module bitwise_not_2(a, b);
  input [1:0] a;
  output [1:0] b;
  assign b = ~a;
endmodule
