//NOTE: no-implementation module stub

module GTECH_MUX4 (
    input wire [1:0] A,
    input wire B,
    input wire D0,
    input wire D1,
    input wire D2,
    input wire D3,
    output wire Z
);

endmodule
