module OptKuznechikEncoder(
  input wire clk,
  input wire [127:0] _block,
  input wire [255:0] key,
  output wire [127:0] out
);
  wire [7:0] arr[256] = '{8'hfc, 8'hee, 8'hdd, 8'h11, 8'hcf, 8'h6e, 8'h31, 8'h16, 8'hfb, 8'hc4, 8'hfa, 8'hda, 8'h23, 8'hc5, 8'h04, 8'h4d, 8'he9, 8'h77, 8'hf0, 8'hdb, 8'h93, 8'h2e, 8'h99, 8'hba, 8'h17, 8'h36, 8'hf1, 8'hbb, 8'h14, 8'hcd, 8'h5f, 8'hc1, 8'hf9, 8'h18, 8'h65, 8'h5a, 8'he2, 8'h5c, 8'hef, 8'h21, 8'h81, 8'h1c, 8'h3c, 8'h42, 8'h8b, 8'h01, 8'h8e, 8'h4f, 8'h05, 8'h84, 8'h02, 8'hae, 8'he3, 8'h6a, 8'h8f, 8'ha0, 8'h06, 8'h0b, 8'hed, 8'h98, 8'h7f, 8'hd4, 8'hd3, 8'h1f, 8'heb, 8'h34, 8'h2c, 8'h51, 8'hea, 8'hc8, 8'h48, 8'hab, 8'hf2, 8'h2a, 8'h68, 8'ha2, 8'hfd, 8'h3a, 8'hce, 8'hcc, 8'hb5, 8'h70, 8'h0e, 8'h56, 8'h08, 8'h0c, 8'h76, 8'h12, 8'hbf, 8'h72, 8'h13, 8'h47, 8'h9c, 8'hb7, 8'h5d, 8'h87, 8'h15, 8'ha1, 8'h96, 8'h29, 8'h10, 8'h7b, 8'h9a, 8'hc7, 8'hf3, 8'h91, 8'h78, 8'h6f, 8'h9d, 8'h9e, 8'hb2, 8'hb1, 8'h32, 8'h75, 8'h19, 8'h3d, 8'hff, 8'h35, 8'h8a, 8'h7e, 8'h6d, 8'h54, 8'hc6, 8'h80, 8'hc3, 8'hbd, 8'h0d, 8'h57, 8'hdf, 8'hf5, 8'h24, 8'ha9, 8'h3e, 8'ha8, 8'h43, 8'hc9, 8'hd7, 8'h79, 8'hd6, 8'hf6, 8'h7c, 8'h22, 8'hb9, 8'h03, 8'he0, 8'h0f, 8'hec, 8'hde, 8'h7a, 8'h94, 8'hb0, 8'hbc, 8'hdc, 8'he8, 8'h28, 8'h50, 8'h4e, 8'h33, 8'h0a, 8'h4a, 8'ha7, 8'h97, 8'h60, 8'h73, 8'h1e, 8'h00, 8'h62, 8'h44, 8'h1a, 8'hb8, 8'h38, 8'h82, 8'h64, 8'h9f, 8'h26, 8'h41, 8'had, 8'h45, 8'h46, 8'h92, 8'h27, 8'h5e, 8'h55, 8'h2f, 8'h8c, 8'ha3, 8'ha5, 8'h7d, 8'h69, 8'hd5, 8'h95, 8'h3b, 8'h07, 8'h58, 8'hb3, 8'h40, 8'h86, 8'hac, 8'h1d, 8'hf7, 8'h30, 8'h37, 8'h6b, 8'he4, 8'h88, 8'hd9, 8'he7, 8'h89, 8'he1, 8'h1b, 8'h83, 8'h49, 8'h4c, 8'h3f, 8'hf8, 8'hfe, 8'h8d, 8'h53, 8'haa, 8'h90, 8'hca, 8'hd8, 8'h85, 8'h61, 8'h20, 8'h71, 8'h67, 8'ha4, 8'h2d, 8'h2b, 8'h09, 8'h5b, 8'hcb, 8'h9b, 8'h25, 8'hd0, 8'hbe, 8'he5, 8'h6c, 8'h52, 8'h59, 8'ha6, 8'h74, 8'hd2, 8'he6, 8'hf4, 8'hb4, 8'hc0, 8'hd1, 8'h66, 8'haf, 8'hc2, 8'h39, 8'h4b, 8'h63, 8'hb6};
  wire [7:0] literal_1076345[256] = '{8'h00, 8'h94, 8'heb, 8'h7f, 8'h15, 8'h81, 8'hfe, 8'h6a, 8'h2a, 8'hbe, 8'hc1, 8'h55, 8'h3f, 8'hab, 8'hd4, 8'h40, 8'h54, 8'hc0, 8'hbf, 8'h2b, 8'h41, 8'hd5, 8'haa, 8'h3e, 8'h7e, 8'hea, 8'h95, 8'h01, 8'h6b, 8'hff, 8'h80, 8'h14, 8'ha8, 8'h3c, 8'h43, 8'hd7, 8'hbd, 8'h29, 8'h56, 8'hc2, 8'h82, 8'h16, 8'h69, 8'hfd, 8'h97, 8'h03, 8'h7c, 8'he8, 8'hfc, 8'h68, 8'h17, 8'h83, 8'he9, 8'h7d, 8'h02, 8'h96, 8'hd6, 8'h42, 8'h3d, 8'ha9, 8'hc3, 8'h57, 8'h28, 8'hbc, 8'h93, 8'h07, 8'h78, 8'hec, 8'h86, 8'h12, 8'h6d, 8'hf9, 8'hb9, 8'h2d, 8'h52, 8'hc6, 8'hac, 8'h38, 8'h47, 8'hd3, 8'hc7, 8'h53, 8'h2c, 8'hb8, 8'hd2, 8'h46, 8'h39, 8'had, 8'hed, 8'h79, 8'h06, 8'h92, 8'hf8, 8'h6c, 8'h13, 8'h87, 8'h3b, 8'haf, 8'hd0, 8'h44, 8'h2e, 8'hba, 8'hc5, 8'h51, 8'h11, 8'h85, 8'hfa, 8'h6e, 8'h04, 8'h90, 8'hef, 8'h7b, 8'h6f, 8'hfb, 8'h84, 8'h10, 8'h7a, 8'hee, 8'h91, 8'h05, 8'h45, 8'hd1, 8'hae, 8'h3a, 8'h50, 8'hc4, 8'hbb, 8'h2f, 8'he5, 8'h71, 8'h0e, 8'h9a, 8'hf0, 8'h64, 8'h1b, 8'h8f, 8'hcf, 8'h5b, 8'h24, 8'hb0, 8'hda, 8'h4e, 8'h31, 8'ha5, 8'hb1, 8'h25, 8'h5a, 8'hce, 8'ha4, 8'h30, 8'h4f, 8'hdb, 8'h9b, 8'h0f, 8'h70, 8'he4, 8'h8e, 8'h1a, 8'h65, 8'hf1, 8'h4d, 8'hd9, 8'ha6, 8'h32, 8'h58, 8'hcc, 8'hb3, 8'h27, 8'h67, 8'hf3, 8'h8c, 8'h18, 8'h72, 8'he6, 8'h99, 8'h0d, 8'h19, 8'h8d, 8'hf2, 8'h66, 8'h0c, 8'h98, 8'he7, 8'h73, 8'h33, 8'ha7, 8'hd8, 8'h4c, 8'h26, 8'hb2, 8'hcd, 8'h59, 8'h76, 8'he2, 8'h9d, 8'h09, 8'h63, 8'hf7, 8'h88, 8'h1c, 8'h5c, 8'hc8, 8'hb7, 8'h23, 8'h49, 8'hdd, 8'ha2, 8'h36, 8'h22, 8'hb6, 8'hc9, 8'h5d, 8'h37, 8'ha3, 8'hdc, 8'h48, 8'h08, 8'h9c, 8'he3, 8'h77, 8'h1d, 8'h89, 8'hf6, 8'h62, 8'hde, 8'h4a, 8'h35, 8'ha1, 8'hcb, 8'h5f, 8'h20, 8'hb4, 8'hf4, 8'h60, 8'h1f, 8'h8b, 8'he1, 8'h75, 8'h0a, 8'h9e, 8'h8a, 8'h1e, 8'h61, 8'hf5, 8'h9f, 8'h0b, 8'h74, 8'he0, 8'ha0, 8'h34, 8'h4b, 8'hdf, 8'hb5, 8'h21, 8'h5e, 8'hca};
  wire [7:0] literal_1076347[256] = '{8'h00, 8'h20, 8'h40, 8'h60, 8'h80, 8'ha0, 8'hc0, 8'he0, 8'hc3, 8'he3, 8'h83, 8'ha3, 8'h43, 8'h63, 8'h03, 8'h23, 8'h45, 8'h65, 8'h05, 8'h25, 8'hc5, 8'he5, 8'h85, 8'ha5, 8'h86, 8'ha6, 8'hc6, 8'he6, 8'h06, 8'h26, 8'h46, 8'h66, 8'h8a, 8'haa, 8'hca, 8'hea, 8'h0a, 8'h2a, 8'h4a, 8'h6a, 8'h49, 8'h69, 8'h09, 8'h29, 8'hc9, 8'he9, 8'h89, 8'ha9, 8'hcf, 8'hef, 8'h8f, 8'haf, 8'h4f, 8'h6f, 8'h0f, 8'h2f, 8'h0c, 8'h2c, 8'h4c, 8'h6c, 8'h8c, 8'hac, 8'hcc, 8'hec, 8'hd7, 8'hf7, 8'h97, 8'hb7, 8'h57, 8'h77, 8'h17, 8'h37, 8'h14, 8'h34, 8'h54, 8'h74, 8'h94, 8'hb4, 8'hd4, 8'hf4, 8'h92, 8'hb2, 8'hd2, 8'hf2, 8'h12, 8'h32, 8'h52, 8'h72, 8'h51, 8'h71, 8'h11, 8'h31, 8'hd1, 8'hf1, 8'h91, 8'hb1, 8'h5d, 8'h7d, 8'h1d, 8'h3d, 8'hdd, 8'hfd, 8'h9d, 8'hbd, 8'h9e, 8'hbe, 8'hde, 8'hfe, 8'h1e, 8'h3e, 8'h5e, 8'h7e, 8'h18, 8'h38, 8'h58, 8'h78, 8'h98, 8'hb8, 8'hd8, 8'hf8, 8'hdb, 8'hfb, 8'h9b, 8'hbb, 8'h5b, 8'h7b, 8'h1b, 8'h3b, 8'h6d, 8'h4d, 8'h2d, 8'h0d, 8'hed, 8'hcd, 8'had, 8'h8d, 8'hae, 8'h8e, 8'hee, 8'hce, 8'h2e, 8'h0e, 8'h6e, 8'h4e, 8'h28, 8'h08, 8'h68, 8'h48, 8'ha8, 8'h88, 8'he8, 8'hc8, 8'heb, 8'hcb, 8'hab, 8'h8b, 8'h6b, 8'h4b, 8'h2b, 8'h0b, 8'he7, 8'hc7, 8'ha7, 8'h87, 8'h67, 8'h47, 8'h27, 8'h07, 8'h24, 8'h04, 8'h64, 8'h44, 8'ha4, 8'h84, 8'he4, 8'hc4, 8'ha2, 8'h82, 8'he2, 8'hc2, 8'h22, 8'h02, 8'h62, 8'h42, 8'h61, 8'h41, 8'h21, 8'h01, 8'he1, 8'hc1, 8'ha1, 8'h81, 8'hba, 8'h9a, 8'hfa, 8'hda, 8'h3a, 8'h1a, 8'h7a, 8'h5a, 8'h79, 8'h59, 8'h39, 8'h19, 8'hf9, 8'hd9, 8'hb9, 8'h99, 8'hff, 8'hdf, 8'hbf, 8'h9f, 8'h7f, 8'h5f, 8'h3f, 8'h1f, 8'h3c, 8'h1c, 8'h7c, 8'h5c, 8'hbc, 8'h9c, 8'hfc, 8'hdc, 8'h30, 8'h10, 8'h70, 8'h50, 8'hb0, 8'h90, 8'hf0, 8'hd0, 8'hf3, 8'hd3, 8'hb3, 8'h93, 8'h73, 8'h53, 8'h33, 8'h13, 8'h75, 8'h55, 8'h35, 8'h15, 8'hf5, 8'hd5, 8'hb5, 8'h95, 8'hb6, 8'h96, 8'hf6, 8'hd6, 8'h36, 8'h16, 8'h76, 8'h56};
  wire [7:0] literal_1076349[256] = '{8'h00, 8'h85, 8'hc9, 8'h4c, 8'h51, 8'hd4, 8'h98, 8'h1d, 8'ha2, 8'h27, 8'h6b, 8'hee, 8'hf3, 8'h76, 8'h3a, 8'hbf, 8'h87, 8'h02, 8'h4e, 8'hcb, 8'hd6, 8'h53, 8'h1f, 8'h9a, 8'h25, 8'ha0, 8'hec, 8'h69, 8'h74, 8'hf1, 8'hbd, 8'h38, 8'hcd, 8'h48, 8'h04, 8'h81, 8'h9c, 8'h19, 8'h55, 8'hd0, 8'h6f, 8'hea, 8'ha6, 8'h23, 8'h3e, 8'hbb, 8'hf7, 8'h72, 8'h4a, 8'hcf, 8'h83, 8'h06, 8'h1b, 8'h9e, 8'hd2, 8'h57, 8'he8, 8'h6d, 8'h21, 8'ha4, 8'hb9, 8'h3c, 8'h70, 8'hf5, 8'h59, 8'hdc, 8'h90, 8'h15, 8'h08, 8'h8d, 8'hc1, 8'h44, 8'hfb, 8'h7e, 8'h32, 8'hb7, 8'haa, 8'h2f, 8'h63, 8'he6, 8'hde, 8'h5b, 8'h17, 8'h92, 8'h8f, 8'h0a, 8'h46, 8'hc3, 8'h7c, 8'hf9, 8'hb5, 8'h30, 8'h2d, 8'ha8, 8'he4, 8'h61, 8'h94, 8'h11, 8'h5d, 8'hd8, 8'hc5, 8'h40, 8'h0c, 8'h89, 8'h36, 8'hb3, 8'hff, 8'h7a, 8'h67, 8'he2, 8'hae, 8'h2b, 8'h13, 8'h96, 8'hda, 8'h5f, 8'h42, 8'hc7, 8'h8b, 8'h0e, 8'hb1, 8'h34, 8'h78, 8'hfd, 8'he0, 8'h65, 8'h29, 8'hac, 8'hb2, 8'h37, 8'h7b, 8'hfe, 8'he3, 8'h66, 8'h2a, 8'haf, 8'h10, 8'h95, 8'hd9, 8'h5c, 8'h41, 8'hc4, 8'h88, 8'h0d, 8'h35, 8'hb0, 8'hfc, 8'h79, 8'h64, 8'he1, 8'had, 8'h28, 8'h97, 8'h12, 8'h5e, 8'hdb, 8'hc6, 8'h43, 8'h0f, 8'h8a, 8'h7f, 8'hfa, 8'hb6, 8'h33, 8'h2e, 8'hab, 8'he7, 8'h62, 8'hdd, 8'h58, 8'h14, 8'h91, 8'h8c, 8'h09, 8'h45, 8'hc0, 8'hf8, 8'h7d, 8'h31, 8'hb4, 8'ha9, 8'h2c, 8'h60, 8'he5, 8'h5a, 8'hdf, 8'h93, 8'h16, 8'h0b, 8'h8e, 8'hc2, 8'h47, 8'heb, 8'h6e, 8'h22, 8'ha7, 8'hba, 8'h3f, 8'h73, 8'hf6, 8'h49, 8'hcc, 8'h80, 8'h05, 8'h18, 8'h9d, 8'hd1, 8'h54, 8'h6c, 8'he9, 8'ha5, 8'h20, 8'h3d, 8'hb8, 8'hf4, 8'h71, 8'hce, 8'h4b, 8'h07, 8'h82, 8'h9f, 8'h1a, 8'h56, 8'hd3, 8'h26, 8'ha3, 8'hef, 8'h6a, 8'h77, 8'hf2, 8'hbe, 8'h3b, 8'h84, 8'h01, 8'h4d, 8'hc8, 8'hd5, 8'h50, 8'h1c, 8'h99, 8'ha1, 8'h24, 8'h68, 8'hed, 8'hf0, 8'h75, 8'h39, 8'hbc, 8'h03, 8'h86, 8'hca, 8'h4f, 8'h52, 8'hd7, 8'h9b, 8'h1e};
  wire [7:0] literal_1076351[256] = '{8'h00, 8'h10, 8'h20, 8'h30, 8'h40, 8'h50, 8'h60, 8'h70, 8'h80, 8'h90, 8'ha0, 8'hb0, 8'hc0, 8'hd0, 8'he0, 8'hf0, 8'hc3, 8'hd3, 8'he3, 8'hf3, 8'h83, 8'h93, 8'ha3, 8'hb3, 8'h43, 8'h53, 8'h63, 8'h73, 8'h03, 8'h13, 8'h23, 8'h33, 8'h45, 8'h55, 8'h65, 8'h75, 8'h05, 8'h15, 8'h25, 8'h35, 8'hc5, 8'hd5, 8'he5, 8'hf5, 8'h85, 8'h95, 8'ha5, 8'hb5, 8'h86, 8'h96, 8'ha6, 8'hb6, 8'hc6, 8'hd6, 8'he6, 8'hf6, 8'h06, 8'h16, 8'h26, 8'h36, 8'h46, 8'h56, 8'h66, 8'h76, 8'h8a, 8'h9a, 8'haa, 8'hba, 8'hca, 8'hda, 8'hea, 8'hfa, 8'h0a, 8'h1a, 8'h2a, 8'h3a, 8'h4a, 8'h5a, 8'h6a, 8'h7a, 8'h49, 8'h59, 8'h69, 8'h79, 8'h09, 8'h19, 8'h29, 8'h39, 8'hc9, 8'hd9, 8'he9, 8'hf9, 8'h89, 8'h99, 8'ha9, 8'hb9, 8'hcf, 8'hdf, 8'hef, 8'hff, 8'h8f, 8'h9f, 8'haf, 8'hbf, 8'h4f, 8'h5f, 8'h6f, 8'h7f, 8'h0f, 8'h1f, 8'h2f, 8'h3f, 8'h0c, 8'h1c, 8'h2c, 8'h3c, 8'h4c, 8'h5c, 8'h6c, 8'h7c, 8'h8c, 8'h9c, 8'hac, 8'hbc, 8'hcc, 8'hdc, 8'hec, 8'hfc, 8'hd7, 8'hc7, 8'hf7, 8'he7, 8'h97, 8'h87, 8'hb7, 8'ha7, 8'h57, 8'h47, 8'h77, 8'h67, 8'h17, 8'h07, 8'h37, 8'h27, 8'h14, 8'h04, 8'h34, 8'h24, 8'h54, 8'h44, 8'h74, 8'h64, 8'h94, 8'h84, 8'hb4, 8'ha4, 8'hd4, 8'hc4, 8'hf4, 8'he4, 8'h92, 8'h82, 8'hb2, 8'ha2, 8'hd2, 8'hc2, 8'hf2, 8'he2, 8'h12, 8'h02, 8'h32, 8'h22, 8'h52, 8'h42, 8'h72, 8'h62, 8'h51, 8'h41, 8'h71, 8'h61, 8'h11, 8'h01, 8'h31, 8'h21, 8'hd1, 8'hc1, 8'hf1, 8'he1, 8'h91, 8'h81, 8'hb1, 8'ha1, 8'h5d, 8'h4d, 8'h7d, 8'h6d, 8'h1d, 8'h0d, 8'h3d, 8'h2d, 8'hdd, 8'hcd, 8'hfd, 8'hed, 8'h9d, 8'h8d, 8'hbd, 8'had, 8'h9e, 8'h8e, 8'hbe, 8'hae, 8'hde, 8'hce, 8'hfe, 8'hee, 8'h1e, 8'h0e, 8'h3e, 8'h2e, 8'h5e, 8'h4e, 8'h7e, 8'h6e, 8'h18, 8'h08, 8'h38, 8'h28, 8'h58, 8'h48, 8'h78, 8'h68, 8'h98, 8'h88, 8'hb8, 8'ha8, 8'hd8, 8'hc8, 8'hf8, 8'he8, 8'hdb, 8'hcb, 8'hfb, 8'heb, 8'h9b, 8'h8b, 8'hbb, 8'hab, 8'h5b, 8'h4b, 8'h7b, 8'h6b, 8'h1b, 8'h0b, 8'h3b, 8'h2b};
  wire [7:0] literal_1076353[256] = '{8'h00, 8'hc2, 8'h47, 8'h85, 8'h8e, 8'h4c, 8'hc9, 8'h0b, 8'hdf, 8'h1d, 8'h98, 8'h5a, 8'h51, 8'h93, 8'h16, 8'hd4, 8'h7d, 8'hbf, 8'h3a, 8'hf8, 8'hf3, 8'h31, 8'hb4, 8'h76, 8'ha2, 8'h60, 8'he5, 8'h27, 8'h2c, 8'hee, 8'h6b, 8'ha9, 8'hfa, 8'h38, 8'hbd, 8'h7f, 8'h74, 8'hb6, 8'h33, 8'hf1, 8'h25, 8'he7, 8'h62, 8'ha0, 8'hab, 8'h69, 8'hec, 8'h2e, 8'h87, 8'h45, 8'hc0, 8'h02, 8'h09, 8'hcb, 8'h4e, 8'h8c, 8'h58, 8'h9a, 8'h1f, 8'hdd, 8'hd6, 8'h14, 8'h91, 8'h53, 8'h37, 8'hf5, 8'h70, 8'hb2, 8'hb9, 8'h7b, 8'hfe, 8'h3c, 8'he8, 8'h2a, 8'haf, 8'h6d, 8'h66, 8'ha4, 8'h21, 8'he3, 8'h4a, 8'h88, 8'h0d, 8'hcf, 8'hc4, 8'h06, 8'h83, 8'h41, 8'h95, 8'h57, 8'hd2, 8'h10, 8'h1b, 8'hd9, 8'h5c, 8'h9e, 8'hcd, 8'h0f, 8'h8a, 8'h48, 8'h43, 8'h81, 8'h04, 8'hc6, 8'h12, 8'hd0, 8'h55, 8'h97, 8'h9c, 8'h5e, 8'hdb, 8'h19, 8'hb0, 8'h72, 8'hf7, 8'h35, 8'h3e, 8'hfc, 8'h79, 8'hbb, 8'h6f, 8'had, 8'h28, 8'hea, 8'he1, 8'h23, 8'ha6, 8'h64, 8'h6e, 8'hac, 8'h29, 8'heb, 8'he0, 8'h22, 8'ha7, 8'h65, 8'hb1, 8'h73, 8'hf6, 8'h34, 8'h3f, 8'hfd, 8'h78, 8'hba, 8'h13, 8'hd1, 8'h54, 8'h96, 8'h9d, 8'h5f, 8'hda, 8'h18, 8'hcc, 8'h0e, 8'h8b, 8'h49, 8'h42, 8'h80, 8'h05, 8'hc7, 8'h94, 8'h56, 8'hd3, 8'h11, 8'h1a, 8'hd8, 8'h5d, 8'h9f, 8'h4b, 8'h89, 8'h0c, 8'hce, 8'hc5, 8'h07, 8'h82, 8'h40, 8'he9, 8'h2b, 8'hae, 8'h6c, 8'h67, 8'ha5, 8'h20, 8'he2, 8'h36, 8'hf4, 8'h71, 8'hb3, 8'hb8, 8'h7a, 8'hff, 8'h3d, 8'h59, 8'h9b, 8'h1e, 8'hdc, 8'hd7, 8'h15, 8'h90, 8'h52, 8'h86, 8'h44, 8'hc1, 8'h03, 8'h08, 8'hca, 8'h4f, 8'h8d, 8'h24, 8'he6, 8'h63, 8'ha1, 8'haa, 8'h68, 8'hed, 8'h2f, 8'hfb, 8'h39, 8'hbc, 8'h7e, 8'h75, 8'hb7, 8'h32, 8'hf0, 8'ha3, 8'h61, 8'he4, 8'h26, 8'h2d, 8'hef, 8'h6a, 8'ha8, 8'h7c, 8'hbe, 8'h3b, 8'hf9, 8'hf2, 8'h30, 8'hb5, 8'h77, 8'hde, 8'h1c, 8'h99, 8'h5b, 8'h50, 8'h92, 8'h17, 8'hd5, 8'h01, 8'hc3, 8'h46, 8'h84, 8'h8f, 8'h4d, 8'hc8, 8'h0a};
  wire [7:0] literal_1076355[256] = '{8'h00, 8'hc0, 8'h43, 8'h83, 8'h86, 8'h46, 8'hc5, 8'h05, 8'hcf, 8'h0f, 8'h8c, 8'h4c, 8'h49, 8'h89, 8'h0a, 8'hca, 8'h5d, 8'h9d, 8'h1e, 8'hde, 8'hdb, 8'h1b, 8'h98, 8'h58, 8'h92, 8'h52, 8'hd1, 8'h11, 8'h14, 8'hd4, 8'h57, 8'h97, 8'hba, 8'h7a, 8'hf9, 8'h39, 8'h3c, 8'hfc, 8'h7f, 8'hbf, 8'h75, 8'hb5, 8'h36, 8'hf6, 8'hf3, 8'h33, 8'hb0, 8'h70, 8'he7, 8'h27, 8'ha4, 8'h64, 8'h61, 8'ha1, 8'h22, 8'he2, 8'h28, 8'he8, 8'h6b, 8'hab, 8'hae, 8'h6e, 8'hed, 8'h2d, 8'hb7, 8'h77, 8'hf4, 8'h34, 8'h31, 8'hf1, 8'h72, 8'hb2, 8'h78, 8'hb8, 8'h3b, 8'hfb, 8'hfe, 8'h3e, 8'hbd, 8'h7d, 8'hea, 8'h2a, 8'ha9, 8'h69, 8'h6c, 8'hac, 8'h2f, 8'hef, 8'h25, 8'he5, 8'h66, 8'ha6, 8'ha3, 8'h63, 8'he0, 8'h20, 8'h0d, 8'hcd, 8'h4e, 8'h8e, 8'h8b, 8'h4b, 8'hc8, 8'h08, 8'hc2, 8'h02, 8'h81, 8'h41, 8'h44, 8'h84, 8'h07, 8'hc7, 8'h50, 8'h90, 8'h13, 8'hd3, 8'hd6, 8'h16, 8'h95, 8'h55, 8'h9f, 8'h5f, 8'hdc, 8'h1c, 8'h19, 8'hd9, 8'h5a, 8'h9a, 8'had, 8'h6d, 8'hee, 8'h2e, 8'h2b, 8'heb, 8'h68, 8'ha8, 8'h62, 8'ha2, 8'h21, 8'he1, 8'he4, 8'h24, 8'ha7, 8'h67, 8'hf0, 8'h30, 8'hb3, 8'h73, 8'h76, 8'hb6, 8'h35, 8'hf5, 8'h3f, 8'hff, 8'h7c, 8'hbc, 8'hb9, 8'h79, 8'hfa, 8'h3a, 8'h17, 8'hd7, 8'h54, 8'h94, 8'h91, 8'h51, 8'hd2, 8'h12, 8'hd8, 8'h18, 8'h9b, 8'h5b, 8'h5e, 8'h9e, 8'h1d, 8'hdd, 8'h4a, 8'h8a, 8'h09, 8'hc9, 8'hcc, 8'h0c, 8'h8f, 8'h4f, 8'h85, 8'h45, 8'hc6, 8'h06, 8'h03, 8'hc3, 8'h40, 8'h80, 8'h1a, 8'hda, 8'h59, 8'h99, 8'h9c, 8'h5c, 8'hdf, 8'h1f, 8'hd5, 8'h15, 8'h96, 8'h56, 8'h53, 8'h93, 8'h10, 8'hd0, 8'h47, 8'h87, 8'h04, 8'hc4, 8'hc1, 8'h01, 8'h82, 8'h42, 8'h88, 8'h48, 8'hcb, 8'h0b, 8'h0e, 8'hce, 8'h4d, 8'h8d, 8'ha0, 8'h60, 8'he3, 8'h23, 8'h26, 8'he6, 8'h65, 8'ha5, 8'h6f, 8'haf, 8'h2c, 8'hec, 8'he9, 8'h29, 8'haa, 8'h6a, 8'hfd, 8'h3d, 8'hbe, 8'h7e, 8'h7b, 8'hbb, 8'h38, 8'hf8, 8'h32, 8'hf2, 8'h71, 8'hb1, 8'hb4, 8'h74, 8'hf7, 8'h37};
  wire [7:0] literal_1076358[256] = '{8'h00, 8'hfb, 8'h35, 8'hce, 8'h6a, 8'h91, 8'h5f, 8'ha4, 8'hd4, 8'h2f, 8'he1, 8'h1a, 8'hbe, 8'h45, 8'h8b, 8'h70, 8'h6b, 8'h90, 8'h5e, 8'ha5, 8'h01, 8'hfa, 8'h34, 8'hcf, 8'hbf, 8'h44, 8'h8a, 8'h71, 8'hd5, 8'h2e, 8'he0, 8'h1b, 8'hd6, 8'h2d, 8'he3, 8'h18, 8'hbc, 8'h47, 8'h89, 8'h72, 8'h02, 8'hf9, 8'h37, 8'hcc, 8'h68, 8'h93, 8'h5d, 8'ha6, 8'hbd, 8'h46, 8'h88, 8'h73, 8'hd7, 8'h2c, 8'he2, 8'h19, 8'h69, 8'h92, 8'h5c, 8'ha7, 8'h03, 8'hf8, 8'h36, 8'hcd, 8'h6f, 8'h94, 8'h5a, 8'ha1, 8'h05, 8'hfe, 8'h30, 8'hcb, 8'hbb, 8'h40, 8'h8e, 8'h75, 8'hd1, 8'h2a, 8'he4, 8'h1f, 8'h04, 8'hff, 8'h31, 8'hca, 8'h6e, 8'h95, 8'h5b, 8'ha0, 8'hd0, 8'h2b, 8'he5, 8'h1e, 8'hba, 8'h41, 8'h8f, 8'h74, 8'hb9, 8'h42, 8'h8c, 8'h77, 8'hd3, 8'h28, 8'he6, 8'h1d, 8'h6d, 8'h96, 8'h58, 8'ha3, 8'h07, 8'hfc, 8'h32, 8'hc9, 8'hd2, 8'h29, 8'he7, 8'h1c, 8'hb8, 8'h43, 8'h8d, 8'h76, 8'h06, 8'hfd, 8'h33, 8'hc8, 8'h6c, 8'h97, 8'h59, 8'ha2, 8'hde, 8'h25, 8'heb, 8'h10, 8'hb4, 8'h4f, 8'h81, 8'h7a, 8'h0a, 8'hf1, 8'h3f, 8'hc4, 8'h60, 8'h9b, 8'h55, 8'hae, 8'hb5, 8'h4e, 8'h80, 8'h7b, 8'hdf, 8'h24, 8'hea, 8'h11, 8'h61, 8'h9a, 8'h54, 8'haf, 8'h0b, 8'hf0, 8'h3e, 8'hc5, 8'h08, 8'hf3, 8'h3d, 8'hc6, 8'h62, 8'h99, 8'h57, 8'hac, 8'hdc, 8'h27, 8'he9, 8'h12, 8'hb6, 8'h4d, 8'h83, 8'h78, 8'h63, 8'h98, 8'h56, 8'had, 8'h09, 8'hf2, 8'h3c, 8'hc7, 8'hb7, 8'h4c, 8'h82, 8'h79, 8'hdd, 8'h26, 8'he8, 8'h13, 8'hb1, 8'h4a, 8'h84, 8'h7f, 8'hdb, 8'h20, 8'hee, 8'h15, 8'h65, 8'h9e, 8'h50, 8'hab, 8'h0f, 8'hf4, 8'h3a, 8'hc1, 8'hda, 8'h21, 8'hef, 8'h14, 8'hb0, 8'h4b, 8'h85, 8'h7e, 8'h0e, 8'hf5, 8'h3b, 8'hc0, 8'h64, 8'h9f, 8'h51, 8'haa, 8'h67, 8'h9c, 8'h52, 8'ha9, 8'h0d, 8'hf6, 8'h38, 8'hc3, 8'hb3, 8'h48, 8'h86, 8'h7d, 8'hd9, 8'h22, 8'hec, 8'h17, 8'h0c, 8'hf7, 8'h39, 8'hc2, 8'h66, 8'h9d, 8'h53, 8'ha8, 8'hd8, 8'h23, 8'hed, 8'h16, 8'hb2, 8'h49, 8'h87, 8'h7c};

  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [127:0] p0__block;
  reg [255:0] p0_key;
  reg [7:0] p1_arr[256];
  reg [7:0] p1_literal_1076345[256];
  reg [7:0] p1_literal_1076347[256];
  reg [7:0] p1_literal_1076349[256];
  reg [7:0] p1_literal_1076351[256];
  reg [7:0] p1_literal_1076353[256];
  reg [7:0] p1_literal_1076355[256];
  reg [7:0] p1_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p0__block <= _block;
    p0_key <= key;
    p1_arr <= arr;
    p1_literal_1076345 <= literal_1076345;
    p1_literal_1076347 <= literal_1076347;
    p1_literal_1076349 <= literal_1076349;
    p1_literal_1076351 <= literal_1076351;
    p1_literal_1076353 <= literal_1076353;
    p1_literal_1076355 <= literal_1076355;
    p1_literal_1076358 <= literal_1076358;
  end

  // ===== Pipe stage 1:
  wire [127:0] p1_addedKey__41_comb;
  wire [7:0] p1_array_index_1076346_comb;
  wire [7:0] p1_array_index_1076348_comb;
  wire [7:0] p1_array_index_1076350_comb;
  wire [7:0] p1_array_index_1076352_comb;
  wire [7:0] p1_array_index_1076354_comb;
  wire [7:0] p1_array_index_1076356_comb;
  wire [7:0] p1_array_index_1076359_comb;
  wire [7:0] p1_array_index_1076361_comb;
  wire [7:0] p1_array_index_1076362_comb;
  wire [7:0] p1_array_index_1076363_comb;
  wire [7:0] p1_array_index_1076364_comb;
  wire [7:0] p1_array_index_1076365_comb;
  wire [7:0] p1_array_index_1076366_comb;
  wire [7:0] p1_array_index_1076368_comb;
  wire [7:0] p1_array_index_1076369_comb;
  wire [7:0] p1_array_index_1076370_comb;
  wire [7:0] p1_array_index_1076371_comb;
  wire [7:0] p1_array_index_1076372_comb;
  wire [7:0] p1_array_index_1076373_comb;
  wire [7:0] p1_array_index_1076374_comb;
  wire [7:0] p1_array_index_1076376_comb;
  wire [7:0] p1_res7_comb;
  wire [7:0] p1_array_index_1076385_comb;
  wire [7:0] p1_array_index_1076386_comb;
  wire [7:0] p1_array_index_1076387_comb;
  wire [7:0] p1_array_index_1076388_comb;
  wire [7:0] p1_array_index_1076389_comb;
  wire [7:0] p1_array_index_1076390_comb;
  wire [7:0] p1_res7__1_comb;
  wire [7:0] p1_array_index_1076400_comb;
  wire [7:0] p1_array_index_1076401_comb;
  wire [7:0] p1_array_index_1076402_comb;
  wire [7:0] p1_array_index_1076403_comb;
  wire [7:0] p1_array_index_1076404_comb;
  wire [7:0] p1_res7__2_comb;
  wire [7:0] p1_array_index_1076414_comb;
  wire [7:0] p1_array_index_1076415_comb;
  wire [7:0] p1_array_index_1076416_comb;
  wire [7:0] p1_array_index_1076417_comb;
  wire [7:0] p1_array_index_1076418_comb;
  wire [7:0] p1_res7__3_comb;
  wire [7:0] p1_array_index_1076429_comb;
  wire [7:0] p1_array_index_1076430_comb;
  wire [7:0] p1_array_index_1076431_comb;
  wire [7:0] p1_array_index_1076432_comb;
  wire [7:0] p1_res7__4_comb;
  wire [7:0] p1_array_index_1076442_comb;
  wire [7:0] p1_array_index_1076443_comb;
  wire [7:0] p1_array_index_1076444_comb;
  wire [7:0] p1_array_index_1076445_comb;
  wire [7:0] p1_res7__5_comb;
  wire [7:0] p1_array_index_1076456_comb;
  wire [7:0] p1_array_index_1076457_comb;
  wire [7:0] p1_array_index_1076458_comb;
  wire [7:0] p1_res7__6_comb;
  wire [7:0] p1_array_index_1076468_comb;
  wire [7:0] p1_array_index_1076469_comb;
  wire [7:0] p1_array_index_1076470_comb;
  wire [7:0] p1_res7__7_comb;
  wire [7:0] p1_array_index_1076481_comb;
  wire [7:0] p1_array_index_1076482_comb;
  wire [7:0] p1_res7__8_comb;
  wire [7:0] p1_array_index_1076492_comb;
  wire [7:0] p1_array_index_1076493_comb;
  wire [7:0] p1_res7__9_comb;
  wire [7:0] p1_array_index_1076504_comb;
  wire [7:0] p1_res7__10_comb;
  wire [7:0] p1_array_index_1076514_comb;
  wire [7:0] p1_res7__11_comb;
  wire [7:0] p1_res7__12_comb;
  wire [7:0] p1_res7__13_comb;
  wire [7:0] p1_res7__14_comb;
  wire [7:0] p1_res7__15_comb;
  wire [127:0] p1_res_comb;
  wire [127:0] p1_xor_1076555_comb;
  wire [127:0] p1_addedKey__42_comb;
  wire [7:0] p1_array_index_1076571_comb;
  wire [7:0] p1_array_index_1076572_comb;
  wire [7:0] p1_array_index_1076573_comb;
  wire [7:0] p1_array_index_1076574_comb;
  wire [7:0] p1_array_index_1076575_comb;
  wire [7:0] p1_array_index_1076576_comb;
  wire [7:0] p1_array_index_1076578_comb;
  wire [7:0] p1_array_index_1076580_comb;
  wire [7:0] p1_array_index_1076581_comb;
  wire [7:0] p1_array_index_1076582_comb;
  wire [7:0] p1_array_index_1076583_comb;
  wire [7:0] p1_array_index_1076584_comb;
  wire [7:0] p1_array_index_1076585_comb;
  wire [7:0] p1_array_index_1076587_comb;
  wire [7:0] p1_array_index_1076588_comb;
  wire [7:0] p1_array_index_1076589_comb;
  wire [7:0] p1_array_index_1076590_comb;
  wire [7:0] p1_array_index_1076591_comb;
  wire [7:0] p1_array_index_1076592_comb;
  wire [7:0] p1_array_index_1076593_comb;
  wire [7:0] p1_array_index_1076595_comb;
  wire [7:0] p1_res7__16_comb;
  wire [7:0] p1_array_index_1076604_comb;
  wire [7:0] p1_array_index_1076605_comb;
  wire [7:0] p1_array_index_1076606_comb;
  wire [7:0] p1_array_index_1076607_comb;
  wire [7:0] p1_array_index_1076608_comb;
  wire [7:0] p1_array_index_1076609_comb;
  wire [7:0] p1_res7__17_comb;
  wire [7:0] p1_array_index_1076619_comb;
  wire [7:0] p1_array_index_1076620_comb;
  wire [7:0] p1_array_index_1076621_comb;
  wire [7:0] p1_array_index_1076622_comb;
  wire [7:0] p1_array_index_1076623_comb;
  wire [7:0] p1_res7__18_comb;
  wire [7:0] p1_array_index_1076633_comb;
  wire [7:0] p1_array_index_1076634_comb;
  wire [7:0] p1_array_index_1076635_comb;
  wire [7:0] p1_array_index_1076636_comb;
  wire [7:0] p1_array_index_1076637_comb;
  wire [7:0] p1_res7__19_comb;
  wire [7:0] p1_array_index_1076648_comb;
  wire [7:0] p1_array_index_1076649_comb;
  wire [7:0] p1_array_index_1076650_comb;
  wire [7:0] p1_array_index_1076651_comb;
  wire [7:0] p1_res7__20_comb;
  wire [7:0] p1_array_index_1076661_comb;
  wire [7:0] p1_array_index_1076662_comb;
  wire [7:0] p1_array_index_1076663_comb;
  wire [7:0] p1_array_index_1076664_comb;
  wire [7:0] p1_res7__21_comb;
  wire [7:0] p1_array_index_1076675_comb;
  wire [7:0] p1_array_index_1076676_comb;
  wire [7:0] p1_array_index_1076677_comb;
  wire [7:0] p1_res7__22_comb;
  wire [7:0] p1_array_index_1076687_comb;
  wire [7:0] p1_array_index_1076688_comb;
  wire [7:0] p1_array_index_1076689_comb;
  wire [7:0] p1_res7__23_comb;
  wire [7:0] p1_array_index_1076700_comb;
  wire [7:0] p1_array_index_1076701_comb;
  wire [7:0] p1_res7__24_comb;
  wire [7:0] p1_array_index_1076711_comb;
  wire [7:0] p1_array_index_1076712_comb;
  wire [7:0] p1_res7__25_comb;
  wire [7:0] p1_array_index_1076723_comb;
  wire [7:0] p1_res7__26_comb;
  wire [7:0] p1_array_index_1076733_comb;
  wire [7:0] p1_res7__27_comb;
  wire [127:0] p1_addedKey__32_comb;
  wire [7:0] p1_res7__28_comb;
  wire [7:0] p1_array_index_1077177_comb;
  wire [7:0] p1_array_index_1077178_comb;
  wire [7:0] p1_array_index_1077179_comb;
  wire [7:0] p1_array_index_1077180_comb;
  wire [7:0] p1_array_index_1077181_comb;
  wire [7:0] p1_array_index_1077182_comb;
  wire [7:0] p1_array_index_1077184_comb;
  wire [7:0] p1_array_index_1077186_comb;
  wire [7:0] p1_array_index_1077187_comb;
  wire [7:0] p1_array_index_1077188_comb;
  wire [7:0] p1_array_index_1077189_comb;
  wire [7:0] p1_array_index_1077190_comb;
  wire [7:0] p1_array_index_1077191_comb;
  wire [7:0] p1_array_index_1077193_comb;
  wire [7:0] p1_array_index_1077194_comb;
  wire [7:0] p1_array_index_1077195_comb;
  wire [7:0] p1_array_index_1077196_comb;
  wire [7:0] p1_array_index_1077197_comb;
  wire [7:0] p1_array_index_1077198_comb;
  wire [7:0] p1_array_index_1077199_comb;
  wire [7:0] p1_array_index_1077201_comb;
  wire [7:0] p1_res7__29_comb;
  wire [7:0] p1_res7__512_comb;
  wire [7:0] p1_array_index_1077210_comb;
  wire [7:0] p1_array_index_1077211_comb;
  wire [7:0] p1_array_index_1077212_comb;
  wire [7:0] p1_array_index_1077213_comb;
  wire [7:0] p1_array_index_1077214_comb;
  wire [7:0] p1_array_index_1077215_comb;
  wire [7:0] p1_res7__30_comb;
  wire [7:0] p1_res7__513_comb;
  wire [7:0] p1_array_index_1077225_comb;
  wire [7:0] p1_array_index_1077226_comb;
  wire [7:0] p1_array_index_1077227_comb;
  wire [7:0] p1_array_index_1077228_comb;
  wire [7:0] p1_array_index_1077229_comb;
  wire [7:0] p1_res7__31_comb;
  wire [7:0] p1_res7__514_comb;
  wire [127:0] p1_res__1_comb;
  wire [7:0] p1_array_index_1077239_comb;
  wire [7:0] p1_array_index_1077240_comb;
  wire [7:0] p1_array_index_1077241_comb;
  wire [7:0] p1_array_index_1077242_comb;
  wire [7:0] p1_array_index_1077243_comb;
  wire [127:0] p1_xor_1076773_comb;
  wire [7:0] p1_res7__515_comb;
  wire [127:0] p1_addedKey__43_comb;
  wire [7:0] p1_array_index_1077254_comb;
  wire [7:0] p1_array_index_1077255_comb;
  wire [7:0] p1_array_index_1077256_comb;
  wire [7:0] p1_array_index_1077257_comb;
  wire [7:0] p1_res7__516_comb;
  wire [7:0] p1_array_index_1076789_comb;
  wire [7:0] p1_array_index_1076790_comb;
  wire [7:0] p1_array_index_1076791_comb;
  wire [7:0] p1_array_index_1076792_comb;
  wire [7:0] p1_array_index_1076793_comb;
  wire [7:0] p1_array_index_1076794_comb;
  wire [7:0] p1_array_index_1076796_comb;
  wire [7:0] p1_array_index_1076798_comb;
  wire [7:0] p1_array_index_1076799_comb;
  wire [7:0] p1_array_index_1076800_comb;
  wire [7:0] p1_array_index_1076801_comb;
  wire [7:0] p1_array_index_1076802_comb;
  wire [7:0] p1_array_index_1076803_comb;
  wire [7:0] p1_array_index_1077267_comb;
  wire [7:0] p1_array_index_1077268_comb;
  wire [7:0] p1_array_index_1077269_comb;
  wire [7:0] p1_array_index_1077270_comb;
  wire [7:0] p1_array_index_1076805_comb;
  wire [7:0] p1_array_index_1076806_comb;
  wire [7:0] p1_array_index_1076807_comb;
  wire [7:0] p1_array_index_1076808_comb;
  wire [7:0] p1_array_index_1076809_comb;
  wire [7:0] p1_array_index_1076810_comb;
  wire [7:0] p1_array_index_1076811_comb;
  wire [7:0] p1_array_index_1076813_comb;
  wire [7:0] p1_res7__517_comb;
  wire [7:0] p1_res7__32_comb;
  wire [7:0] p1_array_index_1077281_comb;
  wire [7:0] p1_array_index_1077282_comb;
  wire [7:0] p1_array_index_1077283_comb;
  wire [7:0] p1_array_index_1076822_comb;
  wire [7:0] p1_array_index_1076823_comb;
  wire [7:0] p1_array_index_1076824_comb;
  wire [7:0] p1_array_index_1076825_comb;
  wire [7:0] p1_array_index_1076826_comb;
  wire [7:0] p1_array_index_1076827_comb;
  wire [7:0] p1_res7__518_comb;
  wire [7:0] p1_res7__33_comb;
  wire [7:0] p1_array_index_1077293_comb;
  wire [7:0] p1_array_index_1077294_comb;
  wire [7:0] p1_array_index_1077295_comb;
  wire [7:0] p1_array_index_1076837_comb;
  wire [7:0] p1_array_index_1076838_comb;
  wire [7:0] p1_array_index_1076839_comb;
  wire [7:0] p1_array_index_1076840_comb;
  wire [7:0] p1_array_index_1076841_comb;
  wire [7:0] p1_res7__519_comb;
  wire [7:0] p1_res7__34_comb;
  wire [7:0] p1_array_index_1077306_comb;
  wire [7:0] p1_array_index_1077307_comb;
  wire [7:0] p1_array_index_1076851_comb;
  wire [7:0] p1_array_index_1076852_comb;
  wire [7:0] p1_array_index_1076853_comb;
  wire [7:0] p1_array_index_1076854_comb;
  wire [7:0] p1_array_index_1076855_comb;
  wire [7:0] p1_res7__520_comb;
  wire [7:0] p1_res7__35_comb;
  wire [7:0] p1_array_index_1077317_comb;
  wire [7:0] p1_array_index_1077318_comb;
  wire [7:0] p1_array_index_1076866_comb;
  wire [7:0] p1_array_index_1076867_comb;
  wire [7:0] p1_array_index_1076868_comb;
  wire [7:0] p1_array_index_1076869_comb;
  wire [7:0] p1_res7__521_comb;
  wire [7:0] p1_res7__36_comb;
  wire [7:0] p1_array_index_1077329_comb;
  wire [7:0] p1_array_index_1076879_comb;
  wire [7:0] p1_array_index_1076880_comb;
  wire [7:0] p1_array_index_1076881_comb;
  wire [7:0] p1_array_index_1076882_comb;
  wire [7:0] p1_res7__522_comb;
  wire [7:0] p1_res7__37_comb;
  wire [7:0] p1_array_index_1077339_comb;
  wire [7:0] p1_array_index_1076893_comb;
  wire [7:0] p1_array_index_1076894_comb;
  wire [7:0] p1_array_index_1076895_comb;
  wire [7:0] p1_res7__523_comb;
  wire [7:0] p1_res7__38_comb;
  wire [7:0] p1_array_index_1076905_comb;
  wire [7:0] p1_array_index_1076906_comb;
  wire [7:0] p1_array_index_1076907_comb;
  wire [7:0] p1_res7__524_comb;
  wire [7:0] p1_res7__39_comb;
  wire [7:0] p1_array_index_1076918_comb;
  wire [7:0] p1_array_index_1076919_comb;
  wire [7:0] p1_res7__525_comb;
  wire [7:0] p1_res7__40_comb;
  wire [7:0] p1_array_index_1076929_comb;
  wire [7:0] p1_array_index_1076930_comb;
  wire [7:0] p1_res7__526_comb;
  wire [7:0] p1_res7__41_comb;
  wire [7:0] p1_array_index_1076941_comb;
  wire [7:0] p1_res7__527_comb;
  wire [7:0] p1_res7__42_comb;
  wire [127:0] p1_res__32_comb;
  wire [7:0] p1_array_index_1076951_comb;
  wire [127:0] p1_addedKey__33_comb;
  wire [7:0] p1_res7__43_comb;
  wire [7:0] p1_array_index_1077393_comb;
  wire [7:0] p1_array_index_1077394_comb;
  wire [7:0] p1_array_index_1077395_comb;
  wire [7:0] p1_array_index_1077396_comb;
  wire [7:0] p1_array_index_1077397_comb;
  wire [7:0] p1_array_index_1077398_comb;
  wire [7:0] p1_array_index_1077400_comb;
  wire [7:0] p1_array_index_1077402_comb;
  wire [7:0] p1_array_index_1077403_comb;
  wire [7:0] p1_array_index_1077404_comb;
  wire [7:0] p1_array_index_1077405_comb;
  wire [7:0] p1_array_index_1077406_comb;
  wire [7:0] p1_array_index_1077407_comb;
  wire [7:0] p1_res7__44_comb;
  wire [7:0] p1_array_index_1077409_comb;
  wire [7:0] p1_array_index_1077410_comb;
  wire [7:0] p1_array_index_1077411_comb;
  wire [7:0] p1_array_index_1077412_comb;
  wire [7:0] p1_array_index_1077413_comb;
  wire [7:0] p1_array_index_1077414_comb;
  wire [7:0] p1_array_index_1077415_comb;
  wire [7:0] p1_array_index_1077417_comb;
  wire [7:0] p1_res7__528_comb;
  wire [7:0] p1_res7__45_comb;
  wire [7:0] p1_array_index_1077426_comb;
  wire [7:0] p1_array_index_1077427_comb;
  wire [7:0] p1_array_index_1077428_comb;
  wire [7:0] p1_array_index_1077429_comb;
  wire [7:0] p1_array_index_1077430_comb;
  wire [7:0] p1_array_index_1077431_comb;
  wire [7:0] p1_res7__529_comb;
  wire [7:0] p1_res7__46_comb;
  wire [7:0] p1_array_index_1077441_comb;
  wire [7:0] p1_array_index_1077442_comb;
  wire [7:0] p1_array_index_1077443_comb;
  wire [7:0] p1_array_index_1077444_comb;
  wire [7:0] p1_array_index_1077445_comb;
  wire [7:0] p1_res7__530_comb;
  wire [7:0] p1_res7__47_comb;
  wire [7:0] p1_array_index_1077455_comb;
  wire [7:0] p1_array_index_1077456_comb;
  wire [7:0] p1_array_index_1077457_comb;
  wire [7:0] p1_array_index_1077458_comb;
  wire [7:0] p1_array_index_1077459_comb;
  wire [127:0] p1_res__2_comb;
  wire [7:0] p1_res7__531_comb;
  wire [127:0] p1_xor_1076991_comb;
  wire [7:0] p1_array_index_1077470_comb;
  wire [7:0] p1_array_index_1077471_comb;
  wire [7:0] p1_array_index_1077472_comb;
  wire [7:0] p1_array_index_1077473_comb;
  wire [127:0] p1_addedKey__44_comb;
  wire [7:0] p1_res7__532_comb;
  wire [7:0] p1_array_index_1077483_comb;
  wire [7:0] p1_array_index_1077484_comb;
  wire [7:0] p1_array_index_1077485_comb;
  wire [7:0] p1_array_index_1077486_comb;
  wire [7:0] p1_array_index_1077007_comb;
  wire [7:0] p1_array_index_1077008_comb;
  wire [7:0] p1_array_index_1077009_comb;
  wire [7:0] p1_array_index_1077010_comb;
  wire [7:0] p1_array_index_1077011_comb;
  wire [7:0] p1_array_index_1077012_comb;
  wire [7:0] p1_array_index_1077014_comb;
  wire [7:0] p1_array_index_1077016_comb;
  wire [7:0] p1_array_index_1077017_comb;
  wire [7:0] p1_array_index_1077018_comb;
  wire [7:0] p1_array_index_1077019_comb;
  wire [7:0] p1_array_index_1077020_comb;
  wire [7:0] p1_array_index_1077021_comb;
  wire [7:0] p1_res7__533_comb;
  wire [7:0] p1_array_index_1077023_comb;
  wire [7:0] p1_array_index_1077024_comb;
  wire [7:0] p1_array_index_1077025_comb;
  wire [7:0] p1_array_index_1077026_comb;
  wire [7:0] p1_array_index_1077027_comb;
  wire [7:0] p1_array_index_1077028_comb;
  wire [7:0] p1_array_index_1077029_comb;
  wire [7:0] p1_array_index_1077031_comb;
  wire [7:0] p1_array_index_1077497_comb;
  wire [7:0] p1_array_index_1077498_comb;
  wire [7:0] p1_array_index_1077499_comb;
  wire [7:0] p1_res7__48_comb;
  wire [7:0] p1_res7__534_comb;
  wire [7:0] p1_array_index_1077040_comb;
  wire [7:0] p1_array_index_1077041_comb;
  wire [7:0] p1_array_index_1077042_comb;
  wire [7:0] p1_array_index_1077043_comb;
  wire [7:0] p1_array_index_1077044_comb;
  wire [7:0] p1_array_index_1077045_comb;
  wire [7:0] p1_array_index_1077509_comb;
  wire [7:0] p1_array_index_1077510_comb;
  wire [7:0] p1_array_index_1077511_comb;
  wire [7:0] p1_res7__49_comb;
  wire [7:0] p1_res7__535_comb;
  wire [7:0] p1_array_index_1077055_comb;
  wire [7:0] p1_array_index_1077056_comb;
  wire [7:0] p1_array_index_1077057_comb;
  wire [7:0] p1_array_index_1077058_comb;
  wire [7:0] p1_array_index_1077059_comb;
  wire [7:0] p1_array_index_1077522_comb;
  wire [7:0] p1_array_index_1077523_comb;
  wire [7:0] p1_res7__50_comb;
  wire [7:0] p1_res7__536_comb;
  wire [7:0] p1_array_index_1077069_comb;
  wire [7:0] p1_array_index_1077070_comb;
  wire [7:0] p1_array_index_1077071_comb;
  wire [7:0] p1_array_index_1077072_comb;
  wire [7:0] p1_array_index_1077073_comb;
  wire [7:0] p1_array_index_1077533_comb;
  wire [7:0] p1_array_index_1077534_comb;
  wire [7:0] p1_res7__51_comb;
  wire [7:0] p1_res7__537_comb;
  wire [7:0] p1_array_index_1077084_comb;
  wire [7:0] p1_array_index_1077085_comb;
  wire [7:0] p1_array_index_1077086_comb;
  wire [7:0] p1_array_index_1077087_comb;
  wire [7:0] p1_array_index_1077545_comb;
  wire [7:0] p1_res7__52_comb;
  wire [7:0] p1_res7__538_comb;
  wire [7:0] p1_array_index_1077097_comb;
  wire [7:0] p1_array_index_1077098_comb;
  wire [7:0] p1_array_index_1077099_comb;
  wire [7:0] p1_array_index_1077100_comb;
  wire [7:0] p1_array_index_1077555_comb;
  wire [7:0] p1_res7__53_comb;
  wire [7:0] p1_res7__539_comb;
  wire [7:0] p1_array_index_1077111_comb;
  wire [7:0] p1_array_index_1077112_comb;
  wire [7:0] p1_array_index_1077113_comb;
  wire [7:0] p1_res7__54_comb;
  wire [7:0] p1_res7__540_comb;
  wire [7:0] p1_array_index_1077123_comb;
  wire [7:0] p1_array_index_1077124_comb;
  wire [7:0] p1_array_index_1077125_comb;
  wire [7:0] p1_res7__55_comb;
  wire [7:0] p1_res7__541_comb;
  wire [7:0] p1_array_index_1077136_comb;
  wire [7:0] p1_array_index_1077137_comb;
  wire [7:0] p1_res7__56_comb;
  wire [7:0] p1_res7__542_comb;
  wire [7:0] p1_array_index_1077147_comb;
  wire [7:0] p1_array_index_1077148_comb;
  wire [7:0] p1_res7__57_comb;
  wire [7:0] p1_res7__543_comb;
  wire [7:0] p1_array_index_1077154_comb;
  wire [7:0] p1_array_index_1077155_comb;
  wire [7:0] p1_array_index_1077156_comb;
  wire [7:0] p1_array_index_1077157_comb;
  wire [7:0] p1_array_index_1077158_comb;
  wire [7:0] p1_array_index_1077159_comb;
  wire [7:0] p1_array_index_1077160_comb;
  wire [7:0] p1_array_index_1077161_comb;
  wire [7:0] p1_array_index_1077162_comb;
  wire [127:0] p1_res__33_comb;
  assign p1_addedKey__41_comb = p0_key[255:128] ^ 128'h6ea2_7672_6c48_7ab8_5d27_bd10_dd84_9401;
  assign p1_array_index_1076346_comb = arr[p1_addedKey__41_comb[127:120]];
  assign p1_array_index_1076348_comb = arr[p1_addedKey__41_comb[119:112]];
  assign p1_array_index_1076350_comb = arr[p1_addedKey__41_comb[111:104]];
  assign p1_array_index_1076352_comb = arr[p1_addedKey__41_comb[103:96]];
  assign p1_array_index_1076354_comb = arr[p1_addedKey__41_comb[95:88]];
  assign p1_array_index_1076356_comb = arr[p1_addedKey__41_comb[87:80]];
  assign p1_array_index_1076359_comb = arr[p1_addedKey__41_comb[71:64]];
  assign p1_array_index_1076361_comb = arr[p1_addedKey__41_comb[55:48]];
  assign p1_array_index_1076362_comb = arr[p1_addedKey__41_comb[47:40]];
  assign p1_array_index_1076363_comb = arr[p1_addedKey__41_comb[39:32]];
  assign p1_array_index_1076364_comb = arr[p1_addedKey__41_comb[31:24]];
  assign p1_array_index_1076365_comb = arr[p1_addedKey__41_comb[23:16]];
  assign p1_array_index_1076366_comb = arr[p1_addedKey__41_comb[15:8]];
  assign p1_array_index_1076368_comb = literal_1076345[p1_array_index_1076346_comb];
  assign p1_array_index_1076369_comb = literal_1076347[p1_array_index_1076348_comb];
  assign p1_array_index_1076370_comb = literal_1076349[p1_array_index_1076350_comb];
  assign p1_array_index_1076371_comb = literal_1076351[p1_array_index_1076352_comb];
  assign p1_array_index_1076372_comb = literal_1076353[p1_array_index_1076354_comb];
  assign p1_array_index_1076373_comb = literal_1076355[p1_array_index_1076356_comb];
  assign p1_array_index_1076374_comb = arr[p1_addedKey__41_comb[79:72]];
  assign p1_array_index_1076376_comb = arr[p1_addedKey__41_comb[63:56]];
  assign p1_res7_comb = p1_array_index_1076368_comb ^ p1_array_index_1076369_comb ^ p1_array_index_1076370_comb ^ p1_array_index_1076371_comb ^ p1_array_index_1076372_comb ^ p1_array_index_1076373_comb ^ p1_array_index_1076374_comb ^ literal_1076358[p1_array_index_1076359_comb] ^ p1_array_index_1076376_comb ^ literal_1076355[p1_array_index_1076361_comb] ^ literal_1076353[p1_array_index_1076362_comb] ^ literal_1076351[p1_array_index_1076363_comb] ^ literal_1076349[p1_array_index_1076364_comb] ^ literal_1076347[p1_array_index_1076365_comb] ^ literal_1076345[p1_array_index_1076366_comb] ^ arr[p1_addedKey__41_comb[7:0]];
  assign p1_array_index_1076385_comb = literal_1076345[p1_res7_comb];
  assign p1_array_index_1076386_comb = literal_1076347[p1_array_index_1076346_comb];
  assign p1_array_index_1076387_comb = literal_1076349[p1_array_index_1076348_comb];
  assign p1_array_index_1076388_comb = literal_1076351[p1_array_index_1076350_comb];
  assign p1_array_index_1076389_comb = literal_1076353[p1_array_index_1076352_comb];
  assign p1_array_index_1076390_comb = literal_1076355[p1_array_index_1076354_comb];
  assign p1_res7__1_comb = p1_array_index_1076385_comb ^ p1_array_index_1076386_comb ^ p1_array_index_1076387_comb ^ p1_array_index_1076388_comb ^ p1_array_index_1076389_comb ^ p1_array_index_1076390_comb ^ p1_array_index_1076356_comb ^ literal_1076358[p1_array_index_1076374_comb] ^ p1_array_index_1076359_comb ^ literal_1076355[p1_array_index_1076376_comb] ^ literal_1076353[p1_array_index_1076361_comb] ^ literal_1076351[p1_array_index_1076362_comb] ^ literal_1076349[p1_array_index_1076363_comb] ^ literal_1076347[p1_array_index_1076364_comb] ^ literal_1076345[p1_array_index_1076365_comb] ^ p1_array_index_1076366_comb;
  assign p1_array_index_1076400_comb = literal_1076347[p1_res7_comb];
  assign p1_array_index_1076401_comb = literal_1076349[p1_array_index_1076346_comb];
  assign p1_array_index_1076402_comb = literal_1076351[p1_array_index_1076348_comb];
  assign p1_array_index_1076403_comb = literal_1076353[p1_array_index_1076350_comb];
  assign p1_array_index_1076404_comb = literal_1076355[p1_array_index_1076352_comb];
  assign p1_res7__2_comb = literal_1076345[p1_res7__1_comb] ^ p1_array_index_1076400_comb ^ p1_array_index_1076401_comb ^ p1_array_index_1076402_comb ^ p1_array_index_1076403_comb ^ p1_array_index_1076404_comb ^ p1_array_index_1076354_comb ^ literal_1076358[p1_array_index_1076356_comb] ^ p1_array_index_1076374_comb ^ literal_1076355[p1_array_index_1076359_comb] ^ literal_1076353[p1_array_index_1076376_comb] ^ literal_1076351[p1_array_index_1076361_comb] ^ literal_1076349[p1_array_index_1076362_comb] ^ literal_1076347[p1_array_index_1076363_comb] ^ literal_1076345[p1_array_index_1076364_comb] ^ p1_array_index_1076365_comb;
  assign p1_array_index_1076414_comb = literal_1076347[p1_res7__1_comb];
  assign p1_array_index_1076415_comb = literal_1076349[p1_res7_comb];
  assign p1_array_index_1076416_comb = literal_1076351[p1_array_index_1076346_comb];
  assign p1_array_index_1076417_comb = literal_1076353[p1_array_index_1076348_comb];
  assign p1_array_index_1076418_comb = literal_1076355[p1_array_index_1076350_comb];
  assign p1_res7__3_comb = literal_1076345[p1_res7__2_comb] ^ p1_array_index_1076414_comb ^ p1_array_index_1076415_comb ^ p1_array_index_1076416_comb ^ p1_array_index_1076417_comb ^ p1_array_index_1076418_comb ^ p1_array_index_1076352_comb ^ literal_1076358[p1_array_index_1076354_comb] ^ p1_array_index_1076356_comb ^ literal_1076355[p1_array_index_1076374_comb] ^ literal_1076353[p1_array_index_1076359_comb] ^ literal_1076351[p1_array_index_1076376_comb] ^ literal_1076349[p1_array_index_1076361_comb] ^ literal_1076347[p1_array_index_1076362_comb] ^ literal_1076345[p1_array_index_1076363_comb] ^ p1_array_index_1076364_comb;
  assign p1_array_index_1076429_comb = literal_1076349[p1_res7__1_comb];
  assign p1_array_index_1076430_comb = literal_1076351[p1_res7_comb];
  assign p1_array_index_1076431_comb = literal_1076353[p1_array_index_1076346_comb];
  assign p1_array_index_1076432_comb = literal_1076355[p1_array_index_1076348_comb];
  assign p1_res7__4_comb = literal_1076345[p1_res7__3_comb] ^ literal_1076347[p1_res7__2_comb] ^ p1_array_index_1076429_comb ^ p1_array_index_1076430_comb ^ p1_array_index_1076431_comb ^ p1_array_index_1076432_comb ^ p1_array_index_1076350_comb ^ literal_1076358[p1_array_index_1076352_comb] ^ p1_array_index_1076354_comb ^ p1_array_index_1076373_comb ^ literal_1076353[p1_array_index_1076374_comb] ^ literal_1076351[p1_array_index_1076359_comb] ^ literal_1076349[p1_array_index_1076376_comb] ^ literal_1076347[p1_array_index_1076361_comb] ^ literal_1076345[p1_array_index_1076362_comb] ^ p1_array_index_1076363_comb;
  assign p1_array_index_1076442_comb = literal_1076349[p1_res7__2_comb];
  assign p1_array_index_1076443_comb = literal_1076351[p1_res7__1_comb];
  assign p1_array_index_1076444_comb = literal_1076353[p1_res7_comb];
  assign p1_array_index_1076445_comb = literal_1076355[p1_array_index_1076346_comb];
  assign p1_res7__5_comb = literal_1076345[p1_res7__4_comb] ^ literal_1076347[p1_res7__3_comb] ^ p1_array_index_1076442_comb ^ p1_array_index_1076443_comb ^ p1_array_index_1076444_comb ^ p1_array_index_1076445_comb ^ p1_array_index_1076348_comb ^ literal_1076358[p1_array_index_1076350_comb] ^ p1_array_index_1076352_comb ^ p1_array_index_1076390_comb ^ literal_1076353[p1_array_index_1076356_comb] ^ literal_1076351[p1_array_index_1076374_comb] ^ literal_1076349[p1_array_index_1076359_comb] ^ literal_1076347[p1_array_index_1076376_comb] ^ literal_1076345[p1_array_index_1076361_comb] ^ p1_array_index_1076362_comb;
  assign p1_array_index_1076456_comb = literal_1076351[p1_res7__2_comb];
  assign p1_array_index_1076457_comb = literal_1076353[p1_res7__1_comb];
  assign p1_array_index_1076458_comb = literal_1076355[p1_res7_comb];
  assign p1_res7__6_comb = literal_1076345[p1_res7__5_comb] ^ literal_1076347[p1_res7__4_comb] ^ literal_1076349[p1_res7__3_comb] ^ p1_array_index_1076456_comb ^ p1_array_index_1076457_comb ^ p1_array_index_1076458_comb ^ p1_array_index_1076346_comb ^ literal_1076358[p1_array_index_1076348_comb] ^ p1_array_index_1076350_comb ^ p1_array_index_1076404_comb ^ p1_array_index_1076372_comb ^ literal_1076351[p1_array_index_1076356_comb] ^ literal_1076349[p1_array_index_1076374_comb] ^ literal_1076347[p1_array_index_1076359_comb] ^ literal_1076345[p1_array_index_1076376_comb] ^ p1_array_index_1076361_comb;
  assign p1_array_index_1076468_comb = literal_1076351[p1_res7__3_comb];
  assign p1_array_index_1076469_comb = literal_1076353[p1_res7__2_comb];
  assign p1_array_index_1076470_comb = literal_1076355[p1_res7__1_comb];
  assign p1_res7__7_comb = literal_1076345[p1_res7__6_comb] ^ literal_1076347[p1_res7__5_comb] ^ literal_1076349[p1_res7__4_comb] ^ p1_array_index_1076468_comb ^ p1_array_index_1076469_comb ^ p1_array_index_1076470_comb ^ p1_res7_comb ^ literal_1076358[p1_array_index_1076346_comb] ^ p1_array_index_1076348_comb ^ p1_array_index_1076418_comb ^ p1_array_index_1076389_comb ^ literal_1076351[p1_array_index_1076354_comb] ^ literal_1076349[p1_array_index_1076356_comb] ^ literal_1076347[p1_array_index_1076374_comb] ^ literal_1076345[p1_array_index_1076359_comb] ^ p1_array_index_1076376_comb;
  assign p1_array_index_1076481_comb = literal_1076353[p1_res7__3_comb];
  assign p1_array_index_1076482_comb = literal_1076355[p1_res7__2_comb];
  assign p1_res7__8_comb = literal_1076345[p1_res7__7_comb] ^ literal_1076347[p1_res7__6_comb] ^ literal_1076349[p1_res7__5_comb] ^ literal_1076351[p1_res7__4_comb] ^ p1_array_index_1076481_comb ^ p1_array_index_1076482_comb ^ p1_res7__1_comb ^ literal_1076358[p1_res7_comb] ^ p1_array_index_1076346_comb ^ p1_array_index_1076432_comb ^ p1_array_index_1076403_comb ^ p1_array_index_1076371_comb ^ literal_1076349[p1_array_index_1076354_comb] ^ literal_1076347[p1_array_index_1076356_comb] ^ literal_1076345[p1_array_index_1076374_comb] ^ p1_array_index_1076359_comb;
  assign p1_array_index_1076492_comb = literal_1076353[p1_res7__4_comb];
  assign p1_array_index_1076493_comb = literal_1076355[p1_res7__3_comb];
  assign p1_res7__9_comb = literal_1076345[p1_res7__8_comb] ^ literal_1076347[p1_res7__7_comb] ^ literal_1076349[p1_res7__6_comb] ^ literal_1076351[p1_res7__5_comb] ^ p1_array_index_1076492_comb ^ p1_array_index_1076493_comb ^ p1_res7__2_comb ^ literal_1076358[p1_res7__1_comb] ^ p1_res7_comb ^ p1_array_index_1076445_comb ^ p1_array_index_1076417_comb ^ p1_array_index_1076388_comb ^ literal_1076349[p1_array_index_1076352_comb] ^ literal_1076347[p1_array_index_1076354_comb] ^ literal_1076345[p1_array_index_1076356_comb] ^ p1_array_index_1076374_comb;
  assign p1_array_index_1076504_comb = literal_1076355[p1_res7__4_comb];
  assign p1_res7__10_comb = literal_1076345[p1_res7__9_comb] ^ literal_1076347[p1_res7__8_comb] ^ literal_1076349[p1_res7__7_comb] ^ literal_1076351[p1_res7__6_comb] ^ literal_1076353[p1_res7__5_comb] ^ p1_array_index_1076504_comb ^ p1_res7__3_comb ^ literal_1076358[p1_res7__2_comb] ^ p1_res7__1_comb ^ p1_array_index_1076458_comb ^ p1_array_index_1076431_comb ^ p1_array_index_1076402_comb ^ p1_array_index_1076370_comb ^ literal_1076347[p1_array_index_1076352_comb] ^ literal_1076345[p1_array_index_1076354_comb] ^ p1_array_index_1076356_comb;
  assign p1_array_index_1076514_comb = literal_1076355[p1_res7__5_comb];
  assign p1_res7__11_comb = literal_1076345[p1_res7__10_comb] ^ literal_1076347[p1_res7__9_comb] ^ literal_1076349[p1_res7__8_comb] ^ literal_1076351[p1_res7__7_comb] ^ literal_1076353[p1_res7__6_comb] ^ p1_array_index_1076514_comb ^ p1_res7__4_comb ^ literal_1076358[p1_res7__3_comb] ^ p1_res7__2_comb ^ p1_array_index_1076470_comb ^ p1_array_index_1076444_comb ^ p1_array_index_1076416_comb ^ p1_array_index_1076387_comb ^ literal_1076347[p1_array_index_1076350_comb] ^ literal_1076345[p1_array_index_1076352_comb] ^ p1_array_index_1076354_comb;
  assign p1_res7__12_comb = literal_1076345[p1_res7__11_comb] ^ literal_1076347[p1_res7__10_comb] ^ literal_1076349[p1_res7__9_comb] ^ literal_1076351[p1_res7__8_comb] ^ literal_1076353[p1_res7__7_comb] ^ literal_1076355[p1_res7__6_comb] ^ p1_res7__5_comb ^ literal_1076358[p1_res7__4_comb] ^ p1_res7__3_comb ^ p1_array_index_1076482_comb ^ p1_array_index_1076457_comb ^ p1_array_index_1076430_comb ^ p1_array_index_1076401_comb ^ p1_array_index_1076369_comb ^ literal_1076345[p1_array_index_1076350_comb] ^ p1_array_index_1076352_comb;
  assign p1_res7__13_comb = literal_1076345[p1_res7__12_comb] ^ literal_1076347[p1_res7__11_comb] ^ literal_1076349[p1_res7__10_comb] ^ literal_1076351[p1_res7__9_comb] ^ literal_1076353[p1_res7__8_comb] ^ literal_1076355[p1_res7__7_comb] ^ p1_res7__6_comb ^ literal_1076358[p1_res7__5_comb] ^ p1_res7__4_comb ^ p1_array_index_1076493_comb ^ p1_array_index_1076469_comb ^ p1_array_index_1076443_comb ^ p1_array_index_1076415_comb ^ p1_array_index_1076386_comb ^ literal_1076345[p1_array_index_1076348_comb] ^ p1_array_index_1076350_comb;
  assign p1_res7__14_comb = literal_1076345[p1_res7__13_comb] ^ literal_1076347[p1_res7__12_comb] ^ literal_1076349[p1_res7__11_comb] ^ literal_1076351[p1_res7__10_comb] ^ literal_1076353[p1_res7__9_comb] ^ literal_1076355[p1_res7__8_comb] ^ p1_res7__7_comb ^ literal_1076358[p1_res7__6_comb] ^ p1_res7__5_comb ^ p1_array_index_1076504_comb ^ p1_array_index_1076481_comb ^ p1_array_index_1076456_comb ^ p1_array_index_1076429_comb ^ p1_array_index_1076400_comb ^ p1_array_index_1076368_comb ^ p1_array_index_1076348_comb;
  assign p1_res7__15_comb = literal_1076345[p1_res7__14_comb] ^ literal_1076347[p1_res7__13_comb] ^ literal_1076349[p1_res7__12_comb] ^ literal_1076351[p1_res7__11_comb] ^ literal_1076353[p1_res7__10_comb] ^ literal_1076355[p1_res7__9_comb] ^ p1_res7__8_comb ^ literal_1076358[p1_res7__7_comb] ^ p1_res7__6_comb ^ p1_array_index_1076514_comb ^ p1_array_index_1076492_comb ^ p1_array_index_1076468_comb ^ p1_array_index_1076442_comb ^ p1_array_index_1076414_comb ^ p1_array_index_1076385_comb ^ p1_array_index_1076346_comb;
  assign p1_res_comb = {p1_res7__15_comb, p1_res7__14_comb, p1_res7__13_comb, p1_res7__12_comb, p1_res7__11_comb, p1_res7__10_comb, p1_res7__9_comb, p1_res7__8_comb, p1_res7__7_comb, p1_res7__6_comb, p1_res7__5_comb, p1_res7__4_comb, p1_res7__3_comb, p1_res7__2_comb, p1_res7__1_comb, p1_res7_comb};
  assign p1_xor_1076555_comb = p1_res_comb ^ p0_key[127:0];
  assign p1_addedKey__42_comb = p1_xor_1076555_comb ^ 128'hdc87_ece4_d890_f4b3_ba4e_b920_79cb_eb02;
  assign p1_array_index_1076571_comb = arr[p1_addedKey__42_comb[127:120]];
  assign p1_array_index_1076572_comb = arr[p1_addedKey__42_comb[119:112]];
  assign p1_array_index_1076573_comb = arr[p1_addedKey__42_comb[111:104]];
  assign p1_array_index_1076574_comb = arr[p1_addedKey__42_comb[103:96]];
  assign p1_array_index_1076575_comb = arr[p1_addedKey__42_comb[95:88]];
  assign p1_array_index_1076576_comb = arr[p1_addedKey__42_comb[87:80]];
  assign p1_array_index_1076578_comb = arr[p1_addedKey__42_comb[71:64]];
  assign p1_array_index_1076580_comb = arr[p1_addedKey__42_comb[55:48]];
  assign p1_array_index_1076581_comb = arr[p1_addedKey__42_comb[47:40]];
  assign p1_array_index_1076582_comb = arr[p1_addedKey__42_comb[39:32]];
  assign p1_array_index_1076583_comb = arr[p1_addedKey__42_comb[31:24]];
  assign p1_array_index_1076584_comb = arr[p1_addedKey__42_comb[23:16]];
  assign p1_array_index_1076585_comb = arr[p1_addedKey__42_comb[15:8]];
  assign p1_array_index_1076587_comb = literal_1076345[p1_array_index_1076571_comb];
  assign p1_array_index_1076588_comb = literal_1076347[p1_array_index_1076572_comb];
  assign p1_array_index_1076589_comb = literal_1076349[p1_array_index_1076573_comb];
  assign p1_array_index_1076590_comb = literal_1076351[p1_array_index_1076574_comb];
  assign p1_array_index_1076591_comb = literal_1076353[p1_array_index_1076575_comb];
  assign p1_array_index_1076592_comb = literal_1076355[p1_array_index_1076576_comb];
  assign p1_array_index_1076593_comb = arr[p1_addedKey__42_comb[79:72]];
  assign p1_array_index_1076595_comb = arr[p1_addedKey__42_comb[63:56]];
  assign p1_res7__16_comb = p1_array_index_1076587_comb ^ p1_array_index_1076588_comb ^ p1_array_index_1076589_comb ^ p1_array_index_1076590_comb ^ p1_array_index_1076591_comb ^ p1_array_index_1076592_comb ^ p1_array_index_1076593_comb ^ literal_1076358[p1_array_index_1076578_comb] ^ p1_array_index_1076595_comb ^ literal_1076355[p1_array_index_1076580_comb] ^ literal_1076353[p1_array_index_1076581_comb] ^ literal_1076351[p1_array_index_1076582_comb] ^ literal_1076349[p1_array_index_1076583_comb] ^ literal_1076347[p1_array_index_1076584_comb] ^ literal_1076345[p1_array_index_1076585_comb] ^ arr[p1_addedKey__42_comb[7:0]];
  assign p1_array_index_1076604_comb = literal_1076345[p1_res7__16_comb];
  assign p1_array_index_1076605_comb = literal_1076347[p1_array_index_1076571_comb];
  assign p1_array_index_1076606_comb = literal_1076349[p1_array_index_1076572_comb];
  assign p1_array_index_1076607_comb = literal_1076351[p1_array_index_1076573_comb];
  assign p1_array_index_1076608_comb = literal_1076353[p1_array_index_1076574_comb];
  assign p1_array_index_1076609_comb = literal_1076355[p1_array_index_1076575_comb];
  assign p1_res7__17_comb = p1_array_index_1076604_comb ^ p1_array_index_1076605_comb ^ p1_array_index_1076606_comb ^ p1_array_index_1076607_comb ^ p1_array_index_1076608_comb ^ p1_array_index_1076609_comb ^ p1_array_index_1076576_comb ^ literal_1076358[p1_array_index_1076593_comb] ^ p1_array_index_1076578_comb ^ literal_1076355[p1_array_index_1076595_comb] ^ literal_1076353[p1_array_index_1076580_comb] ^ literal_1076351[p1_array_index_1076581_comb] ^ literal_1076349[p1_array_index_1076582_comb] ^ literal_1076347[p1_array_index_1076583_comb] ^ literal_1076345[p1_array_index_1076584_comb] ^ p1_array_index_1076585_comb;
  assign p1_array_index_1076619_comb = literal_1076347[p1_res7__16_comb];
  assign p1_array_index_1076620_comb = literal_1076349[p1_array_index_1076571_comb];
  assign p1_array_index_1076621_comb = literal_1076351[p1_array_index_1076572_comb];
  assign p1_array_index_1076622_comb = literal_1076353[p1_array_index_1076573_comb];
  assign p1_array_index_1076623_comb = literal_1076355[p1_array_index_1076574_comb];
  assign p1_res7__18_comb = literal_1076345[p1_res7__17_comb] ^ p1_array_index_1076619_comb ^ p1_array_index_1076620_comb ^ p1_array_index_1076621_comb ^ p1_array_index_1076622_comb ^ p1_array_index_1076623_comb ^ p1_array_index_1076575_comb ^ literal_1076358[p1_array_index_1076576_comb] ^ p1_array_index_1076593_comb ^ literal_1076355[p1_array_index_1076578_comb] ^ literal_1076353[p1_array_index_1076595_comb] ^ literal_1076351[p1_array_index_1076580_comb] ^ literal_1076349[p1_array_index_1076581_comb] ^ literal_1076347[p1_array_index_1076582_comb] ^ literal_1076345[p1_array_index_1076583_comb] ^ p1_array_index_1076584_comb;
  assign p1_array_index_1076633_comb = literal_1076347[p1_res7__17_comb];
  assign p1_array_index_1076634_comb = literal_1076349[p1_res7__16_comb];
  assign p1_array_index_1076635_comb = literal_1076351[p1_array_index_1076571_comb];
  assign p1_array_index_1076636_comb = literal_1076353[p1_array_index_1076572_comb];
  assign p1_array_index_1076637_comb = literal_1076355[p1_array_index_1076573_comb];
  assign p1_res7__19_comb = literal_1076345[p1_res7__18_comb] ^ p1_array_index_1076633_comb ^ p1_array_index_1076634_comb ^ p1_array_index_1076635_comb ^ p1_array_index_1076636_comb ^ p1_array_index_1076637_comb ^ p1_array_index_1076574_comb ^ literal_1076358[p1_array_index_1076575_comb] ^ p1_array_index_1076576_comb ^ literal_1076355[p1_array_index_1076593_comb] ^ literal_1076353[p1_array_index_1076578_comb] ^ literal_1076351[p1_array_index_1076595_comb] ^ literal_1076349[p1_array_index_1076580_comb] ^ literal_1076347[p1_array_index_1076581_comb] ^ literal_1076345[p1_array_index_1076582_comb] ^ p1_array_index_1076583_comb;
  assign p1_array_index_1076648_comb = literal_1076349[p1_res7__17_comb];
  assign p1_array_index_1076649_comb = literal_1076351[p1_res7__16_comb];
  assign p1_array_index_1076650_comb = literal_1076353[p1_array_index_1076571_comb];
  assign p1_array_index_1076651_comb = literal_1076355[p1_array_index_1076572_comb];
  assign p1_res7__20_comb = literal_1076345[p1_res7__19_comb] ^ literal_1076347[p1_res7__18_comb] ^ p1_array_index_1076648_comb ^ p1_array_index_1076649_comb ^ p1_array_index_1076650_comb ^ p1_array_index_1076651_comb ^ p1_array_index_1076573_comb ^ literal_1076358[p1_array_index_1076574_comb] ^ p1_array_index_1076575_comb ^ p1_array_index_1076592_comb ^ literal_1076353[p1_array_index_1076593_comb] ^ literal_1076351[p1_array_index_1076578_comb] ^ literal_1076349[p1_array_index_1076595_comb] ^ literal_1076347[p1_array_index_1076580_comb] ^ literal_1076345[p1_array_index_1076581_comb] ^ p1_array_index_1076582_comb;
  assign p1_array_index_1076661_comb = literal_1076349[p1_res7__18_comb];
  assign p1_array_index_1076662_comb = literal_1076351[p1_res7__17_comb];
  assign p1_array_index_1076663_comb = literal_1076353[p1_res7__16_comb];
  assign p1_array_index_1076664_comb = literal_1076355[p1_array_index_1076571_comb];
  assign p1_res7__21_comb = literal_1076345[p1_res7__20_comb] ^ literal_1076347[p1_res7__19_comb] ^ p1_array_index_1076661_comb ^ p1_array_index_1076662_comb ^ p1_array_index_1076663_comb ^ p1_array_index_1076664_comb ^ p1_array_index_1076572_comb ^ literal_1076358[p1_array_index_1076573_comb] ^ p1_array_index_1076574_comb ^ p1_array_index_1076609_comb ^ literal_1076353[p1_array_index_1076576_comb] ^ literal_1076351[p1_array_index_1076593_comb] ^ literal_1076349[p1_array_index_1076578_comb] ^ literal_1076347[p1_array_index_1076595_comb] ^ literal_1076345[p1_array_index_1076580_comb] ^ p1_array_index_1076581_comb;
  assign p1_array_index_1076675_comb = literal_1076351[p1_res7__18_comb];
  assign p1_array_index_1076676_comb = literal_1076353[p1_res7__17_comb];
  assign p1_array_index_1076677_comb = literal_1076355[p1_res7__16_comb];
  assign p1_res7__22_comb = literal_1076345[p1_res7__21_comb] ^ literal_1076347[p1_res7__20_comb] ^ literal_1076349[p1_res7__19_comb] ^ p1_array_index_1076675_comb ^ p1_array_index_1076676_comb ^ p1_array_index_1076677_comb ^ p1_array_index_1076571_comb ^ literal_1076358[p1_array_index_1076572_comb] ^ p1_array_index_1076573_comb ^ p1_array_index_1076623_comb ^ p1_array_index_1076591_comb ^ literal_1076351[p1_array_index_1076576_comb] ^ literal_1076349[p1_array_index_1076593_comb] ^ literal_1076347[p1_array_index_1076578_comb] ^ literal_1076345[p1_array_index_1076595_comb] ^ p1_array_index_1076580_comb;
  assign p1_array_index_1076687_comb = literal_1076351[p1_res7__19_comb];
  assign p1_array_index_1076688_comb = literal_1076353[p1_res7__18_comb];
  assign p1_array_index_1076689_comb = literal_1076355[p1_res7__17_comb];
  assign p1_res7__23_comb = literal_1076345[p1_res7__22_comb] ^ literal_1076347[p1_res7__21_comb] ^ literal_1076349[p1_res7__20_comb] ^ p1_array_index_1076687_comb ^ p1_array_index_1076688_comb ^ p1_array_index_1076689_comb ^ p1_res7__16_comb ^ literal_1076358[p1_array_index_1076571_comb] ^ p1_array_index_1076572_comb ^ p1_array_index_1076637_comb ^ p1_array_index_1076608_comb ^ literal_1076351[p1_array_index_1076575_comb] ^ literal_1076349[p1_array_index_1076576_comb] ^ literal_1076347[p1_array_index_1076593_comb] ^ literal_1076345[p1_array_index_1076578_comb] ^ p1_array_index_1076595_comb;
  assign p1_array_index_1076700_comb = literal_1076353[p1_res7__19_comb];
  assign p1_array_index_1076701_comb = literal_1076355[p1_res7__18_comb];
  assign p1_res7__24_comb = literal_1076345[p1_res7__23_comb] ^ literal_1076347[p1_res7__22_comb] ^ literal_1076349[p1_res7__21_comb] ^ literal_1076351[p1_res7__20_comb] ^ p1_array_index_1076700_comb ^ p1_array_index_1076701_comb ^ p1_res7__17_comb ^ literal_1076358[p1_res7__16_comb] ^ p1_array_index_1076571_comb ^ p1_array_index_1076651_comb ^ p1_array_index_1076622_comb ^ p1_array_index_1076590_comb ^ literal_1076349[p1_array_index_1076575_comb] ^ literal_1076347[p1_array_index_1076576_comb] ^ literal_1076345[p1_array_index_1076593_comb] ^ p1_array_index_1076578_comb;
  assign p1_array_index_1076711_comb = literal_1076353[p1_res7__20_comb];
  assign p1_array_index_1076712_comb = literal_1076355[p1_res7__19_comb];
  assign p1_res7__25_comb = literal_1076345[p1_res7__24_comb] ^ literal_1076347[p1_res7__23_comb] ^ literal_1076349[p1_res7__22_comb] ^ literal_1076351[p1_res7__21_comb] ^ p1_array_index_1076711_comb ^ p1_array_index_1076712_comb ^ p1_res7__18_comb ^ literal_1076358[p1_res7__17_comb] ^ p1_res7__16_comb ^ p1_array_index_1076664_comb ^ p1_array_index_1076636_comb ^ p1_array_index_1076607_comb ^ literal_1076349[p1_array_index_1076574_comb] ^ literal_1076347[p1_array_index_1076575_comb] ^ literal_1076345[p1_array_index_1076576_comb] ^ p1_array_index_1076593_comb;
  assign p1_array_index_1076723_comb = literal_1076355[p1_res7__20_comb];
  assign p1_res7__26_comb = literal_1076345[p1_res7__25_comb] ^ literal_1076347[p1_res7__24_comb] ^ literal_1076349[p1_res7__23_comb] ^ literal_1076351[p1_res7__22_comb] ^ literal_1076353[p1_res7__21_comb] ^ p1_array_index_1076723_comb ^ p1_res7__19_comb ^ literal_1076358[p1_res7__18_comb] ^ p1_res7__17_comb ^ p1_array_index_1076677_comb ^ p1_array_index_1076650_comb ^ p1_array_index_1076621_comb ^ p1_array_index_1076589_comb ^ literal_1076347[p1_array_index_1076574_comb] ^ literal_1076345[p1_array_index_1076575_comb] ^ p1_array_index_1076576_comb;
  assign p1_array_index_1076733_comb = literal_1076355[p1_res7__21_comb];
  assign p1_res7__27_comb = literal_1076345[p1_res7__26_comb] ^ literal_1076347[p1_res7__25_comb] ^ literal_1076349[p1_res7__24_comb] ^ literal_1076351[p1_res7__23_comb] ^ literal_1076353[p1_res7__22_comb] ^ p1_array_index_1076733_comb ^ p1_res7__20_comb ^ literal_1076358[p1_res7__19_comb] ^ p1_res7__18_comb ^ p1_array_index_1076689_comb ^ p1_array_index_1076663_comb ^ p1_array_index_1076635_comb ^ p1_array_index_1076606_comb ^ literal_1076347[p1_array_index_1076573_comb] ^ literal_1076345[p1_array_index_1076574_comb] ^ p1_array_index_1076575_comb;
  assign p1_addedKey__32_comb = p0_key[255:128] ^ p0__block;
  assign p1_res7__28_comb = literal_1076345[p1_res7__27_comb] ^ literal_1076347[p1_res7__26_comb] ^ literal_1076349[p1_res7__25_comb] ^ literal_1076351[p1_res7__24_comb] ^ literal_1076353[p1_res7__23_comb] ^ literal_1076355[p1_res7__22_comb] ^ p1_res7__21_comb ^ literal_1076358[p1_res7__20_comb] ^ p1_res7__19_comb ^ p1_array_index_1076701_comb ^ p1_array_index_1076676_comb ^ p1_array_index_1076649_comb ^ p1_array_index_1076620_comb ^ p1_array_index_1076588_comb ^ literal_1076345[p1_array_index_1076573_comb] ^ p1_array_index_1076574_comb;
  assign p1_array_index_1077177_comb = arr[p1_addedKey__32_comb[127:120]];
  assign p1_array_index_1077178_comb = arr[p1_addedKey__32_comb[119:112]];
  assign p1_array_index_1077179_comb = arr[p1_addedKey__32_comb[111:104]];
  assign p1_array_index_1077180_comb = arr[p1_addedKey__32_comb[103:96]];
  assign p1_array_index_1077181_comb = arr[p1_addedKey__32_comb[95:88]];
  assign p1_array_index_1077182_comb = arr[p1_addedKey__32_comb[87:80]];
  assign p1_array_index_1077184_comb = arr[p1_addedKey__32_comb[71:64]];
  assign p1_array_index_1077186_comb = arr[p1_addedKey__32_comb[55:48]];
  assign p1_array_index_1077187_comb = arr[p1_addedKey__32_comb[47:40]];
  assign p1_array_index_1077188_comb = arr[p1_addedKey__32_comb[39:32]];
  assign p1_array_index_1077189_comb = arr[p1_addedKey__32_comb[31:24]];
  assign p1_array_index_1077190_comb = arr[p1_addedKey__32_comb[23:16]];
  assign p1_array_index_1077191_comb = arr[p1_addedKey__32_comb[15:8]];
  assign p1_array_index_1077193_comb = literal_1076345[p1_array_index_1077177_comb];
  assign p1_array_index_1077194_comb = literal_1076347[p1_array_index_1077178_comb];
  assign p1_array_index_1077195_comb = literal_1076349[p1_array_index_1077179_comb];
  assign p1_array_index_1077196_comb = literal_1076351[p1_array_index_1077180_comb];
  assign p1_array_index_1077197_comb = literal_1076353[p1_array_index_1077181_comb];
  assign p1_array_index_1077198_comb = literal_1076355[p1_array_index_1077182_comb];
  assign p1_array_index_1077199_comb = arr[p1_addedKey__32_comb[79:72]];
  assign p1_array_index_1077201_comb = arr[p1_addedKey__32_comb[63:56]];
  assign p1_res7__29_comb = literal_1076345[p1_res7__28_comb] ^ literal_1076347[p1_res7__27_comb] ^ literal_1076349[p1_res7__26_comb] ^ literal_1076351[p1_res7__25_comb] ^ literal_1076353[p1_res7__24_comb] ^ literal_1076355[p1_res7__23_comb] ^ p1_res7__22_comb ^ literal_1076358[p1_res7__21_comb] ^ p1_res7__20_comb ^ p1_array_index_1076712_comb ^ p1_array_index_1076688_comb ^ p1_array_index_1076662_comb ^ p1_array_index_1076634_comb ^ p1_array_index_1076605_comb ^ literal_1076345[p1_array_index_1076572_comb] ^ p1_array_index_1076573_comb;
  assign p1_res7__512_comb = p1_array_index_1077193_comb ^ p1_array_index_1077194_comb ^ p1_array_index_1077195_comb ^ p1_array_index_1077196_comb ^ p1_array_index_1077197_comb ^ p1_array_index_1077198_comb ^ p1_array_index_1077199_comb ^ literal_1076358[p1_array_index_1077184_comb] ^ p1_array_index_1077201_comb ^ literal_1076355[p1_array_index_1077186_comb] ^ literal_1076353[p1_array_index_1077187_comb] ^ literal_1076351[p1_array_index_1077188_comb] ^ literal_1076349[p1_array_index_1077189_comb] ^ literal_1076347[p1_array_index_1077190_comb] ^ literal_1076345[p1_array_index_1077191_comb] ^ arr[p1_addedKey__32_comb[7:0]];
  assign p1_array_index_1077210_comb = literal_1076345[p1_res7__512_comb];
  assign p1_array_index_1077211_comb = literal_1076347[p1_array_index_1077177_comb];
  assign p1_array_index_1077212_comb = literal_1076349[p1_array_index_1077178_comb];
  assign p1_array_index_1077213_comb = literal_1076351[p1_array_index_1077179_comb];
  assign p1_array_index_1077214_comb = literal_1076353[p1_array_index_1077180_comb];
  assign p1_array_index_1077215_comb = literal_1076355[p1_array_index_1077181_comb];
  assign p1_res7__30_comb = literal_1076345[p1_res7__29_comb] ^ literal_1076347[p1_res7__28_comb] ^ literal_1076349[p1_res7__27_comb] ^ literal_1076351[p1_res7__26_comb] ^ literal_1076353[p1_res7__25_comb] ^ literal_1076355[p1_res7__24_comb] ^ p1_res7__23_comb ^ literal_1076358[p1_res7__22_comb] ^ p1_res7__21_comb ^ p1_array_index_1076723_comb ^ p1_array_index_1076700_comb ^ p1_array_index_1076675_comb ^ p1_array_index_1076648_comb ^ p1_array_index_1076619_comb ^ p1_array_index_1076587_comb ^ p1_array_index_1076572_comb;
  assign p1_res7__513_comb = p1_array_index_1077210_comb ^ p1_array_index_1077211_comb ^ p1_array_index_1077212_comb ^ p1_array_index_1077213_comb ^ p1_array_index_1077214_comb ^ p1_array_index_1077215_comb ^ p1_array_index_1077182_comb ^ literal_1076358[p1_array_index_1077199_comb] ^ p1_array_index_1077184_comb ^ literal_1076355[p1_array_index_1077201_comb] ^ literal_1076353[p1_array_index_1077186_comb] ^ literal_1076351[p1_array_index_1077187_comb] ^ literal_1076349[p1_array_index_1077188_comb] ^ literal_1076347[p1_array_index_1077189_comb] ^ literal_1076345[p1_array_index_1077190_comb] ^ p1_array_index_1077191_comb;
  assign p1_array_index_1077225_comb = literal_1076347[p1_res7__512_comb];
  assign p1_array_index_1077226_comb = literal_1076349[p1_array_index_1077177_comb];
  assign p1_array_index_1077227_comb = literal_1076351[p1_array_index_1077178_comb];
  assign p1_array_index_1077228_comb = literal_1076353[p1_array_index_1077179_comb];
  assign p1_array_index_1077229_comb = literal_1076355[p1_array_index_1077180_comb];
  assign p1_res7__31_comb = literal_1076345[p1_res7__30_comb] ^ literal_1076347[p1_res7__29_comb] ^ literal_1076349[p1_res7__28_comb] ^ literal_1076351[p1_res7__27_comb] ^ literal_1076353[p1_res7__26_comb] ^ literal_1076355[p1_res7__25_comb] ^ p1_res7__24_comb ^ literal_1076358[p1_res7__23_comb] ^ p1_res7__22_comb ^ p1_array_index_1076733_comb ^ p1_array_index_1076711_comb ^ p1_array_index_1076687_comb ^ p1_array_index_1076661_comb ^ p1_array_index_1076633_comb ^ p1_array_index_1076604_comb ^ p1_array_index_1076571_comb;
  assign p1_res7__514_comb = literal_1076345[p1_res7__513_comb] ^ p1_array_index_1077225_comb ^ p1_array_index_1077226_comb ^ p1_array_index_1077227_comb ^ p1_array_index_1077228_comb ^ p1_array_index_1077229_comb ^ p1_array_index_1077181_comb ^ literal_1076358[p1_array_index_1077182_comb] ^ p1_array_index_1077199_comb ^ literal_1076355[p1_array_index_1077184_comb] ^ literal_1076353[p1_array_index_1077201_comb] ^ literal_1076351[p1_array_index_1077186_comb] ^ literal_1076349[p1_array_index_1077187_comb] ^ literal_1076347[p1_array_index_1077188_comb] ^ literal_1076345[p1_array_index_1077189_comb] ^ p1_array_index_1077190_comb;
  assign p1_res__1_comb = {p1_res7__31_comb, p1_res7__30_comb, p1_res7__29_comb, p1_res7__28_comb, p1_res7__27_comb, p1_res7__26_comb, p1_res7__25_comb, p1_res7__24_comb, p1_res7__23_comb, p1_res7__22_comb, p1_res7__21_comb, p1_res7__20_comb, p1_res7__19_comb, p1_res7__18_comb, p1_res7__17_comb, p1_res7__16_comb};
  assign p1_array_index_1077239_comb = literal_1076347[p1_res7__513_comb];
  assign p1_array_index_1077240_comb = literal_1076349[p1_res7__512_comb];
  assign p1_array_index_1077241_comb = literal_1076351[p1_array_index_1077177_comb];
  assign p1_array_index_1077242_comb = literal_1076353[p1_array_index_1077178_comb];
  assign p1_array_index_1077243_comb = literal_1076355[p1_array_index_1077179_comb];
  assign p1_xor_1076773_comb = p1_res__1_comb ^ p0_key[255:128];
  assign p1_res7__515_comb = literal_1076345[p1_res7__514_comb] ^ p1_array_index_1077239_comb ^ p1_array_index_1077240_comb ^ p1_array_index_1077241_comb ^ p1_array_index_1077242_comb ^ p1_array_index_1077243_comb ^ p1_array_index_1077180_comb ^ literal_1076358[p1_array_index_1077181_comb] ^ p1_array_index_1077182_comb ^ literal_1076355[p1_array_index_1077199_comb] ^ literal_1076353[p1_array_index_1077184_comb] ^ literal_1076351[p1_array_index_1077201_comb] ^ literal_1076349[p1_array_index_1077186_comb] ^ literal_1076347[p1_array_index_1077187_comb] ^ literal_1076345[p1_array_index_1077188_comb] ^ p1_array_index_1077189_comb;
  assign p1_addedKey__43_comb = p1_xor_1076773_comb ^ 128'hb225_9a96_b4d8_8e0b_e769_0430_a44f_7f03;
  assign p1_array_index_1077254_comb = literal_1076349[p1_res7__513_comb];
  assign p1_array_index_1077255_comb = literal_1076351[p1_res7__512_comb];
  assign p1_array_index_1077256_comb = literal_1076353[p1_array_index_1077177_comb];
  assign p1_array_index_1077257_comb = literal_1076355[p1_array_index_1077178_comb];
  assign p1_res7__516_comb = literal_1076345[p1_res7__515_comb] ^ literal_1076347[p1_res7__514_comb] ^ p1_array_index_1077254_comb ^ p1_array_index_1077255_comb ^ p1_array_index_1077256_comb ^ p1_array_index_1077257_comb ^ p1_array_index_1077179_comb ^ literal_1076358[p1_array_index_1077180_comb] ^ p1_array_index_1077181_comb ^ p1_array_index_1077198_comb ^ literal_1076353[p1_array_index_1077199_comb] ^ literal_1076351[p1_array_index_1077184_comb] ^ literal_1076349[p1_array_index_1077201_comb] ^ literal_1076347[p1_array_index_1077186_comb] ^ literal_1076345[p1_array_index_1077187_comb] ^ p1_array_index_1077188_comb;
  assign p1_array_index_1076789_comb = arr[p1_addedKey__43_comb[127:120]];
  assign p1_array_index_1076790_comb = arr[p1_addedKey__43_comb[119:112]];
  assign p1_array_index_1076791_comb = arr[p1_addedKey__43_comb[111:104]];
  assign p1_array_index_1076792_comb = arr[p1_addedKey__43_comb[103:96]];
  assign p1_array_index_1076793_comb = arr[p1_addedKey__43_comb[95:88]];
  assign p1_array_index_1076794_comb = arr[p1_addedKey__43_comb[87:80]];
  assign p1_array_index_1076796_comb = arr[p1_addedKey__43_comb[71:64]];
  assign p1_array_index_1076798_comb = arr[p1_addedKey__43_comb[55:48]];
  assign p1_array_index_1076799_comb = arr[p1_addedKey__43_comb[47:40]];
  assign p1_array_index_1076800_comb = arr[p1_addedKey__43_comb[39:32]];
  assign p1_array_index_1076801_comb = arr[p1_addedKey__43_comb[31:24]];
  assign p1_array_index_1076802_comb = arr[p1_addedKey__43_comb[23:16]];
  assign p1_array_index_1076803_comb = arr[p1_addedKey__43_comb[15:8]];
  assign p1_array_index_1077267_comb = literal_1076349[p1_res7__514_comb];
  assign p1_array_index_1077268_comb = literal_1076351[p1_res7__513_comb];
  assign p1_array_index_1077269_comb = literal_1076353[p1_res7__512_comb];
  assign p1_array_index_1077270_comb = literal_1076355[p1_array_index_1077177_comb];
  assign p1_array_index_1076805_comb = literal_1076345[p1_array_index_1076789_comb];
  assign p1_array_index_1076806_comb = literal_1076347[p1_array_index_1076790_comb];
  assign p1_array_index_1076807_comb = literal_1076349[p1_array_index_1076791_comb];
  assign p1_array_index_1076808_comb = literal_1076351[p1_array_index_1076792_comb];
  assign p1_array_index_1076809_comb = literal_1076353[p1_array_index_1076793_comb];
  assign p1_array_index_1076810_comb = literal_1076355[p1_array_index_1076794_comb];
  assign p1_array_index_1076811_comb = arr[p1_addedKey__43_comb[79:72]];
  assign p1_array_index_1076813_comb = arr[p1_addedKey__43_comb[63:56]];
  assign p1_res7__517_comb = literal_1076345[p1_res7__516_comb] ^ literal_1076347[p1_res7__515_comb] ^ p1_array_index_1077267_comb ^ p1_array_index_1077268_comb ^ p1_array_index_1077269_comb ^ p1_array_index_1077270_comb ^ p1_array_index_1077178_comb ^ literal_1076358[p1_array_index_1077179_comb] ^ p1_array_index_1077180_comb ^ p1_array_index_1077215_comb ^ literal_1076353[p1_array_index_1077182_comb] ^ literal_1076351[p1_array_index_1077199_comb] ^ literal_1076349[p1_array_index_1077184_comb] ^ literal_1076347[p1_array_index_1077201_comb] ^ literal_1076345[p1_array_index_1077186_comb] ^ p1_array_index_1077187_comb;
  assign p1_res7__32_comb = p1_array_index_1076805_comb ^ p1_array_index_1076806_comb ^ p1_array_index_1076807_comb ^ p1_array_index_1076808_comb ^ p1_array_index_1076809_comb ^ p1_array_index_1076810_comb ^ p1_array_index_1076811_comb ^ literal_1076358[p1_array_index_1076796_comb] ^ p1_array_index_1076813_comb ^ literal_1076355[p1_array_index_1076798_comb] ^ literal_1076353[p1_array_index_1076799_comb] ^ literal_1076351[p1_array_index_1076800_comb] ^ literal_1076349[p1_array_index_1076801_comb] ^ literal_1076347[p1_array_index_1076802_comb] ^ literal_1076345[p1_array_index_1076803_comb] ^ arr[p1_addedKey__43_comb[7:0]];
  assign p1_array_index_1077281_comb = literal_1076351[p1_res7__514_comb];
  assign p1_array_index_1077282_comb = literal_1076353[p1_res7__513_comb];
  assign p1_array_index_1077283_comb = literal_1076355[p1_res7__512_comb];
  assign p1_array_index_1076822_comb = literal_1076345[p1_res7__32_comb];
  assign p1_array_index_1076823_comb = literal_1076347[p1_array_index_1076789_comb];
  assign p1_array_index_1076824_comb = literal_1076349[p1_array_index_1076790_comb];
  assign p1_array_index_1076825_comb = literal_1076351[p1_array_index_1076791_comb];
  assign p1_array_index_1076826_comb = literal_1076353[p1_array_index_1076792_comb];
  assign p1_array_index_1076827_comb = literal_1076355[p1_array_index_1076793_comb];
  assign p1_res7__518_comb = literal_1076345[p1_res7__517_comb] ^ literal_1076347[p1_res7__516_comb] ^ literal_1076349[p1_res7__515_comb] ^ p1_array_index_1077281_comb ^ p1_array_index_1077282_comb ^ p1_array_index_1077283_comb ^ p1_array_index_1077177_comb ^ literal_1076358[p1_array_index_1077178_comb] ^ p1_array_index_1077179_comb ^ p1_array_index_1077229_comb ^ p1_array_index_1077197_comb ^ literal_1076351[p1_array_index_1077182_comb] ^ literal_1076349[p1_array_index_1077199_comb] ^ literal_1076347[p1_array_index_1077184_comb] ^ literal_1076345[p1_array_index_1077201_comb] ^ p1_array_index_1077186_comb;
  assign p1_res7__33_comb = p1_array_index_1076822_comb ^ p1_array_index_1076823_comb ^ p1_array_index_1076824_comb ^ p1_array_index_1076825_comb ^ p1_array_index_1076826_comb ^ p1_array_index_1076827_comb ^ p1_array_index_1076794_comb ^ literal_1076358[p1_array_index_1076811_comb] ^ p1_array_index_1076796_comb ^ literal_1076355[p1_array_index_1076813_comb] ^ literal_1076353[p1_array_index_1076798_comb] ^ literal_1076351[p1_array_index_1076799_comb] ^ literal_1076349[p1_array_index_1076800_comb] ^ literal_1076347[p1_array_index_1076801_comb] ^ literal_1076345[p1_array_index_1076802_comb] ^ p1_array_index_1076803_comb;
  assign p1_array_index_1077293_comb = literal_1076351[p1_res7__515_comb];
  assign p1_array_index_1077294_comb = literal_1076353[p1_res7__514_comb];
  assign p1_array_index_1077295_comb = literal_1076355[p1_res7__513_comb];
  assign p1_array_index_1076837_comb = literal_1076347[p1_res7__32_comb];
  assign p1_array_index_1076838_comb = literal_1076349[p1_array_index_1076789_comb];
  assign p1_array_index_1076839_comb = literal_1076351[p1_array_index_1076790_comb];
  assign p1_array_index_1076840_comb = literal_1076353[p1_array_index_1076791_comb];
  assign p1_array_index_1076841_comb = literal_1076355[p1_array_index_1076792_comb];
  assign p1_res7__519_comb = literal_1076345[p1_res7__518_comb] ^ literal_1076347[p1_res7__517_comb] ^ literal_1076349[p1_res7__516_comb] ^ p1_array_index_1077293_comb ^ p1_array_index_1077294_comb ^ p1_array_index_1077295_comb ^ p1_res7__512_comb ^ literal_1076358[p1_array_index_1077177_comb] ^ p1_array_index_1077178_comb ^ p1_array_index_1077243_comb ^ p1_array_index_1077214_comb ^ literal_1076351[p1_array_index_1077181_comb] ^ literal_1076349[p1_array_index_1077182_comb] ^ literal_1076347[p1_array_index_1077199_comb] ^ literal_1076345[p1_array_index_1077184_comb] ^ p1_array_index_1077201_comb;
  assign p1_res7__34_comb = literal_1076345[p1_res7__33_comb] ^ p1_array_index_1076837_comb ^ p1_array_index_1076838_comb ^ p1_array_index_1076839_comb ^ p1_array_index_1076840_comb ^ p1_array_index_1076841_comb ^ p1_array_index_1076793_comb ^ literal_1076358[p1_array_index_1076794_comb] ^ p1_array_index_1076811_comb ^ literal_1076355[p1_array_index_1076796_comb] ^ literal_1076353[p1_array_index_1076813_comb] ^ literal_1076351[p1_array_index_1076798_comb] ^ literal_1076349[p1_array_index_1076799_comb] ^ literal_1076347[p1_array_index_1076800_comb] ^ literal_1076345[p1_array_index_1076801_comb] ^ p1_array_index_1076802_comb;
  assign p1_array_index_1077306_comb = literal_1076353[p1_res7__515_comb];
  assign p1_array_index_1077307_comb = literal_1076355[p1_res7__514_comb];
  assign p1_array_index_1076851_comb = literal_1076347[p1_res7__33_comb];
  assign p1_array_index_1076852_comb = literal_1076349[p1_res7__32_comb];
  assign p1_array_index_1076853_comb = literal_1076351[p1_array_index_1076789_comb];
  assign p1_array_index_1076854_comb = literal_1076353[p1_array_index_1076790_comb];
  assign p1_array_index_1076855_comb = literal_1076355[p1_array_index_1076791_comb];
  assign p1_res7__520_comb = literal_1076345[p1_res7__519_comb] ^ literal_1076347[p1_res7__518_comb] ^ literal_1076349[p1_res7__517_comb] ^ literal_1076351[p1_res7__516_comb] ^ p1_array_index_1077306_comb ^ p1_array_index_1077307_comb ^ p1_res7__513_comb ^ literal_1076358[p1_res7__512_comb] ^ p1_array_index_1077177_comb ^ p1_array_index_1077257_comb ^ p1_array_index_1077228_comb ^ p1_array_index_1077196_comb ^ literal_1076349[p1_array_index_1077181_comb] ^ literal_1076347[p1_array_index_1077182_comb] ^ literal_1076345[p1_array_index_1077199_comb] ^ p1_array_index_1077184_comb;
  assign p1_res7__35_comb = literal_1076345[p1_res7__34_comb] ^ p1_array_index_1076851_comb ^ p1_array_index_1076852_comb ^ p1_array_index_1076853_comb ^ p1_array_index_1076854_comb ^ p1_array_index_1076855_comb ^ p1_array_index_1076792_comb ^ literal_1076358[p1_array_index_1076793_comb] ^ p1_array_index_1076794_comb ^ literal_1076355[p1_array_index_1076811_comb] ^ literal_1076353[p1_array_index_1076796_comb] ^ literal_1076351[p1_array_index_1076813_comb] ^ literal_1076349[p1_array_index_1076798_comb] ^ literal_1076347[p1_array_index_1076799_comb] ^ literal_1076345[p1_array_index_1076800_comb] ^ p1_array_index_1076801_comb;
  assign p1_array_index_1077317_comb = literal_1076353[p1_res7__516_comb];
  assign p1_array_index_1077318_comb = literal_1076355[p1_res7__515_comb];
  assign p1_array_index_1076866_comb = literal_1076349[p1_res7__33_comb];
  assign p1_array_index_1076867_comb = literal_1076351[p1_res7__32_comb];
  assign p1_array_index_1076868_comb = literal_1076353[p1_array_index_1076789_comb];
  assign p1_array_index_1076869_comb = literal_1076355[p1_array_index_1076790_comb];
  assign p1_res7__521_comb = literal_1076345[p1_res7__520_comb] ^ literal_1076347[p1_res7__519_comb] ^ literal_1076349[p1_res7__518_comb] ^ literal_1076351[p1_res7__517_comb] ^ p1_array_index_1077317_comb ^ p1_array_index_1077318_comb ^ p1_res7__514_comb ^ literal_1076358[p1_res7__513_comb] ^ p1_res7__512_comb ^ p1_array_index_1077270_comb ^ p1_array_index_1077242_comb ^ p1_array_index_1077213_comb ^ literal_1076349[p1_array_index_1077180_comb] ^ literal_1076347[p1_array_index_1077181_comb] ^ literal_1076345[p1_array_index_1077182_comb] ^ p1_array_index_1077199_comb;
  assign p1_res7__36_comb = literal_1076345[p1_res7__35_comb] ^ literal_1076347[p1_res7__34_comb] ^ p1_array_index_1076866_comb ^ p1_array_index_1076867_comb ^ p1_array_index_1076868_comb ^ p1_array_index_1076869_comb ^ p1_array_index_1076791_comb ^ literal_1076358[p1_array_index_1076792_comb] ^ p1_array_index_1076793_comb ^ p1_array_index_1076810_comb ^ literal_1076353[p1_array_index_1076811_comb] ^ literal_1076351[p1_array_index_1076796_comb] ^ literal_1076349[p1_array_index_1076813_comb] ^ literal_1076347[p1_array_index_1076798_comb] ^ literal_1076345[p1_array_index_1076799_comb] ^ p1_array_index_1076800_comb;
  assign p1_array_index_1077329_comb = literal_1076355[p1_res7__516_comb];
  assign p1_array_index_1076879_comb = literal_1076349[p1_res7__34_comb];
  assign p1_array_index_1076880_comb = literal_1076351[p1_res7__33_comb];
  assign p1_array_index_1076881_comb = literal_1076353[p1_res7__32_comb];
  assign p1_array_index_1076882_comb = literal_1076355[p1_array_index_1076789_comb];
  assign p1_res7__522_comb = literal_1076345[p1_res7__521_comb] ^ literal_1076347[p1_res7__520_comb] ^ literal_1076349[p1_res7__519_comb] ^ literal_1076351[p1_res7__518_comb] ^ literal_1076353[p1_res7__517_comb] ^ p1_array_index_1077329_comb ^ p1_res7__515_comb ^ literal_1076358[p1_res7__514_comb] ^ p1_res7__513_comb ^ p1_array_index_1077283_comb ^ p1_array_index_1077256_comb ^ p1_array_index_1077227_comb ^ p1_array_index_1077195_comb ^ literal_1076347[p1_array_index_1077180_comb] ^ literal_1076345[p1_array_index_1077181_comb] ^ p1_array_index_1077182_comb;
  assign p1_res7__37_comb = literal_1076345[p1_res7__36_comb] ^ literal_1076347[p1_res7__35_comb] ^ p1_array_index_1076879_comb ^ p1_array_index_1076880_comb ^ p1_array_index_1076881_comb ^ p1_array_index_1076882_comb ^ p1_array_index_1076790_comb ^ literal_1076358[p1_array_index_1076791_comb] ^ p1_array_index_1076792_comb ^ p1_array_index_1076827_comb ^ literal_1076353[p1_array_index_1076794_comb] ^ literal_1076351[p1_array_index_1076811_comb] ^ literal_1076349[p1_array_index_1076796_comb] ^ literal_1076347[p1_array_index_1076813_comb] ^ literal_1076345[p1_array_index_1076798_comb] ^ p1_array_index_1076799_comb;
  assign p1_array_index_1077339_comb = literal_1076355[p1_res7__517_comb];
  assign p1_array_index_1076893_comb = literal_1076351[p1_res7__34_comb];
  assign p1_array_index_1076894_comb = literal_1076353[p1_res7__33_comb];
  assign p1_array_index_1076895_comb = literal_1076355[p1_res7__32_comb];
  assign p1_res7__523_comb = literal_1076345[p1_res7__522_comb] ^ literal_1076347[p1_res7__521_comb] ^ literal_1076349[p1_res7__520_comb] ^ literal_1076351[p1_res7__519_comb] ^ literal_1076353[p1_res7__518_comb] ^ p1_array_index_1077339_comb ^ p1_res7__516_comb ^ literal_1076358[p1_res7__515_comb] ^ p1_res7__514_comb ^ p1_array_index_1077295_comb ^ p1_array_index_1077269_comb ^ p1_array_index_1077241_comb ^ p1_array_index_1077212_comb ^ literal_1076347[p1_array_index_1077179_comb] ^ literal_1076345[p1_array_index_1077180_comb] ^ p1_array_index_1077181_comb;
  assign p1_res7__38_comb = literal_1076345[p1_res7__37_comb] ^ literal_1076347[p1_res7__36_comb] ^ literal_1076349[p1_res7__35_comb] ^ p1_array_index_1076893_comb ^ p1_array_index_1076894_comb ^ p1_array_index_1076895_comb ^ p1_array_index_1076789_comb ^ literal_1076358[p1_array_index_1076790_comb] ^ p1_array_index_1076791_comb ^ p1_array_index_1076841_comb ^ p1_array_index_1076809_comb ^ literal_1076351[p1_array_index_1076794_comb] ^ literal_1076349[p1_array_index_1076811_comb] ^ literal_1076347[p1_array_index_1076796_comb] ^ literal_1076345[p1_array_index_1076813_comb] ^ p1_array_index_1076798_comb;
  assign p1_array_index_1076905_comb = literal_1076351[p1_res7__35_comb];
  assign p1_array_index_1076906_comb = literal_1076353[p1_res7__34_comb];
  assign p1_array_index_1076907_comb = literal_1076355[p1_res7__33_comb];
  assign p1_res7__524_comb = literal_1076345[p1_res7__523_comb] ^ literal_1076347[p1_res7__522_comb] ^ literal_1076349[p1_res7__521_comb] ^ literal_1076351[p1_res7__520_comb] ^ literal_1076353[p1_res7__519_comb] ^ literal_1076355[p1_res7__518_comb] ^ p1_res7__517_comb ^ literal_1076358[p1_res7__516_comb] ^ p1_res7__515_comb ^ p1_array_index_1077307_comb ^ p1_array_index_1077282_comb ^ p1_array_index_1077255_comb ^ p1_array_index_1077226_comb ^ p1_array_index_1077194_comb ^ literal_1076345[p1_array_index_1077179_comb] ^ p1_array_index_1077180_comb;
  assign p1_res7__39_comb = literal_1076345[p1_res7__38_comb] ^ literal_1076347[p1_res7__37_comb] ^ literal_1076349[p1_res7__36_comb] ^ p1_array_index_1076905_comb ^ p1_array_index_1076906_comb ^ p1_array_index_1076907_comb ^ p1_res7__32_comb ^ literal_1076358[p1_array_index_1076789_comb] ^ p1_array_index_1076790_comb ^ p1_array_index_1076855_comb ^ p1_array_index_1076826_comb ^ literal_1076351[p1_array_index_1076793_comb] ^ literal_1076349[p1_array_index_1076794_comb] ^ literal_1076347[p1_array_index_1076811_comb] ^ literal_1076345[p1_array_index_1076796_comb] ^ p1_array_index_1076813_comb;
  assign p1_array_index_1076918_comb = literal_1076353[p1_res7__35_comb];
  assign p1_array_index_1076919_comb = literal_1076355[p1_res7__34_comb];
  assign p1_res7__525_comb = literal_1076345[p1_res7__524_comb] ^ literal_1076347[p1_res7__523_comb] ^ literal_1076349[p1_res7__522_comb] ^ literal_1076351[p1_res7__521_comb] ^ literal_1076353[p1_res7__520_comb] ^ literal_1076355[p1_res7__519_comb] ^ p1_res7__518_comb ^ literal_1076358[p1_res7__517_comb] ^ p1_res7__516_comb ^ p1_array_index_1077318_comb ^ p1_array_index_1077294_comb ^ p1_array_index_1077268_comb ^ p1_array_index_1077240_comb ^ p1_array_index_1077211_comb ^ literal_1076345[p1_array_index_1077178_comb] ^ p1_array_index_1077179_comb;
  assign p1_res7__40_comb = literal_1076345[p1_res7__39_comb] ^ literal_1076347[p1_res7__38_comb] ^ literal_1076349[p1_res7__37_comb] ^ literal_1076351[p1_res7__36_comb] ^ p1_array_index_1076918_comb ^ p1_array_index_1076919_comb ^ p1_res7__33_comb ^ literal_1076358[p1_res7__32_comb] ^ p1_array_index_1076789_comb ^ p1_array_index_1076869_comb ^ p1_array_index_1076840_comb ^ p1_array_index_1076808_comb ^ literal_1076349[p1_array_index_1076793_comb] ^ literal_1076347[p1_array_index_1076794_comb] ^ literal_1076345[p1_array_index_1076811_comb] ^ p1_array_index_1076796_comb;
  assign p1_array_index_1076929_comb = literal_1076353[p1_res7__36_comb];
  assign p1_array_index_1076930_comb = literal_1076355[p1_res7__35_comb];
  assign p1_res7__526_comb = literal_1076345[p1_res7__525_comb] ^ literal_1076347[p1_res7__524_comb] ^ literal_1076349[p1_res7__523_comb] ^ literal_1076351[p1_res7__522_comb] ^ literal_1076353[p1_res7__521_comb] ^ literal_1076355[p1_res7__520_comb] ^ p1_res7__519_comb ^ literal_1076358[p1_res7__518_comb] ^ p1_res7__517_comb ^ p1_array_index_1077329_comb ^ p1_array_index_1077306_comb ^ p1_array_index_1077281_comb ^ p1_array_index_1077254_comb ^ p1_array_index_1077225_comb ^ p1_array_index_1077193_comb ^ p1_array_index_1077178_comb;
  assign p1_res7__41_comb = literal_1076345[p1_res7__40_comb] ^ literal_1076347[p1_res7__39_comb] ^ literal_1076349[p1_res7__38_comb] ^ literal_1076351[p1_res7__37_comb] ^ p1_array_index_1076929_comb ^ p1_array_index_1076930_comb ^ p1_res7__34_comb ^ literal_1076358[p1_res7__33_comb] ^ p1_res7__32_comb ^ p1_array_index_1076882_comb ^ p1_array_index_1076854_comb ^ p1_array_index_1076825_comb ^ literal_1076349[p1_array_index_1076792_comb] ^ literal_1076347[p1_array_index_1076793_comb] ^ literal_1076345[p1_array_index_1076794_comb] ^ p1_array_index_1076811_comb;
  assign p1_array_index_1076941_comb = literal_1076355[p1_res7__36_comb];
  assign p1_res7__527_comb = literal_1076345[p1_res7__526_comb] ^ literal_1076347[p1_res7__525_comb] ^ literal_1076349[p1_res7__524_comb] ^ literal_1076351[p1_res7__523_comb] ^ literal_1076353[p1_res7__522_comb] ^ literal_1076355[p1_res7__521_comb] ^ p1_res7__520_comb ^ literal_1076358[p1_res7__519_comb] ^ p1_res7__518_comb ^ p1_array_index_1077339_comb ^ p1_array_index_1077317_comb ^ p1_array_index_1077293_comb ^ p1_array_index_1077267_comb ^ p1_array_index_1077239_comb ^ p1_array_index_1077210_comb ^ p1_array_index_1077177_comb;
  assign p1_res7__42_comb = literal_1076345[p1_res7__41_comb] ^ literal_1076347[p1_res7__40_comb] ^ literal_1076349[p1_res7__39_comb] ^ literal_1076351[p1_res7__38_comb] ^ literal_1076353[p1_res7__37_comb] ^ p1_array_index_1076941_comb ^ p1_res7__35_comb ^ literal_1076358[p1_res7__34_comb] ^ p1_res7__33_comb ^ p1_array_index_1076895_comb ^ p1_array_index_1076868_comb ^ p1_array_index_1076839_comb ^ p1_array_index_1076807_comb ^ literal_1076347[p1_array_index_1076792_comb] ^ literal_1076345[p1_array_index_1076793_comb] ^ p1_array_index_1076794_comb;
  assign p1_res__32_comb = {p1_res7__527_comb, p1_res7__526_comb, p1_res7__525_comb, p1_res7__524_comb, p1_res7__523_comb, p1_res7__522_comb, p1_res7__521_comb, p1_res7__520_comb, p1_res7__519_comb, p1_res7__518_comb, p1_res7__517_comb, p1_res7__516_comb, p1_res7__515_comb, p1_res7__514_comb, p1_res7__513_comb, p1_res7__512_comb};
  assign p1_array_index_1076951_comb = literal_1076355[p1_res7__37_comb];
  assign p1_addedKey__33_comb = p0_key[127:0] ^ p1_res__32_comb;
  assign p1_res7__43_comb = literal_1076345[p1_res7__42_comb] ^ literal_1076347[p1_res7__41_comb] ^ literal_1076349[p1_res7__40_comb] ^ literal_1076351[p1_res7__39_comb] ^ literal_1076353[p1_res7__38_comb] ^ p1_array_index_1076951_comb ^ p1_res7__36_comb ^ literal_1076358[p1_res7__35_comb] ^ p1_res7__34_comb ^ p1_array_index_1076907_comb ^ p1_array_index_1076881_comb ^ p1_array_index_1076853_comb ^ p1_array_index_1076824_comb ^ literal_1076347[p1_array_index_1076791_comb] ^ literal_1076345[p1_array_index_1076792_comb] ^ p1_array_index_1076793_comb;
  assign p1_array_index_1077393_comb = arr[p1_addedKey__33_comb[127:120]];
  assign p1_array_index_1077394_comb = arr[p1_addedKey__33_comb[119:112]];
  assign p1_array_index_1077395_comb = arr[p1_addedKey__33_comb[111:104]];
  assign p1_array_index_1077396_comb = arr[p1_addedKey__33_comb[103:96]];
  assign p1_array_index_1077397_comb = arr[p1_addedKey__33_comb[95:88]];
  assign p1_array_index_1077398_comb = arr[p1_addedKey__33_comb[87:80]];
  assign p1_array_index_1077400_comb = arr[p1_addedKey__33_comb[71:64]];
  assign p1_array_index_1077402_comb = arr[p1_addedKey__33_comb[55:48]];
  assign p1_array_index_1077403_comb = arr[p1_addedKey__33_comb[47:40]];
  assign p1_array_index_1077404_comb = arr[p1_addedKey__33_comb[39:32]];
  assign p1_array_index_1077405_comb = arr[p1_addedKey__33_comb[31:24]];
  assign p1_array_index_1077406_comb = arr[p1_addedKey__33_comb[23:16]];
  assign p1_array_index_1077407_comb = arr[p1_addedKey__33_comb[15:8]];
  assign p1_res7__44_comb = literal_1076345[p1_res7__43_comb] ^ literal_1076347[p1_res7__42_comb] ^ literal_1076349[p1_res7__41_comb] ^ literal_1076351[p1_res7__40_comb] ^ literal_1076353[p1_res7__39_comb] ^ literal_1076355[p1_res7__38_comb] ^ p1_res7__37_comb ^ literal_1076358[p1_res7__36_comb] ^ p1_res7__35_comb ^ p1_array_index_1076919_comb ^ p1_array_index_1076894_comb ^ p1_array_index_1076867_comb ^ p1_array_index_1076838_comb ^ p1_array_index_1076806_comb ^ literal_1076345[p1_array_index_1076791_comb] ^ p1_array_index_1076792_comb;
  assign p1_array_index_1077409_comb = literal_1076345[p1_array_index_1077393_comb];
  assign p1_array_index_1077410_comb = literal_1076347[p1_array_index_1077394_comb];
  assign p1_array_index_1077411_comb = literal_1076349[p1_array_index_1077395_comb];
  assign p1_array_index_1077412_comb = literal_1076351[p1_array_index_1077396_comb];
  assign p1_array_index_1077413_comb = literal_1076353[p1_array_index_1077397_comb];
  assign p1_array_index_1077414_comb = literal_1076355[p1_array_index_1077398_comb];
  assign p1_array_index_1077415_comb = arr[p1_addedKey__33_comb[79:72]];
  assign p1_array_index_1077417_comb = arr[p1_addedKey__33_comb[63:56]];
  assign p1_res7__528_comb = p1_array_index_1077409_comb ^ p1_array_index_1077410_comb ^ p1_array_index_1077411_comb ^ p1_array_index_1077412_comb ^ p1_array_index_1077413_comb ^ p1_array_index_1077414_comb ^ p1_array_index_1077415_comb ^ literal_1076358[p1_array_index_1077400_comb] ^ p1_array_index_1077417_comb ^ literal_1076355[p1_array_index_1077402_comb] ^ literal_1076353[p1_array_index_1077403_comb] ^ literal_1076351[p1_array_index_1077404_comb] ^ literal_1076349[p1_array_index_1077405_comb] ^ literal_1076347[p1_array_index_1077406_comb] ^ literal_1076345[p1_array_index_1077407_comb] ^ arr[p1_addedKey__33_comb[7:0]];
  assign p1_res7__45_comb = literal_1076345[p1_res7__44_comb] ^ literal_1076347[p1_res7__43_comb] ^ literal_1076349[p1_res7__42_comb] ^ literal_1076351[p1_res7__41_comb] ^ literal_1076353[p1_res7__40_comb] ^ literal_1076355[p1_res7__39_comb] ^ p1_res7__38_comb ^ literal_1076358[p1_res7__37_comb] ^ p1_res7__36_comb ^ p1_array_index_1076930_comb ^ p1_array_index_1076906_comb ^ p1_array_index_1076880_comb ^ p1_array_index_1076852_comb ^ p1_array_index_1076823_comb ^ literal_1076345[p1_array_index_1076790_comb] ^ p1_array_index_1076791_comb;
  assign p1_array_index_1077426_comb = literal_1076345[p1_res7__528_comb];
  assign p1_array_index_1077427_comb = literal_1076347[p1_array_index_1077393_comb];
  assign p1_array_index_1077428_comb = literal_1076349[p1_array_index_1077394_comb];
  assign p1_array_index_1077429_comb = literal_1076351[p1_array_index_1077395_comb];
  assign p1_array_index_1077430_comb = literal_1076353[p1_array_index_1077396_comb];
  assign p1_array_index_1077431_comb = literal_1076355[p1_array_index_1077397_comb];
  assign p1_res7__529_comb = p1_array_index_1077426_comb ^ p1_array_index_1077427_comb ^ p1_array_index_1077428_comb ^ p1_array_index_1077429_comb ^ p1_array_index_1077430_comb ^ p1_array_index_1077431_comb ^ p1_array_index_1077398_comb ^ literal_1076358[p1_array_index_1077415_comb] ^ p1_array_index_1077400_comb ^ literal_1076355[p1_array_index_1077417_comb] ^ literal_1076353[p1_array_index_1077402_comb] ^ literal_1076351[p1_array_index_1077403_comb] ^ literal_1076349[p1_array_index_1077404_comb] ^ literal_1076347[p1_array_index_1077405_comb] ^ literal_1076345[p1_array_index_1077406_comb] ^ p1_array_index_1077407_comb;
  assign p1_res7__46_comb = literal_1076345[p1_res7__45_comb] ^ literal_1076347[p1_res7__44_comb] ^ literal_1076349[p1_res7__43_comb] ^ literal_1076351[p1_res7__42_comb] ^ literal_1076353[p1_res7__41_comb] ^ literal_1076355[p1_res7__40_comb] ^ p1_res7__39_comb ^ literal_1076358[p1_res7__38_comb] ^ p1_res7__37_comb ^ p1_array_index_1076941_comb ^ p1_array_index_1076918_comb ^ p1_array_index_1076893_comb ^ p1_array_index_1076866_comb ^ p1_array_index_1076837_comb ^ p1_array_index_1076805_comb ^ p1_array_index_1076790_comb;
  assign p1_array_index_1077441_comb = literal_1076347[p1_res7__528_comb];
  assign p1_array_index_1077442_comb = literal_1076349[p1_array_index_1077393_comb];
  assign p1_array_index_1077443_comb = literal_1076351[p1_array_index_1077394_comb];
  assign p1_array_index_1077444_comb = literal_1076353[p1_array_index_1077395_comb];
  assign p1_array_index_1077445_comb = literal_1076355[p1_array_index_1077396_comb];
  assign p1_res7__530_comb = literal_1076345[p1_res7__529_comb] ^ p1_array_index_1077441_comb ^ p1_array_index_1077442_comb ^ p1_array_index_1077443_comb ^ p1_array_index_1077444_comb ^ p1_array_index_1077445_comb ^ p1_array_index_1077397_comb ^ literal_1076358[p1_array_index_1077398_comb] ^ p1_array_index_1077415_comb ^ literal_1076355[p1_array_index_1077400_comb] ^ literal_1076353[p1_array_index_1077417_comb] ^ literal_1076351[p1_array_index_1077402_comb] ^ literal_1076349[p1_array_index_1077403_comb] ^ literal_1076347[p1_array_index_1077404_comb] ^ literal_1076345[p1_array_index_1077405_comb] ^ p1_array_index_1077406_comb;
  assign p1_res7__47_comb = literal_1076345[p1_res7__46_comb] ^ literal_1076347[p1_res7__45_comb] ^ literal_1076349[p1_res7__44_comb] ^ literal_1076351[p1_res7__43_comb] ^ literal_1076353[p1_res7__42_comb] ^ literal_1076355[p1_res7__41_comb] ^ p1_res7__40_comb ^ literal_1076358[p1_res7__39_comb] ^ p1_res7__38_comb ^ p1_array_index_1076951_comb ^ p1_array_index_1076929_comb ^ p1_array_index_1076905_comb ^ p1_array_index_1076879_comb ^ p1_array_index_1076851_comb ^ p1_array_index_1076822_comb ^ p1_array_index_1076789_comb;
  assign p1_array_index_1077455_comb = literal_1076347[p1_res7__529_comb];
  assign p1_array_index_1077456_comb = literal_1076349[p1_res7__528_comb];
  assign p1_array_index_1077457_comb = literal_1076351[p1_array_index_1077393_comb];
  assign p1_array_index_1077458_comb = literal_1076353[p1_array_index_1077394_comb];
  assign p1_array_index_1077459_comb = literal_1076355[p1_array_index_1077395_comb];
  assign p1_res__2_comb = {p1_res7__47_comb, p1_res7__46_comb, p1_res7__45_comb, p1_res7__44_comb, p1_res7__43_comb, p1_res7__42_comb, p1_res7__41_comb, p1_res7__40_comb, p1_res7__39_comb, p1_res7__38_comb, p1_res7__37_comb, p1_res7__36_comb, p1_res7__35_comb, p1_res7__34_comb, p1_res7__33_comb, p1_res7__32_comb};
  assign p1_res7__531_comb = literal_1076345[p1_res7__530_comb] ^ p1_array_index_1077455_comb ^ p1_array_index_1077456_comb ^ p1_array_index_1077457_comb ^ p1_array_index_1077458_comb ^ p1_array_index_1077459_comb ^ p1_array_index_1077396_comb ^ literal_1076358[p1_array_index_1077397_comb] ^ p1_array_index_1077398_comb ^ literal_1076355[p1_array_index_1077415_comb] ^ literal_1076353[p1_array_index_1077400_comb] ^ literal_1076351[p1_array_index_1077417_comb] ^ literal_1076349[p1_array_index_1077402_comb] ^ literal_1076347[p1_array_index_1077403_comb] ^ literal_1076345[p1_array_index_1077404_comb] ^ p1_array_index_1077405_comb;
  assign p1_xor_1076991_comb = p1_res__2_comb ^ p1_xor_1076555_comb;
  assign p1_array_index_1077470_comb = literal_1076349[p1_res7__529_comb];
  assign p1_array_index_1077471_comb = literal_1076351[p1_res7__528_comb];
  assign p1_array_index_1077472_comb = literal_1076353[p1_array_index_1077393_comb];
  assign p1_array_index_1077473_comb = literal_1076355[p1_array_index_1077394_comb];
  assign p1_addedKey__44_comb = p1_xor_1076991_comb ^ 128'h7bcd_1b0b_73e3_2ba5_b79c_b140_f255_1504;
  assign p1_res7__532_comb = literal_1076345[p1_res7__531_comb] ^ literal_1076347[p1_res7__530_comb] ^ p1_array_index_1077470_comb ^ p1_array_index_1077471_comb ^ p1_array_index_1077472_comb ^ p1_array_index_1077473_comb ^ p1_array_index_1077395_comb ^ literal_1076358[p1_array_index_1077396_comb] ^ p1_array_index_1077397_comb ^ p1_array_index_1077414_comb ^ literal_1076353[p1_array_index_1077415_comb] ^ literal_1076351[p1_array_index_1077400_comb] ^ literal_1076349[p1_array_index_1077417_comb] ^ literal_1076347[p1_array_index_1077402_comb] ^ literal_1076345[p1_array_index_1077403_comb] ^ p1_array_index_1077404_comb;
  assign p1_array_index_1077483_comb = literal_1076349[p1_res7__530_comb];
  assign p1_array_index_1077484_comb = literal_1076351[p1_res7__529_comb];
  assign p1_array_index_1077485_comb = literal_1076353[p1_res7__528_comb];
  assign p1_array_index_1077486_comb = literal_1076355[p1_array_index_1077393_comb];
  assign p1_array_index_1077007_comb = arr[p1_addedKey__44_comb[127:120]];
  assign p1_array_index_1077008_comb = arr[p1_addedKey__44_comb[119:112]];
  assign p1_array_index_1077009_comb = arr[p1_addedKey__44_comb[111:104]];
  assign p1_array_index_1077010_comb = arr[p1_addedKey__44_comb[103:96]];
  assign p1_array_index_1077011_comb = arr[p1_addedKey__44_comb[95:88]];
  assign p1_array_index_1077012_comb = arr[p1_addedKey__44_comb[87:80]];
  assign p1_array_index_1077014_comb = arr[p1_addedKey__44_comb[71:64]];
  assign p1_array_index_1077016_comb = arr[p1_addedKey__44_comb[55:48]];
  assign p1_array_index_1077017_comb = arr[p1_addedKey__44_comb[47:40]];
  assign p1_array_index_1077018_comb = arr[p1_addedKey__44_comb[39:32]];
  assign p1_array_index_1077019_comb = arr[p1_addedKey__44_comb[31:24]];
  assign p1_array_index_1077020_comb = arr[p1_addedKey__44_comb[23:16]];
  assign p1_array_index_1077021_comb = arr[p1_addedKey__44_comb[15:8]];
  assign p1_res7__533_comb = literal_1076345[p1_res7__532_comb] ^ literal_1076347[p1_res7__531_comb] ^ p1_array_index_1077483_comb ^ p1_array_index_1077484_comb ^ p1_array_index_1077485_comb ^ p1_array_index_1077486_comb ^ p1_array_index_1077394_comb ^ literal_1076358[p1_array_index_1077395_comb] ^ p1_array_index_1077396_comb ^ p1_array_index_1077431_comb ^ literal_1076353[p1_array_index_1077398_comb] ^ literal_1076351[p1_array_index_1077415_comb] ^ literal_1076349[p1_array_index_1077400_comb] ^ literal_1076347[p1_array_index_1077417_comb] ^ literal_1076345[p1_array_index_1077402_comb] ^ p1_array_index_1077403_comb;
  assign p1_array_index_1077023_comb = literal_1076345[p1_array_index_1077007_comb];
  assign p1_array_index_1077024_comb = literal_1076347[p1_array_index_1077008_comb];
  assign p1_array_index_1077025_comb = literal_1076349[p1_array_index_1077009_comb];
  assign p1_array_index_1077026_comb = literal_1076351[p1_array_index_1077010_comb];
  assign p1_array_index_1077027_comb = literal_1076353[p1_array_index_1077011_comb];
  assign p1_array_index_1077028_comb = literal_1076355[p1_array_index_1077012_comb];
  assign p1_array_index_1077029_comb = arr[p1_addedKey__44_comb[79:72]];
  assign p1_array_index_1077031_comb = arr[p1_addedKey__44_comb[63:56]];
  assign p1_array_index_1077497_comb = literal_1076351[p1_res7__530_comb];
  assign p1_array_index_1077498_comb = literal_1076353[p1_res7__529_comb];
  assign p1_array_index_1077499_comb = literal_1076355[p1_res7__528_comb];
  assign p1_res7__48_comb = p1_array_index_1077023_comb ^ p1_array_index_1077024_comb ^ p1_array_index_1077025_comb ^ p1_array_index_1077026_comb ^ p1_array_index_1077027_comb ^ p1_array_index_1077028_comb ^ p1_array_index_1077029_comb ^ literal_1076358[p1_array_index_1077014_comb] ^ p1_array_index_1077031_comb ^ literal_1076355[p1_array_index_1077016_comb] ^ literal_1076353[p1_array_index_1077017_comb] ^ literal_1076351[p1_array_index_1077018_comb] ^ literal_1076349[p1_array_index_1077019_comb] ^ literal_1076347[p1_array_index_1077020_comb] ^ literal_1076345[p1_array_index_1077021_comb] ^ arr[p1_addedKey__44_comb[7:0]];
  assign p1_res7__534_comb = literal_1076345[p1_res7__533_comb] ^ literal_1076347[p1_res7__532_comb] ^ literal_1076349[p1_res7__531_comb] ^ p1_array_index_1077497_comb ^ p1_array_index_1077498_comb ^ p1_array_index_1077499_comb ^ p1_array_index_1077393_comb ^ literal_1076358[p1_array_index_1077394_comb] ^ p1_array_index_1077395_comb ^ p1_array_index_1077445_comb ^ p1_array_index_1077413_comb ^ literal_1076351[p1_array_index_1077398_comb] ^ literal_1076349[p1_array_index_1077415_comb] ^ literal_1076347[p1_array_index_1077400_comb] ^ literal_1076345[p1_array_index_1077417_comb] ^ p1_array_index_1077402_comb;
  assign p1_array_index_1077040_comb = literal_1076345[p1_res7__48_comb];
  assign p1_array_index_1077041_comb = literal_1076347[p1_array_index_1077007_comb];
  assign p1_array_index_1077042_comb = literal_1076349[p1_array_index_1077008_comb];
  assign p1_array_index_1077043_comb = literal_1076351[p1_array_index_1077009_comb];
  assign p1_array_index_1077044_comb = literal_1076353[p1_array_index_1077010_comb];
  assign p1_array_index_1077045_comb = literal_1076355[p1_array_index_1077011_comb];
  assign p1_array_index_1077509_comb = literal_1076351[p1_res7__531_comb];
  assign p1_array_index_1077510_comb = literal_1076353[p1_res7__530_comb];
  assign p1_array_index_1077511_comb = literal_1076355[p1_res7__529_comb];
  assign p1_res7__49_comb = p1_array_index_1077040_comb ^ p1_array_index_1077041_comb ^ p1_array_index_1077042_comb ^ p1_array_index_1077043_comb ^ p1_array_index_1077044_comb ^ p1_array_index_1077045_comb ^ p1_array_index_1077012_comb ^ literal_1076358[p1_array_index_1077029_comb] ^ p1_array_index_1077014_comb ^ literal_1076355[p1_array_index_1077031_comb] ^ literal_1076353[p1_array_index_1077016_comb] ^ literal_1076351[p1_array_index_1077017_comb] ^ literal_1076349[p1_array_index_1077018_comb] ^ literal_1076347[p1_array_index_1077019_comb] ^ literal_1076345[p1_array_index_1077020_comb] ^ p1_array_index_1077021_comb;
  assign p1_res7__535_comb = literal_1076345[p1_res7__534_comb] ^ literal_1076347[p1_res7__533_comb] ^ literal_1076349[p1_res7__532_comb] ^ p1_array_index_1077509_comb ^ p1_array_index_1077510_comb ^ p1_array_index_1077511_comb ^ p1_res7__528_comb ^ literal_1076358[p1_array_index_1077393_comb] ^ p1_array_index_1077394_comb ^ p1_array_index_1077459_comb ^ p1_array_index_1077430_comb ^ literal_1076351[p1_array_index_1077397_comb] ^ literal_1076349[p1_array_index_1077398_comb] ^ literal_1076347[p1_array_index_1077415_comb] ^ literal_1076345[p1_array_index_1077400_comb] ^ p1_array_index_1077417_comb;
  assign p1_array_index_1077055_comb = literal_1076347[p1_res7__48_comb];
  assign p1_array_index_1077056_comb = literal_1076349[p1_array_index_1077007_comb];
  assign p1_array_index_1077057_comb = literal_1076351[p1_array_index_1077008_comb];
  assign p1_array_index_1077058_comb = literal_1076353[p1_array_index_1077009_comb];
  assign p1_array_index_1077059_comb = literal_1076355[p1_array_index_1077010_comb];
  assign p1_array_index_1077522_comb = literal_1076353[p1_res7__531_comb];
  assign p1_array_index_1077523_comb = literal_1076355[p1_res7__530_comb];
  assign p1_res7__50_comb = literal_1076345[p1_res7__49_comb] ^ p1_array_index_1077055_comb ^ p1_array_index_1077056_comb ^ p1_array_index_1077057_comb ^ p1_array_index_1077058_comb ^ p1_array_index_1077059_comb ^ p1_array_index_1077011_comb ^ literal_1076358[p1_array_index_1077012_comb] ^ p1_array_index_1077029_comb ^ literal_1076355[p1_array_index_1077014_comb] ^ literal_1076353[p1_array_index_1077031_comb] ^ literal_1076351[p1_array_index_1077016_comb] ^ literal_1076349[p1_array_index_1077017_comb] ^ literal_1076347[p1_array_index_1077018_comb] ^ literal_1076345[p1_array_index_1077019_comb] ^ p1_array_index_1077020_comb;
  assign p1_res7__536_comb = literal_1076345[p1_res7__535_comb] ^ literal_1076347[p1_res7__534_comb] ^ literal_1076349[p1_res7__533_comb] ^ literal_1076351[p1_res7__532_comb] ^ p1_array_index_1077522_comb ^ p1_array_index_1077523_comb ^ p1_res7__529_comb ^ literal_1076358[p1_res7__528_comb] ^ p1_array_index_1077393_comb ^ p1_array_index_1077473_comb ^ p1_array_index_1077444_comb ^ p1_array_index_1077412_comb ^ literal_1076349[p1_array_index_1077397_comb] ^ literal_1076347[p1_array_index_1077398_comb] ^ literal_1076345[p1_array_index_1077415_comb] ^ p1_array_index_1077400_comb;
  assign p1_array_index_1077069_comb = literal_1076347[p1_res7__49_comb];
  assign p1_array_index_1077070_comb = literal_1076349[p1_res7__48_comb];
  assign p1_array_index_1077071_comb = literal_1076351[p1_array_index_1077007_comb];
  assign p1_array_index_1077072_comb = literal_1076353[p1_array_index_1077008_comb];
  assign p1_array_index_1077073_comb = literal_1076355[p1_array_index_1077009_comb];
  assign p1_array_index_1077533_comb = literal_1076353[p1_res7__532_comb];
  assign p1_array_index_1077534_comb = literal_1076355[p1_res7__531_comb];
  assign p1_res7__51_comb = literal_1076345[p1_res7__50_comb] ^ p1_array_index_1077069_comb ^ p1_array_index_1077070_comb ^ p1_array_index_1077071_comb ^ p1_array_index_1077072_comb ^ p1_array_index_1077073_comb ^ p1_array_index_1077010_comb ^ literal_1076358[p1_array_index_1077011_comb] ^ p1_array_index_1077012_comb ^ literal_1076355[p1_array_index_1077029_comb] ^ literal_1076353[p1_array_index_1077014_comb] ^ literal_1076351[p1_array_index_1077031_comb] ^ literal_1076349[p1_array_index_1077016_comb] ^ literal_1076347[p1_array_index_1077017_comb] ^ literal_1076345[p1_array_index_1077018_comb] ^ p1_array_index_1077019_comb;
  assign p1_res7__537_comb = literal_1076345[p1_res7__536_comb] ^ literal_1076347[p1_res7__535_comb] ^ literal_1076349[p1_res7__534_comb] ^ literal_1076351[p1_res7__533_comb] ^ p1_array_index_1077533_comb ^ p1_array_index_1077534_comb ^ p1_res7__530_comb ^ literal_1076358[p1_res7__529_comb] ^ p1_res7__528_comb ^ p1_array_index_1077486_comb ^ p1_array_index_1077458_comb ^ p1_array_index_1077429_comb ^ literal_1076349[p1_array_index_1077396_comb] ^ literal_1076347[p1_array_index_1077397_comb] ^ literal_1076345[p1_array_index_1077398_comb] ^ p1_array_index_1077415_comb;
  assign p1_array_index_1077084_comb = literal_1076349[p1_res7__49_comb];
  assign p1_array_index_1077085_comb = literal_1076351[p1_res7__48_comb];
  assign p1_array_index_1077086_comb = literal_1076353[p1_array_index_1077007_comb];
  assign p1_array_index_1077087_comb = literal_1076355[p1_array_index_1077008_comb];
  assign p1_array_index_1077545_comb = literal_1076355[p1_res7__532_comb];
  assign p1_res7__52_comb = literal_1076345[p1_res7__51_comb] ^ literal_1076347[p1_res7__50_comb] ^ p1_array_index_1077084_comb ^ p1_array_index_1077085_comb ^ p1_array_index_1077086_comb ^ p1_array_index_1077087_comb ^ p1_array_index_1077009_comb ^ literal_1076358[p1_array_index_1077010_comb] ^ p1_array_index_1077011_comb ^ p1_array_index_1077028_comb ^ literal_1076353[p1_array_index_1077029_comb] ^ literal_1076351[p1_array_index_1077014_comb] ^ literal_1076349[p1_array_index_1077031_comb] ^ literal_1076347[p1_array_index_1077016_comb] ^ literal_1076345[p1_array_index_1077017_comb] ^ p1_array_index_1077018_comb;
  assign p1_res7__538_comb = literal_1076345[p1_res7__537_comb] ^ literal_1076347[p1_res7__536_comb] ^ literal_1076349[p1_res7__535_comb] ^ literal_1076351[p1_res7__534_comb] ^ literal_1076353[p1_res7__533_comb] ^ p1_array_index_1077545_comb ^ p1_res7__531_comb ^ literal_1076358[p1_res7__530_comb] ^ p1_res7__529_comb ^ p1_array_index_1077499_comb ^ p1_array_index_1077472_comb ^ p1_array_index_1077443_comb ^ p1_array_index_1077411_comb ^ literal_1076347[p1_array_index_1077396_comb] ^ literal_1076345[p1_array_index_1077397_comb] ^ p1_array_index_1077398_comb;
  assign p1_array_index_1077097_comb = literal_1076349[p1_res7__50_comb];
  assign p1_array_index_1077098_comb = literal_1076351[p1_res7__49_comb];
  assign p1_array_index_1077099_comb = literal_1076353[p1_res7__48_comb];
  assign p1_array_index_1077100_comb = literal_1076355[p1_array_index_1077007_comb];
  assign p1_array_index_1077555_comb = literal_1076355[p1_res7__533_comb];
  assign p1_res7__53_comb = literal_1076345[p1_res7__52_comb] ^ literal_1076347[p1_res7__51_comb] ^ p1_array_index_1077097_comb ^ p1_array_index_1077098_comb ^ p1_array_index_1077099_comb ^ p1_array_index_1077100_comb ^ p1_array_index_1077008_comb ^ literal_1076358[p1_array_index_1077009_comb] ^ p1_array_index_1077010_comb ^ p1_array_index_1077045_comb ^ literal_1076353[p1_array_index_1077012_comb] ^ literal_1076351[p1_array_index_1077029_comb] ^ literal_1076349[p1_array_index_1077014_comb] ^ literal_1076347[p1_array_index_1077031_comb] ^ literal_1076345[p1_array_index_1077016_comb] ^ p1_array_index_1077017_comb;
  assign p1_res7__539_comb = literal_1076345[p1_res7__538_comb] ^ literal_1076347[p1_res7__537_comb] ^ literal_1076349[p1_res7__536_comb] ^ literal_1076351[p1_res7__535_comb] ^ literal_1076353[p1_res7__534_comb] ^ p1_array_index_1077555_comb ^ p1_res7__532_comb ^ literal_1076358[p1_res7__531_comb] ^ p1_res7__530_comb ^ p1_array_index_1077511_comb ^ p1_array_index_1077485_comb ^ p1_array_index_1077457_comb ^ p1_array_index_1077428_comb ^ literal_1076347[p1_array_index_1077395_comb] ^ literal_1076345[p1_array_index_1077396_comb] ^ p1_array_index_1077397_comb;
  assign p1_array_index_1077111_comb = literal_1076351[p1_res7__50_comb];
  assign p1_array_index_1077112_comb = literal_1076353[p1_res7__49_comb];
  assign p1_array_index_1077113_comb = literal_1076355[p1_res7__48_comb];
  assign p1_res7__54_comb = literal_1076345[p1_res7__53_comb] ^ literal_1076347[p1_res7__52_comb] ^ literal_1076349[p1_res7__51_comb] ^ p1_array_index_1077111_comb ^ p1_array_index_1077112_comb ^ p1_array_index_1077113_comb ^ p1_array_index_1077007_comb ^ literal_1076358[p1_array_index_1077008_comb] ^ p1_array_index_1077009_comb ^ p1_array_index_1077059_comb ^ p1_array_index_1077027_comb ^ literal_1076351[p1_array_index_1077012_comb] ^ literal_1076349[p1_array_index_1077029_comb] ^ literal_1076347[p1_array_index_1077014_comb] ^ literal_1076345[p1_array_index_1077031_comb] ^ p1_array_index_1077016_comb;
  assign p1_res7__540_comb = literal_1076345[p1_res7__539_comb] ^ literal_1076347[p1_res7__538_comb] ^ literal_1076349[p1_res7__537_comb] ^ literal_1076351[p1_res7__536_comb] ^ literal_1076353[p1_res7__535_comb] ^ literal_1076355[p1_res7__534_comb] ^ p1_res7__533_comb ^ literal_1076358[p1_res7__532_comb] ^ p1_res7__531_comb ^ p1_array_index_1077523_comb ^ p1_array_index_1077498_comb ^ p1_array_index_1077471_comb ^ p1_array_index_1077442_comb ^ p1_array_index_1077410_comb ^ literal_1076345[p1_array_index_1077395_comb] ^ p1_array_index_1077396_comb;
  assign p1_array_index_1077123_comb = literal_1076351[p1_res7__51_comb];
  assign p1_array_index_1077124_comb = literal_1076353[p1_res7__50_comb];
  assign p1_array_index_1077125_comb = literal_1076355[p1_res7__49_comb];
  assign p1_res7__55_comb = literal_1076345[p1_res7__54_comb] ^ literal_1076347[p1_res7__53_comb] ^ literal_1076349[p1_res7__52_comb] ^ p1_array_index_1077123_comb ^ p1_array_index_1077124_comb ^ p1_array_index_1077125_comb ^ p1_res7__48_comb ^ literal_1076358[p1_array_index_1077007_comb] ^ p1_array_index_1077008_comb ^ p1_array_index_1077073_comb ^ p1_array_index_1077044_comb ^ literal_1076351[p1_array_index_1077011_comb] ^ literal_1076349[p1_array_index_1077012_comb] ^ literal_1076347[p1_array_index_1077029_comb] ^ literal_1076345[p1_array_index_1077014_comb] ^ p1_array_index_1077031_comb;
  assign p1_res7__541_comb = literal_1076345[p1_res7__540_comb] ^ literal_1076347[p1_res7__539_comb] ^ literal_1076349[p1_res7__538_comb] ^ literal_1076351[p1_res7__537_comb] ^ literal_1076353[p1_res7__536_comb] ^ literal_1076355[p1_res7__535_comb] ^ p1_res7__534_comb ^ literal_1076358[p1_res7__533_comb] ^ p1_res7__532_comb ^ p1_array_index_1077534_comb ^ p1_array_index_1077510_comb ^ p1_array_index_1077484_comb ^ p1_array_index_1077456_comb ^ p1_array_index_1077427_comb ^ literal_1076345[p1_array_index_1077394_comb] ^ p1_array_index_1077395_comb;
  assign p1_array_index_1077136_comb = literal_1076353[p1_res7__51_comb];
  assign p1_array_index_1077137_comb = literal_1076355[p1_res7__50_comb];
  assign p1_res7__56_comb = literal_1076345[p1_res7__55_comb] ^ literal_1076347[p1_res7__54_comb] ^ literal_1076349[p1_res7__53_comb] ^ literal_1076351[p1_res7__52_comb] ^ p1_array_index_1077136_comb ^ p1_array_index_1077137_comb ^ p1_res7__49_comb ^ literal_1076358[p1_res7__48_comb] ^ p1_array_index_1077007_comb ^ p1_array_index_1077087_comb ^ p1_array_index_1077058_comb ^ p1_array_index_1077026_comb ^ literal_1076349[p1_array_index_1077011_comb] ^ literal_1076347[p1_array_index_1077012_comb] ^ literal_1076345[p1_array_index_1077029_comb] ^ p1_array_index_1077014_comb;
  assign p1_res7__542_comb = literal_1076345[p1_res7__541_comb] ^ literal_1076347[p1_res7__540_comb] ^ literal_1076349[p1_res7__539_comb] ^ literal_1076351[p1_res7__538_comb] ^ literal_1076353[p1_res7__537_comb] ^ literal_1076355[p1_res7__536_comb] ^ p1_res7__535_comb ^ literal_1076358[p1_res7__534_comb] ^ p1_res7__533_comb ^ p1_array_index_1077545_comb ^ p1_array_index_1077522_comb ^ p1_array_index_1077497_comb ^ p1_array_index_1077470_comb ^ p1_array_index_1077441_comb ^ p1_array_index_1077409_comb ^ p1_array_index_1077394_comb;
  assign p1_array_index_1077147_comb = literal_1076353[p1_res7__52_comb];
  assign p1_array_index_1077148_comb = literal_1076355[p1_res7__51_comb];
  assign p1_res7__57_comb = literal_1076345[p1_res7__56_comb] ^ literal_1076347[p1_res7__55_comb] ^ literal_1076349[p1_res7__54_comb] ^ literal_1076351[p1_res7__53_comb] ^ p1_array_index_1077147_comb ^ p1_array_index_1077148_comb ^ p1_res7__50_comb ^ literal_1076358[p1_res7__49_comb] ^ p1_res7__48_comb ^ p1_array_index_1077100_comb ^ p1_array_index_1077072_comb ^ p1_array_index_1077043_comb ^ literal_1076349[p1_array_index_1077010_comb] ^ literal_1076347[p1_array_index_1077011_comb] ^ literal_1076345[p1_array_index_1077012_comb] ^ p1_array_index_1077029_comb;
  assign p1_res7__543_comb = literal_1076345[p1_res7__542_comb] ^ literal_1076347[p1_res7__541_comb] ^ literal_1076349[p1_res7__540_comb] ^ literal_1076351[p1_res7__539_comb] ^ literal_1076353[p1_res7__538_comb] ^ literal_1076355[p1_res7__537_comb] ^ p1_res7__536_comb ^ literal_1076358[p1_res7__535_comb] ^ p1_res7__534_comb ^ p1_array_index_1077555_comb ^ p1_array_index_1077533_comb ^ p1_array_index_1077509_comb ^ p1_array_index_1077483_comb ^ p1_array_index_1077455_comb ^ p1_array_index_1077426_comb ^ p1_array_index_1077393_comb;
  assign p1_array_index_1077154_comb = literal_1076345[p1_res7__57_comb];
  assign p1_array_index_1077155_comb = literal_1076347[p1_res7__56_comb];
  assign p1_array_index_1077156_comb = literal_1076349[p1_res7__55_comb];
  assign p1_array_index_1077157_comb = literal_1076351[p1_res7__54_comb];
  assign p1_array_index_1077158_comb = literal_1076353[p1_res7__53_comb];
  assign p1_array_index_1077159_comb = literal_1076355[p1_res7__52_comb];
  assign p1_array_index_1077160_comb = literal_1076358[p1_res7__50_comb];
  assign p1_array_index_1077161_comb = literal_1076347[p1_array_index_1077010_comb];
  assign p1_array_index_1077162_comb = literal_1076345[p1_array_index_1077011_comb];
  assign p1_res__33_comb = {p1_res7__543_comb, p1_res7__542_comb, p1_res7__541_comb, p1_res7__540_comb, p1_res7__539_comb, p1_res7__538_comb, p1_res7__537_comb, p1_res7__536_comb, p1_res7__535_comb, p1_res7__534_comb, p1_res7__533_comb, p1_res7__532_comb, p1_res7__531_comb, p1_res7__530_comb, p1_res7__529_comb, p1_res7__528_comb};

  // Registers for pipe stage 1:
  reg [127:0] p1_xor_1076773;
  reg [127:0] p1_xor_1076991;
  reg [7:0] p1_array_index_1077007;
  reg [7:0] p1_array_index_1077008;
  reg [7:0] p1_array_index_1077009;
  reg [7:0] p1_array_index_1077010;
  reg [7:0] p1_array_index_1077011;
  reg [7:0] p1_array_index_1077012;
  reg [7:0] p1_array_index_1077023;
  reg [7:0] p1_array_index_1077024;
  reg [7:0] p1_array_index_1077025;
  reg [7:0] p1_res7__48;
  reg [7:0] p1_array_index_1077040;
  reg [7:0] p1_array_index_1077041;
  reg [7:0] p1_array_index_1077042;
  reg [7:0] p1_res7__49;
  reg [7:0] p1_array_index_1077055;
  reg [7:0] p1_array_index_1077056;
  reg [7:0] p1_array_index_1077057;
  reg [7:0] p1_res7__50;
  reg [7:0] p1_array_index_1077069;
  reg [7:0] p1_array_index_1077070;
  reg [7:0] p1_array_index_1077071;
  reg [7:0] p1_res7__51;
  reg [7:0] p1_array_index_1077084;
  reg [7:0] p1_array_index_1077085;
  reg [7:0] p1_array_index_1077086;
  reg [7:0] p1_res7__52;
  reg [7:0] p1_array_index_1077097;
  reg [7:0] p1_array_index_1077098;
  reg [7:0] p1_array_index_1077099;
  reg [7:0] p1_res7__53;
  reg [7:0] p1_array_index_1077111;
  reg [7:0] p1_array_index_1077112;
  reg [7:0] p1_array_index_1077113;
  reg [7:0] p1_res7__54;
  reg [7:0] p1_array_index_1077123;
  reg [7:0] p1_array_index_1077124;
  reg [7:0] p1_array_index_1077125;
  reg [7:0] p1_res7__55;
  reg [7:0] p1_array_index_1077136;
  reg [7:0] p1_array_index_1077137;
  reg [7:0] p1_res7__56;
  reg [7:0] p1_array_index_1077147;
  reg [7:0] p1_array_index_1077148;
  reg [7:0] p1_res7__57;
  reg [7:0] p1_array_index_1077154;
  reg [7:0] p1_array_index_1077155;
  reg [7:0] p1_array_index_1077156;
  reg [7:0] p1_array_index_1077157;
  reg [7:0] p1_array_index_1077158;
  reg [7:0] p1_array_index_1077159;
  reg [7:0] p1_array_index_1077160;
  reg [7:0] p1_array_index_1077161;
  reg [7:0] p1_array_index_1077162;
  reg [127:0] p1_res__33;
  reg [7:0] p2_arr[256];
  reg [7:0] p2_literal_1076345[256];
  reg [7:0] p2_literal_1076347[256];
  reg [7:0] p2_literal_1076349[256];
  reg [7:0] p2_literal_1076351[256];
  reg [7:0] p2_literal_1076353[256];
  reg [7:0] p2_literal_1076355[256];
  reg [7:0] p2_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p1_xor_1076773 <= p1_xor_1076773_comb;
    p1_xor_1076991 <= p1_xor_1076991_comb;
    p1_array_index_1077007 <= p1_array_index_1077007_comb;
    p1_array_index_1077008 <= p1_array_index_1077008_comb;
    p1_array_index_1077009 <= p1_array_index_1077009_comb;
    p1_array_index_1077010 <= p1_array_index_1077010_comb;
    p1_array_index_1077011 <= p1_array_index_1077011_comb;
    p1_array_index_1077012 <= p1_array_index_1077012_comb;
    p1_array_index_1077023 <= p1_array_index_1077023_comb;
    p1_array_index_1077024 <= p1_array_index_1077024_comb;
    p1_array_index_1077025 <= p1_array_index_1077025_comb;
    p1_res7__48 <= p1_res7__48_comb;
    p1_array_index_1077040 <= p1_array_index_1077040_comb;
    p1_array_index_1077041 <= p1_array_index_1077041_comb;
    p1_array_index_1077042 <= p1_array_index_1077042_comb;
    p1_res7__49 <= p1_res7__49_comb;
    p1_array_index_1077055 <= p1_array_index_1077055_comb;
    p1_array_index_1077056 <= p1_array_index_1077056_comb;
    p1_array_index_1077057 <= p1_array_index_1077057_comb;
    p1_res7__50 <= p1_res7__50_comb;
    p1_array_index_1077069 <= p1_array_index_1077069_comb;
    p1_array_index_1077070 <= p1_array_index_1077070_comb;
    p1_array_index_1077071 <= p1_array_index_1077071_comb;
    p1_res7__51 <= p1_res7__51_comb;
    p1_array_index_1077084 <= p1_array_index_1077084_comb;
    p1_array_index_1077085 <= p1_array_index_1077085_comb;
    p1_array_index_1077086 <= p1_array_index_1077086_comb;
    p1_res7__52 <= p1_res7__52_comb;
    p1_array_index_1077097 <= p1_array_index_1077097_comb;
    p1_array_index_1077098 <= p1_array_index_1077098_comb;
    p1_array_index_1077099 <= p1_array_index_1077099_comb;
    p1_res7__53 <= p1_res7__53_comb;
    p1_array_index_1077111 <= p1_array_index_1077111_comb;
    p1_array_index_1077112 <= p1_array_index_1077112_comb;
    p1_array_index_1077113 <= p1_array_index_1077113_comb;
    p1_res7__54 <= p1_res7__54_comb;
    p1_array_index_1077123 <= p1_array_index_1077123_comb;
    p1_array_index_1077124 <= p1_array_index_1077124_comb;
    p1_array_index_1077125 <= p1_array_index_1077125_comb;
    p1_res7__55 <= p1_res7__55_comb;
    p1_array_index_1077136 <= p1_array_index_1077136_comb;
    p1_array_index_1077137 <= p1_array_index_1077137_comb;
    p1_res7__56 <= p1_res7__56_comb;
    p1_array_index_1077147 <= p1_array_index_1077147_comb;
    p1_array_index_1077148 <= p1_array_index_1077148_comb;
    p1_res7__57 <= p1_res7__57_comb;
    p1_array_index_1077154 <= p1_array_index_1077154_comb;
    p1_array_index_1077155 <= p1_array_index_1077155_comb;
    p1_array_index_1077156 <= p1_array_index_1077156_comb;
    p1_array_index_1077157 <= p1_array_index_1077157_comb;
    p1_array_index_1077158 <= p1_array_index_1077158_comb;
    p1_array_index_1077159 <= p1_array_index_1077159_comb;
    p1_array_index_1077160 <= p1_array_index_1077160_comb;
    p1_array_index_1077161 <= p1_array_index_1077161_comb;
    p1_array_index_1077162 <= p1_array_index_1077162_comb;
    p1_res__33 <= p1_res__33_comb;
    p2_arr <= p1_arr;
    p2_literal_1076345 <= p1_literal_1076345;
    p2_literal_1076347 <= p1_literal_1076347;
    p2_literal_1076349 <= p1_literal_1076349;
    p2_literal_1076351 <= p1_literal_1076351;
    p2_literal_1076353 <= p1_literal_1076353;
    p2_literal_1076355 <= p1_literal_1076355;
    p2_literal_1076358 <= p1_literal_1076358;
  end

  // ===== Pipe stage 2:
  wire [7:0] p2_res7__58_comb;
  wire [7:0] p2_array_index_1077729_comb;
  wire [7:0] p2_res7__59_comb;
  wire [7:0] p2_res7__60_comb;
  wire [7:0] p2_res7__61_comb;
  wire [7:0] p2_res7__62_comb;
  wire [7:0] p2_res7__63_comb;
  wire [127:0] p2_res__3_comb;
  wire [127:0] p2_xor_1077769_comb;
  wire [127:0] p2_addedKey__45_comb;
  wire [7:0] p2_array_index_1077785_comb;
  wire [7:0] p2_array_index_1077786_comb;
  wire [7:0] p2_array_index_1077787_comb;
  wire [7:0] p2_array_index_1077788_comb;
  wire [7:0] p2_array_index_1077789_comb;
  wire [7:0] p2_array_index_1077790_comb;
  wire [7:0] p2_array_index_1077792_comb;
  wire [7:0] p2_array_index_1077794_comb;
  wire [7:0] p2_array_index_1077795_comb;
  wire [7:0] p2_array_index_1077796_comb;
  wire [7:0] p2_array_index_1077797_comb;
  wire [7:0] p2_array_index_1077798_comb;
  wire [7:0] p2_array_index_1077799_comb;
  wire [7:0] p2_array_index_1077801_comb;
  wire [7:0] p2_array_index_1077802_comb;
  wire [7:0] p2_array_index_1077803_comb;
  wire [7:0] p2_array_index_1077804_comb;
  wire [7:0] p2_array_index_1077805_comb;
  wire [7:0] p2_array_index_1077806_comb;
  wire [7:0] p2_array_index_1077807_comb;
  wire [7:0] p2_array_index_1077809_comb;
  wire [7:0] p2_res7__64_comb;
  wire [7:0] p2_array_index_1077818_comb;
  wire [7:0] p2_array_index_1077819_comb;
  wire [7:0] p2_array_index_1077820_comb;
  wire [7:0] p2_array_index_1077821_comb;
  wire [7:0] p2_array_index_1077822_comb;
  wire [7:0] p2_array_index_1077823_comb;
  wire [7:0] p2_res7__65_comb;
  wire [7:0] p2_array_index_1077833_comb;
  wire [7:0] p2_array_index_1077834_comb;
  wire [7:0] p2_array_index_1077835_comb;
  wire [7:0] p2_array_index_1077836_comb;
  wire [7:0] p2_array_index_1077837_comb;
  wire [7:0] p2_res7__66_comb;
  wire [7:0] p2_array_index_1077847_comb;
  wire [7:0] p2_array_index_1077848_comb;
  wire [7:0] p2_array_index_1077849_comb;
  wire [7:0] p2_array_index_1077850_comb;
  wire [7:0] p2_array_index_1077851_comb;
  wire [7:0] p2_res7__67_comb;
  wire [7:0] p2_array_index_1077862_comb;
  wire [7:0] p2_array_index_1077863_comb;
  wire [7:0] p2_array_index_1077864_comb;
  wire [7:0] p2_array_index_1077865_comb;
  wire [7:0] p2_res7__68_comb;
  wire [7:0] p2_array_index_1077875_comb;
  wire [7:0] p2_array_index_1077876_comb;
  wire [7:0] p2_array_index_1077877_comb;
  wire [7:0] p2_array_index_1077878_comb;
  wire [7:0] p2_res7__69_comb;
  wire [7:0] p2_array_index_1077889_comb;
  wire [7:0] p2_array_index_1077890_comb;
  wire [7:0] p2_array_index_1077891_comb;
  wire [7:0] p2_res7__70_comb;
  wire [7:0] p2_array_index_1077901_comb;
  wire [7:0] p2_array_index_1077902_comb;
  wire [7:0] p2_array_index_1077903_comb;
  wire [7:0] p2_res7__71_comb;
  wire [7:0] p2_array_index_1077914_comb;
  wire [7:0] p2_array_index_1077915_comb;
  wire [7:0] p2_res7__72_comb;
  wire [7:0] p2_array_index_1077925_comb;
  wire [7:0] p2_array_index_1077926_comb;
  wire [7:0] p2_res7__73_comb;
  wire [7:0] p2_array_index_1077937_comb;
  wire [7:0] p2_res7__74_comb;
  wire [7:0] p2_array_index_1077947_comb;
  wire [7:0] p2_res7__75_comb;
  wire [7:0] p2_res7__76_comb;
  wire [7:0] p2_res7__77_comb;
  wire [7:0] p2_res7__78_comb;
  wire [7:0] p2_res7__79_comb;
  wire [127:0] p2_res__4_comb;
  wire [127:0] p2_xor_1077987_comb;
  wire [127:0] p2_addedKey__46_comb;
  wire [7:0] p2_array_index_1078003_comb;
  wire [7:0] p2_array_index_1078004_comb;
  wire [7:0] p2_array_index_1078005_comb;
  wire [7:0] p2_array_index_1078006_comb;
  wire [7:0] p2_array_index_1078007_comb;
  wire [7:0] p2_array_index_1078008_comb;
  wire [7:0] p2_array_index_1078010_comb;
  wire [7:0] p2_array_index_1078012_comb;
  wire [7:0] p2_array_index_1078013_comb;
  wire [7:0] p2_array_index_1078014_comb;
  wire [7:0] p2_array_index_1078015_comb;
  wire [7:0] p2_array_index_1078016_comb;
  wire [7:0] p2_array_index_1078017_comb;
  wire [7:0] p2_array_index_1078019_comb;
  wire [7:0] p2_array_index_1078020_comb;
  wire [7:0] p2_array_index_1078021_comb;
  wire [7:0] p2_array_index_1078022_comb;
  wire [7:0] p2_array_index_1078023_comb;
  wire [7:0] p2_array_index_1078024_comb;
  wire [7:0] p2_array_index_1078025_comb;
  wire [7:0] p2_array_index_1078027_comb;
  wire [7:0] p2_res7__80_comb;
  wire [7:0] p2_array_index_1078036_comb;
  wire [7:0] p2_array_index_1078037_comb;
  wire [7:0] p2_array_index_1078038_comb;
  wire [7:0] p2_array_index_1078039_comb;
  wire [7:0] p2_array_index_1078040_comb;
  wire [7:0] p2_array_index_1078041_comb;
  wire [7:0] p2_res7__81_comb;
  wire [7:0] p2_array_index_1078051_comb;
  wire [7:0] p2_array_index_1078052_comb;
  wire [7:0] p2_array_index_1078053_comb;
  wire [7:0] p2_array_index_1078054_comb;
  wire [7:0] p2_array_index_1078055_comb;
  wire [7:0] p2_res7__82_comb;
  wire [7:0] p2_array_index_1078065_comb;
  wire [7:0] p2_array_index_1078066_comb;
  wire [7:0] p2_array_index_1078067_comb;
  wire [7:0] p2_array_index_1078068_comb;
  wire [7:0] p2_array_index_1078069_comb;
  wire [7:0] p2_res7__83_comb;
  wire [7:0] p2_array_index_1078080_comb;
  wire [7:0] p2_array_index_1078081_comb;
  wire [7:0] p2_array_index_1078082_comb;
  wire [7:0] p2_array_index_1078083_comb;
  wire [7:0] p2_res7__84_comb;
  wire [7:0] p2_array_index_1078093_comb;
  wire [7:0] p2_array_index_1078094_comb;
  wire [7:0] p2_array_index_1078095_comb;
  wire [7:0] p2_array_index_1078096_comb;
  wire [7:0] p2_res7__85_comb;
  wire [7:0] p2_array_index_1078107_comb;
  wire [7:0] p2_array_index_1078108_comb;
  wire [7:0] p2_array_index_1078109_comb;
  wire [7:0] p2_res7__86_comb;
  wire [7:0] p2_array_index_1078119_comb;
  wire [7:0] p2_array_index_1078120_comb;
  wire [7:0] p2_array_index_1078121_comb;
  wire [7:0] p2_res7__87_comb;
  wire [7:0] p2_array_index_1078132_comb;
  wire [7:0] p2_array_index_1078133_comb;
  wire [7:0] p2_res7__88_comb;
  wire [7:0] p2_array_index_1078143_comb;
  wire [7:0] p2_array_index_1078144_comb;
  wire [7:0] p2_res7__89_comb;
  wire [7:0] p2_array_index_1078155_comb;
  wire [7:0] p2_res7__90_comb;
  wire [7:0] p2_array_index_1078165_comb;
  wire [7:0] p2_res7__91_comb;
  wire [7:0] p2_res7__92_comb;
  wire [7:0] p2_res7__93_comb;
  wire [7:0] p2_res7__94_comb;
  wire [7:0] p2_res7__95_comb;
  wire [127:0] p2_res__5_comb;
  wire [127:0] p2_xor_1078205_comb;
  wire [127:0] p2_addedKey__47_comb;
  wire [7:0] p2_array_index_1078221_comb;
  wire [7:0] p2_array_index_1078222_comb;
  wire [7:0] p2_array_index_1078223_comb;
  wire [7:0] p2_array_index_1078224_comb;
  wire [7:0] p2_array_index_1078225_comb;
  wire [7:0] p2_array_index_1078226_comb;
  wire [7:0] p2_array_index_1078228_comb;
  wire [7:0] p2_array_index_1078230_comb;
  wire [7:0] p2_array_index_1078231_comb;
  wire [7:0] p2_array_index_1078232_comb;
  wire [7:0] p2_array_index_1078233_comb;
  wire [7:0] p2_array_index_1078234_comb;
  wire [7:0] p2_array_index_1078235_comb;
  wire [7:0] p2_array_index_1078237_comb;
  wire [7:0] p2_array_index_1078238_comb;
  wire [7:0] p2_array_index_1078239_comb;
  wire [7:0] p2_array_index_1078240_comb;
  wire [7:0] p2_array_index_1078241_comb;
  wire [7:0] p2_array_index_1078242_comb;
  wire [7:0] p2_array_index_1078243_comb;
  wire [7:0] p2_array_index_1078245_comb;
  wire [7:0] p2_res7__96_comb;
  wire [7:0] p2_array_index_1078254_comb;
  wire [7:0] p2_array_index_1078255_comb;
  wire [7:0] p2_array_index_1078256_comb;
  wire [7:0] p2_array_index_1078257_comb;
  wire [7:0] p2_array_index_1078258_comb;
  wire [7:0] p2_array_index_1078259_comb;
  wire [7:0] p2_res7__97_comb;
  wire [7:0] p2_array_index_1078269_comb;
  wire [7:0] p2_array_index_1078270_comb;
  wire [7:0] p2_array_index_1078271_comb;
  wire [7:0] p2_array_index_1078272_comb;
  wire [7:0] p2_array_index_1078273_comb;
  wire [7:0] p2_res7__98_comb;
  wire [7:0] p2_array_index_1078283_comb;
  wire [7:0] p2_array_index_1078284_comb;
  wire [7:0] p2_array_index_1078285_comb;
  wire [7:0] p2_array_index_1078286_comb;
  wire [7:0] p2_array_index_1078287_comb;
  wire [7:0] p2_res7__99_comb;
  wire [7:0] p2_array_index_1078298_comb;
  wire [7:0] p2_array_index_1078299_comb;
  wire [7:0] p2_array_index_1078300_comb;
  wire [7:0] p2_array_index_1078301_comb;
  wire [7:0] p2_res7__100_comb;
  wire [7:0] p2_array_index_1078311_comb;
  wire [7:0] p2_array_index_1078312_comb;
  wire [7:0] p2_array_index_1078313_comb;
  wire [7:0] p2_array_index_1078314_comb;
  wire [7:0] p2_res7__101_comb;
  wire [7:0] p2_array_index_1078325_comb;
  wire [7:0] p2_array_index_1078326_comb;
  wire [7:0] p2_array_index_1078327_comb;
  wire [7:0] p2_res7__102_comb;
  wire [7:0] p2_array_index_1078337_comb;
  wire [7:0] p2_array_index_1078338_comb;
  wire [7:0] p2_array_index_1078339_comb;
  wire [7:0] p2_res7__103_comb;
  wire [7:0] p2_array_index_1078350_comb;
  wire [7:0] p2_array_index_1078351_comb;
  wire [7:0] p2_res7__104_comb;
  wire [7:0] p2_array_index_1078361_comb;
  wire [7:0] p2_array_index_1078362_comb;
  wire [7:0] p2_res7__105_comb;
  wire [7:0] p2_array_index_1078373_comb;
  wire [7:0] p2_res7__106_comb;
  wire [7:0] p2_array_index_1078383_comb;
  wire [7:0] p2_res7__107_comb;
  wire [7:0] p2_res7__108_comb;
  wire [7:0] p2_res7__109_comb;
  wire [7:0] p2_res7__110_comb;
  wire [7:0] p2_res7__111_comb;
  wire [127:0] p2_res__6_comb;
  wire [127:0] p2_k3_comb;
  wire [127:0] p2_addedKey__48_comb;
  wire [7:0] p2_array_index_1078439_comb;
  wire [7:0] p2_array_index_1078440_comb;
  wire [7:0] p2_array_index_1078441_comb;
  wire [7:0] p2_array_index_1078442_comb;
  wire [7:0] p2_array_index_1078443_comb;
  wire [7:0] p2_array_index_1078444_comb;
  wire [7:0] p2_array_index_1078446_comb;
  wire [7:0] p2_array_index_1078448_comb;
  wire [7:0] p2_array_index_1078449_comb;
  wire [7:0] p2_array_index_1078450_comb;
  wire [7:0] p2_array_index_1078451_comb;
  wire [7:0] p2_array_index_1078452_comb;
  wire [7:0] p2_array_index_1078453_comb;
  wire [7:0] p2_array_index_1078455_comb;
  wire [7:0] p2_array_index_1078456_comb;
  wire [7:0] p2_array_index_1078457_comb;
  wire [7:0] p2_array_index_1078458_comb;
  wire [7:0] p2_array_index_1078459_comb;
  wire [7:0] p2_array_index_1078460_comb;
  wire [7:0] p2_array_index_1078461_comb;
  wire [7:0] p2_array_index_1078463_comb;
  wire [7:0] p2_res7__112_comb;
  wire [7:0] p2_array_index_1078472_comb;
  wire [7:0] p2_array_index_1078473_comb;
  wire [7:0] p2_array_index_1078474_comb;
  wire [7:0] p2_array_index_1078475_comb;
  wire [7:0] p2_array_index_1078476_comb;
  wire [7:0] p2_array_index_1078477_comb;
  wire [7:0] p2_res7__113_comb;
  wire [7:0] p2_array_index_1078487_comb;
  wire [7:0] p2_array_index_1078488_comb;
  wire [7:0] p2_array_index_1078489_comb;
  wire [7:0] p2_array_index_1078490_comb;
  wire [7:0] p2_array_index_1078491_comb;
  wire [7:0] p2_res7__114_comb;
  wire [7:0] p2_array_index_1078501_comb;
  wire [7:0] p2_array_index_1078502_comb;
  wire [7:0] p2_array_index_1078503_comb;
  wire [7:0] p2_array_index_1078504_comb;
  wire [7:0] p2_array_index_1078505_comb;
  wire [7:0] p2_res7__115_comb;
  wire [7:0] p2_array_index_1078516_comb;
  wire [7:0] p2_array_index_1078517_comb;
  wire [7:0] p2_array_index_1078518_comb;
  wire [7:0] p2_array_index_1078519_comb;
  wire [7:0] p2_res7__116_comb;
  assign p2_res7__58_comb = p1_array_index_1077154 ^ p1_array_index_1077155 ^ p1_array_index_1077156 ^ p1_array_index_1077157 ^ p1_array_index_1077158 ^ p1_array_index_1077159 ^ p1_res7__51 ^ p1_array_index_1077160 ^ p1_res7__49 ^ p1_array_index_1077113 ^ p1_array_index_1077086 ^ p1_array_index_1077057 ^ p1_array_index_1077025 ^ p1_array_index_1077161 ^ p1_array_index_1077162 ^ p1_array_index_1077012;
  assign p2_array_index_1077729_comb = p1_literal_1076355[p1_res7__53];
  assign p2_res7__59_comb = p1_literal_1076345[p2_res7__58_comb] ^ p1_literal_1076347[p1_res7__57] ^ p1_literal_1076349[p1_res7__56] ^ p1_literal_1076351[p1_res7__55] ^ p1_literal_1076353[p1_res7__54] ^ p2_array_index_1077729_comb ^ p1_res7__52 ^ p1_literal_1076358[p1_res7__51] ^ p1_res7__50 ^ p1_array_index_1077125 ^ p1_array_index_1077099 ^ p1_array_index_1077071 ^ p1_array_index_1077042 ^ p1_literal_1076347[p1_array_index_1077009] ^ p1_literal_1076345[p1_array_index_1077010] ^ p1_array_index_1077011;
  assign p2_res7__60_comb = p1_literal_1076345[p2_res7__59_comb] ^ p1_literal_1076347[p2_res7__58_comb] ^ p1_literal_1076349[p1_res7__57] ^ p1_literal_1076351[p1_res7__56] ^ p1_literal_1076353[p1_res7__55] ^ p1_literal_1076355[p1_res7__54] ^ p1_res7__53 ^ p1_literal_1076358[p1_res7__52] ^ p1_res7__51 ^ p1_array_index_1077137 ^ p1_array_index_1077112 ^ p1_array_index_1077085 ^ p1_array_index_1077056 ^ p1_array_index_1077024 ^ p1_literal_1076345[p1_array_index_1077009] ^ p1_array_index_1077010;
  assign p2_res7__61_comb = p1_literal_1076345[p2_res7__60_comb] ^ p1_literal_1076347[p2_res7__59_comb] ^ p1_literal_1076349[p2_res7__58_comb] ^ p1_literal_1076351[p1_res7__57] ^ p1_literal_1076353[p1_res7__56] ^ p1_literal_1076355[p1_res7__55] ^ p1_res7__54 ^ p1_literal_1076358[p1_res7__53] ^ p1_res7__52 ^ p1_array_index_1077148 ^ p1_array_index_1077124 ^ p1_array_index_1077098 ^ p1_array_index_1077070 ^ p1_array_index_1077041 ^ p1_literal_1076345[p1_array_index_1077008] ^ p1_array_index_1077009;
  assign p2_res7__62_comb = p1_literal_1076345[p2_res7__61_comb] ^ p1_literal_1076347[p2_res7__60_comb] ^ p1_literal_1076349[p2_res7__59_comb] ^ p1_literal_1076351[p2_res7__58_comb] ^ p1_literal_1076353[p1_res7__57] ^ p1_literal_1076355[p1_res7__56] ^ p1_res7__55 ^ p1_literal_1076358[p1_res7__54] ^ p1_res7__53 ^ p1_array_index_1077159 ^ p1_array_index_1077136 ^ p1_array_index_1077111 ^ p1_array_index_1077084 ^ p1_array_index_1077055 ^ p1_array_index_1077023 ^ p1_array_index_1077008;
  assign p2_res7__63_comb = p1_literal_1076345[p2_res7__62_comb] ^ p1_literal_1076347[p2_res7__61_comb] ^ p1_literal_1076349[p2_res7__60_comb] ^ p1_literal_1076351[p2_res7__59_comb] ^ p1_literal_1076353[p2_res7__58_comb] ^ p1_literal_1076355[p1_res7__57] ^ p1_res7__56 ^ p1_literal_1076358[p1_res7__55] ^ p1_res7__54 ^ p2_array_index_1077729_comb ^ p1_array_index_1077147 ^ p1_array_index_1077123 ^ p1_array_index_1077097 ^ p1_array_index_1077069 ^ p1_array_index_1077040 ^ p1_array_index_1077007;
  assign p2_res__3_comb = {p2_res7__63_comb, p2_res7__62_comb, p2_res7__61_comb, p2_res7__60_comb, p2_res7__59_comb, p2_res7__58_comb, p1_res7__57, p1_res7__56, p1_res7__55, p1_res7__54, p1_res7__53, p1_res7__52, p1_res7__51, p1_res7__50, p1_res7__49, p1_res7__48};
  assign p2_xor_1077769_comb = p2_res__3_comb ^ p1_xor_1076773;
  assign p2_addedKey__45_comb = p2_xor_1077769_comb ^ 128'h156f_6d79_1fab_511d_eabb_0c50_2fd1_8105;
  assign p2_array_index_1077785_comb = p1_arr[p2_addedKey__45_comb[127:120]];
  assign p2_array_index_1077786_comb = p1_arr[p2_addedKey__45_comb[119:112]];
  assign p2_array_index_1077787_comb = p1_arr[p2_addedKey__45_comb[111:104]];
  assign p2_array_index_1077788_comb = p1_arr[p2_addedKey__45_comb[103:96]];
  assign p2_array_index_1077789_comb = p1_arr[p2_addedKey__45_comb[95:88]];
  assign p2_array_index_1077790_comb = p1_arr[p2_addedKey__45_comb[87:80]];
  assign p2_array_index_1077792_comb = p1_arr[p2_addedKey__45_comb[71:64]];
  assign p2_array_index_1077794_comb = p1_arr[p2_addedKey__45_comb[55:48]];
  assign p2_array_index_1077795_comb = p1_arr[p2_addedKey__45_comb[47:40]];
  assign p2_array_index_1077796_comb = p1_arr[p2_addedKey__45_comb[39:32]];
  assign p2_array_index_1077797_comb = p1_arr[p2_addedKey__45_comb[31:24]];
  assign p2_array_index_1077798_comb = p1_arr[p2_addedKey__45_comb[23:16]];
  assign p2_array_index_1077799_comb = p1_arr[p2_addedKey__45_comb[15:8]];
  assign p2_array_index_1077801_comb = p1_literal_1076345[p2_array_index_1077785_comb];
  assign p2_array_index_1077802_comb = p1_literal_1076347[p2_array_index_1077786_comb];
  assign p2_array_index_1077803_comb = p1_literal_1076349[p2_array_index_1077787_comb];
  assign p2_array_index_1077804_comb = p1_literal_1076351[p2_array_index_1077788_comb];
  assign p2_array_index_1077805_comb = p1_literal_1076353[p2_array_index_1077789_comb];
  assign p2_array_index_1077806_comb = p1_literal_1076355[p2_array_index_1077790_comb];
  assign p2_array_index_1077807_comb = p1_arr[p2_addedKey__45_comb[79:72]];
  assign p2_array_index_1077809_comb = p1_arr[p2_addedKey__45_comb[63:56]];
  assign p2_res7__64_comb = p2_array_index_1077801_comb ^ p2_array_index_1077802_comb ^ p2_array_index_1077803_comb ^ p2_array_index_1077804_comb ^ p2_array_index_1077805_comb ^ p2_array_index_1077806_comb ^ p2_array_index_1077807_comb ^ p1_literal_1076358[p2_array_index_1077792_comb] ^ p2_array_index_1077809_comb ^ p1_literal_1076355[p2_array_index_1077794_comb] ^ p1_literal_1076353[p2_array_index_1077795_comb] ^ p1_literal_1076351[p2_array_index_1077796_comb] ^ p1_literal_1076349[p2_array_index_1077797_comb] ^ p1_literal_1076347[p2_array_index_1077798_comb] ^ p1_literal_1076345[p2_array_index_1077799_comb] ^ p1_arr[p2_addedKey__45_comb[7:0]];
  assign p2_array_index_1077818_comb = p1_literal_1076345[p2_res7__64_comb];
  assign p2_array_index_1077819_comb = p1_literal_1076347[p2_array_index_1077785_comb];
  assign p2_array_index_1077820_comb = p1_literal_1076349[p2_array_index_1077786_comb];
  assign p2_array_index_1077821_comb = p1_literal_1076351[p2_array_index_1077787_comb];
  assign p2_array_index_1077822_comb = p1_literal_1076353[p2_array_index_1077788_comb];
  assign p2_array_index_1077823_comb = p1_literal_1076355[p2_array_index_1077789_comb];
  assign p2_res7__65_comb = p2_array_index_1077818_comb ^ p2_array_index_1077819_comb ^ p2_array_index_1077820_comb ^ p2_array_index_1077821_comb ^ p2_array_index_1077822_comb ^ p2_array_index_1077823_comb ^ p2_array_index_1077790_comb ^ p1_literal_1076358[p2_array_index_1077807_comb] ^ p2_array_index_1077792_comb ^ p1_literal_1076355[p2_array_index_1077809_comb] ^ p1_literal_1076353[p2_array_index_1077794_comb] ^ p1_literal_1076351[p2_array_index_1077795_comb] ^ p1_literal_1076349[p2_array_index_1077796_comb] ^ p1_literal_1076347[p2_array_index_1077797_comb] ^ p1_literal_1076345[p2_array_index_1077798_comb] ^ p2_array_index_1077799_comb;
  assign p2_array_index_1077833_comb = p1_literal_1076347[p2_res7__64_comb];
  assign p2_array_index_1077834_comb = p1_literal_1076349[p2_array_index_1077785_comb];
  assign p2_array_index_1077835_comb = p1_literal_1076351[p2_array_index_1077786_comb];
  assign p2_array_index_1077836_comb = p1_literal_1076353[p2_array_index_1077787_comb];
  assign p2_array_index_1077837_comb = p1_literal_1076355[p2_array_index_1077788_comb];
  assign p2_res7__66_comb = p1_literal_1076345[p2_res7__65_comb] ^ p2_array_index_1077833_comb ^ p2_array_index_1077834_comb ^ p2_array_index_1077835_comb ^ p2_array_index_1077836_comb ^ p2_array_index_1077837_comb ^ p2_array_index_1077789_comb ^ p1_literal_1076358[p2_array_index_1077790_comb] ^ p2_array_index_1077807_comb ^ p1_literal_1076355[p2_array_index_1077792_comb] ^ p1_literal_1076353[p2_array_index_1077809_comb] ^ p1_literal_1076351[p2_array_index_1077794_comb] ^ p1_literal_1076349[p2_array_index_1077795_comb] ^ p1_literal_1076347[p2_array_index_1077796_comb] ^ p1_literal_1076345[p2_array_index_1077797_comb] ^ p2_array_index_1077798_comb;
  assign p2_array_index_1077847_comb = p1_literal_1076347[p2_res7__65_comb];
  assign p2_array_index_1077848_comb = p1_literal_1076349[p2_res7__64_comb];
  assign p2_array_index_1077849_comb = p1_literal_1076351[p2_array_index_1077785_comb];
  assign p2_array_index_1077850_comb = p1_literal_1076353[p2_array_index_1077786_comb];
  assign p2_array_index_1077851_comb = p1_literal_1076355[p2_array_index_1077787_comb];
  assign p2_res7__67_comb = p1_literal_1076345[p2_res7__66_comb] ^ p2_array_index_1077847_comb ^ p2_array_index_1077848_comb ^ p2_array_index_1077849_comb ^ p2_array_index_1077850_comb ^ p2_array_index_1077851_comb ^ p2_array_index_1077788_comb ^ p1_literal_1076358[p2_array_index_1077789_comb] ^ p2_array_index_1077790_comb ^ p1_literal_1076355[p2_array_index_1077807_comb] ^ p1_literal_1076353[p2_array_index_1077792_comb] ^ p1_literal_1076351[p2_array_index_1077809_comb] ^ p1_literal_1076349[p2_array_index_1077794_comb] ^ p1_literal_1076347[p2_array_index_1077795_comb] ^ p1_literal_1076345[p2_array_index_1077796_comb] ^ p2_array_index_1077797_comb;
  assign p2_array_index_1077862_comb = p1_literal_1076349[p2_res7__65_comb];
  assign p2_array_index_1077863_comb = p1_literal_1076351[p2_res7__64_comb];
  assign p2_array_index_1077864_comb = p1_literal_1076353[p2_array_index_1077785_comb];
  assign p2_array_index_1077865_comb = p1_literal_1076355[p2_array_index_1077786_comb];
  assign p2_res7__68_comb = p1_literal_1076345[p2_res7__67_comb] ^ p1_literal_1076347[p2_res7__66_comb] ^ p2_array_index_1077862_comb ^ p2_array_index_1077863_comb ^ p2_array_index_1077864_comb ^ p2_array_index_1077865_comb ^ p2_array_index_1077787_comb ^ p1_literal_1076358[p2_array_index_1077788_comb] ^ p2_array_index_1077789_comb ^ p2_array_index_1077806_comb ^ p1_literal_1076353[p2_array_index_1077807_comb] ^ p1_literal_1076351[p2_array_index_1077792_comb] ^ p1_literal_1076349[p2_array_index_1077809_comb] ^ p1_literal_1076347[p2_array_index_1077794_comb] ^ p1_literal_1076345[p2_array_index_1077795_comb] ^ p2_array_index_1077796_comb;
  assign p2_array_index_1077875_comb = p1_literal_1076349[p2_res7__66_comb];
  assign p2_array_index_1077876_comb = p1_literal_1076351[p2_res7__65_comb];
  assign p2_array_index_1077877_comb = p1_literal_1076353[p2_res7__64_comb];
  assign p2_array_index_1077878_comb = p1_literal_1076355[p2_array_index_1077785_comb];
  assign p2_res7__69_comb = p1_literal_1076345[p2_res7__68_comb] ^ p1_literal_1076347[p2_res7__67_comb] ^ p2_array_index_1077875_comb ^ p2_array_index_1077876_comb ^ p2_array_index_1077877_comb ^ p2_array_index_1077878_comb ^ p2_array_index_1077786_comb ^ p1_literal_1076358[p2_array_index_1077787_comb] ^ p2_array_index_1077788_comb ^ p2_array_index_1077823_comb ^ p1_literal_1076353[p2_array_index_1077790_comb] ^ p1_literal_1076351[p2_array_index_1077807_comb] ^ p1_literal_1076349[p2_array_index_1077792_comb] ^ p1_literal_1076347[p2_array_index_1077809_comb] ^ p1_literal_1076345[p2_array_index_1077794_comb] ^ p2_array_index_1077795_comb;
  assign p2_array_index_1077889_comb = p1_literal_1076351[p2_res7__66_comb];
  assign p2_array_index_1077890_comb = p1_literal_1076353[p2_res7__65_comb];
  assign p2_array_index_1077891_comb = p1_literal_1076355[p2_res7__64_comb];
  assign p2_res7__70_comb = p1_literal_1076345[p2_res7__69_comb] ^ p1_literal_1076347[p2_res7__68_comb] ^ p1_literal_1076349[p2_res7__67_comb] ^ p2_array_index_1077889_comb ^ p2_array_index_1077890_comb ^ p2_array_index_1077891_comb ^ p2_array_index_1077785_comb ^ p1_literal_1076358[p2_array_index_1077786_comb] ^ p2_array_index_1077787_comb ^ p2_array_index_1077837_comb ^ p2_array_index_1077805_comb ^ p1_literal_1076351[p2_array_index_1077790_comb] ^ p1_literal_1076349[p2_array_index_1077807_comb] ^ p1_literal_1076347[p2_array_index_1077792_comb] ^ p1_literal_1076345[p2_array_index_1077809_comb] ^ p2_array_index_1077794_comb;
  assign p2_array_index_1077901_comb = p1_literal_1076351[p2_res7__67_comb];
  assign p2_array_index_1077902_comb = p1_literal_1076353[p2_res7__66_comb];
  assign p2_array_index_1077903_comb = p1_literal_1076355[p2_res7__65_comb];
  assign p2_res7__71_comb = p1_literal_1076345[p2_res7__70_comb] ^ p1_literal_1076347[p2_res7__69_comb] ^ p1_literal_1076349[p2_res7__68_comb] ^ p2_array_index_1077901_comb ^ p2_array_index_1077902_comb ^ p2_array_index_1077903_comb ^ p2_res7__64_comb ^ p1_literal_1076358[p2_array_index_1077785_comb] ^ p2_array_index_1077786_comb ^ p2_array_index_1077851_comb ^ p2_array_index_1077822_comb ^ p1_literal_1076351[p2_array_index_1077789_comb] ^ p1_literal_1076349[p2_array_index_1077790_comb] ^ p1_literal_1076347[p2_array_index_1077807_comb] ^ p1_literal_1076345[p2_array_index_1077792_comb] ^ p2_array_index_1077809_comb;
  assign p2_array_index_1077914_comb = p1_literal_1076353[p2_res7__67_comb];
  assign p2_array_index_1077915_comb = p1_literal_1076355[p2_res7__66_comb];
  assign p2_res7__72_comb = p1_literal_1076345[p2_res7__71_comb] ^ p1_literal_1076347[p2_res7__70_comb] ^ p1_literal_1076349[p2_res7__69_comb] ^ p1_literal_1076351[p2_res7__68_comb] ^ p2_array_index_1077914_comb ^ p2_array_index_1077915_comb ^ p2_res7__65_comb ^ p1_literal_1076358[p2_res7__64_comb] ^ p2_array_index_1077785_comb ^ p2_array_index_1077865_comb ^ p2_array_index_1077836_comb ^ p2_array_index_1077804_comb ^ p1_literal_1076349[p2_array_index_1077789_comb] ^ p1_literal_1076347[p2_array_index_1077790_comb] ^ p1_literal_1076345[p2_array_index_1077807_comb] ^ p2_array_index_1077792_comb;
  assign p2_array_index_1077925_comb = p1_literal_1076353[p2_res7__68_comb];
  assign p2_array_index_1077926_comb = p1_literal_1076355[p2_res7__67_comb];
  assign p2_res7__73_comb = p1_literal_1076345[p2_res7__72_comb] ^ p1_literal_1076347[p2_res7__71_comb] ^ p1_literal_1076349[p2_res7__70_comb] ^ p1_literal_1076351[p2_res7__69_comb] ^ p2_array_index_1077925_comb ^ p2_array_index_1077926_comb ^ p2_res7__66_comb ^ p1_literal_1076358[p2_res7__65_comb] ^ p2_res7__64_comb ^ p2_array_index_1077878_comb ^ p2_array_index_1077850_comb ^ p2_array_index_1077821_comb ^ p1_literal_1076349[p2_array_index_1077788_comb] ^ p1_literal_1076347[p2_array_index_1077789_comb] ^ p1_literal_1076345[p2_array_index_1077790_comb] ^ p2_array_index_1077807_comb;
  assign p2_array_index_1077937_comb = p1_literal_1076355[p2_res7__68_comb];
  assign p2_res7__74_comb = p1_literal_1076345[p2_res7__73_comb] ^ p1_literal_1076347[p2_res7__72_comb] ^ p1_literal_1076349[p2_res7__71_comb] ^ p1_literal_1076351[p2_res7__70_comb] ^ p1_literal_1076353[p2_res7__69_comb] ^ p2_array_index_1077937_comb ^ p2_res7__67_comb ^ p1_literal_1076358[p2_res7__66_comb] ^ p2_res7__65_comb ^ p2_array_index_1077891_comb ^ p2_array_index_1077864_comb ^ p2_array_index_1077835_comb ^ p2_array_index_1077803_comb ^ p1_literal_1076347[p2_array_index_1077788_comb] ^ p1_literal_1076345[p2_array_index_1077789_comb] ^ p2_array_index_1077790_comb;
  assign p2_array_index_1077947_comb = p1_literal_1076355[p2_res7__69_comb];
  assign p2_res7__75_comb = p1_literal_1076345[p2_res7__74_comb] ^ p1_literal_1076347[p2_res7__73_comb] ^ p1_literal_1076349[p2_res7__72_comb] ^ p1_literal_1076351[p2_res7__71_comb] ^ p1_literal_1076353[p2_res7__70_comb] ^ p2_array_index_1077947_comb ^ p2_res7__68_comb ^ p1_literal_1076358[p2_res7__67_comb] ^ p2_res7__66_comb ^ p2_array_index_1077903_comb ^ p2_array_index_1077877_comb ^ p2_array_index_1077849_comb ^ p2_array_index_1077820_comb ^ p1_literal_1076347[p2_array_index_1077787_comb] ^ p1_literal_1076345[p2_array_index_1077788_comb] ^ p2_array_index_1077789_comb;
  assign p2_res7__76_comb = p1_literal_1076345[p2_res7__75_comb] ^ p1_literal_1076347[p2_res7__74_comb] ^ p1_literal_1076349[p2_res7__73_comb] ^ p1_literal_1076351[p2_res7__72_comb] ^ p1_literal_1076353[p2_res7__71_comb] ^ p1_literal_1076355[p2_res7__70_comb] ^ p2_res7__69_comb ^ p1_literal_1076358[p2_res7__68_comb] ^ p2_res7__67_comb ^ p2_array_index_1077915_comb ^ p2_array_index_1077890_comb ^ p2_array_index_1077863_comb ^ p2_array_index_1077834_comb ^ p2_array_index_1077802_comb ^ p1_literal_1076345[p2_array_index_1077787_comb] ^ p2_array_index_1077788_comb;
  assign p2_res7__77_comb = p1_literal_1076345[p2_res7__76_comb] ^ p1_literal_1076347[p2_res7__75_comb] ^ p1_literal_1076349[p2_res7__74_comb] ^ p1_literal_1076351[p2_res7__73_comb] ^ p1_literal_1076353[p2_res7__72_comb] ^ p1_literal_1076355[p2_res7__71_comb] ^ p2_res7__70_comb ^ p1_literal_1076358[p2_res7__69_comb] ^ p2_res7__68_comb ^ p2_array_index_1077926_comb ^ p2_array_index_1077902_comb ^ p2_array_index_1077876_comb ^ p2_array_index_1077848_comb ^ p2_array_index_1077819_comb ^ p1_literal_1076345[p2_array_index_1077786_comb] ^ p2_array_index_1077787_comb;
  assign p2_res7__78_comb = p1_literal_1076345[p2_res7__77_comb] ^ p1_literal_1076347[p2_res7__76_comb] ^ p1_literal_1076349[p2_res7__75_comb] ^ p1_literal_1076351[p2_res7__74_comb] ^ p1_literal_1076353[p2_res7__73_comb] ^ p1_literal_1076355[p2_res7__72_comb] ^ p2_res7__71_comb ^ p1_literal_1076358[p2_res7__70_comb] ^ p2_res7__69_comb ^ p2_array_index_1077937_comb ^ p2_array_index_1077914_comb ^ p2_array_index_1077889_comb ^ p2_array_index_1077862_comb ^ p2_array_index_1077833_comb ^ p2_array_index_1077801_comb ^ p2_array_index_1077786_comb;
  assign p2_res7__79_comb = p1_literal_1076345[p2_res7__78_comb] ^ p1_literal_1076347[p2_res7__77_comb] ^ p1_literal_1076349[p2_res7__76_comb] ^ p1_literal_1076351[p2_res7__75_comb] ^ p1_literal_1076353[p2_res7__74_comb] ^ p1_literal_1076355[p2_res7__73_comb] ^ p2_res7__72_comb ^ p1_literal_1076358[p2_res7__71_comb] ^ p2_res7__70_comb ^ p2_array_index_1077947_comb ^ p2_array_index_1077925_comb ^ p2_array_index_1077901_comb ^ p2_array_index_1077875_comb ^ p2_array_index_1077847_comb ^ p2_array_index_1077818_comb ^ p2_array_index_1077785_comb;
  assign p2_res__4_comb = {p2_res7__79_comb, p2_res7__78_comb, p2_res7__77_comb, p2_res7__76_comb, p2_res7__75_comb, p2_res7__74_comb, p2_res7__73_comb, p2_res7__72_comb, p2_res7__71_comb, p2_res7__70_comb, p2_res7__69_comb, p2_res7__68_comb, p2_res7__67_comb, p2_res7__66_comb, p2_res7__65_comb, p2_res7__64_comb};
  assign p2_xor_1077987_comb = p2_res__4_comb ^ p1_xor_1076991;
  assign p2_addedKey__46_comb = p2_xor_1077987_comb ^ 128'ha74a_f7ef_ab73_df16_0dd2_0860_8b9e_fe06;
  assign p2_array_index_1078003_comb = p1_arr[p2_addedKey__46_comb[127:120]];
  assign p2_array_index_1078004_comb = p1_arr[p2_addedKey__46_comb[119:112]];
  assign p2_array_index_1078005_comb = p1_arr[p2_addedKey__46_comb[111:104]];
  assign p2_array_index_1078006_comb = p1_arr[p2_addedKey__46_comb[103:96]];
  assign p2_array_index_1078007_comb = p1_arr[p2_addedKey__46_comb[95:88]];
  assign p2_array_index_1078008_comb = p1_arr[p2_addedKey__46_comb[87:80]];
  assign p2_array_index_1078010_comb = p1_arr[p2_addedKey__46_comb[71:64]];
  assign p2_array_index_1078012_comb = p1_arr[p2_addedKey__46_comb[55:48]];
  assign p2_array_index_1078013_comb = p1_arr[p2_addedKey__46_comb[47:40]];
  assign p2_array_index_1078014_comb = p1_arr[p2_addedKey__46_comb[39:32]];
  assign p2_array_index_1078015_comb = p1_arr[p2_addedKey__46_comb[31:24]];
  assign p2_array_index_1078016_comb = p1_arr[p2_addedKey__46_comb[23:16]];
  assign p2_array_index_1078017_comb = p1_arr[p2_addedKey__46_comb[15:8]];
  assign p2_array_index_1078019_comb = p1_literal_1076345[p2_array_index_1078003_comb];
  assign p2_array_index_1078020_comb = p1_literal_1076347[p2_array_index_1078004_comb];
  assign p2_array_index_1078021_comb = p1_literal_1076349[p2_array_index_1078005_comb];
  assign p2_array_index_1078022_comb = p1_literal_1076351[p2_array_index_1078006_comb];
  assign p2_array_index_1078023_comb = p1_literal_1076353[p2_array_index_1078007_comb];
  assign p2_array_index_1078024_comb = p1_literal_1076355[p2_array_index_1078008_comb];
  assign p2_array_index_1078025_comb = p1_arr[p2_addedKey__46_comb[79:72]];
  assign p2_array_index_1078027_comb = p1_arr[p2_addedKey__46_comb[63:56]];
  assign p2_res7__80_comb = p2_array_index_1078019_comb ^ p2_array_index_1078020_comb ^ p2_array_index_1078021_comb ^ p2_array_index_1078022_comb ^ p2_array_index_1078023_comb ^ p2_array_index_1078024_comb ^ p2_array_index_1078025_comb ^ p1_literal_1076358[p2_array_index_1078010_comb] ^ p2_array_index_1078027_comb ^ p1_literal_1076355[p2_array_index_1078012_comb] ^ p1_literal_1076353[p2_array_index_1078013_comb] ^ p1_literal_1076351[p2_array_index_1078014_comb] ^ p1_literal_1076349[p2_array_index_1078015_comb] ^ p1_literal_1076347[p2_array_index_1078016_comb] ^ p1_literal_1076345[p2_array_index_1078017_comb] ^ p1_arr[p2_addedKey__46_comb[7:0]];
  assign p2_array_index_1078036_comb = p1_literal_1076345[p2_res7__80_comb];
  assign p2_array_index_1078037_comb = p1_literal_1076347[p2_array_index_1078003_comb];
  assign p2_array_index_1078038_comb = p1_literal_1076349[p2_array_index_1078004_comb];
  assign p2_array_index_1078039_comb = p1_literal_1076351[p2_array_index_1078005_comb];
  assign p2_array_index_1078040_comb = p1_literal_1076353[p2_array_index_1078006_comb];
  assign p2_array_index_1078041_comb = p1_literal_1076355[p2_array_index_1078007_comb];
  assign p2_res7__81_comb = p2_array_index_1078036_comb ^ p2_array_index_1078037_comb ^ p2_array_index_1078038_comb ^ p2_array_index_1078039_comb ^ p2_array_index_1078040_comb ^ p2_array_index_1078041_comb ^ p2_array_index_1078008_comb ^ p1_literal_1076358[p2_array_index_1078025_comb] ^ p2_array_index_1078010_comb ^ p1_literal_1076355[p2_array_index_1078027_comb] ^ p1_literal_1076353[p2_array_index_1078012_comb] ^ p1_literal_1076351[p2_array_index_1078013_comb] ^ p1_literal_1076349[p2_array_index_1078014_comb] ^ p1_literal_1076347[p2_array_index_1078015_comb] ^ p1_literal_1076345[p2_array_index_1078016_comb] ^ p2_array_index_1078017_comb;
  assign p2_array_index_1078051_comb = p1_literal_1076347[p2_res7__80_comb];
  assign p2_array_index_1078052_comb = p1_literal_1076349[p2_array_index_1078003_comb];
  assign p2_array_index_1078053_comb = p1_literal_1076351[p2_array_index_1078004_comb];
  assign p2_array_index_1078054_comb = p1_literal_1076353[p2_array_index_1078005_comb];
  assign p2_array_index_1078055_comb = p1_literal_1076355[p2_array_index_1078006_comb];
  assign p2_res7__82_comb = p1_literal_1076345[p2_res7__81_comb] ^ p2_array_index_1078051_comb ^ p2_array_index_1078052_comb ^ p2_array_index_1078053_comb ^ p2_array_index_1078054_comb ^ p2_array_index_1078055_comb ^ p2_array_index_1078007_comb ^ p1_literal_1076358[p2_array_index_1078008_comb] ^ p2_array_index_1078025_comb ^ p1_literal_1076355[p2_array_index_1078010_comb] ^ p1_literal_1076353[p2_array_index_1078027_comb] ^ p1_literal_1076351[p2_array_index_1078012_comb] ^ p1_literal_1076349[p2_array_index_1078013_comb] ^ p1_literal_1076347[p2_array_index_1078014_comb] ^ p1_literal_1076345[p2_array_index_1078015_comb] ^ p2_array_index_1078016_comb;
  assign p2_array_index_1078065_comb = p1_literal_1076347[p2_res7__81_comb];
  assign p2_array_index_1078066_comb = p1_literal_1076349[p2_res7__80_comb];
  assign p2_array_index_1078067_comb = p1_literal_1076351[p2_array_index_1078003_comb];
  assign p2_array_index_1078068_comb = p1_literal_1076353[p2_array_index_1078004_comb];
  assign p2_array_index_1078069_comb = p1_literal_1076355[p2_array_index_1078005_comb];
  assign p2_res7__83_comb = p1_literal_1076345[p2_res7__82_comb] ^ p2_array_index_1078065_comb ^ p2_array_index_1078066_comb ^ p2_array_index_1078067_comb ^ p2_array_index_1078068_comb ^ p2_array_index_1078069_comb ^ p2_array_index_1078006_comb ^ p1_literal_1076358[p2_array_index_1078007_comb] ^ p2_array_index_1078008_comb ^ p1_literal_1076355[p2_array_index_1078025_comb] ^ p1_literal_1076353[p2_array_index_1078010_comb] ^ p1_literal_1076351[p2_array_index_1078027_comb] ^ p1_literal_1076349[p2_array_index_1078012_comb] ^ p1_literal_1076347[p2_array_index_1078013_comb] ^ p1_literal_1076345[p2_array_index_1078014_comb] ^ p2_array_index_1078015_comb;
  assign p2_array_index_1078080_comb = p1_literal_1076349[p2_res7__81_comb];
  assign p2_array_index_1078081_comb = p1_literal_1076351[p2_res7__80_comb];
  assign p2_array_index_1078082_comb = p1_literal_1076353[p2_array_index_1078003_comb];
  assign p2_array_index_1078083_comb = p1_literal_1076355[p2_array_index_1078004_comb];
  assign p2_res7__84_comb = p1_literal_1076345[p2_res7__83_comb] ^ p1_literal_1076347[p2_res7__82_comb] ^ p2_array_index_1078080_comb ^ p2_array_index_1078081_comb ^ p2_array_index_1078082_comb ^ p2_array_index_1078083_comb ^ p2_array_index_1078005_comb ^ p1_literal_1076358[p2_array_index_1078006_comb] ^ p2_array_index_1078007_comb ^ p2_array_index_1078024_comb ^ p1_literal_1076353[p2_array_index_1078025_comb] ^ p1_literal_1076351[p2_array_index_1078010_comb] ^ p1_literal_1076349[p2_array_index_1078027_comb] ^ p1_literal_1076347[p2_array_index_1078012_comb] ^ p1_literal_1076345[p2_array_index_1078013_comb] ^ p2_array_index_1078014_comb;
  assign p2_array_index_1078093_comb = p1_literal_1076349[p2_res7__82_comb];
  assign p2_array_index_1078094_comb = p1_literal_1076351[p2_res7__81_comb];
  assign p2_array_index_1078095_comb = p1_literal_1076353[p2_res7__80_comb];
  assign p2_array_index_1078096_comb = p1_literal_1076355[p2_array_index_1078003_comb];
  assign p2_res7__85_comb = p1_literal_1076345[p2_res7__84_comb] ^ p1_literal_1076347[p2_res7__83_comb] ^ p2_array_index_1078093_comb ^ p2_array_index_1078094_comb ^ p2_array_index_1078095_comb ^ p2_array_index_1078096_comb ^ p2_array_index_1078004_comb ^ p1_literal_1076358[p2_array_index_1078005_comb] ^ p2_array_index_1078006_comb ^ p2_array_index_1078041_comb ^ p1_literal_1076353[p2_array_index_1078008_comb] ^ p1_literal_1076351[p2_array_index_1078025_comb] ^ p1_literal_1076349[p2_array_index_1078010_comb] ^ p1_literal_1076347[p2_array_index_1078027_comb] ^ p1_literal_1076345[p2_array_index_1078012_comb] ^ p2_array_index_1078013_comb;
  assign p2_array_index_1078107_comb = p1_literal_1076351[p2_res7__82_comb];
  assign p2_array_index_1078108_comb = p1_literal_1076353[p2_res7__81_comb];
  assign p2_array_index_1078109_comb = p1_literal_1076355[p2_res7__80_comb];
  assign p2_res7__86_comb = p1_literal_1076345[p2_res7__85_comb] ^ p1_literal_1076347[p2_res7__84_comb] ^ p1_literal_1076349[p2_res7__83_comb] ^ p2_array_index_1078107_comb ^ p2_array_index_1078108_comb ^ p2_array_index_1078109_comb ^ p2_array_index_1078003_comb ^ p1_literal_1076358[p2_array_index_1078004_comb] ^ p2_array_index_1078005_comb ^ p2_array_index_1078055_comb ^ p2_array_index_1078023_comb ^ p1_literal_1076351[p2_array_index_1078008_comb] ^ p1_literal_1076349[p2_array_index_1078025_comb] ^ p1_literal_1076347[p2_array_index_1078010_comb] ^ p1_literal_1076345[p2_array_index_1078027_comb] ^ p2_array_index_1078012_comb;
  assign p2_array_index_1078119_comb = p1_literal_1076351[p2_res7__83_comb];
  assign p2_array_index_1078120_comb = p1_literal_1076353[p2_res7__82_comb];
  assign p2_array_index_1078121_comb = p1_literal_1076355[p2_res7__81_comb];
  assign p2_res7__87_comb = p1_literal_1076345[p2_res7__86_comb] ^ p1_literal_1076347[p2_res7__85_comb] ^ p1_literal_1076349[p2_res7__84_comb] ^ p2_array_index_1078119_comb ^ p2_array_index_1078120_comb ^ p2_array_index_1078121_comb ^ p2_res7__80_comb ^ p1_literal_1076358[p2_array_index_1078003_comb] ^ p2_array_index_1078004_comb ^ p2_array_index_1078069_comb ^ p2_array_index_1078040_comb ^ p1_literal_1076351[p2_array_index_1078007_comb] ^ p1_literal_1076349[p2_array_index_1078008_comb] ^ p1_literal_1076347[p2_array_index_1078025_comb] ^ p1_literal_1076345[p2_array_index_1078010_comb] ^ p2_array_index_1078027_comb;
  assign p2_array_index_1078132_comb = p1_literal_1076353[p2_res7__83_comb];
  assign p2_array_index_1078133_comb = p1_literal_1076355[p2_res7__82_comb];
  assign p2_res7__88_comb = p1_literal_1076345[p2_res7__87_comb] ^ p1_literal_1076347[p2_res7__86_comb] ^ p1_literal_1076349[p2_res7__85_comb] ^ p1_literal_1076351[p2_res7__84_comb] ^ p2_array_index_1078132_comb ^ p2_array_index_1078133_comb ^ p2_res7__81_comb ^ p1_literal_1076358[p2_res7__80_comb] ^ p2_array_index_1078003_comb ^ p2_array_index_1078083_comb ^ p2_array_index_1078054_comb ^ p2_array_index_1078022_comb ^ p1_literal_1076349[p2_array_index_1078007_comb] ^ p1_literal_1076347[p2_array_index_1078008_comb] ^ p1_literal_1076345[p2_array_index_1078025_comb] ^ p2_array_index_1078010_comb;
  assign p2_array_index_1078143_comb = p1_literal_1076353[p2_res7__84_comb];
  assign p2_array_index_1078144_comb = p1_literal_1076355[p2_res7__83_comb];
  assign p2_res7__89_comb = p1_literal_1076345[p2_res7__88_comb] ^ p1_literal_1076347[p2_res7__87_comb] ^ p1_literal_1076349[p2_res7__86_comb] ^ p1_literal_1076351[p2_res7__85_comb] ^ p2_array_index_1078143_comb ^ p2_array_index_1078144_comb ^ p2_res7__82_comb ^ p1_literal_1076358[p2_res7__81_comb] ^ p2_res7__80_comb ^ p2_array_index_1078096_comb ^ p2_array_index_1078068_comb ^ p2_array_index_1078039_comb ^ p1_literal_1076349[p2_array_index_1078006_comb] ^ p1_literal_1076347[p2_array_index_1078007_comb] ^ p1_literal_1076345[p2_array_index_1078008_comb] ^ p2_array_index_1078025_comb;
  assign p2_array_index_1078155_comb = p1_literal_1076355[p2_res7__84_comb];
  assign p2_res7__90_comb = p1_literal_1076345[p2_res7__89_comb] ^ p1_literal_1076347[p2_res7__88_comb] ^ p1_literal_1076349[p2_res7__87_comb] ^ p1_literal_1076351[p2_res7__86_comb] ^ p1_literal_1076353[p2_res7__85_comb] ^ p2_array_index_1078155_comb ^ p2_res7__83_comb ^ p1_literal_1076358[p2_res7__82_comb] ^ p2_res7__81_comb ^ p2_array_index_1078109_comb ^ p2_array_index_1078082_comb ^ p2_array_index_1078053_comb ^ p2_array_index_1078021_comb ^ p1_literal_1076347[p2_array_index_1078006_comb] ^ p1_literal_1076345[p2_array_index_1078007_comb] ^ p2_array_index_1078008_comb;
  assign p2_array_index_1078165_comb = p1_literal_1076355[p2_res7__85_comb];
  assign p2_res7__91_comb = p1_literal_1076345[p2_res7__90_comb] ^ p1_literal_1076347[p2_res7__89_comb] ^ p1_literal_1076349[p2_res7__88_comb] ^ p1_literal_1076351[p2_res7__87_comb] ^ p1_literal_1076353[p2_res7__86_comb] ^ p2_array_index_1078165_comb ^ p2_res7__84_comb ^ p1_literal_1076358[p2_res7__83_comb] ^ p2_res7__82_comb ^ p2_array_index_1078121_comb ^ p2_array_index_1078095_comb ^ p2_array_index_1078067_comb ^ p2_array_index_1078038_comb ^ p1_literal_1076347[p2_array_index_1078005_comb] ^ p1_literal_1076345[p2_array_index_1078006_comb] ^ p2_array_index_1078007_comb;
  assign p2_res7__92_comb = p1_literal_1076345[p2_res7__91_comb] ^ p1_literal_1076347[p2_res7__90_comb] ^ p1_literal_1076349[p2_res7__89_comb] ^ p1_literal_1076351[p2_res7__88_comb] ^ p1_literal_1076353[p2_res7__87_comb] ^ p1_literal_1076355[p2_res7__86_comb] ^ p2_res7__85_comb ^ p1_literal_1076358[p2_res7__84_comb] ^ p2_res7__83_comb ^ p2_array_index_1078133_comb ^ p2_array_index_1078108_comb ^ p2_array_index_1078081_comb ^ p2_array_index_1078052_comb ^ p2_array_index_1078020_comb ^ p1_literal_1076345[p2_array_index_1078005_comb] ^ p2_array_index_1078006_comb;
  assign p2_res7__93_comb = p1_literal_1076345[p2_res7__92_comb] ^ p1_literal_1076347[p2_res7__91_comb] ^ p1_literal_1076349[p2_res7__90_comb] ^ p1_literal_1076351[p2_res7__89_comb] ^ p1_literal_1076353[p2_res7__88_comb] ^ p1_literal_1076355[p2_res7__87_comb] ^ p2_res7__86_comb ^ p1_literal_1076358[p2_res7__85_comb] ^ p2_res7__84_comb ^ p2_array_index_1078144_comb ^ p2_array_index_1078120_comb ^ p2_array_index_1078094_comb ^ p2_array_index_1078066_comb ^ p2_array_index_1078037_comb ^ p1_literal_1076345[p2_array_index_1078004_comb] ^ p2_array_index_1078005_comb;
  assign p2_res7__94_comb = p1_literal_1076345[p2_res7__93_comb] ^ p1_literal_1076347[p2_res7__92_comb] ^ p1_literal_1076349[p2_res7__91_comb] ^ p1_literal_1076351[p2_res7__90_comb] ^ p1_literal_1076353[p2_res7__89_comb] ^ p1_literal_1076355[p2_res7__88_comb] ^ p2_res7__87_comb ^ p1_literal_1076358[p2_res7__86_comb] ^ p2_res7__85_comb ^ p2_array_index_1078155_comb ^ p2_array_index_1078132_comb ^ p2_array_index_1078107_comb ^ p2_array_index_1078080_comb ^ p2_array_index_1078051_comb ^ p2_array_index_1078019_comb ^ p2_array_index_1078004_comb;
  assign p2_res7__95_comb = p1_literal_1076345[p2_res7__94_comb] ^ p1_literal_1076347[p2_res7__93_comb] ^ p1_literal_1076349[p2_res7__92_comb] ^ p1_literal_1076351[p2_res7__91_comb] ^ p1_literal_1076353[p2_res7__90_comb] ^ p1_literal_1076355[p2_res7__89_comb] ^ p2_res7__88_comb ^ p1_literal_1076358[p2_res7__87_comb] ^ p2_res7__86_comb ^ p2_array_index_1078165_comb ^ p2_array_index_1078143_comb ^ p2_array_index_1078119_comb ^ p2_array_index_1078093_comb ^ p2_array_index_1078065_comb ^ p2_array_index_1078036_comb ^ p2_array_index_1078003_comb;
  assign p2_res__5_comb = {p2_res7__95_comb, p2_res7__94_comb, p2_res7__93_comb, p2_res7__92_comb, p2_res7__91_comb, p2_res7__90_comb, p2_res7__89_comb, p2_res7__88_comb, p2_res7__87_comb, p2_res7__86_comb, p2_res7__85_comb, p2_res7__84_comb, p2_res7__83_comb, p2_res7__82_comb, p2_res7__81_comb, p2_res7__80_comb};
  assign p2_xor_1078205_comb = p2_res__5_comb ^ p2_xor_1077769_comb;
  assign p2_addedKey__47_comb = p2_xor_1078205_comb ^ 128'hc9e8_819d_c73b_a5ae_50f5_b570_561a_6a07;
  assign p2_array_index_1078221_comb = p1_arr[p2_addedKey__47_comb[127:120]];
  assign p2_array_index_1078222_comb = p1_arr[p2_addedKey__47_comb[119:112]];
  assign p2_array_index_1078223_comb = p1_arr[p2_addedKey__47_comb[111:104]];
  assign p2_array_index_1078224_comb = p1_arr[p2_addedKey__47_comb[103:96]];
  assign p2_array_index_1078225_comb = p1_arr[p2_addedKey__47_comb[95:88]];
  assign p2_array_index_1078226_comb = p1_arr[p2_addedKey__47_comb[87:80]];
  assign p2_array_index_1078228_comb = p1_arr[p2_addedKey__47_comb[71:64]];
  assign p2_array_index_1078230_comb = p1_arr[p2_addedKey__47_comb[55:48]];
  assign p2_array_index_1078231_comb = p1_arr[p2_addedKey__47_comb[47:40]];
  assign p2_array_index_1078232_comb = p1_arr[p2_addedKey__47_comb[39:32]];
  assign p2_array_index_1078233_comb = p1_arr[p2_addedKey__47_comb[31:24]];
  assign p2_array_index_1078234_comb = p1_arr[p2_addedKey__47_comb[23:16]];
  assign p2_array_index_1078235_comb = p1_arr[p2_addedKey__47_comb[15:8]];
  assign p2_array_index_1078237_comb = p1_literal_1076345[p2_array_index_1078221_comb];
  assign p2_array_index_1078238_comb = p1_literal_1076347[p2_array_index_1078222_comb];
  assign p2_array_index_1078239_comb = p1_literal_1076349[p2_array_index_1078223_comb];
  assign p2_array_index_1078240_comb = p1_literal_1076351[p2_array_index_1078224_comb];
  assign p2_array_index_1078241_comb = p1_literal_1076353[p2_array_index_1078225_comb];
  assign p2_array_index_1078242_comb = p1_literal_1076355[p2_array_index_1078226_comb];
  assign p2_array_index_1078243_comb = p1_arr[p2_addedKey__47_comb[79:72]];
  assign p2_array_index_1078245_comb = p1_arr[p2_addedKey__47_comb[63:56]];
  assign p2_res7__96_comb = p2_array_index_1078237_comb ^ p2_array_index_1078238_comb ^ p2_array_index_1078239_comb ^ p2_array_index_1078240_comb ^ p2_array_index_1078241_comb ^ p2_array_index_1078242_comb ^ p2_array_index_1078243_comb ^ p1_literal_1076358[p2_array_index_1078228_comb] ^ p2_array_index_1078245_comb ^ p1_literal_1076355[p2_array_index_1078230_comb] ^ p1_literal_1076353[p2_array_index_1078231_comb] ^ p1_literal_1076351[p2_array_index_1078232_comb] ^ p1_literal_1076349[p2_array_index_1078233_comb] ^ p1_literal_1076347[p2_array_index_1078234_comb] ^ p1_literal_1076345[p2_array_index_1078235_comb] ^ p1_arr[p2_addedKey__47_comb[7:0]];
  assign p2_array_index_1078254_comb = p1_literal_1076345[p2_res7__96_comb];
  assign p2_array_index_1078255_comb = p1_literal_1076347[p2_array_index_1078221_comb];
  assign p2_array_index_1078256_comb = p1_literal_1076349[p2_array_index_1078222_comb];
  assign p2_array_index_1078257_comb = p1_literal_1076351[p2_array_index_1078223_comb];
  assign p2_array_index_1078258_comb = p1_literal_1076353[p2_array_index_1078224_comb];
  assign p2_array_index_1078259_comb = p1_literal_1076355[p2_array_index_1078225_comb];
  assign p2_res7__97_comb = p2_array_index_1078254_comb ^ p2_array_index_1078255_comb ^ p2_array_index_1078256_comb ^ p2_array_index_1078257_comb ^ p2_array_index_1078258_comb ^ p2_array_index_1078259_comb ^ p2_array_index_1078226_comb ^ p1_literal_1076358[p2_array_index_1078243_comb] ^ p2_array_index_1078228_comb ^ p1_literal_1076355[p2_array_index_1078245_comb] ^ p1_literal_1076353[p2_array_index_1078230_comb] ^ p1_literal_1076351[p2_array_index_1078231_comb] ^ p1_literal_1076349[p2_array_index_1078232_comb] ^ p1_literal_1076347[p2_array_index_1078233_comb] ^ p1_literal_1076345[p2_array_index_1078234_comb] ^ p2_array_index_1078235_comb;
  assign p2_array_index_1078269_comb = p1_literal_1076347[p2_res7__96_comb];
  assign p2_array_index_1078270_comb = p1_literal_1076349[p2_array_index_1078221_comb];
  assign p2_array_index_1078271_comb = p1_literal_1076351[p2_array_index_1078222_comb];
  assign p2_array_index_1078272_comb = p1_literal_1076353[p2_array_index_1078223_comb];
  assign p2_array_index_1078273_comb = p1_literal_1076355[p2_array_index_1078224_comb];
  assign p2_res7__98_comb = p1_literal_1076345[p2_res7__97_comb] ^ p2_array_index_1078269_comb ^ p2_array_index_1078270_comb ^ p2_array_index_1078271_comb ^ p2_array_index_1078272_comb ^ p2_array_index_1078273_comb ^ p2_array_index_1078225_comb ^ p1_literal_1076358[p2_array_index_1078226_comb] ^ p2_array_index_1078243_comb ^ p1_literal_1076355[p2_array_index_1078228_comb] ^ p1_literal_1076353[p2_array_index_1078245_comb] ^ p1_literal_1076351[p2_array_index_1078230_comb] ^ p1_literal_1076349[p2_array_index_1078231_comb] ^ p1_literal_1076347[p2_array_index_1078232_comb] ^ p1_literal_1076345[p2_array_index_1078233_comb] ^ p2_array_index_1078234_comb;
  assign p2_array_index_1078283_comb = p1_literal_1076347[p2_res7__97_comb];
  assign p2_array_index_1078284_comb = p1_literal_1076349[p2_res7__96_comb];
  assign p2_array_index_1078285_comb = p1_literal_1076351[p2_array_index_1078221_comb];
  assign p2_array_index_1078286_comb = p1_literal_1076353[p2_array_index_1078222_comb];
  assign p2_array_index_1078287_comb = p1_literal_1076355[p2_array_index_1078223_comb];
  assign p2_res7__99_comb = p1_literal_1076345[p2_res7__98_comb] ^ p2_array_index_1078283_comb ^ p2_array_index_1078284_comb ^ p2_array_index_1078285_comb ^ p2_array_index_1078286_comb ^ p2_array_index_1078287_comb ^ p2_array_index_1078224_comb ^ p1_literal_1076358[p2_array_index_1078225_comb] ^ p2_array_index_1078226_comb ^ p1_literal_1076355[p2_array_index_1078243_comb] ^ p1_literal_1076353[p2_array_index_1078228_comb] ^ p1_literal_1076351[p2_array_index_1078245_comb] ^ p1_literal_1076349[p2_array_index_1078230_comb] ^ p1_literal_1076347[p2_array_index_1078231_comb] ^ p1_literal_1076345[p2_array_index_1078232_comb] ^ p2_array_index_1078233_comb;
  assign p2_array_index_1078298_comb = p1_literal_1076349[p2_res7__97_comb];
  assign p2_array_index_1078299_comb = p1_literal_1076351[p2_res7__96_comb];
  assign p2_array_index_1078300_comb = p1_literal_1076353[p2_array_index_1078221_comb];
  assign p2_array_index_1078301_comb = p1_literal_1076355[p2_array_index_1078222_comb];
  assign p2_res7__100_comb = p1_literal_1076345[p2_res7__99_comb] ^ p1_literal_1076347[p2_res7__98_comb] ^ p2_array_index_1078298_comb ^ p2_array_index_1078299_comb ^ p2_array_index_1078300_comb ^ p2_array_index_1078301_comb ^ p2_array_index_1078223_comb ^ p1_literal_1076358[p2_array_index_1078224_comb] ^ p2_array_index_1078225_comb ^ p2_array_index_1078242_comb ^ p1_literal_1076353[p2_array_index_1078243_comb] ^ p1_literal_1076351[p2_array_index_1078228_comb] ^ p1_literal_1076349[p2_array_index_1078245_comb] ^ p1_literal_1076347[p2_array_index_1078230_comb] ^ p1_literal_1076345[p2_array_index_1078231_comb] ^ p2_array_index_1078232_comb;
  assign p2_array_index_1078311_comb = p1_literal_1076349[p2_res7__98_comb];
  assign p2_array_index_1078312_comb = p1_literal_1076351[p2_res7__97_comb];
  assign p2_array_index_1078313_comb = p1_literal_1076353[p2_res7__96_comb];
  assign p2_array_index_1078314_comb = p1_literal_1076355[p2_array_index_1078221_comb];
  assign p2_res7__101_comb = p1_literal_1076345[p2_res7__100_comb] ^ p1_literal_1076347[p2_res7__99_comb] ^ p2_array_index_1078311_comb ^ p2_array_index_1078312_comb ^ p2_array_index_1078313_comb ^ p2_array_index_1078314_comb ^ p2_array_index_1078222_comb ^ p1_literal_1076358[p2_array_index_1078223_comb] ^ p2_array_index_1078224_comb ^ p2_array_index_1078259_comb ^ p1_literal_1076353[p2_array_index_1078226_comb] ^ p1_literal_1076351[p2_array_index_1078243_comb] ^ p1_literal_1076349[p2_array_index_1078228_comb] ^ p1_literal_1076347[p2_array_index_1078245_comb] ^ p1_literal_1076345[p2_array_index_1078230_comb] ^ p2_array_index_1078231_comb;
  assign p2_array_index_1078325_comb = p1_literal_1076351[p2_res7__98_comb];
  assign p2_array_index_1078326_comb = p1_literal_1076353[p2_res7__97_comb];
  assign p2_array_index_1078327_comb = p1_literal_1076355[p2_res7__96_comb];
  assign p2_res7__102_comb = p1_literal_1076345[p2_res7__101_comb] ^ p1_literal_1076347[p2_res7__100_comb] ^ p1_literal_1076349[p2_res7__99_comb] ^ p2_array_index_1078325_comb ^ p2_array_index_1078326_comb ^ p2_array_index_1078327_comb ^ p2_array_index_1078221_comb ^ p1_literal_1076358[p2_array_index_1078222_comb] ^ p2_array_index_1078223_comb ^ p2_array_index_1078273_comb ^ p2_array_index_1078241_comb ^ p1_literal_1076351[p2_array_index_1078226_comb] ^ p1_literal_1076349[p2_array_index_1078243_comb] ^ p1_literal_1076347[p2_array_index_1078228_comb] ^ p1_literal_1076345[p2_array_index_1078245_comb] ^ p2_array_index_1078230_comb;
  assign p2_array_index_1078337_comb = p1_literal_1076351[p2_res7__99_comb];
  assign p2_array_index_1078338_comb = p1_literal_1076353[p2_res7__98_comb];
  assign p2_array_index_1078339_comb = p1_literal_1076355[p2_res7__97_comb];
  assign p2_res7__103_comb = p1_literal_1076345[p2_res7__102_comb] ^ p1_literal_1076347[p2_res7__101_comb] ^ p1_literal_1076349[p2_res7__100_comb] ^ p2_array_index_1078337_comb ^ p2_array_index_1078338_comb ^ p2_array_index_1078339_comb ^ p2_res7__96_comb ^ p1_literal_1076358[p2_array_index_1078221_comb] ^ p2_array_index_1078222_comb ^ p2_array_index_1078287_comb ^ p2_array_index_1078258_comb ^ p1_literal_1076351[p2_array_index_1078225_comb] ^ p1_literal_1076349[p2_array_index_1078226_comb] ^ p1_literal_1076347[p2_array_index_1078243_comb] ^ p1_literal_1076345[p2_array_index_1078228_comb] ^ p2_array_index_1078245_comb;
  assign p2_array_index_1078350_comb = p1_literal_1076353[p2_res7__99_comb];
  assign p2_array_index_1078351_comb = p1_literal_1076355[p2_res7__98_comb];
  assign p2_res7__104_comb = p1_literal_1076345[p2_res7__103_comb] ^ p1_literal_1076347[p2_res7__102_comb] ^ p1_literal_1076349[p2_res7__101_comb] ^ p1_literal_1076351[p2_res7__100_comb] ^ p2_array_index_1078350_comb ^ p2_array_index_1078351_comb ^ p2_res7__97_comb ^ p1_literal_1076358[p2_res7__96_comb] ^ p2_array_index_1078221_comb ^ p2_array_index_1078301_comb ^ p2_array_index_1078272_comb ^ p2_array_index_1078240_comb ^ p1_literal_1076349[p2_array_index_1078225_comb] ^ p1_literal_1076347[p2_array_index_1078226_comb] ^ p1_literal_1076345[p2_array_index_1078243_comb] ^ p2_array_index_1078228_comb;
  assign p2_array_index_1078361_comb = p1_literal_1076353[p2_res7__100_comb];
  assign p2_array_index_1078362_comb = p1_literal_1076355[p2_res7__99_comb];
  assign p2_res7__105_comb = p1_literal_1076345[p2_res7__104_comb] ^ p1_literal_1076347[p2_res7__103_comb] ^ p1_literal_1076349[p2_res7__102_comb] ^ p1_literal_1076351[p2_res7__101_comb] ^ p2_array_index_1078361_comb ^ p2_array_index_1078362_comb ^ p2_res7__98_comb ^ p1_literal_1076358[p2_res7__97_comb] ^ p2_res7__96_comb ^ p2_array_index_1078314_comb ^ p2_array_index_1078286_comb ^ p2_array_index_1078257_comb ^ p1_literal_1076349[p2_array_index_1078224_comb] ^ p1_literal_1076347[p2_array_index_1078225_comb] ^ p1_literal_1076345[p2_array_index_1078226_comb] ^ p2_array_index_1078243_comb;
  assign p2_array_index_1078373_comb = p1_literal_1076355[p2_res7__100_comb];
  assign p2_res7__106_comb = p1_literal_1076345[p2_res7__105_comb] ^ p1_literal_1076347[p2_res7__104_comb] ^ p1_literal_1076349[p2_res7__103_comb] ^ p1_literal_1076351[p2_res7__102_comb] ^ p1_literal_1076353[p2_res7__101_comb] ^ p2_array_index_1078373_comb ^ p2_res7__99_comb ^ p1_literal_1076358[p2_res7__98_comb] ^ p2_res7__97_comb ^ p2_array_index_1078327_comb ^ p2_array_index_1078300_comb ^ p2_array_index_1078271_comb ^ p2_array_index_1078239_comb ^ p1_literal_1076347[p2_array_index_1078224_comb] ^ p1_literal_1076345[p2_array_index_1078225_comb] ^ p2_array_index_1078226_comb;
  assign p2_array_index_1078383_comb = p1_literal_1076355[p2_res7__101_comb];
  assign p2_res7__107_comb = p1_literal_1076345[p2_res7__106_comb] ^ p1_literal_1076347[p2_res7__105_comb] ^ p1_literal_1076349[p2_res7__104_comb] ^ p1_literal_1076351[p2_res7__103_comb] ^ p1_literal_1076353[p2_res7__102_comb] ^ p2_array_index_1078383_comb ^ p2_res7__100_comb ^ p1_literal_1076358[p2_res7__99_comb] ^ p2_res7__98_comb ^ p2_array_index_1078339_comb ^ p2_array_index_1078313_comb ^ p2_array_index_1078285_comb ^ p2_array_index_1078256_comb ^ p1_literal_1076347[p2_array_index_1078223_comb] ^ p1_literal_1076345[p2_array_index_1078224_comb] ^ p2_array_index_1078225_comb;
  assign p2_res7__108_comb = p1_literal_1076345[p2_res7__107_comb] ^ p1_literal_1076347[p2_res7__106_comb] ^ p1_literal_1076349[p2_res7__105_comb] ^ p1_literal_1076351[p2_res7__104_comb] ^ p1_literal_1076353[p2_res7__103_comb] ^ p1_literal_1076355[p2_res7__102_comb] ^ p2_res7__101_comb ^ p1_literal_1076358[p2_res7__100_comb] ^ p2_res7__99_comb ^ p2_array_index_1078351_comb ^ p2_array_index_1078326_comb ^ p2_array_index_1078299_comb ^ p2_array_index_1078270_comb ^ p2_array_index_1078238_comb ^ p1_literal_1076345[p2_array_index_1078223_comb] ^ p2_array_index_1078224_comb;
  assign p2_res7__109_comb = p1_literal_1076345[p2_res7__108_comb] ^ p1_literal_1076347[p2_res7__107_comb] ^ p1_literal_1076349[p2_res7__106_comb] ^ p1_literal_1076351[p2_res7__105_comb] ^ p1_literal_1076353[p2_res7__104_comb] ^ p1_literal_1076355[p2_res7__103_comb] ^ p2_res7__102_comb ^ p1_literal_1076358[p2_res7__101_comb] ^ p2_res7__100_comb ^ p2_array_index_1078362_comb ^ p2_array_index_1078338_comb ^ p2_array_index_1078312_comb ^ p2_array_index_1078284_comb ^ p2_array_index_1078255_comb ^ p1_literal_1076345[p2_array_index_1078222_comb] ^ p2_array_index_1078223_comb;
  assign p2_res7__110_comb = p1_literal_1076345[p2_res7__109_comb] ^ p1_literal_1076347[p2_res7__108_comb] ^ p1_literal_1076349[p2_res7__107_comb] ^ p1_literal_1076351[p2_res7__106_comb] ^ p1_literal_1076353[p2_res7__105_comb] ^ p1_literal_1076355[p2_res7__104_comb] ^ p2_res7__103_comb ^ p1_literal_1076358[p2_res7__102_comb] ^ p2_res7__101_comb ^ p2_array_index_1078373_comb ^ p2_array_index_1078350_comb ^ p2_array_index_1078325_comb ^ p2_array_index_1078298_comb ^ p2_array_index_1078269_comb ^ p2_array_index_1078237_comb ^ p2_array_index_1078222_comb;
  assign p2_res7__111_comb = p1_literal_1076345[p2_res7__110_comb] ^ p1_literal_1076347[p2_res7__109_comb] ^ p1_literal_1076349[p2_res7__108_comb] ^ p1_literal_1076351[p2_res7__107_comb] ^ p1_literal_1076353[p2_res7__106_comb] ^ p1_literal_1076355[p2_res7__105_comb] ^ p2_res7__104_comb ^ p1_literal_1076358[p2_res7__103_comb] ^ p2_res7__102_comb ^ p2_array_index_1078383_comb ^ p2_array_index_1078361_comb ^ p2_array_index_1078337_comb ^ p2_array_index_1078311_comb ^ p2_array_index_1078283_comb ^ p2_array_index_1078254_comb ^ p2_array_index_1078221_comb;
  assign p2_res__6_comb = {p2_res7__111_comb, p2_res7__110_comb, p2_res7__109_comb, p2_res7__108_comb, p2_res7__107_comb, p2_res7__106_comb, p2_res7__105_comb, p2_res7__104_comb, p2_res7__103_comb, p2_res7__102_comb, p2_res7__101_comb, p2_res7__100_comb, p2_res7__99_comb, p2_res7__98_comb, p2_res7__97_comb, p2_res7__96_comb};
  assign p2_k3_comb = p2_res__6_comb ^ p2_xor_1077987_comb;
  assign p2_addedKey__48_comb = p2_k3_comb ^ 128'hf659_3616_e605_5689_adfb_a180_27aa_2a08;
  assign p2_array_index_1078439_comb = p1_arr[p2_addedKey__48_comb[127:120]];
  assign p2_array_index_1078440_comb = p1_arr[p2_addedKey__48_comb[119:112]];
  assign p2_array_index_1078441_comb = p1_arr[p2_addedKey__48_comb[111:104]];
  assign p2_array_index_1078442_comb = p1_arr[p2_addedKey__48_comb[103:96]];
  assign p2_array_index_1078443_comb = p1_arr[p2_addedKey__48_comb[95:88]];
  assign p2_array_index_1078444_comb = p1_arr[p2_addedKey__48_comb[87:80]];
  assign p2_array_index_1078446_comb = p1_arr[p2_addedKey__48_comb[71:64]];
  assign p2_array_index_1078448_comb = p1_arr[p2_addedKey__48_comb[55:48]];
  assign p2_array_index_1078449_comb = p1_arr[p2_addedKey__48_comb[47:40]];
  assign p2_array_index_1078450_comb = p1_arr[p2_addedKey__48_comb[39:32]];
  assign p2_array_index_1078451_comb = p1_arr[p2_addedKey__48_comb[31:24]];
  assign p2_array_index_1078452_comb = p1_arr[p2_addedKey__48_comb[23:16]];
  assign p2_array_index_1078453_comb = p1_arr[p2_addedKey__48_comb[15:8]];
  assign p2_array_index_1078455_comb = p1_literal_1076345[p2_array_index_1078439_comb];
  assign p2_array_index_1078456_comb = p1_literal_1076347[p2_array_index_1078440_comb];
  assign p2_array_index_1078457_comb = p1_literal_1076349[p2_array_index_1078441_comb];
  assign p2_array_index_1078458_comb = p1_literal_1076351[p2_array_index_1078442_comb];
  assign p2_array_index_1078459_comb = p1_literal_1076353[p2_array_index_1078443_comb];
  assign p2_array_index_1078460_comb = p1_literal_1076355[p2_array_index_1078444_comb];
  assign p2_array_index_1078461_comb = p1_arr[p2_addedKey__48_comb[79:72]];
  assign p2_array_index_1078463_comb = p1_arr[p2_addedKey__48_comb[63:56]];
  assign p2_res7__112_comb = p2_array_index_1078455_comb ^ p2_array_index_1078456_comb ^ p2_array_index_1078457_comb ^ p2_array_index_1078458_comb ^ p2_array_index_1078459_comb ^ p2_array_index_1078460_comb ^ p2_array_index_1078461_comb ^ p1_literal_1076358[p2_array_index_1078446_comb] ^ p2_array_index_1078463_comb ^ p1_literal_1076355[p2_array_index_1078448_comb] ^ p1_literal_1076353[p2_array_index_1078449_comb] ^ p1_literal_1076351[p2_array_index_1078450_comb] ^ p1_literal_1076349[p2_array_index_1078451_comb] ^ p1_literal_1076347[p2_array_index_1078452_comb] ^ p1_literal_1076345[p2_array_index_1078453_comb] ^ p1_arr[p2_addedKey__48_comb[7:0]];
  assign p2_array_index_1078472_comb = p1_literal_1076345[p2_res7__112_comb];
  assign p2_array_index_1078473_comb = p1_literal_1076347[p2_array_index_1078439_comb];
  assign p2_array_index_1078474_comb = p1_literal_1076349[p2_array_index_1078440_comb];
  assign p2_array_index_1078475_comb = p1_literal_1076351[p2_array_index_1078441_comb];
  assign p2_array_index_1078476_comb = p1_literal_1076353[p2_array_index_1078442_comb];
  assign p2_array_index_1078477_comb = p1_literal_1076355[p2_array_index_1078443_comb];
  assign p2_res7__113_comb = p2_array_index_1078472_comb ^ p2_array_index_1078473_comb ^ p2_array_index_1078474_comb ^ p2_array_index_1078475_comb ^ p2_array_index_1078476_comb ^ p2_array_index_1078477_comb ^ p2_array_index_1078444_comb ^ p1_literal_1076358[p2_array_index_1078461_comb] ^ p2_array_index_1078446_comb ^ p1_literal_1076355[p2_array_index_1078463_comb] ^ p1_literal_1076353[p2_array_index_1078448_comb] ^ p1_literal_1076351[p2_array_index_1078449_comb] ^ p1_literal_1076349[p2_array_index_1078450_comb] ^ p1_literal_1076347[p2_array_index_1078451_comb] ^ p1_literal_1076345[p2_array_index_1078452_comb] ^ p2_array_index_1078453_comb;
  assign p2_array_index_1078487_comb = p1_literal_1076347[p2_res7__112_comb];
  assign p2_array_index_1078488_comb = p1_literal_1076349[p2_array_index_1078439_comb];
  assign p2_array_index_1078489_comb = p1_literal_1076351[p2_array_index_1078440_comb];
  assign p2_array_index_1078490_comb = p1_literal_1076353[p2_array_index_1078441_comb];
  assign p2_array_index_1078491_comb = p1_literal_1076355[p2_array_index_1078442_comb];
  assign p2_res7__114_comb = p1_literal_1076345[p2_res7__113_comb] ^ p2_array_index_1078487_comb ^ p2_array_index_1078488_comb ^ p2_array_index_1078489_comb ^ p2_array_index_1078490_comb ^ p2_array_index_1078491_comb ^ p2_array_index_1078443_comb ^ p1_literal_1076358[p2_array_index_1078444_comb] ^ p2_array_index_1078461_comb ^ p1_literal_1076355[p2_array_index_1078446_comb] ^ p1_literal_1076353[p2_array_index_1078463_comb] ^ p1_literal_1076351[p2_array_index_1078448_comb] ^ p1_literal_1076349[p2_array_index_1078449_comb] ^ p1_literal_1076347[p2_array_index_1078450_comb] ^ p1_literal_1076345[p2_array_index_1078451_comb] ^ p2_array_index_1078452_comb;
  assign p2_array_index_1078501_comb = p1_literal_1076347[p2_res7__113_comb];
  assign p2_array_index_1078502_comb = p1_literal_1076349[p2_res7__112_comb];
  assign p2_array_index_1078503_comb = p1_literal_1076351[p2_array_index_1078439_comb];
  assign p2_array_index_1078504_comb = p1_literal_1076353[p2_array_index_1078440_comb];
  assign p2_array_index_1078505_comb = p1_literal_1076355[p2_array_index_1078441_comb];
  assign p2_res7__115_comb = p1_literal_1076345[p2_res7__114_comb] ^ p2_array_index_1078501_comb ^ p2_array_index_1078502_comb ^ p2_array_index_1078503_comb ^ p2_array_index_1078504_comb ^ p2_array_index_1078505_comb ^ p2_array_index_1078442_comb ^ p1_literal_1076358[p2_array_index_1078443_comb] ^ p2_array_index_1078444_comb ^ p1_literal_1076355[p2_array_index_1078461_comb] ^ p1_literal_1076353[p2_array_index_1078446_comb] ^ p1_literal_1076351[p2_array_index_1078463_comb] ^ p1_literal_1076349[p2_array_index_1078448_comb] ^ p1_literal_1076347[p2_array_index_1078449_comb] ^ p1_literal_1076345[p2_array_index_1078450_comb] ^ p2_array_index_1078451_comb;
  assign p2_array_index_1078516_comb = p1_literal_1076349[p2_res7__113_comb];
  assign p2_array_index_1078517_comb = p1_literal_1076351[p2_res7__112_comb];
  assign p2_array_index_1078518_comb = p1_literal_1076353[p2_array_index_1078439_comb];
  assign p2_array_index_1078519_comb = p1_literal_1076355[p2_array_index_1078440_comb];
  assign p2_res7__116_comb = p1_literal_1076345[p2_res7__115_comb] ^ p1_literal_1076347[p2_res7__114_comb] ^ p2_array_index_1078516_comb ^ p2_array_index_1078517_comb ^ p2_array_index_1078518_comb ^ p2_array_index_1078519_comb ^ p2_array_index_1078441_comb ^ p1_literal_1076358[p2_array_index_1078442_comb] ^ p2_array_index_1078443_comb ^ p2_array_index_1078460_comb ^ p1_literal_1076353[p2_array_index_1078461_comb] ^ p1_literal_1076351[p2_array_index_1078446_comb] ^ p1_literal_1076349[p2_array_index_1078463_comb] ^ p1_literal_1076347[p2_array_index_1078448_comb] ^ p1_literal_1076345[p2_array_index_1078449_comb] ^ p2_array_index_1078450_comb;

  // Registers for pipe stage 2:
  reg [127:0] p2_xor_1078205;
  reg [127:0] p2_k3;
  reg [7:0] p2_array_index_1078439;
  reg [7:0] p2_array_index_1078440;
  reg [7:0] p2_array_index_1078441;
  reg [7:0] p2_array_index_1078442;
  reg [7:0] p2_array_index_1078443;
  reg [7:0] p2_array_index_1078444;
  reg [7:0] p2_array_index_1078446;
  reg [7:0] p2_array_index_1078448;
  reg [7:0] p2_array_index_1078449;
  reg [7:0] p2_array_index_1078455;
  reg [7:0] p2_array_index_1078456;
  reg [7:0] p2_array_index_1078457;
  reg [7:0] p2_array_index_1078458;
  reg [7:0] p2_array_index_1078459;
  reg [7:0] p2_array_index_1078461;
  reg [7:0] p2_array_index_1078463;
  reg [7:0] p2_res7__112;
  reg [7:0] p2_array_index_1078472;
  reg [7:0] p2_array_index_1078473;
  reg [7:0] p2_array_index_1078474;
  reg [7:0] p2_array_index_1078475;
  reg [7:0] p2_array_index_1078476;
  reg [7:0] p2_array_index_1078477;
  reg [7:0] p2_res7__113;
  reg [7:0] p2_array_index_1078487;
  reg [7:0] p2_array_index_1078488;
  reg [7:0] p2_array_index_1078489;
  reg [7:0] p2_array_index_1078490;
  reg [7:0] p2_array_index_1078491;
  reg [7:0] p2_res7__114;
  reg [7:0] p2_array_index_1078501;
  reg [7:0] p2_array_index_1078502;
  reg [7:0] p2_array_index_1078503;
  reg [7:0] p2_array_index_1078504;
  reg [7:0] p2_array_index_1078505;
  reg [7:0] p2_res7__115;
  reg [7:0] p2_array_index_1078516;
  reg [7:0] p2_array_index_1078517;
  reg [7:0] p2_array_index_1078518;
  reg [7:0] p2_array_index_1078519;
  reg [7:0] p2_res7__116;
  reg [127:0] p2_res__33;
  reg [7:0] p3_arr[256];
  reg [7:0] p3_literal_1076345[256];
  reg [7:0] p3_literal_1076347[256];
  reg [7:0] p3_literal_1076349[256];
  reg [7:0] p3_literal_1076351[256];
  reg [7:0] p3_literal_1076353[256];
  reg [7:0] p3_literal_1076355[256];
  reg [7:0] p3_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p2_xor_1078205 <= p2_xor_1078205_comb;
    p2_k3 <= p2_k3_comb;
    p2_array_index_1078439 <= p2_array_index_1078439_comb;
    p2_array_index_1078440 <= p2_array_index_1078440_comb;
    p2_array_index_1078441 <= p2_array_index_1078441_comb;
    p2_array_index_1078442 <= p2_array_index_1078442_comb;
    p2_array_index_1078443 <= p2_array_index_1078443_comb;
    p2_array_index_1078444 <= p2_array_index_1078444_comb;
    p2_array_index_1078446 <= p2_array_index_1078446_comb;
    p2_array_index_1078448 <= p2_array_index_1078448_comb;
    p2_array_index_1078449 <= p2_array_index_1078449_comb;
    p2_array_index_1078455 <= p2_array_index_1078455_comb;
    p2_array_index_1078456 <= p2_array_index_1078456_comb;
    p2_array_index_1078457 <= p2_array_index_1078457_comb;
    p2_array_index_1078458 <= p2_array_index_1078458_comb;
    p2_array_index_1078459 <= p2_array_index_1078459_comb;
    p2_array_index_1078461 <= p2_array_index_1078461_comb;
    p2_array_index_1078463 <= p2_array_index_1078463_comb;
    p2_res7__112 <= p2_res7__112_comb;
    p2_array_index_1078472 <= p2_array_index_1078472_comb;
    p2_array_index_1078473 <= p2_array_index_1078473_comb;
    p2_array_index_1078474 <= p2_array_index_1078474_comb;
    p2_array_index_1078475 <= p2_array_index_1078475_comb;
    p2_array_index_1078476 <= p2_array_index_1078476_comb;
    p2_array_index_1078477 <= p2_array_index_1078477_comb;
    p2_res7__113 <= p2_res7__113_comb;
    p2_array_index_1078487 <= p2_array_index_1078487_comb;
    p2_array_index_1078488 <= p2_array_index_1078488_comb;
    p2_array_index_1078489 <= p2_array_index_1078489_comb;
    p2_array_index_1078490 <= p2_array_index_1078490_comb;
    p2_array_index_1078491 <= p2_array_index_1078491_comb;
    p2_res7__114 <= p2_res7__114_comb;
    p2_array_index_1078501 <= p2_array_index_1078501_comb;
    p2_array_index_1078502 <= p2_array_index_1078502_comb;
    p2_array_index_1078503 <= p2_array_index_1078503_comb;
    p2_array_index_1078504 <= p2_array_index_1078504_comb;
    p2_array_index_1078505 <= p2_array_index_1078505_comb;
    p2_res7__115 <= p2_res7__115_comb;
    p2_array_index_1078516 <= p2_array_index_1078516_comb;
    p2_array_index_1078517 <= p2_array_index_1078517_comb;
    p2_array_index_1078518 <= p2_array_index_1078518_comb;
    p2_array_index_1078519 <= p2_array_index_1078519_comb;
    p2_res7__116 <= p2_res7__116_comb;
    p2_res__33 <= p1_res__33;
    p3_arr <= p2_arr;
    p3_literal_1076345 <= p2_literal_1076345;
    p3_literal_1076347 <= p2_literal_1076347;
    p3_literal_1076349 <= p2_literal_1076349;
    p3_literal_1076351 <= p2_literal_1076351;
    p3_literal_1076353 <= p2_literal_1076353;
    p3_literal_1076355 <= p2_literal_1076355;
    p3_literal_1076358 <= p2_literal_1076358;
  end

  // ===== Pipe stage 3:
  wire [7:0] p3_array_index_1078633_comb;
  wire [7:0] p3_array_index_1078634_comb;
  wire [7:0] p3_array_index_1078635_comb;
  wire [7:0] p3_array_index_1078636_comb;
  wire [7:0] p3_res7__117_comb;
  wire [7:0] p3_array_index_1078647_comb;
  wire [7:0] p3_array_index_1078648_comb;
  wire [7:0] p3_array_index_1078649_comb;
  wire [7:0] p3_res7__118_comb;
  wire [7:0] p3_array_index_1078659_comb;
  wire [7:0] p3_array_index_1078660_comb;
  wire [7:0] p3_array_index_1078661_comb;
  wire [7:0] p3_res7__119_comb;
  wire [7:0] p3_array_index_1078672_comb;
  wire [7:0] p3_array_index_1078673_comb;
  wire [7:0] p3_res7__120_comb;
  wire [7:0] p3_array_index_1078683_comb;
  wire [7:0] p3_array_index_1078684_comb;
  wire [7:0] p3_res7__121_comb;
  wire [7:0] p3_array_index_1078695_comb;
  wire [7:0] p3_res7__122_comb;
  wire [7:0] p3_array_index_1078705_comb;
  wire [7:0] p3_res7__123_comb;
  wire [7:0] p3_res7__124_comb;
  wire [7:0] p3_res7__125_comb;
  wire [7:0] p3_res7__126_comb;
  wire [7:0] p3_res7__127_comb;
  wire [127:0] p3_res__7_comb;
  wire [127:0] p3_k2_comb;
  wire [127:0] p3_addedKey__49_comb;
  wire [7:0] p3_array_index_1078761_comb;
  wire [7:0] p3_array_index_1078762_comb;
  wire [7:0] p3_array_index_1078763_comb;
  wire [7:0] p3_array_index_1078764_comb;
  wire [7:0] p3_array_index_1078765_comb;
  wire [7:0] p3_array_index_1078766_comb;
  wire [7:0] p3_array_index_1078768_comb;
  wire [7:0] p3_array_index_1078770_comb;
  wire [7:0] p3_array_index_1078771_comb;
  wire [7:0] p3_array_index_1078772_comb;
  wire [7:0] p3_array_index_1078773_comb;
  wire [7:0] p3_array_index_1078774_comb;
  wire [7:0] p3_array_index_1078775_comb;
  wire [7:0] p3_array_index_1078777_comb;
  wire [7:0] p3_array_index_1078778_comb;
  wire [7:0] p3_array_index_1078779_comb;
  wire [7:0] p3_array_index_1078780_comb;
  wire [7:0] p3_array_index_1078781_comb;
  wire [7:0] p3_array_index_1078782_comb;
  wire [7:0] p3_array_index_1078783_comb;
  wire [7:0] p3_array_index_1078785_comb;
  wire [7:0] p3_res7__128_comb;
  wire [7:0] p3_array_index_1078794_comb;
  wire [7:0] p3_array_index_1078795_comb;
  wire [7:0] p3_array_index_1078796_comb;
  wire [7:0] p3_array_index_1078797_comb;
  wire [7:0] p3_array_index_1078798_comb;
  wire [7:0] p3_array_index_1078799_comb;
  wire [7:0] p3_res7__129_comb;
  wire [7:0] p3_array_index_1078809_comb;
  wire [7:0] p3_array_index_1078810_comb;
  wire [7:0] p3_array_index_1078811_comb;
  wire [7:0] p3_array_index_1078812_comb;
  wire [7:0] p3_array_index_1078813_comb;
  wire [7:0] p3_res7__130_comb;
  wire [7:0] p3_array_index_1078823_comb;
  wire [7:0] p3_array_index_1078824_comb;
  wire [7:0] p3_array_index_1078825_comb;
  wire [7:0] p3_array_index_1078826_comb;
  wire [7:0] p3_array_index_1078827_comb;
  wire [7:0] p3_res7__131_comb;
  wire [7:0] p3_array_index_1078838_comb;
  wire [7:0] p3_array_index_1078839_comb;
  wire [7:0] p3_array_index_1078840_comb;
  wire [7:0] p3_array_index_1078841_comb;
  wire [7:0] p3_res7__132_comb;
  wire [7:0] p3_array_index_1078851_comb;
  wire [7:0] p3_array_index_1078852_comb;
  wire [7:0] p3_array_index_1078853_comb;
  wire [7:0] p3_array_index_1078854_comb;
  wire [7:0] p3_res7__133_comb;
  wire [7:0] p3_array_index_1078865_comb;
  wire [7:0] p3_array_index_1078866_comb;
  wire [7:0] p3_array_index_1078867_comb;
  wire [7:0] p3_res7__134_comb;
  wire [7:0] p3_array_index_1078877_comb;
  wire [7:0] p3_array_index_1078878_comb;
  wire [7:0] p3_array_index_1078879_comb;
  wire [7:0] p3_res7__135_comb;
  wire [7:0] p3_array_index_1078890_comb;
  wire [7:0] p3_array_index_1078891_comb;
  wire [7:0] p3_res7__136_comb;
  wire [7:0] p3_array_index_1078901_comb;
  wire [7:0] p3_array_index_1078902_comb;
  wire [7:0] p3_res7__137_comb;
  wire [7:0] p3_array_index_1078913_comb;
  wire [7:0] p3_res7__138_comb;
  wire [7:0] p3_array_index_1078923_comb;
  wire [7:0] p3_res7__139_comb;
  wire [7:0] p3_res7__140_comb;
  wire [7:0] p3_res7__141_comb;
  wire [7:0] p3_res7__142_comb;
  wire [7:0] p3_res7__143_comb;
  wire [127:0] p3_res__8_comb;
  wire [127:0] p3_xor_1078963_comb;
  wire [127:0] p3_addedKey__50_comb;
  wire [7:0] p3_array_index_1078979_comb;
  wire [7:0] p3_array_index_1078980_comb;
  wire [7:0] p3_array_index_1078981_comb;
  wire [7:0] p3_array_index_1078982_comb;
  wire [7:0] p3_array_index_1078983_comb;
  wire [7:0] p3_array_index_1078984_comb;
  wire [7:0] p3_array_index_1078986_comb;
  wire [7:0] p3_array_index_1078988_comb;
  wire [7:0] p3_array_index_1078989_comb;
  wire [7:0] p3_array_index_1078990_comb;
  wire [7:0] p3_array_index_1078991_comb;
  wire [7:0] p3_array_index_1078992_comb;
  wire [7:0] p3_array_index_1078993_comb;
  wire [127:0] p3_addedKey__34_comb;
  wire [7:0] p3_array_index_1078995_comb;
  wire [7:0] p3_array_index_1078996_comb;
  wire [7:0] p3_array_index_1078997_comb;
  wire [7:0] p3_array_index_1078998_comb;
  wire [7:0] p3_array_index_1078999_comb;
  wire [7:0] p3_array_index_1079000_comb;
  wire [7:0] p3_array_index_1079001_comb;
  wire [7:0] p3_array_index_1079003_comb;
  wire [7:0] p3_res7__144_comb;
  wire [7:0] p3_array_index_1079414_comb;
  wire [7:0] p3_array_index_1079415_comb;
  wire [7:0] p3_array_index_1079416_comb;
  wire [7:0] p3_array_index_1079417_comb;
  wire [7:0] p3_array_index_1079418_comb;
  wire [7:0] p3_array_index_1079419_comb;
  wire [7:0] p3_array_index_1079421_comb;
  wire [7:0] p3_array_index_1079423_comb;
  wire [7:0] p3_array_index_1079424_comb;
  wire [7:0] p3_array_index_1079425_comb;
  wire [7:0] p3_array_index_1079426_comb;
  wire [7:0] p3_array_index_1079427_comb;
  wire [7:0] p3_array_index_1079428_comb;
  wire [7:0] p3_array_index_1079012_comb;
  wire [7:0] p3_array_index_1079013_comb;
  wire [7:0] p3_array_index_1079014_comb;
  wire [7:0] p3_array_index_1079015_comb;
  wire [7:0] p3_array_index_1079016_comb;
  wire [7:0] p3_array_index_1079017_comb;
  wire [7:0] p3_array_index_1079430_comb;
  wire [7:0] p3_array_index_1079431_comb;
  wire [7:0] p3_array_index_1079432_comb;
  wire [7:0] p3_array_index_1079433_comb;
  wire [7:0] p3_array_index_1079434_comb;
  wire [7:0] p3_array_index_1079435_comb;
  wire [7:0] p3_array_index_1079436_comb;
  wire [7:0] p3_array_index_1079438_comb;
  wire [7:0] p3_res7__145_comb;
  wire [7:0] p3_res7__544_comb;
  wire [7:0] p3_array_index_1079027_comb;
  wire [7:0] p3_array_index_1079028_comb;
  wire [7:0] p3_array_index_1079029_comb;
  wire [7:0] p3_array_index_1079030_comb;
  wire [7:0] p3_array_index_1079031_comb;
  wire [7:0] p3_array_index_1079447_comb;
  wire [7:0] p3_array_index_1079448_comb;
  wire [7:0] p3_array_index_1079449_comb;
  wire [7:0] p3_array_index_1079450_comb;
  wire [7:0] p3_array_index_1079451_comb;
  wire [7:0] p3_array_index_1079452_comb;
  wire [7:0] p3_res7__146_comb;
  wire [7:0] p3_res7__545_comb;
  wire [7:0] p3_array_index_1079041_comb;
  wire [7:0] p3_array_index_1079042_comb;
  wire [7:0] p3_array_index_1079043_comb;
  wire [7:0] p3_array_index_1079044_comb;
  wire [7:0] p3_array_index_1079045_comb;
  wire [7:0] p3_array_index_1079462_comb;
  wire [7:0] p3_array_index_1079463_comb;
  wire [7:0] p3_array_index_1079464_comb;
  wire [7:0] p3_array_index_1079465_comb;
  wire [7:0] p3_array_index_1079466_comb;
  wire [7:0] p3_res7__147_comb;
  wire [7:0] p3_res7__546_comb;
  wire [7:0] p3_array_index_1079056_comb;
  wire [7:0] p3_array_index_1079057_comb;
  wire [7:0] p3_array_index_1079058_comb;
  wire [7:0] p3_array_index_1079059_comb;
  wire [7:0] p3_array_index_1079476_comb;
  wire [7:0] p3_array_index_1079477_comb;
  wire [7:0] p3_array_index_1079478_comb;
  wire [7:0] p3_array_index_1079479_comb;
  wire [7:0] p3_array_index_1079480_comb;
  wire [7:0] p3_res7__148_comb;
  wire [7:0] p3_res7__547_comb;
  wire [7:0] p3_array_index_1079069_comb;
  wire [7:0] p3_array_index_1079070_comb;
  wire [7:0] p3_array_index_1079071_comb;
  wire [7:0] p3_array_index_1079072_comb;
  wire [7:0] p3_array_index_1079491_comb;
  wire [7:0] p3_array_index_1079492_comb;
  wire [7:0] p3_array_index_1079493_comb;
  wire [7:0] p3_array_index_1079494_comb;
  wire [7:0] p3_res7__149_comb;
  wire [7:0] p3_res7__548_comb;
  wire [7:0] p3_array_index_1079083_comb;
  wire [7:0] p3_array_index_1079084_comb;
  wire [7:0] p3_array_index_1079085_comb;
  wire [7:0] p3_array_index_1079504_comb;
  wire [7:0] p3_array_index_1079505_comb;
  wire [7:0] p3_array_index_1079506_comb;
  wire [7:0] p3_array_index_1079507_comb;
  wire [7:0] p3_res7__150_comb;
  wire [7:0] p3_res7__549_comb;
  wire [7:0] p3_array_index_1079095_comb;
  wire [7:0] p3_array_index_1079096_comb;
  wire [7:0] p3_array_index_1079097_comb;
  wire [7:0] p3_array_index_1079518_comb;
  wire [7:0] p3_array_index_1079519_comb;
  wire [7:0] p3_array_index_1079520_comb;
  wire [7:0] p3_res7__151_comb;
  wire [7:0] p3_res7__550_comb;
  wire [7:0] p3_array_index_1079108_comb;
  wire [7:0] p3_array_index_1079109_comb;
  wire [7:0] p3_array_index_1079530_comb;
  wire [7:0] p3_array_index_1079531_comb;
  wire [7:0] p3_array_index_1079532_comb;
  wire [7:0] p3_res7__152_comb;
  wire [7:0] p3_res7__551_comb;
  wire [7:0] p3_array_index_1079119_comb;
  wire [7:0] p3_array_index_1079120_comb;
  wire [7:0] p3_array_index_1079543_comb;
  wire [7:0] p3_array_index_1079544_comb;
  wire [7:0] p3_res7__153_comb;
  wire [7:0] p3_res7__552_comb;
  wire [7:0] p3_array_index_1079131_comb;
  wire [7:0] p3_array_index_1079554_comb;
  wire [7:0] p3_array_index_1079555_comb;
  wire [7:0] p3_res7__154_comb;
  wire [7:0] p3_res7__553_comb;
  wire [7:0] p3_array_index_1079141_comb;
  wire [7:0] p3_array_index_1079566_comb;
  wire [7:0] p3_res7__155_comb;
  wire [7:0] p3_res7__554_comb;
  wire [7:0] p3_array_index_1079576_comb;
  wire [7:0] p3_res7__156_comb;
  wire [7:0] p3_res7__555_comb;
  wire [7:0] p3_res7__157_comb;
  wire [7:0] p3_res7__556_comb;
  wire [7:0] p3_res7__158_comb;
  wire [7:0] p3_res7__557_comb;
  wire [7:0] p3_res7__159_comb;
  wire [7:0] p3_res7__558_comb;
  wire [127:0] p3_res__9_comb;
  wire [127:0] p3_xor_1079181_comb;
  wire [7:0] p3_res7__559_comb;
  wire [127:0] p3_addedKey__51_comb;
  wire [127:0] p3_res__34_comb;
  wire [127:0] p3_addedKey__35_comb;
  wire [7:0] p3_array_index_1079197_comb;
  wire [7:0] p3_array_index_1079198_comb;
  wire [7:0] p3_array_index_1079199_comb;
  wire [7:0] p3_array_index_1079200_comb;
  wire [7:0] p3_array_index_1079201_comb;
  wire [7:0] p3_array_index_1079202_comb;
  wire [7:0] p3_array_index_1079204_comb;
  wire [7:0] p3_array_index_1079206_comb;
  wire [7:0] p3_array_index_1079207_comb;
  wire [7:0] p3_array_index_1079208_comb;
  wire [7:0] p3_array_index_1079209_comb;
  wire [7:0] p3_array_index_1079210_comb;
  wire [7:0] p3_array_index_1079211_comb;
  wire [7:0] p3_array_index_1079213_comb;
  wire [7:0] p3_array_index_1079214_comb;
  wire [7:0] p3_array_index_1079215_comb;
  wire [7:0] p3_array_index_1079216_comb;
  wire [7:0] p3_array_index_1079217_comb;
  wire [7:0] p3_array_index_1079218_comb;
  wire [7:0] p3_array_index_1079219_comb;
  wire [7:0] p3_array_index_1079221_comb;
  wire [7:0] p3_array_index_1079630_comb;
  wire [7:0] p3_array_index_1079631_comb;
  wire [7:0] p3_array_index_1079632_comb;
  wire [7:0] p3_array_index_1079633_comb;
  wire [7:0] p3_array_index_1079634_comb;
  wire [7:0] p3_array_index_1079635_comb;
  wire [7:0] p3_array_index_1079637_comb;
  wire [7:0] p3_array_index_1079639_comb;
  wire [7:0] p3_array_index_1079640_comb;
  wire [7:0] p3_array_index_1079641_comb;
  wire [7:0] p3_array_index_1079642_comb;
  wire [7:0] p3_array_index_1079643_comb;
  wire [7:0] p3_array_index_1079644_comb;
  wire [7:0] p3_res7__160_comb;
  wire [7:0] p3_array_index_1079646_comb;
  wire [7:0] p3_array_index_1079647_comb;
  wire [7:0] p3_array_index_1079648_comb;
  wire [7:0] p3_array_index_1079649_comb;
  wire [7:0] p3_array_index_1079650_comb;
  wire [7:0] p3_array_index_1079651_comb;
  wire [7:0] p3_array_index_1079652_comb;
  wire [7:0] p3_array_index_1079654_comb;
  wire [7:0] p3_array_index_1079230_comb;
  wire [7:0] p3_array_index_1079231_comb;
  wire [7:0] p3_array_index_1079232_comb;
  wire [7:0] p3_array_index_1079233_comb;
  wire [7:0] p3_array_index_1079234_comb;
  wire [7:0] p3_array_index_1079235_comb;
  wire [7:0] p3_res7__560_comb;
  wire [7:0] p3_res7__161_comb;
  wire [7:0] p3_array_index_1079663_comb;
  wire [7:0] p3_array_index_1079664_comb;
  wire [7:0] p3_array_index_1079665_comb;
  wire [7:0] p3_array_index_1079666_comb;
  wire [7:0] p3_array_index_1079667_comb;
  wire [7:0] p3_array_index_1079668_comb;
  wire [7:0] p3_array_index_1079245_comb;
  wire [7:0] p3_array_index_1079246_comb;
  wire [7:0] p3_array_index_1079247_comb;
  wire [7:0] p3_array_index_1079248_comb;
  wire [7:0] p3_array_index_1079249_comb;
  wire [7:0] p3_res7__561_comb;
  wire [7:0] p3_res7__162_comb;
  wire [7:0] p3_array_index_1079678_comb;
  wire [7:0] p3_array_index_1079679_comb;
  wire [7:0] p3_array_index_1079680_comb;
  wire [7:0] p3_array_index_1079681_comb;
  wire [7:0] p3_array_index_1079682_comb;
  wire [7:0] p3_array_index_1079259_comb;
  wire [7:0] p3_array_index_1079260_comb;
  wire [7:0] p3_array_index_1079261_comb;
  wire [7:0] p3_array_index_1079262_comb;
  wire [7:0] p3_array_index_1079263_comb;
  wire [7:0] p3_res7__562_comb;
  wire [7:0] p3_res7__163_comb;
  wire [7:0] p3_array_index_1079692_comb;
  wire [7:0] p3_array_index_1079693_comb;
  wire [7:0] p3_array_index_1079694_comb;
  wire [7:0] p3_array_index_1079695_comb;
  wire [7:0] p3_array_index_1079696_comb;
  wire [7:0] p3_array_index_1079274_comb;
  wire [7:0] p3_array_index_1079275_comb;
  wire [7:0] p3_array_index_1079276_comb;
  wire [7:0] p3_array_index_1079277_comb;
  wire [7:0] p3_res7__563_comb;
  wire [7:0] p3_res7__164_comb;
  wire [7:0] p3_array_index_1079707_comb;
  wire [7:0] p3_array_index_1079708_comb;
  wire [7:0] p3_array_index_1079709_comb;
  wire [7:0] p3_array_index_1079710_comb;
  wire [7:0] p3_array_index_1079287_comb;
  wire [7:0] p3_array_index_1079288_comb;
  wire [7:0] p3_array_index_1079289_comb;
  wire [7:0] p3_array_index_1079290_comb;
  wire [7:0] p3_res7__564_comb;
  wire [7:0] p3_res7__165_comb;
  wire [7:0] p3_array_index_1079720_comb;
  wire [7:0] p3_array_index_1079721_comb;
  wire [7:0] p3_array_index_1079722_comb;
  wire [7:0] p3_array_index_1079723_comb;
  wire [7:0] p3_array_index_1079301_comb;
  wire [7:0] p3_array_index_1079302_comb;
  wire [7:0] p3_array_index_1079303_comb;
  wire [7:0] p3_res7__565_comb;
  wire [7:0] p3_res7__166_comb;
  wire [7:0] p3_array_index_1079734_comb;
  wire [7:0] p3_array_index_1079735_comb;
  wire [7:0] p3_array_index_1079736_comb;
  wire [7:0] p3_array_index_1079313_comb;
  wire [7:0] p3_array_index_1079314_comb;
  wire [7:0] p3_array_index_1079315_comb;
  wire [7:0] p3_res7__566_comb;
  wire [7:0] p3_res7__167_comb;
  wire [7:0] p3_array_index_1079746_comb;
  wire [7:0] p3_array_index_1079747_comb;
  wire [7:0] p3_array_index_1079748_comb;
  wire [7:0] p3_array_index_1079326_comb;
  wire [7:0] p3_array_index_1079327_comb;
  wire [7:0] p3_res7__567_comb;
  wire [7:0] p3_res7__168_comb;
  wire [7:0] p3_array_index_1079759_comb;
  wire [7:0] p3_array_index_1079760_comb;
  wire [7:0] p3_array_index_1079337_comb;
  wire [7:0] p3_array_index_1079338_comb;
  wire [7:0] p3_res7__568_comb;
  wire [7:0] p3_res7__169_comb;
  wire [7:0] p3_array_index_1079770_comb;
  wire [7:0] p3_array_index_1079771_comb;
  wire [7:0] p3_array_index_1079349_comb;
  wire [7:0] p3_res7__569_comb;
  wire [7:0] p3_res7__170_comb;
  wire [7:0] p3_array_index_1079782_comb;
  wire [7:0] p3_array_index_1079359_comb;
  wire [7:0] p3_res7__570_comb;
  wire [7:0] p3_res7__171_comb;
  wire [7:0] p3_array_index_1079792_comb;
  wire [7:0] p3_res7__571_comb;
  wire [7:0] p3_res7__172_comb;
  wire [7:0] p3_res7__572_comb;
  wire [7:0] p3_res7__173_comb;
  wire [7:0] p3_res7__573_comb;
  wire [7:0] p3_res7__174_comb;
  wire [7:0] p3_res7__574_comb;
  wire [7:0] p3_res7__175_comb;
  wire [127:0] p3_res__10_comb;
  wire [7:0] p3_res7__575_comb;
  wire [127:0] p3_xor_1079399_comb;
  wire [127:0] p3_res__35_comb;
  assign p3_array_index_1078633_comb = p2_literal_1076349[p2_res7__114];
  assign p3_array_index_1078634_comb = p2_literal_1076351[p2_res7__113];
  assign p3_array_index_1078635_comb = p2_literal_1076353[p2_res7__112];
  assign p3_array_index_1078636_comb = p2_literal_1076355[p2_array_index_1078439];
  assign p3_res7__117_comb = p2_literal_1076345[p2_res7__116] ^ p2_literal_1076347[p2_res7__115] ^ p3_array_index_1078633_comb ^ p3_array_index_1078634_comb ^ p3_array_index_1078635_comb ^ p3_array_index_1078636_comb ^ p2_array_index_1078440 ^ p2_literal_1076358[p2_array_index_1078441] ^ p2_array_index_1078442 ^ p2_array_index_1078477 ^ p2_literal_1076353[p2_array_index_1078444] ^ p2_literal_1076351[p2_array_index_1078461] ^ p2_literal_1076349[p2_array_index_1078446] ^ p2_literal_1076347[p2_array_index_1078463] ^ p2_literal_1076345[p2_array_index_1078448] ^ p2_array_index_1078449;
  assign p3_array_index_1078647_comb = p2_literal_1076351[p2_res7__114];
  assign p3_array_index_1078648_comb = p2_literal_1076353[p2_res7__113];
  assign p3_array_index_1078649_comb = p2_literal_1076355[p2_res7__112];
  assign p3_res7__118_comb = p2_literal_1076345[p3_res7__117_comb] ^ p2_literal_1076347[p2_res7__116] ^ p2_literal_1076349[p2_res7__115] ^ p3_array_index_1078647_comb ^ p3_array_index_1078648_comb ^ p3_array_index_1078649_comb ^ p2_array_index_1078439 ^ p2_literal_1076358[p2_array_index_1078440] ^ p2_array_index_1078441 ^ p2_array_index_1078491 ^ p2_array_index_1078459 ^ p2_literal_1076351[p2_array_index_1078444] ^ p2_literal_1076349[p2_array_index_1078461] ^ p2_literal_1076347[p2_array_index_1078446] ^ p2_literal_1076345[p2_array_index_1078463] ^ p2_array_index_1078448;
  assign p3_array_index_1078659_comb = p2_literal_1076351[p2_res7__115];
  assign p3_array_index_1078660_comb = p2_literal_1076353[p2_res7__114];
  assign p3_array_index_1078661_comb = p2_literal_1076355[p2_res7__113];
  assign p3_res7__119_comb = p2_literal_1076345[p3_res7__118_comb] ^ p2_literal_1076347[p3_res7__117_comb] ^ p2_literal_1076349[p2_res7__116] ^ p3_array_index_1078659_comb ^ p3_array_index_1078660_comb ^ p3_array_index_1078661_comb ^ p2_res7__112 ^ p2_literal_1076358[p2_array_index_1078439] ^ p2_array_index_1078440 ^ p2_array_index_1078505 ^ p2_array_index_1078476 ^ p2_literal_1076351[p2_array_index_1078443] ^ p2_literal_1076349[p2_array_index_1078444] ^ p2_literal_1076347[p2_array_index_1078461] ^ p2_literal_1076345[p2_array_index_1078446] ^ p2_array_index_1078463;
  assign p3_array_index_1078672_comb = p2_literal_1076353[p2_res7__115];
  assign p3_array_index_1078673_comb = p2_literal_1076355[p2_res7__114];
  assign p3_res7__120_comb = p2_literal_1076345[p3_res7__119_comb] ^ p2_literal_1076347[p3_res7__118_comb] ^ p2_literal_1076349[p3_res7__117_comb] ^ p2_literal_1076351[p2_res7__116] ^ p3_array_index_1078672_comb ^ p3_array_index_1078673_comb ^ p2_res7__113 ^ p2_literal_1076358[p2_res7__112] ^ p2_array_index_1078439 ^ p2_array_index_1078519 ^ p2_array_index_1078490 ^ p2_array_index_1078458 ^ p2_literal_1076349[p2_array_index_1078443] ^ p2_literal_1076347[p2_array_index_1078444] ^ p2_literal_1076345[p2_array_index_1078461] ^ p2_array_index_1078446;
  assign p3_array_index_1078683_comb = p2_literal_1076353[p2_res7__116];
  assign p3_array_index_1078684_comb = p2_literal_1076355[p2_res7__115];
  assign p3_res7__121_comb = p2_literal_1076345[p3_res7__120_comb] ^ p2_literal_1076347[p3_res7__119_comb] ^ p2_literal_1076349[p3_res7__118_comb] ^ p2_literal_1076351[p3_res7__117_comb] ^ p3_array_index_1078683_comb ^ p3_array_index_1078684_comb ^ p2_res7__114 ^ p2_literal_1076358[p2_res7__113] ^ p2_res7__112 ^ p3_array_index_1078636_comb ^ p2_array_index_1078504 ^ p2_array_index_1078475 ^ p2_literal_1076349[p2_array_index_1078442] ^ p2_literal_1076347[p2_array_index_1078443] ^ p2_literal_1076345[p2_array_index_1078444] ^ p2_array_index_1078461;
  assign p3_array_index_1078695_comb = p2_literal_1076355[p2_res7__116];
  assign p3_res7__122_comb = p2_literal_1076345[p3_res7__121_comb] ^ p2_literal_1076347[p3_res7__120_comb] ^ p2_literal_1076349[p3_res7__119_comb] ^ p2_literal_1076351[p3_res7__118_comb] ^ p2_literal_1076353[p3_res7__117_comb] ^ p3_array_index_1078695_comb ^ p2_res7__115 ^ p2_literal_1076358[p2_res7__114] ^ p2_res7__113 ^ p3_array_index_1078649_comb ^ p2_array_index_1078518 ^ p2_array_index_1078489 ^ p2_array_index_1078457 ^ p2_literal_1076347[p2_array_index_1078442] ^ p2_literal_1076345[p2_array_index_1078443] ^ p2_array_index_1078444;
  assign p3_array_index_1078705_comb = p2_literal_1076355[p3_res7__117_comb];
  assign p3_res7__123_comb = p2_literal_1076345[p3_res7__122_comb] ^ p2_literal_1076347[p3_res7__121_comb] ^ p2_literal_1076349[p3_res7__120_comb] ^ p2_literal_1076351[p3_res7__119_comb] ^ p2_literal_1076353[p3_res7__118_comb] ^ p3_array_index_1078705_comb ^ p2_res7__116 ^ p2_literal_1076358[p2_res7__115] ^ p2_res7__114 ^ p3_array_index_1078661_comb ^ p3_array_index_1078635_comb ^ p2_array_index_1078503 ^ p2_array_index_1078474 ^ p2_literal_1076347[p2_array_index_1078441] ^ p2_literal_1076345[p2_array_index_1078442] ^ p2_array_index_1078443;
  assign p3_res7__124_comb = p2_literal_1076345[p3_res7__123_comb] ^ p2_literal_1076347[p3_res7__122_comb] ^ p2_literal_1076349[p3_res7__121_comb] ^ p2_literal_1076351[p3_res7__120_comb] ^ p2_literal_1076353[p3_res7__119_comb] ^ p2_literal_1076355[p3_res7__118_comb] ^ p3_res7__117_comb ^ p2_literal_1076358[p2_res7__116] ^ p2_res7__115 ^ p3_array_index_1078673_comb ^ p3_array_index_1078648_comb ^ p2_array_index_1078517 ^ p2_array_index_1078488 ^ p2_array_index_1078456 ^ p2_literal_1076345[p2_array_index_1078441] ^ p2_array_index_1078442;
  assign p3_res7__125_comb = p2_literal_1076345[p3_res7__124_comb] ^ p2_literal_1076347[p3_res7__123_comb] ^ p2_literal_1076349[p3_res7__122_comb] ^ p2_literal_1076351[p3_res7__121_comb] ^ p2_literal_1076353[p3_res7__120_comb] ^ p2_literal_1076355[p3_res7__119_comb] ^ p3_res7__118_comb ^ p2_literal_1076358[p3_res7__117_comb] ^ p2_res7__116 ^ p3_array_index_1078684_comb ^ p3_array_index_1078660_comb ^ p3_array_index_1078634_comb ^ p2_array_index_1078502 ^ p2_array_index_1078473 ^ p2_literal_1076345[p2_array_index_1078440] ^ p2_array_index_1078441;
  assign p3_res7__126_comb = p2_literal_1076345[p3_res7__125_comb] ^ p2_literal_1076347[p3_res7__124_comb] ^ p2_literal_1076349[p3_res7__123_comb] ^ p2_literal_1076351[p3_res7__122_comb] ^ p2_literal_1076353[p3_res7__121_comb] ^ p2_literal_1076355[p3_res7__120_comb] ^ p3_res7__119_comb ^ p2_literal_1076358[p3_res7__118_comb] ^ p3_res7__117_comb ^ p3_array_index_1078695_comb ^ p3_array_index_1078672_comb ^ p3_array_index_1078647_comb ^ p2_array_index_1078516 ^ p2_array_index_1078487 ^ p2_array_index_1078455 ^ p2_array_index_1078440;
  assign p3_res7__127_comb = p2_literal_1076345[p3_res7__126_comb] ^ p2_literal_1076347[p3_res7__125_comb] ^ p2_literal_1076349[p3_res7__124_comb] ^ p2_literal_1076351[p3_res7__123_comb] ^ p2_literal_1076353[p3_res7__122_comb] ^ p2_literal_1076355[p3_res7__121_comb] ^ p3_res7__120_comb ^ p2_literal_1076358[p3_res7__119_comb] ^ p3_res7__118_comb ^ p3_array_index_1078705_comb ^ p3_array_index_1078683_comb ^ p3_array_index_1078659_comb ^ p3_array_index_1078633_comb ^ p2_array_index_1078501 ^ p2_array_index_1078472 ^ p2_array_index_1078439;
  assign p3_res__7_comb = {p3_res7__127_comb, p3_res7__126_comb, p3_res7__125_comb, p3_res7__124_comb, p3_res7__123_comb, p3_res7__122_comb, p3_res7__121_comb, p3_res7__120_comb, p3_res7__119_comb, p3_res7__118_comb, p3_res7__117_comb, p2_res7__116, p2_res7__115, p2_res7__114, p2_res7__113, p2_res7__112};
  assign p3_k2_comb = p3_res__7_comb ^ p2_xor_1078205;
  assign p3_addedKey__49_comb = p3_k2_comb ^ 128'h98fb_4064_8a4d_2c31_f0dc_1c90_fa2e_be09;
  assign p3_array_index_1078761_comb = p2_arr[p3_addedKey__49_comb[127:120]];
  assign p3_array_index_1078762_comb = p2_arr[p3_addedKey__49_comb[119:112]];
  assign p3_array_index_1078763_comb = p2_arr[p3_addedKey__49_comb[111:104]];
  assign p3_array_index_1078764_comb = p2_arr[p3_addedKey__49_comb[103:96]];
  assign p3_array_index_1078765_comb = p2_arr[p3_addedKey__49_comb[95:88]];
  assign p3_array_index_1078766_comb = p2_arr[p3_addedKey__49_comb[87:80]];
  assign p3_array_index_1078768_comb = p2_arr[p3_addedKey__49_comb[71:64]];
  assign p3_array_index_1078770_comb = p2_arr[p3_addedKey__49_comb[55:48]];
  assign p3_array_index_1078771_comb = p2_arr[p3_addedKey__49_comb[47:40]];
  assign p3_array_index_1078772_comb = p2_arr[p3_addedKey__49_comb[39:32]];
  assign p3_array_index_1078773_comb = p2_arr[p3_addedKey__49_comb[31:24]];
  assign p3_array_index_1078774_comb = p2_arr[p3_addedKey__49_comb[23:16]];
  assign p3_array_index_1078775_comb = p2_arr[p3_addedKey__49_comb[15:8]];
  assign p3_array_index_1078777_comb = p2_literal_1076345[p3_array_index_1078761_comb];
  assign p3_array_index_1078778_comb = p2_literal_1076347[p3_array_index_1078762_comb];
  assign p3_array_index_1078779_comb = p2_literal_1076349[p3_array_index_1078763_comb];
  assign p3_array_index_1078780_comb = p2_literal_1076351[p3_array_index_1078764_comb];
  assign p3_array_index_1078781_comb = p2_literal_1076353[p3_array_index_1078765_comb];
  assign p3_array_index_1078782_comb = p2_literal_1076355[p3_array_index_1078766_comb];
  assign p3_array_index_1078783_comb = p2_arr[p3_addedKey__49_comb[79:72]];
  assign p3_array_index_1078785_comb = p2_arr[p3_addedKey__49_comb[63:56]];
  assign p3_res7__128_comb = p3_array_index_1078777_comb ^ p3_array_index_1078778_comb ^ p3_array_index_1078779_comb ^ p3_array_index_1078780_comb ^ p3_array_index_1078781_comb ^ p3_array_index_1078782_comb ^ p3_array_index_1078783_comb ^ p2_literal_1076358[p3_array_index_1078768_comb] ^ p3_array_index_1078785_comb ^ p2_literal_1076355[p3_array_index_1078770_comb] ^ p2_literal_1076353[p3_array_index_1078771_comb] ^ p2_literal_1076351[p3_array_index_1078772_comb] ^ p2_literal_1076349[p3_array_index_1078773_comb] ^ p2_literal_1076347[p3_array_index_1078774_comb] ^ p2_literal_1076345[p3_array_index_1078775_comb] ^ p2_arr[p3_addedKey__49_comb[7:0]];
  assign p3_array_index_1078794_comb = p2_literal_1076345[p3_res7__128_comb];
  assign p3_array_index_1078795_comb = p2_literal_1076347[p3_array_index_1078761_comb];
  assign p3_array_index_1078796_comb = p2_literal_1076349[p3_array_index_1078762_comb];
  assign p3_array_index_1078797_comb = p2_literal_1076351[p3_array_index_1078763_comb];
  assign p3_array_index_1078798_comb = p2_literal_1076353[p3_array_index_1078764_comb];
  assign p3_array_index_1078799_comb = p2_literal_1076355[p3_array_index_1078765_comb];
  assign p3_res7__129_comb = p3_array_index_1078794_comb ^ p3_array_index_1078795_comb ^ p3_array_index_1078796_comb ^ p3_array_index_1078797_comb ^ p3_array_index_1078798_comb ^ p3_array_index_1078799_comb ^ p3_array_index_1078766_comb ^ p2_literal_1076358[p3_array_index_1078783_comb] ^ p3_array_index_1078768_comb ^ p2_literal_1076355[p3_array_index_1078785_comb] ^ p2_literal_1076353[p3_array_index_1078770_comb] ^ p2_literal_1076351[p3_array_index_1078771_comb] ^ p2_literal_1076349[p3_array_index_1078772_comb] ^ p2_literal_1076347[p3_array_index_1078773_comb] ^ p2_literal_1076345[p3_array_index_1078774_comb] ^ p3_array_index_1078775_comb;
  assign p3_array_index_1078809_comb = p2_literal_1076347[p3_res7__128_comb];
  assign p3_array_index_1078810_comb = p2_literal_1076349[p3_array_index_1078761_comb];
  assign p3_array_index_1078811_comb = p2_literal_1076351[p3_array_index_1078762_comb];
  assign p3_array_index_1078812_comb = p2_literal_1076353[p3_array_index_1078763_comb];
  assign p3_array_index_1078813_comb = p2_literal_1076355[p3_array_index_1078764_comb];
  assign p3_res7__130_comb = p2_literal_1076345[p3_res7__129_comb] ^ p3_array_index_1078809_comb ^ p3_array_index_1078810_comb ^ p3_array_index_1078811_comb ^ p3_array_index_1078812_comb ^ p3_array_index_1078813_comb ^ p3_array_index_1078765_comb ^ p2_literal_1076358[p3_array_index_1078766_comb] ^ p3_array_index_1078783_comb ^ p2_literal_1076355[p3_array_index_1078768_comb] ^ p2_literal_1076353[p3_array_index_1078785_comb] ^ p2_literal_1076351[p3_array_index_1078770_comb] ^ p2_literal_1076349[p3_array_index_1078771_comb] ^ p2_literal_1076347[p3_array_index_1078772_comb] ^ p2_literal_1076345[p3_array_index_1078773_comb] ^ p3_array_index_1078774_comb;
  assign p3_array_index_1078823_comb = p2_literal_1076347[p3_res7__129_comb];
  assign p3_array_index_1078824_comb = p2_literal_1076349[p3_res7__128_comb];
  assign p3_array_index_1078825_comb = p2_literal_1076351[p3_array_index_1078761_comb];
  assign p3_array_index_1078826_comb = p2_literal_1076353[p3_array_index_1078762_comb];
  assign p3_array_index_1078827_comb = p2_literal_1076355[p3_array_index_1078763_comb];
  assign p3_res7__131_comb = p2_literal_1076345[p3_res7__130_comb] ^ p3_array_index_1078823_comb ^ p3_array_index_1078824_comb ^ p3_array_index_1078825_comb ^ p3_array_index_1078826_comb ^ p3_array_index_1078827_comb ^ p3_array_index_1078764_comb ^ p2_literal_1076358[p3_array_index_1078765_comb] ^ p3_array_index_1078766_comb ^ p2_literal_1076355[p3_array_index_1078783_comb] ^ p2_literal_1076353[p3_array_index_1078768_comb] ^ p2_literal_1076351[p3_array_index_1078785_comb] ^ p2_literal_1076349[p3_array_index_1078770_comb] ^ p2_literal_1076347[p3_array_index_1078771_comb] ^ p2_literal_1076345[p3_array_index_1078772_comb] ^ p3_array_index_1078773_comb;
  assign p3_array_index_1078838_comb = p2_literal_1076349[p3_res7__129_comb];
  assign p3_array_index_1078839_comb = p2_literal_1076351[p3_res7__128_comb];
  assign p3_array_index_1078840_comb = p2_literal_1076353[p3_array_index_1078761_comb];
  assign p3_array_index_1078841_comb = p2_literal_1076355[p3_array_index_1078762_comb];
  assign p3_res7__132_comb = p2_literal_1076345[p3_res7__131_comb] ^ p2_literal_1076347[p3_res7__130_comb] ^ p3_array_index_1078838_comb ^ p3_array_index_1078839_comb ^ p3_array_index_1078840_comb ^ p3_array_index_1078841_comb ^ p3_array_index_1078763_comb ^ p2_literal_1076358[p3_array_index_1078764_comb] ^ p3_array_index_1078765_comb ^ p3_array_index_1078782_comb ^ p2_literal_1076353[p3_array_index_1078783_comb] ^ p2_literal_1076351[p3_array_index_1078768_comb] ^ p2_literal_1076349[p3_array_index_1078785_comb] ^ p2_literal_1076347[p3_array_index_1078770_comb] ^ p2_literal_1076345[p3_array_index_1078771_comb] ^ p3_array_index_1078772_comb;
  assign p3_array_index_1078851_comb = p2_literal_1076349[p3_res7__130_comb];
  assign p3_array_index_1078852_comb = p2_literal_1076351[p3_res7__129_comb];
  assign p3_array_index_1078853_comb = p2_literal_1076353[p3_res7__128_comb];
  assign p3_array_index_1078854_comb = p2_literal_1076355[p3_array_index_1078761_comb];
  assign p3_res7__133_comb = p2_literal_1076345[p3_res7__132_comb] ^ p2_literal_1076347[p3_res7__131_comb] ^ p3_array_index_1078851_comb ^ p3_array_index_1078852_comb ^ p3_array_index_1078853_comb ^ p3_array_index_1078854_comb ^ p3_array_index_1078762_comb ^ p2_literal_1076358[p3_array_index_1078763_comb] ^ p3_array_index_1078764_comb ^ p3_array_index_1078799_comb ^ p2_literal_1076353[p3_array_index_1078766_comb] ^ p2_literal_1076351[p3_array_index_1078783_comb] ^ p2_literal_1076349[p3_array_index_1078768_comb] ^ p2_literal_1076347[p3_array_index_1078785_comb] ^ p2_literal_1076345[p3_array_index_1078770_comb] ^ p3_array_index_1078771_comb;
  assign p3_array_index_1078865_comb = p2_literal_1076351[p3_res7__130_comb];
  assign p3_array_index_1078866_comb = p2_literal_1076353[p3_res7__129_comb];
  assign p3_array_index_1078867_comb = p2_literal_1076355[p3_res7__128_comb];
  assign p3_res7__134_comb = p2_literal_1076345[p3_res7__133_comb] ^ p2_literal_1076347[p3_res7__132_comb] ^ p2_literal_1076349[p3_res7__131_comb] ^ p3_array_index_1078865_comb ^ p3_array_index_1078866_comb ^ p3_array_index_1078867_comb ^ p3_array_index_1078761_comb ^ p2_literal_1076358[p3_array_index_1078762_comb] ^ p3_array_index_1078763_comb ^ p3_array_index_1078813_comb ^ p3_array_index_1078781_comb ^ p2_literal_1076351[p3_array_index_1078766_comb] ^ p2_literal_1076349[p3_array_index_1078783_comb] ^ p2_literal_1076347[p3_array_index_1078768_comb] ^ p2_literal_1076345[p3_array_index_1078785_comb] ^ p3_array_index_1078770_comb;
  assign p3_array_index_1078877_comb = p2_literal_1076351[p3_res7__131_comb];
  assign p3_array_index_1078878_comb = p2_literal_1076353[p3_res7__130_comb];
  assign p3_array_index_1078879_comb = p2_literal_1076355[p3_res7__129_comb];
  assign p3_res7__135_comb = p2_literal_1076345[p3_res7__134_comb] ^ p2_literal_1076347[p3_res7__133_comb] ^ p2_literal_1076349[p3_res7__132_comb] ^ p3_array_index_1078877_comb ^ p3_array_index_1078878_comb ^ p3_array_index_1078879_comb ^ p3_res7__128_comb ^ p2_literal_1076358[p3_array_index_1078761_comb] ^ p3_array_index_1078762_comb ^ p3_array_index_1078827_comb ^ p3_array_index_1078798_comb ^ p2_literal_1076351[p3_array_index_1078765_comb] ^ p2_literal_1076349[p3_array_index_1078766_comb] ^ p2_literal_1076347[p3_array_index_1078783_comb] ^ p2_literal_1076345[p3_array_index_1078768_comb] ^ p3_array_index_1078785_comb;
  assign p3_array_index_1078890_comb = p2_literal_1076353[p3_res7__131_comb];
  assign p3_array_index_1078891_comb = p2_literal_1076355[p3_res7__130_comb];
  assign p3_res7__136_comb = p2_literal_1076345[p3_res7__135_comb] ^ p2_literal_1076347[p3_res7__134_comb] ^ p2_literal_1076349[p3_res7__133_comb] ^ p2_literal_1076351[p3_res7__132_comb] ^ p3_array_index_1078890_comb ^ p3_array_index_1078891_comb ^ p3_res7__129_comb ^ p2_literal_1076358[p3_res7__128_comb] ^ p3_array_index_1078761_comb ^ p3_array_index_1078841_comb ^ p3_array_index_1078812_comb ^ p3_array_index_1078780_comb ^ p2_literal_1076349[p3_array_index_1078765_comb] ^ p2_literal_1076347[p3_array_index_1078766_comb] ^ p2_literal_1076345[p3_array_index_1078783_comb] ^ p3_array_index_1078768_comb;
  assign p3_array_index_1078901_comb = p2_literal_1076353[p3_res7__132_comb];
  assign p3_array_index_1078902_comb = p2_literal_1076355[p3_res7__131_comb];
  assign p3_res7__137_comb = p2_literal_1076345[p3_res7__136_comb] ^ p2_literal_1076347[p3_res7__135_comb] ^ p2_literal_1076349[p3_res7__134_comb] ^ p2_literal_1076351[p3_res7__133_comb] ^ p3_array_index_1078901_comb ^ p3_array_index_1078902_comb ^ p3_res7__130_comb ^ p2_literal_1076358[p3_res7__129_comb] ^ p3_res7__128_comb ^ p3_array_index_1078854_comb ^ p3_array_index_1078826_comb ^ p3_array_index_1078797_comb ^ p2_literal_1076349[p3_array_index_1078764_comb] ^ p2_literal_1076347[p3_array_index_1078765_comb] ^ p2_literal_1076345[p3_array_index_1078766_comb] ^ p3_array_index_1078783_comb;
  assign p3_array_index_1078913_comb = p2_literal_1076355[p3_res7__132_comb];
  assign p3_res7__138_comb = p2_literal_1076345[p3_res7__137_comb] ^ p2_literal_1076347[p3_res7__136_comb] ^ p2_literal_1076349[p3_res7__135_comb] ^ p2_literal_1076351[p3_res7__134_comb] ^ p2_literal_1076353[p3_res7__133_comb] ^ p3_array_index_1078913_comb ^ p3_res7__131_comb ^ p2_literal_1076358[p3_res7__130_comb] ^ p3_res7__129_comb ^ p3_array_index_1078867_comb ^ p3_array_index_1078840_comb ^ p3_array_index_1078811_comb ^ p3_array_index_1078779_comb ^ p2_literal_1076347[p3_array_index_1078764_comb] ^ p2_literal_1076345[p3_array_index_1078765_comb] ^ p3_array_index_1078766_comb;
  assign p3_array_index_1078923_comb = p2_literal_1076355[p3_res7__133_comb];
  assign p3_res7__139_comb = p2_literal_1076345[p3_res7__138_comb] ^ p2_literal_1076347[p3_res7__137_comb] ^ p2_literal_1076349[p3_res7__136_comb] ^ p2_literal_1076351[p3_res7__135_comb] ^ p2_literal_1076353[p3_res7__134_comb] ^ p3_array_index_1078923_comb ^ p3_res7__132_comb ^ p2_literal_1076358[p3_res7__131_comb] ^ p3_res7__130_comb ^ p3_array_index_1078879_comb ^ p3_array_index_1078853_comb ^ p3_array_index_1078825_comb ^ p3_array_index_1078796_comb ^ p2_literal_1076347[p3_array_index_1078763_comb] ^ p2_literal_1076345[p3_array_index_1078764_comb] ^ p3_array_index_1078765_comb;
  assign p3_res7__140_comb = p2_literal_1076345[p3_res7__139_comb] ^ p2_literal_1076347[p3_res7__138_comb] ^ p2_literal_1076349[p3_res7__137_comb] ^ p2_literal_1076351[p3_res7__136_comb] ^ p2_literal_1076353[p3_res7__135_comb] ^ p2_literal_1076355[p3_res7__134_comb] ^ p3_res7__133_comb ^ p2_literal_1076358[p3_res7__132_comb] ^ p3_res7__131_comb ^ p3_array_index_1078891_comb ^ p3_array_index_1078866_comb ^ p3_array_index_1078839_comb ^ p3_array_index_1078810_comb ^ p3_array_index_1078778_comb ^ p2_literal_1076345[p3_array_index_1078763_comb] ^ p3_array_index_1078764_comb;
  assign p3_res7__141_comb = p2_literal_1076345[p3_res7__140_comb] ^ p2_literal_1076347[p3_res7__139_comb] ^ p2_literal_1076349[p3_res7__138_comb] ^ p2_literal_1076351[p3_res7__137_comb] ^ p2_literal_1076353[p3_res7__136_comb] ^ p2_literal_1076355[p3_res7__135_comb] ^ p3_res7__134_comb ^ p2_literal_1076358[p3_res7__133_comb] ^ p3_res7__132_comb ^ p3_array_index_1078902_comb ^ p3_array_index_1078878_comb ^ p3_array_index_1078852_comb ^ p3_array_index_1078824_comb ^ p3_array_index_1078795_comb ^ p2_literal_1076345[p3_array_index_1078762_comb] ^ p3_array_index_1078763_comb;
  assign p3_res7__142_comb = p2_literal_1076345[p3_res7__141_comb] ^ p2_literal_1076347[p3_res7__140_comb] ^ p2_literal_1076349[p3_res7__139_comb] ^ p2_literal_1076351[p3_res7__138_comb] ^ p2_literal_1076353[p3_res7__137_comb] ^ p2_literal_1076355[p3_res7__136_comb] ^ p3_res7__135_comb ^ p2_literal_1076358[p3_res7__134_comb] ^ p3_res7__133_comb ^ p3_array_index_1078913_comb ^ p3_array_index_1078890_comb ^ p3_array_index_1078865_comb ^ p3_array_index_1078838_comb ^ p3_array_index_1078809_comb ^ p3_array_index_1078777_comb ^ p3_array_index_1078762_comb;
  assign p3_res7__143_comb = p2_literal_1076345[p3_res7__142_comb] ^ p2_literal_1076347[p3_res7__141_comb] ^ p2_literal_1076349[p3_res7__140_comb] ^ p2_literal_1076351[p3_res7__139_comb] ^ p2_literal_1076353[p3_res7__138_comb] ^ p2_literal_1076355[p3_res7__137_comb] ^ p3_res7__136_comb ^ p2_literal_1076358[p3_res7__135_comb] ^ p3_res7__134_comb ^ p3_array_index_1078923_comb ^ p3_array_index_1078901_comb ^ p3_array_index_1078877_comb ^ p3_array_index_1078851_comb ^ p3_array_index_1078823_comb ^ p3_array_index_1078794_comb ^ p3_array_index_1078761_comb;
  assign p3_res__8_comb = {p3_res7__143_comb, p3_res7__142_comb, p3_res7__141_comb, p3_res7__140_comb, p3_res7__139_comb, p3_res7__138_comb, p3_res7__137_comb, p3_res7__136_comb, p3_res7__135_comb, p3_res7__134_comb, p3_res7__133_comb, p3_res7__132_comb, p3_res7__131_comb, p3_res7__130_comb, p3_res7__129_comb, p3_res7__128_comb};
  assign p3_xor_1078963_comb = p3_res__8_comb ^ p2_k3;
  assign p3_addedKey__50_comb = p3_xor_1078963_comb ^ 128'h2ade_daf2_3e95_a23a_17b5_18a0_5e61_c10a;
  assign p3_array_index_1078979_comb = p2_arr[p3_addedKey__50_comb[127:120]];
  assign p3_array_index_1078980_comb = p2_arr[p3_addedKey__50_comb[119:112]];
  assign p3_array_index_1078981_comb = p2_arr[p3_addedKey__50_comb[111:104]];
  assign p3_array_index_1078982_comb = p2_arr[p3_addedKey__50_comb[103:96]];
  assign p3_array_index_1078983_comb = p2_arr[p3_addedKey__50_comb[95:88]];
  assign p3_array_index_1078984_comb = p2_arr[p3_addedKey__50_comb[87:80]];
  assign p3_array_index_1078986_comb = p2_arr[p3_addedKey__50_comb[71:64]];
  assign p3_array_index_1078988_comb = p2_arr[p3_addedKey__50_comb[55:48]];
  assign p3_array_index_1078989_comb = p2_arr[p3_addedKey__50_comb[47:40]];
  assign p3_array_index_1078990_comb = p2_arr[p3_addedKey__50_comb[39:32]];
  assign p3_array_index_1078991_comb = p2_arr[p3_addedKey__50_comb[31:24]];
  assign p3_array_index_1078992_comb = p2_arr[p3_addedKey__50_comb[23:16]];
  assign p3_array_index_1078993_comb = p2_arr[p3_addedKey__50_comb[15:8]];
  assign p3_addedKey__34_comb = p3_k2_comb ^ p2_res__33;
  assign p3_array_index_1078995_comb = p2_literal_1076345[p3_array_index_1078979_comb];
  assign p3_array_index_1078996_comb = p2_literal_1076347[p3_array_index_1078980_comb];
  assign p3_array_index_1078997_comb = p2_literal_1076349[p3_array_index_1078981_comb];
  assign p3_array_index_1078998_comb = p2_literal_1076351[p3_array_index_1078982_comb];
  assign p3_array_index_1078999_comb = p2_literal_1076353[p3_array_index_1078983_comb];
  assign p3_array_index_1079000_comb = p2_literal_1076355[p3_array_index_1078984_comb];
  assign p3_array_index_1079001_comb = p2_arr[p3_addedKey__50_comb[79:72]];
  assign p3_array_index_1079003_comb = p2_arr[p3_addedKey__50_comb[63:56]];
  assign p3_res7__144_comb = p3_array_index_1078995_comb ^ p3_array_index_1078996_comb ^ p3_array_index_1078997_comb ^ p3_array_index_1078998_comb ^ p3_array_index_1078999_comb ^ p3_array_index_1079000_comb ^ p3_array_index_1079001_comb ^ p2_literal_1076358[p3_array_index_1078986_comb] ^ p3_array_index_1079003_comb ^ p2_literal_1076355[p3_array_index_1078988_comb] ^ p2_literal_1076353[p3_array_index_1078989_comb] ^ p2_literal_1076351[p3_array_index_1078990_comb] ^ p2_literal_1076349[p3_array_index_1078991_comb] ^ p2_literal_1076347[p3_array_index_1078992_comb] ^ p2_literal_1076345[p3_array_index_1078993_comb] ^ p2_arr[p3_addedKey__50_comb[7:0]];
  assign p3_array_index_1079414_comb = p2_arr[p3_addedKey__34_comb[127:120]];
  assign p3_array_index_1079415_comb = p2_arr[p3_addedKey__34_comb[119:112]];
  assign p3_array_index_1079416_comb = p2_arr[p3_addedKey__34_comb[111:104]];
  assign p3_array_index_1079417_comb = p2_arr[p3_addedKey__34_comb[103:96]];
  assign p3_array_index_1079418_comb = p2_arr[p3_addedKey__34_comb[95:88]];
  assign p3_array_index_1079419_comb = p2_arr[p3_addedKey__34_comb[87:80]];
  assign p3_array_index_1079421_comb = p2_arr[p3_addedKey__34_comb[71:64]];
  assign p3_array_index_1079423_comb = p2_arr[p3_addedKey__34_comb[55:48]];
  assign p3_array_index_1079424_comb = p2_arr[p3_addedKey__34_comb[47:40]];
  assign p3_array_index_1079425_comb = p2_arr[p3_addedKey__34_comb[39:32]];
  assign p3_array_index_1079426_comb = p2_arr[p3_addedKey__34_comb[31:24]];
  assign p3_array_index_1079427_comb = p2_arr[p3_addedKey__34_comb[23:16]];
  assign p3_array_index_1079428_comb = p2_arr[p3_addedKey__34_comb[15:8]];
  assign p3_array_index_1079012_comb = p2_literal_1076345[p3_res7__144_comb];
  assign p3_array_index_1079013_comb = p2_literal_1076347[p3_array_index_1078979_comb];
  assign p3_array_index_1079014_comb = p2_literal_1076349[p3_array_index_1078980_comb];
  assign p3_array_index_1079015_comb = p2_literal_1076351[p3_array_index_1078981_comb];
  assign p3_array_index_1079016_comb = p2_literal_1076353[p3_array_index_1078982_comb];
  assign p3_array_index_1079017_comb = p2_literal_1076355[p3_array_index_1078983_comb];
  assign p3_array_index_1079430_comb = p2_literal_1076345[p3_array_index_1079414_comb];
  assign p3_array_index_1079431_comb = p2_literal_1076347[p3_array_index_1079415_comb];
  assign p3_array_index_1079432_comb = p2_literal_1076349[p3_array_index_1079416_comb];
  assign p3_array_index_1079433_comb = p2_literal_1076351[p3_array_index_1079417_comb];
  assign p3_array_index_1079434_comb = p2_literal_1076353[p3_array_index_1079418_comb];
  assign p3_array_index_1079435_comb = p2_literal_1076355[p3_array_index_1079419_comb];
  assign p3_array_index_1079436_comb = p2_arr[p3_addedKey__34_comb[79:72]];
  assign p3_array_index_1079438_comb = p2_arr[p3_addedKey__34_comb[63:56]];
  assign p3_res7__145_comb = p3_array_index_1079012_comb ^ p3_array_index_1079013_comb ^ p3_array_index_1079014_comb ^ p3_array_index_1079015_comb ^ p3_array_index_1079016_comb ^ p3_array_index_1079017_comb ^ p3_array_index_1078984_comb ^ p2_literal_1076358[p3_array_index_1079001_comb] ^ p3_array_index_1078986_comb ^ p2_literal_1076355[p3_array_index_1079003_comb] ^ p2_literal_1076353[p3_array_index_1078988_comb] ^ p2_literal_1076351[p3_array_index_1078989_comb] ^ p2_literal_1076349[p3_array_index_1078990_comb] ^ p2_literal_1076347[p3_array_index_1078991_comb] ^ p2_literal_1076345[p3_array_index_1078992_comb] ^ p3_array_index_1078993_comb;
  assign p3_res7__544_comb = p3_array_index_1079430_comb ^ p3_array_index_1079431_comb ^ p3_array_index_1079432_comb ^ p3_array_index_1079433_comb ^ p3_array_index_1079434_comb ^ p3_array_index_1079435_comb ^ p3_array_index_1079436_comb ^ p2_literal_1076358[p3_array_index_1079421_comb] ^ p3_array_index_1079438_comb ^ p2_literal_1076355[p3_array_index_1079423_comb] ^ p2_literal_1076353[p3_array_index_1079424_comb] ^ p2_literal_1076351[p3_array_index_1079425_comb] ^ p2_literal_1076349[p3_array_index_1079426_comb] ^ p2_literal_1076347[p3_array_index_1079427_comb] ^ p2_literal_1076345[p3_array_index_1079428_comb] ^ p2_arr[p3_addedKey__34_comb[7:0]];
  assign p3_array_index_1079027_comb = p2_literal_1076347[p3_res7__144_comb];
  assign p3_array_index_1079028_comb = p2_literal_1076349[p3_array_index_1078979_comb];
  assign p3_array_index_1079029_comb = p2_literal_1076351[p3_array_index_1078980_comb];
  assign p3_array_index_1079030_comb = p2_literal_1076353[p3_array_index_1078981_comb];
  assign p3_array_index_1079031_comb = p2_literal_1076355[p3_array_index_1078982_comb];
  assign p3_array_index_1079447_comb = p2_literal_1076345[p3_res7__544_comb];
  assign p3_array_index_1079448_comb = p2_literal_1076347[p3_array_index_1079414_comb];
  assign p3_array_index_1079449_comb = p2_literal_1076349[p3_array_index_1079415_comb];
  assign p3_array_index_1079450_comb = p2_literal_1076351[p3_array_index_1079416_comb];
  assign p3_array_index_1079451_comb = p2_literal_1076353[p3_array_index_1079417_comb];
  assign p3_array_index_1079452_comb = p2_literal_1076355[p3_array_index_1079418_comb];
  assign p3_res7__146_comb = p2_literal_1076345[p3_res7__145_comb] ^ p3_array_index_1079027_comb ^ p3_array_index_1079028_comb ^ p3_array_index_1079029_comb ^ p3_array_index_1079030_comb ^ p3_array_index_1079031_comb ^ p3_array_index_1078983_comb ^ p2_literal_1076358[p3_array_index_1078984_comb] ^ p3_array_index_1079001_comb ^ p2_literal_1076355[p3_array_index_1078986_comb] ^ p2_literal_1076353[p3_array_index_1079003_comb] ^ p2_literal_1076351[p3_array_index_1078988_comb] ^ p2_literal_1076349[p3_array_index_1078989_comb] ^ p2_literal_1076347[p3_array_index_1078990_comb] ^ p2_literal_1076345[p3_array_index_1078991_comb] ^ p3_array_index_1078992_comb;
  assign p3_res7__545_comb = p3_array_index_1079447_comb ^ p3_array_index_1079448_comb ^ p3_array_index_1079449_comb ^ p3_array_index_1079450_comb ^ p3_array_index_1079451_comb ^ p3_array_index_1079452_comb ^ p3_array_index_1079419_comb ^ p2_literal_1076358[p3_array_index_1079436_comb] ^ p3_array_index_1079421_comb ^ p2_literal_1076355[p3_array_index_1079438_comb] ^ p2_literal_1076353[p3_array_index_1079423_comb] ^ p2_literal_1076351[p3_array_index_1079424_comb] ^ p2_literal_1076349[p3_array_index_1079425_comb] ^ p2_literal_1076347[p3_array_index_1079426_comb] ^ p2_literal_1076345[p3_array_index_1079427_comb] ^ p3_array_index_1079428_comb;
  assign p3_array_index_1079041_comb = p2_literal_1076347[p3_res7__145_comb];
  assign p3_array_index_1079042_comb = p2_literal_1076349[p3_res7__144_comb];
  assign p3_array_index_1079043_comb = p2_literal_1076351[p3_array_index_1078979_comb];
  assign p3_array_index_1079044_comb = p2_literal_1076353[p3_array_index_1078980_comb];
  assign p3_array_index_1079045_comb = p2_literal_1076355[p3_array_index_1078981_comb];
  assign p3_array_index_1079462_comb = p2_literal_1076347[p3_res7__544_comb];
  assign p3_array_index_1079463_comb = p2_literal_1076349[p3_array_index_1079414_comb];
  assign p3_array_index_1079464_comb = p2_literal_1076351[p3_array_index_1079415_comb];
  assign p3_array_index_1079465_comb = p2_literal_1076353[p3_array_index_1079416_comb];
  assign p3_array_index_1079466_comb = p2_literal_1076355[p3_array_index_1079417_comb];
  assign p3_res7__147_comb = p2_literal_1076345[p3_res7__146_comb] ^ p3_array_index_1079041_comb ^ p3_array_index_1079042_comb ^ p3_array_index_1079043_comb ^ p3_array_index_1079044_comb ^ p3_array_index_1079045_comb ^ p3_array_index_1078982_comb ^ p2_literal_1076358[p3_array_index_1078983_comb] ^ p3_array_index_1078984_comb ^ p2_literal_1076355[p3_array_index_1079001_comb] ^ p2_literal_1076353[p3_array_index_1078986_comb] ^ p2_literal_1076351[p3_array_index_1079003_comb] ^ p2_literal_1076349[p3_array_index_1078988_comb] ^ p2_literal_1076347[p3_array_index_1078989_comb] ^ p2_literal_1076345[p3_array_index_1078990_comb] ^ p3_array_index_1078991_comb;
  assign p3_res7__546_comb = p2_literal_1076345[p3_res7__545_comb] ^ p3_array_index_1079462_comb ^ p3_array_index_1079463_comb ^ p3_array_index_1079464_comb ^ p3_array_index_1079465_comb ^ p3_array_index_1079466_comb ^ p3_array_index_1079418_comb ^ p2_literal_1076358[p3_array_index_1079419_comb] ^ p3_array_index_1079436_comb ^ p2_literal_1076355[p3_array_index_1079421_comb] ^ p2_literal_1076353[p3_array_index_1079438_comb] ^ p2_literal_1076351[p3_array_index_1079423_comb] ^ p2_literal_1076349[p3_array_index_1079424_comb] ^ p2_literal_1076347[p3_array_index_1079425_comb] ^ p2_literal_1076345[p3_array_index_1079426_comb] ^ p3_array_index_1079427_comb;
  assign p3_array_index_1079056_comb = p2_literal_1076349[p3_res7__145_comb];
  assign p3_array_index_1079057_comb = p2_literal_1076351[p3_res7__144_comb];
  assign p3_array_index_1079058_comb = p2_literal_1076353[p3_array_index_1078979_comb];
  assign p3_array_index_1079059_comb = p2_literal_1076355[p3_array_index_1078980_comb];
  assign p3_array_index_1079476_comb = p2_literal_1076347[p3_res7__545_comb];
  assign p3_array_index_1079477_comb = p2_literal_1076349[p3_res7__544_comb];
  assign p3_array_index_1079478_comb = p2_literal_1076351[p3_array_index_1079414_comb];
  assign p3_array_index_1079479_comb = p2_literal_1076353[p3_array_index_1079415_comb];
  assign p3_array_index_1079480_comb = p2_literal_1076355[p3_array_index_1079416_comb];
  assign p3_res7__148_comb = p2_literal_1076345[p3_res7__147_comb] ^ p2_literal_1076347[p3_res7__146_comb] ^ p3_array_index_1079056_comb ^ p3_array_index_1079057_comb ^ p3_array_index_1079058_comb ^ p3_array_index_1079059_comb ^ p3_array_index_1078981_comb ^ p2_literal_1076358[p3_array_index_1078982_comb] ^ p3_array_index_1078983_comb ^ p3_array_index_1079000_comb ^ p2_literal_1076353[p3_array_index_1079001_comb] ^ p2_literal_1076351[p3_array_index_1078986_comb] ^ p2_literal_1076349[p3_array_index_1079003_comb] ^ p2_literal_1076347[p3_array_index_1078988_comb] ^ p2_literal_1076345[p3_array_index_1078989_comb] ^ p3_array_index_1078990_comb;
  assign p3_res7__547_comb = p2_literal_1076345[p3_res7__546_comb] ^ p3_array_index_1079476_comb ^ p3_array_index_1079477_comb ^ p3_array_index_1079478_comb ^ p3_array_index_1079479_comb ^ p3_array_index_1079480_comb ^ p3_array_index_1079417_comb ^ p2_literal_1076358[p3_array_index_1079418_comb] ^ p3_array_index_1079419_comb ^ p2_literal_1076355[p3_array_index_1079436_comb] ^ p2_literal_1076353[p3_array_index_1079421_comb] ^ p2_literal_1076351[p3_array_index_1079438_comb] ^ p2_literal_1076349[p3_array_index_1079423_comb] ^ p2_literal_1076347[p3_array_index_1079424_comb] ^ p2_literal_1076345[p3_array_index_1079425_comb] ^ p3_array_index_1079426_comb;
  assign p3_array_index_1079069_comb = p2_literal_1076349[p3_res7__146_comb];
  assign p3_array_index_1079070_comb = p2_literal_1076351[p3_res7__145_comb];
  assign p3_array_index_1079071_comb = p2_literal_1076353[p3_res7__144_comb];
  assign p3_array_index_1079072_comb = p2_literal_1076355[p3_array_index_1078979_comb];
  assign p3_array_index_1079491_comb = p2_literal_1076349[p3_res7__545_comb];
  assign p3_array_index_1079492_comb = p2_literal_1076351[p3_res7__544_comb];
  assign p3_array_index_1079493_comb = p2_literal_1076353[p3_array_index_1079414_comb];
  assign p3_array_index_1079494_comb = p2_literal_1076355[p3_array_index_1079415_comb];
  assign p3_res7__149_comb = p2_literal_1076345[p3_res7__148_comb] ^ p2_literal_1076347[p3_res7__147_comb] ^ p3_array_index_1079069_comb ^ p3_array_index_1079070_comb ^ p3_array_index_1079071_comb ^ p3_array_index_1079072_comb ^ p3_array_index_1078980_comb ^ p2_literal_1076358[p3_array_index_1078981_comb] ^ p3_array_index_1078982_comb ^ p3_array_index_1079017_comb ^ p2_literal_1076353[p3_array_index_1078984_comb] ^ p2_literal_1076351[p3_array_index_1079001_comb] ^ p2_literal_1076349[p3_array_index_1078986_comb] ^ p2_literal_1076347[p3_array_index_1079003_comb] ^ p2_literal_1076345[p3_array_index_1078988_comb] ^ p3_array_index_1078989_comb;
  assign p3_res7__548_comb = p2_literal_1076345[p3_res7__547_comb] ^ p2_literal_1076347[p3_res7__546_comb] ^ p3_array_index_1079491_comb ^ p3_array_index_1079492_comb ^ p3_array_index_1079493_comb ^ p3_array_index_1079494_comb ^ p3_array_index_1079416_comb ^ p2_literal_1076358[p3_array_index_1079417_comb] ^ p3_array_index_1079418_comb ^ p3_array_index_1079435_comb ^ p2_literal_1076353[p3_array_index_1079436_comb] ^ p2_literal_1076351[p3_array_index_1079421_comb] ^ p2_literal_1076349[p3_array_index_1079438_comb] ^ p2_literal_1076347[p3_array_index_1079423_comb] ^ p2_literal_1076345[p3_array_index_1079424_comb] ^ p3_array_index_1079425_comb;
  assign p3_array_index_1079083_comb = p2_literal_1076351[p3_res7__146_comb];
  assign p3_array_index_1079084_comb = p2_literal_1076353[p3_res7__145_comb];
  assign p3_array_index_1079085_comb = p2_literal_1076355[p3_res7__144_comb];
  assign p3_array_index_1079504_comb = p2_literal_1076349[p3_res7__546_comb];
  assign p3_array_index_1079505_comb = p2_literal_1076351[p3_res7__545_comb];
  assign p3_array_index_1079506_comb = p2_literal_1076353[p3_res7__544_comb];
  assign p3_array_index_1079507_comb = p2_literal_1076355[p3_array_index_1079414_comb];
  assign p3_res7__150_comb = p2_literal_1076345[p3_res7__149_comb] ^ p2_literal_1076347[p3_res7__148_comb] ^ p2_literal_1076349[p3_res7__147_comb] ^ p3_array_index_1079083_comb ^ p3_array_index_1079084_comb ^ p3_array_index_1079085_comb ^ p3_array_index_1078979_comb ^ p2_literal_1076358[p3_array_index_1078980_comb] ^ p3_array_index_1078981_comb ^ p3_array_index_1079031_comb ^ p3_array_index_1078999_comb ^ p2_literal_1076351[p3_array_index_1078984_comb] ^ p2_literal_1076349[p3_array_index_1079001_comb] ^ p2_literal_1076347[p3_array_index_1078986_comb] ^ p2_literal_1076345[p3_array_index_1079003_comb] ^ p3_array_index_1078988_comb;
  assign p3_res7__549_comb = p2_literal_1076345[p3_res7__548_comb] ^ p2_literal_1076347[p3_res7__547_comb] ^ p3_array_index_1079504_comb ^ p3_array_index_1079505_comb ^ p3_array_index_1079506_comb ^ p3_array_index_1079507_comb ^ p3_array_index_1079415_comb ^ p2_literal_1076358[p3_array_index_1079416_comb] ^ p3_array_index_1079417_comb ^ p3_array_index_1079452_comb ^ p2_literal_1076353[p3_array_index_1079419_comb] ^ p2_literal_1076351[p3_array_index_1079436_comb] ^ p2_literal_1076349[p3_array_index_1079421_comb] ^ p2_literal_1076347[p3_array_index_1079438_comb] ^ p2_literal_1076345[p3_array_index_1079423_comb] ^ p3_array_index_1079424_comb;
  assign p3_array_index_1079095_comb = p2_literal_1076351[p3_res7__147_comb];
  assign p3_array_index_1079096_comb = p2_literal_1076353[p3_res7__146_comb];
  assign p3_array_index_1079097_comb = p2_literal_1076355[p3_res7__145_comb];
  assign p3_array_index_1079518_comb = p2_literal_1076351[p3_res7__546_comb];
  assign p3_array_index_1079519_comb = p2_literal_1076353[p3_res7__545_comb];
  assign p3_array_index_1079520_comb = p2_literal_1076355[p3_res7__544_comb];
  assign p3_res7__151_comb = p2_literal_1076345[p3_res7__150_comb] ^ p2_literal_1076347[p3_res7__149_comb] ^ p2_literal_1076349[p3_res7__148_comb] ^ p3_array_index_1079095_comb ^ p3_array_index_1079096_comb ^ p3_array_index_1079097_comb ^ p3_res7__144_comb ^ p2_literal_1076358[p3_array_index_1078979_comb] ^ p3_array_index_1078980_comb ^ p3_array_index_1079045_comb ^ p3_array_index_1079016_comb ^ p2_literal_1076351[p3_array_index_1078983_comb] ^ p2_literal_1076349[p3_array_index_1078984_comb] ^ p2_literal_1076347[p3_array_index_1079001_comb] ^ p2_literal_1076345[p3_array_index_1078986_comb] ^ p3_array_index_1079003_comb;
  assign p3_res7__550_comb = p2_literal_1076345[p3_res7__549_comb] ^ p2_literal_1076347[p3_res7__548_comb] ^ p2_literal_1076349[p3_res7__547_comb] ^ p3_array_index_1079518_comb ^ p3_array_index_1079519_comb ^ p3_array_index_1079520_comb ^ p3_array_index_1079414_comb ^ p2_literal_1076358[p3_array_index_1079415_comb] ^ p3_array_index_1079416_comb ^ p3_array_index_1079466_comb ^ p3_array_index_1079434_comb ^ p2_literal_1076351[p3_array_index_1079419_comb] ^ p2_literal_1076349[p3_array_index_1079436_comb] ^ p2_literal_1076347[p3_array_index_1079421_comb] ^ p2_literal_1076345[p3_array_index_1079438_comb] ^ p3_array_index_1079423_comb;
  assign p3_array_index_1079108_comb = p2_literal_1076353[p3_res7__147_comb];
  assign p3_array_index_1079109_comb = p2_literal_1076355[p3_res7__146_comb];
  assign p3_array_index_1079530_comb = p2_literal_1076351[p3_res7__547_comb];
  assign p3_array_index_1079531_comb = p2_literal_1076353[p3_res7__546_comb];
  assign p3_array_index_1079532_comb = p2_literal_1076355[p3_res7__545_comb];
  assign p3_res7__152_comb = p2_literal_1076345[p3_res7__151_comb] ^ p2_literal_1076347[p3_res7__150_comb] ^ p2_literal_1076349[p3_res7__149_comb] ^ p2_literal_1076351[p3_res7__148_comb] ^ p3_array_index_1079108_comb ^ p3_array_index_1079109_comb ^ p3_res7__145_comb ^ p2_literal_1076358[p3_res7__144_comb] ^ p3_array_index_1078979_comb ^ p3_array_index_1079059_comb ^ p3_array_index_1079030_comb ^ p3_array_index_1078998_comb ^ p2_literal_1076349[p3_array_index_1078983_comb] ^ p2_literal_1076347[p3_array_index_1078984_comb] ^ p2_literal_1076345[p3_array_index_1079001_comb] ^ p3_array_index_1078986_comb;
  assign p3_res7__551_comb = p2_literal_1076345[p3_res7__550_comb] ^ p2_literal_1076347[p3_res7__549_comb] ^ p2_literal_1076349[p3_res7__548_comb] ^ p3_array_index_1079530_comb ^ p3_array_index_1079531_comb ^ p3_array_index_1079532_comb ^ p3_res7__544_comb ^ p2_literal_1076358[p3_array_index_1079414_comb] ^ p3_array_index_1079415_comb ^ p3_array_index_1079480_comb ^ p3_array_index_1079451_comb ^ p2_literal_1076351[p3_array_index_1079418_comb] ^ p2_literal_1076349[p3_array_index_1079419_comb] ^ p2_literal_1076347[p3_array_index_1079436_comb] ^ p2_literal_1076345[p3_array_index_1079421_comb] ^ p3_array_index_1079438_comb;
  assign p3_array_index_1079119_comb = p2_literal_1076353[p3_res7__148_comb];
  assign p3_array_index_1079120_comb = p2_literal_1076355[p3_res7__147_comb];
  assign p3_array_index_1079543_comb = p2_literal_1076353[p3_res7__547_comb];
  assign p3_array_index_1079544_comb = p2_literal_1076355[p3_res7__546_comb];
  assign p3_res7__153_comb = p2_literal_1076345[p3_res7__152_comb] ^ p2_literal_1076347[p3_res7__151_comb] ^ p2_literal_1076349[p3_res7__150_comb] ^ p2_literal_1076351[p3_res7__149_comb] ^ p3_array_index_1079119_comb ^ p3_array_index_1079120_comb ^ p3_res7__146_comb ^ p2_literal_1076358[p3_res7__145_comb] ^ p3_res7__144_comb ^ p3_array_index_1079072_comb ^ p3_array_index_1079044_comb ^ p3_array_index_1079015_comb ^ p2_literal_1076349[p3_array_index_1078982_comb] ^ p2_literal_1076347[p3_array_index_1078983_comb] ^ p2_literal_1076345[p3_array_index_1078984_comb] ^ p3_array_index_1079001_comb;
  assign p3_res7__552_comb = p2_literal_1076345[p3_res7__551_comb] ^ p2_literal_1076347[p3_res7__550_comb] ^ p2_literal_1076349[p3_res7__549_comb] ^ p2_literal_1076351[p3_res7__548_comb] ^ p3_array_index_1079543_comb ^ p3_array_index_1079544_comb ^ p3_res7__545_comb ^ p2_literal_1076358[p3_res7__544_comb] ^ p3_array_index_1079414_comb ^ p3_array_index_1079494_comb ^ p3_array_index_1079465_comb ^ p3_array_index_1079433_comb ^ p2_literal_1076349[p3_array_index_1079418_comb] ^ p2_literal_1076347[p3_array_index_1079419_comb] ^ p2_literal_1076345[p3_array_index_1079436_comb] ^ p3_array_index_1079421_comb;
  assign p3_array_index_1079131_comb = p2_literal_1076355[p3_res7__148_comb];
  assign p3_array_index_1079554_comb = p2_literal_1076353[p3_res7__548_comb];
  assign p3_array_index_1079555_comb = p2_literal_1076355[p3_res7__547_comb];
  assign p3_res7__154_comb = p2_literal_1076345[p3_res7__153_comb] ^ p2_literal_1076347[p3_res7__152_comb] ^ p2_literal_1076349[p3_res7__151_comb] ^ p2_literal_1076351[p3_res7__150_comb] ^ p2_literal_1076353[p3_res7__149_comb] ^ p3_array_index_1079131_comb ^ p3_res7__147_comb ^ p2_literal_1076358[p3_res7__146_comb] ^ p3_res7__145_comb ^ p3_array_index_1079085_comb ^ p3_array_index_1079058_comb ^ p3_array_index_1079029_comb ^ p3_array_index_1078997_comb ^ p2_literal_1076347[p3_array_index_1078982_comb] ^ p2_literal_1076345[p3_array_index_1078983_comb] ^ p3_array_index_1078984_comb;
  assign p3_res7__553_comb = p2_literal_1076345[p3_res7__552_comb] ^ p2_literal_1076347[p3_res7__551_comb] ^ p2_literal_1076349[p3_res7__550_comb] ^ p2_literal_1076351[p3_res7__549_comb] ^ p3_array_index_1079554_comb ^ p3_array_index_1079555_comb ^ p3_res7__546_comb ^ p2_literal_1076358[p3_res7__545_comb] ^ p3_res7__544_comb ^ p3_array_index_1079507_comb ^ p3_array_index_1079479_comb ^ p3_array_index_1079450_comb ^ p2_literal_1076349[p3_array_index_1079417_comb] ^ p2_literal_1076347[p3_array_index_1079418_comb] ^ p2_literal_1076345[p3_array_index_1079419_comb] ^ p3_array_index_1079436_comb;
  assign p3_array_index_1079141_comb = p2_literal_1076355[p3_res7__149_comb];
  assign p3_array_index_1079566_comb = p2_literal_1076355[p3_res7__548_comb];
  assign p3_res7__155_comb = p2_literal_1076345[p3_res7__154_comb] ^ p2_literal_1076347[p3_res7__153_comb] ^ p2_literal_1076349[p3_res7__152_comb] ^ p2_literal_1076351[p3_res7__151_comb] ^ p2_literal_1076353[p3_res7__150_comb] ^ p3_array_index_1079141_comb ^ p3_res7__148_comb ^ p2_literal_1076358[p3_res7__147_comb] ^ p3_res7__146_comb ^ p3_array_index_1079097_comb ^ p3_array_index_1079071_comb ^ p3_array_index_1079043_comb ^ p3_array_index_1079014_comb ^ p2_literal_1076347[p3_array_index_1078981_comb] ^ p2_literal_1076345[p3_array_index_1078982_comb] ^ p3_array_index_1078983_comb;
  assign p3_res7__554_comb = p2_literal_1076345[p3_res7__553_comb] ^ p2_literal_1076347[p3_res7__552_comb] ^ p2_literal_1076349[p3_res7__551_comb] ^ p2_literal_1076351[p3_res7__550_comb] ^ p2_literal_1076353[p3_res7__549_comb] ^ p3_array_index_1079566_comb ^ p3_res7__547_comb ^ p2_literal_1076358[p3_res7__546_comb] ^ p3_res7__545_comb ^ p3_array_index_1079520_comb ^ p3_array_index_1079493_comb ^ p3_array_index_1079464_comb ^ p3_array_index_1079432_comb ^ p2_literal_1076347[p3_array_index_1079417_comb] ^ p2_literal_1076345[p3_array_index_1079418_comb] ^ p3_array_index_1079419_comb;
  assign p3_array_index_1079576_comb = p2_literal_1076355[p3_res7__549_comb];
  assign p3_res7__156_comb = p2_literal_1076345[p3_res7__155_comb] ^ p2_literal_1076347[p3_res7__154_comb] ^ p2_literal_1076349[p3_res7__153_comb] ^ p2_literal_1076351[p3_res7__152_comb] ^ p2_literal_1076353[p3_res7__151_comb] ^ p2_literal_1076355[p3_res7__150_comb] ^ p3_res7__149_comb ^ p2_literal_1076358[p3_res7__148_comb] ^ p3_res7__147_comb ^ p3_array_index_1079109_comb ^ p3_array_index_1079084_comb ^ p3_array_index_1079057_comb ^ p3_array_index_1079028_comb ^ p3_array_index_1078996_comb ^ p2_literal_1076345[p3_array_index_1078981_comb] ^ p3_array_index_1078982_comb;
  assign p3_res7__555_comb = p2_literal_1076345[p3_res7__554_comb] ^ p2_literal_1076347[p3_res7__553_comb] ^ p2_literal_1076349[p3_res7__552_comb] ^ p2_literal_1076351[p3_res7__551_comb] ^ p2_literal_1076353[p3_res7__550_comb] ^ p3_array_index_1079576_comb ^ p3_res7__548_comb ^ p2_literal_1076358[p3_res7__547_comb] ^ p3_res7__546_comb ^ p3_array_index_1079532_comb ^ p3_array_index_1079506_comb ^ p3_array_index_1079478_comb ^ p3_array_index_1079449_comb ^ p2_literal_1076347[p3_array_index_1079416_comb] ^ p2_literal_1076345[p3_array_index_1079417_comb] ^ p3_array_index_1079418_comb;
  assign p3_res7__157_comb = p2_literal_1076345[p3_res7__156_comb] ^ p2_literal_1076347[p3_res7__155_comb] ^ p2_literal_1076349[p3_res7__154_comb] ^ p2_literal_1076351[p3_res7__153_comb] ^ p2_literal_1076353[p3_res7__152_comb] ^ p2_literal_1076355[p3_res7__151_comb] ^ p3_res7__150_comb ^ p2_literal_1076358[p3_res7__149_comb] ^ p3_res7__148_comb ^ p3_array_index_1079120_comb ^ p3_array_index_1079096_comb ^ p3_array_index_1079070_comb ^ p3_array_index_1079042_comb ^ p3_array_index_1079013_comb ^ p2_literal_1076345[p3_array_index_1078980_comb] ^ p3_array_index_1078981_comb;
  assign p3_res7__556_comb = p2_literal_1076345[p3_res7__555_comb] ^ p2_literal_1076347[p3_res7__554_comb] ^ p2_literal_1076349[p3_res7__553_comb] ^ p2_literal_1076351[p3_res7__552_comb] ^ p2_literal_1076353[p3_res7__551_comb] ^ p2_literal_1076355[p3_res7__550_comb] ^ p3_res7__549_comb ^ p2_literal_1076358[p3_res7__548_comb] ^ p3_res7__547_comb ^ p3_array_index_1079544_comb ^ p3_array_index_1079519_comb ^ p3_array_index_1079492_comb ^ p3_array_index_1079463_comb ^ p3_array_index_1079431_comb ^ p2_literal_1076345[p3_array_index_1079416_comb] ^ p3_array_index_1079417_comb;
  assign p3_res7__158_comb = p2_literal_1076345[p3_res7__157_comb] ^ p2_literal_1076347[p3_res7__156_comb] ^ p2_literal_1076349[p3_res7__155_comb] ^ p2_literal_1076351[p3_res7__154_comb] ^ p2_literal_1076353[p3_res7__153_comb] ^ p2_literal_1076355[p3_res7__152_comb] ^ p3_res7__151_comb ^ p2_literal_1076358[p3_res7__150_comb] ^ p3_res7__149_comb ^ p3_array_index_1079131_comb ^ p3_array_index_1079108_comb ^ p3_array_index_1079083_comb ^ p3_array_index_1079056_comb ^ p3_array_index_1079027_comb ^ p3_array_index_1078995_comb ^ p3_array_index_1078980_comb;
  assign p3_res7__557_comb = p2_literal_1076345[p3_res7__556_comb] ^ p2_literal_1076347[p3_res7__555_comb] ^ p2_literal_1076349[p3_res7__554_comb] ^ p2_literal_1076351[p3_res7__553_comb] ^ p2_literal_1076353[p3_res7__552_comb] ^ p2_literal_1076355[p3_res7__551_comb] ^ p3_res7__550_comb ^ p2_literal_1076358[p3_res7__549_comb] ^ p3_res7__548_comb ^ p3_array_index_1079555_comb ^ p3_array_index_1079531_comb ^ p3_array_index_1079505_comb ^ p3_array_index_1079477_comb ^ p3_array_index_1079448_comb ^ p2_literal_1076345[p3_array_index_1079415_comb] ^ p3_array_index_1079416_comb;
  assign p3_res7__159_comb = p2_literal_1076345[p3_res7__158_comb] ^ p2_literal_1076347[p3_res7__157_comb] ^ p2_literal_1076349[p3_res7__156_comb] ^ p2_literal_1076351[p3_res7__155_comb] ^ p2_literal_1076353[p3_res7__154_comb] ^ p2_literal_1076355[p3_res7__153_comb] ^ p3_res7__152_comb ^ p2_literal_1076358[p3_res7__151_comb] ^ p3_res7__150_comb ^ p3_array_index_1079141_comb ^ p3_array_index_1079119_comb ^ p3_array_index_1079095_comb ^ p3_array_index_1079069_comb ^ p3_array_index_1079041_comb ^ p3_array_index_1079012_comb ^ p3_array_index_1078979_comb;
  assign p3_res7__558_comb = p2_literal_1076345[p3_res7__557_comb] ^ p2_literal_1076347[p3_res7__556_comb] ^ p2_literal_1076349[p3_res7__555_comb] ^ p2_literal_1076351[p3_res7__554_comb] ^ p2_literal_1076353[p3_res7__553_comb] ^ p2_literal_1076355[p3_res7__552_comb] ^ p3_res7__551_comb ^ p2_literal_1076358[p3_res7__550_comb] ^ p3_res7__549_comb ^ p3_array_index_1079566_comb ^ p3_array_index_1079543_comb ^ p3_array_index_1079518_comb ^ p3_array_index_1079491_comb ^ p3_array_index_1079462_comb ^ p3_array_index_1079430_comb ^ p3_array_index_1079415_comb;
  assign p3_res__9_comb = {p3_res7__159_comb, p3_res7__158_comb, p3_res7__157_comb, p3_res7__156_comb, p3_res7__155_comb, p3_res7__154_comb, p3_res7__153_comb, p3_res7__152_comb, p3_res7__151_comb, p3_res7__150_comb, p3_res7__149_comb, p3_res7__148_comb, p3_res7__147_comb, p3_res7__146_comb, p3_res7__145_comb, p3_res7__144_comb};
  assign p3_xor_1079181_comb = p3_res__9_comb ^ p3_k2_comb;
  assign p3_res7__559_comb = p2_literal_1076345[p3_res7__558_comb] ^ p2_literal_1076347[p3_res7__557_comb] ^ p2_literal_1076349[p3_res7__556_comb] ^ p2_literal_1076351[p3_res7__555_comb] ^ p2_literal_1076353[p3_res7__554_comb] ^ p2_literal_1076355[p3_res7__553_comb] ^ p3_res7__552_comb ^ p2_literal_1076358[p3_res7__551_comb] ^ p3_res7__550_comb ^ p3_array_index_1079576_comb ^ p3_array_index_1079554_comb ^ p3_array_index_1079530_comb ^ p3_array_index_1079504_comb ^ p3_array_index_1079476_comb ^ p3_array_index_1079447_comb ^ p3_array_index_1079414_comb;
  assign p3_addedKey__51_comb = p3_xor_1079181_comb ^ 128'h447c_ac80_52dd_d882_4a92_a5b0_83e5_550b;
  assign p3_res__34_comb = {p3_res7__559_comb, p3_res7__558_comb, p3_res7__557_comb, p3_res7__556_comb, p3_res7__555_comb, p3_res7__554_comb, p3_res7__553_comb, p3_res7__552_comb, p3_res7__551_comb, p3_res7__550_comb, p3_res7__549_comb, p3_res7__548_comb, p3_res7__547_comb, p3_res7__546_comb, p3_res7__545_comb, p3_res7__544_comb};
  assign p3_addedKey__35_comb = p2_k3 ^ p3_res__34_comb;
  assign p3_array_index_1079197_comb = p2_arr[p3_addedKey__51_comb[127:120]];
  assign p3_array_index_1079198_comb = p2_arr[p3_addedKey__51_comb[119:112]];
  assign p3_array_index_1079199_comb = p2_arr[p3_addedKey__51_comb[111:104]];
  assign p3_array_index_1079200_comb = p2_arr[p3_addedKey__51_comb[103:96]];
  assign p3_array_index_1079201_comb = p2_arr[p3_addedKey__51_comb[95:88]];
  assign p3_array_index_1079202_comb = p2_arr[p3_addedKey__51_comb[87:80]];
  assign p3_array_index_1079204_comb = p2_arr[p3_addedKey__51_comb[71:64]];
  assign p3_array_index_1079206_comb = p2_arr[p3_addedKey__51_comb[55:48]];
  assign p3_array_index_1079207_comb = p2_arr[p3_addedKey__51_comb[47:40]];
  assign p3_array_index_1079208_comb = p2_arr[p3_addedKey__51_comb[39:32]];
  assign p3_array_index_1079209_comb = p2_arr[p3_addedKey__51_comb[31:24]];
  assign p3_array_index_1079210_comb = p2_arr[p3_addedKey__51_comb[23:16]];
  assign p3_array_index_1079211_comb = p2_arr[p3_addedKey__51_comb[15:8]];
  assign p3_array_index_1079213_comb = p2_literal_1076345[p3_array_index_1079197_comb];
  assign p3_array_index_1079214_comb = p2_literal_1076347[p3_array_index_1079198_comb];
  assign p3_array_index_1079215_comb = p2_literal_1076349[p3_array_index_1079199_comb];
  assign p3_array_index_1079216_comb = p2_literal_1076351[p3_array_index_1079200_comb];
  assign p3_array_index_1079217_comb = p2_literal_1076353[p3_array_index_1079201_comb];
  assign p3_array_index_1079218_comb = p2_literal_1076355[p3_array_index_1079202_comb];
  assign p3_array_index_1079219_comb = p2_arr[p3_addedKey__51_comb[79:72]];
  assign p3_array_index_1079221_comb = p2_arr[p3_addedKey__51_comb[63:56]];
  assign p3_array_index_1079630_comb = p2_arr[p3_addedKey__35_comb[127:120]];
  assign p3_array_index_1079631_comb = p2_arr[p3_addedKey__35_comb[119:112]];
  assign p3_array_index_1079632_comb = p2_arr[p3_addedKey__35_comb[111:104]];
  assign p3_array_index_1079633_comb = p2_arr[p3_addedKey__35_comb[103:96]];
  assign p3_array_index_1079634_comb = p2_arr[p3_addedKey__35_comb[95:88]];
  assign p3_array_index_1079635_comb = p2_arr[p3_addedKey__35_comb[87:80]];
  assign p3_array_index_1079637_comb = p2_arr[p3_addedKey__35_comb[71:64]];
  assign p3_array_index_1079639_comb = p2_arr[p3_addedKey__35_comb[55:48]];
  assign p3_array_index_1079640_comb = p2_arr[p3_addedKey__35_comb[47:40]];
  assign p3_array_index_1079641_comb = p2_arr[p3_addedKey__35_comb[39:32]];
  assign p3_array_index_1079642_comb = p2_arr[p3_addedKey__35_comb[31:24]];
  assign p3_array_index_1079643_comb = p2_arr[p3_addedKey__35_comb[23:16]];
  assign p3_array_index_1079644_comb = p2_arr[p3_addedKey__35_comb[15:8]];
  assign p3_res7__160_comb = p3_array_index_1079213_comb ^ p3_array_index_1079214_comb ^ p3_array_index_1079215_comb ^ p3_array_index_1079216_comb ^ p3_array_index_1079217_comb ^ p3_array_index_1079218_comb ^ p3_array_index_1079219_comb ^ p2_literal_1076358[p3_array_index_1079204_comb] ^ p3_array_index_1079221_comb ^ p2_literal_1076355[p3_array_index_1079206_comb] ^ p2_literal_1076353[p3_array_index_1079207_comb] ^ p2_literal_1076351[p3_array_index_1079208_comb] ^ p2_literal_1076349[p3_array_index_1079209_comb] ^ p2_literal_1076347[p3_array_index_1079210_comb] ^ p2_literal_1076345[p3_array_index_1079211_comb] ^ p2_arr[p3_addedKey__51_comb[7:0]];
  assign p3_array_index_1079646_comb = p2_literal_1076345[p3_array_index_1079630_comb];
  assign p3_array_index_1079647_comb = p2_literal_1076347[p3_array_index_1079631_comb];
  assign p3_array_index_1079648_comb = p2_literal_1076349[p3_array_index_1079632_comb];
  assign p3_array_index_1079649_comb = p2_literal_1076351[p3_array_index_1079633_comb];
  assign p3_array_index_1079650_comb = p2_literal_1076353[p3_array_index_1079634_comb];
  assign p3_array_index_1079651_comb = p2_literal_1076355[p3_array_index_1079635_comb];
  assign p3_array_index_1079652_comb = p2_arr[p3_addedKey__35_comb[79:72]];
  assign p3_array_index_1079654_comb = p2_arr[p3_addedKey__35_comb[63:56]];
  assign p3_array_index_1079230_comb = p2_literal_1076345[p3_res7__160_comb];
  assign p3_array_index_1079231_comb = p2_literal_1076347[p3_array_index_1079197_comb];
  assign p3_array_index_1079232_comb = p2_literal_1076349[p3_array_index_1079198_comb];
  assign p3_array_index_1079233_comb = p2_literal_1076351[p3_array_index_1079199_comb];
  assign p3_array_index_1079234_comb = p2_literal_1076353[p3_array_index_1079200_comb];
  assign p3_array_index_1079235_comb = p2_literal_1076355[p3_array_index_1079201_comb];
  assign p3_res7__560_comb = p3_array_index_1079646_comb ^ p3_array_index_1079647_comb ^ p3_array_index_1079648_comb ^ p3_array_index_1079649_comb ^ p3_array_index_1079650_comb ^ p3_array_index_1079651_comb ^ p3_array_index_1079652_comb ^ p2_literal_1076358[p3_array_index_1079637_comb] ^ p3_array_index_1079654_comb ^ p2_literal_1076355[p3_array_index_1079639_comb] ^ p2_literal_1076353[p3_array_index_1079640_comb] ^ p2_literal_1076351[p3_array_index_1079641_comb] ^ p2_literal_1076349[p3_array_index_1079642_comb] ^ p2_literal_1076347[p3_array_index_1079643_comb] ^ p2_literal_1076345[p3_array_index_1079644_comb] ^ p2_arr[p3_addedKey__35_comb[7:0]];
  assign p3_res7__161_comb = p3_array_index_1079230_comb ^ p3_array_index_1079231_comb ^ p3_array_index_1079232_comb ^ p3_array_index_1079233_comb ^ p3_array_index_1079234_comb ^ p3_array_index_1079235_comb ^ p3_array_index_1079202_comb ^ p2_literal_1076358[p3_array_index_1079219_comb] ^ p3_array_index_1079204_comb ^ p2_literal_1076355[p3_array_index_1079221_comb] ^ p2_literal_1076353[p3_array_index_1079206_comb] ^ p2_literal_1076351[p3_array_index_1079207_comb] ^ p2_literal_1076349[p3_array_index_1079208_comb] ^ p2_literal_1076347[p3_array_index_1079209_comb] ^ p2_literal_1076345[p3_array_index_1079210_comb] ^ p3_array_index_1079211_comb;
  assign p3_array_index_1079663_comb = p2_literal_1076345[p3_res7__560_comb];
  assign p3_array_index_1079664_comb = p2_literal_1076347[p3_array_index_1079630_comb];
  assign p3_array_index_1079665_comb = p2_literal_1076349[p3_array_index_1079631_comb];
  assign p3_array_index_1079666_comb = p2_literal_1076351[p3_array_index_1079632_comb];
  assign p3_array_index_1079667_comb = p2_literal_1076353[p3_array_index_1079633_comb];
  assign p3_array_index_1079668_comb = p2_literal_1076355[p3_array_index_1079634_comb];
  assign p3_array_index_1079245_comb = p2_literal_1076347[p3_res7__160_comb];
  assign p3_array_index_1079246_comb = p2_literal_1076349[p3_array_index_1079197_comb];
  assign p3_array_index_1079247_comb = p2_literal_1076351[p3_array_index_1079198_comb];
  assign p3_array_index_1079248_comb = p2_literal_1076353[p3_array_index_1079199_comb];
  assign p3_array_index_1079249_comb = p2_literal_1076355[p3_array_index_1079200_comb];
  assign p3_res7__561_comb = p3_array_index_1079663_comb ^ p3_array_index_1079664_comb ^ p3_array_index_1079665_comb ^ p3_array_index_1079666_comb ^ p3_array_index_1079667_comb ^ p3_array_index_1079668_comb ^ p3_array_index_1079635_comb ^ p2_literal_1076358[p3_array_index_1079652_comb] ^ p3_array_index_1079637_comb ^ p2_literal_1076355[p3_array_index_1079654_comb] ^ p2_literal_1076353[p3_array_index_1079639_comb] ^ p2_literal_1076351[p3_array_index_1079640_comb] ^ p2_literal_1076349[p3_array_index_1079641_comb] ^ p2_literal_1076347[p3_array_index_1079642_comb] ^ p2_literal_1076345[p3_array_index_1079643_comb] ^ p3_array_index_1079644_comb;
  assign p3_res7__162_comb = p2_literal_1076345[p3_res7__161_comb] ^ p3_array_index_1079245_comb ^ p3_array_index_1079246_comb ^ p3_array_index_1079247_comb ^ p3_array_index_1079248_comb ^ p3_array_index_1079249_comb ^ p3_array_index_1079201_comb ^ p2_literal_1076358[p3_array_index_1079202_comb] ^ p3_array_index_1079219_comb ^ p2_literal_1076355[p3_array_index_1079204_comb] ^ p2_literal_1076353[p3_array_index_1079221_comb] ^ p2_literal_1076351[p3_array_index_1079206_comb] ^ p2_literal_1076349[p3_array_index_1079207_comb] ^ p2_literal_1076347[p3_array_index_1079208_comb] ^ p2_literal_1076345[p3_array_index_1079209_comb] ^ p3_array_index_1079210_comb;
  assign p3_array_index_1079678_comb = p2_literal_1076347[p3_res7__560_comb];
  assign p3_array_index_1079679_comb = p2_literal_1076349[p3_array_index_1079630_comb];
  assign p3_array_index_1079680_comb = p2_literal_1076351[p3_array_index_1079631_comb];
  assign p3_array_index_1079681_comb = p2_literal_1076353[p3_array_index_1079632_comb];
  assign p3_array_index_1079682_comb = p2_literal_1076355[p3_array_index_1079633_comb];
  assign p3_array_index_1079259_comb = p2_literal_1076347[p3_res7__161_comb];
  assign p3_array_index_1079260_comb = p2_literal_1076349[p3_res7__160_comb];
  assign p3_array_index_1079261_comb = p2_literal_1076351[p3_array_index_1079197_comb];
  assign p3_array_index_1079262_comb = p2_literal_1076353[p3_array_index_1079198_comb];
  assign p3_array_index_1079263_comb = p2_literal_1076355[p3_array_index_1079199_comb];
  assign p3_res7__562_comb = p2_literal_1076345[p3_res7__561_comb] ^ p3_array_index_1079678_comb ^ p3_array_index_1079679_comb ^ p3_array_index_1079680_comb ^ p3_array_index_1079681_comb ^ p3_array_index_1079682_comb ^ p3_array_index_1079634_comb ^ p2_literal_1076358[p3_array_index_1079635_comb] ^ p3_array_index_1079652_comb ^ p2_literal_1076355[p3_array_index_1079637_comb] ^ p2_literal_1076353[p3_array_index_1079654_comb] ^ p2_literal_1076351[p3_array_index_1079639_comb] ^ p2_literal_1076349[p3_array_index_1079640_comb] ^ p2_literal_1076347[p3_array_index_1079641_comb] ^ p2_literal_1076345[p3_array_index_1079642_comb] ^ p3_array_index_1079643_comb;
  assign p3_res7__163_comb = p2_literal_1076345[p3_res7__162_comb] ^ p3_array_index_1079259_comb ^ p3_array_index_1079260_comb ^ p3_array_index_1079261_comb ^ p3_array_index_1079262_comb ^ p3_array_index_1079263_comb ^ p3_array_index_1079200_comb ^ p2_literal_1076358[p3_array_index_1079201_comb] ^ p3_array_index_1079202_comb ^ p2_literal_1076355[p3_array_index_1079219_comb] ^ p2_literal_1076353[p3_array_index_1079204_comb] ^ p2_literal_1076351[p3_array_index_1079221_comb] ^ p2_literal_1076349[p3_array_index_1079206_comb] ^ p2_literal_1076347[p3_array_index_1079207_comb] ^ p2_literal_1076345[p3_array_index_1079208_comb] ^ p3_array_index_1079209_comb;
  assign p3_array_index_1079692_comb = p2_literal_1076347[p3_res7__561_comb];
  assign p3_array_index_1079693_comb = p2_literal_1076349[p3_res7__560_comb];
  assign p3_array_index_1079694_comb = p2_literal_1076351[p3_array_index_1079630_comb];
  assign p3_array_index_1079695_comb = p2_literal_1076353[p3_array_index_1079631_comb];
  assign p3_array_index_1079696_comb = p2_literal_1076355[p3_array_index_1079632_comb];
  assign p3_array_index_1079274_comb = p2_literal_1076349[p3_res7__161_comb];
  assign p3_array_index_1079275_comb = p2_literal_1076351[p3_res7__160_comb];
  assign p3_array_index_1079276_comb = p2_literal_1076353[p3_array_index_1079197_comb];
  assign p3_array_index_1079277_comb = p2_literal_1076355[p3_array_index_1079198_comb];
  assign p3_res7__563_comb = p2_literal_1076345[p3_res7__562_comb] ^ p3_array_index_1079692_comb ^ p3_array_index_1079693_comb ^ p3_array_index_1079694_comb ^ p3_array_index_1079695_comb ^ p3_array_index_1079696_comb ^ p3_array_index_1079633_comb ^ p2_literal_1076358[p3_array_index_1079634_comb] ^ p3_array_index_1079635_comb ^ p2_literal_1076355[p3_array_index_1079652_comb] ^ p2_literal_1076353[p3_array_index_1079637_comb] ^ p2_literal_1076351[p3_array_index_1079654_comb] ^ p2_literal_1076349[p3_array_index_1079639_comb] ^ p2_literal_1076347[p3_array_index_1079640_comb] ^ p2_literal_1076345[p3_array_index_1079641_comb] ^ p3_array_index_1079642_comb;
  assign p3_res7__164_comb = p2_literal_1076345[p3_res7__163_comb] ^ p2_literal_1076347[p3_res7__162_comb] ^ p3_array_index_1079274_comb ^ p3_array_index_1079275_comb ^ p3_array_index_1079276_comb ^ p3_array_index_1079277_comb ^ p3_array_index_1079199_comb ^ p2_literal_1076358[p3_array_index_1079200_comb] ^ p3_array_index_1079201_comb ^ p3_array_index_1079218_comb ^ p2_literal_1076353[p3_array_index_1079219_comb] ^ p2_literal_1076351[p3_array_index_1079204_comb] ^ p2_literal_1076349[p3_array_index_1079221_comb] ^ p2_literal_1076347[p3_array_index_1079206_comb] ^ p2_literal_1076345[p3_array_index_1079207_comb] ^ p3_array_index_1079208_comb;
  assign p3_array_index_1079707_comb = p2_literal_1076349[p3_res7__561_comb];
  assign p3_array_index_1079708_comb = p2_literal_1076351[p3_res7__560_comb];
  assign p3_array_index_1079709_comb = p2_literal_1076353[p3_array_index_1079630_comb];
  assign p3_array_index_1079710_comb = p2_literal_1076355[p3_array_index_1079631_comb];
  assign p3_array_index_1079287_comb = p2_literal_1076349[p3_res7__162_comb];
  assign p3_array_index_1079288_comb = p2_literal_1076351[p3_res7__161_comb];
  assign p3_array_index_1079289_comb = p2_literal_1076353[p3_res7__160_comb];
  assign p3_array_index_1079290_comb = p2_literal_1076355[p3_array_index_1079197_comb];
  assign p3_res7__564_comb = p2_literal_1076345[p3_res7__563_comb] ^ p2_literal_1076347[p3_res7__562_comb] ^ p3_array_index_1079707_comb ^ p3_array_index_1079708_comb ^ p3_array_index_1079709_comb ^ p3_array_index_1079710_comb ^ p3_array_index_1079632_comb ^ p2_literal_1076358[p3_array_index_1079633_comb] ^ p3_array_index_1079634_comb ^ p3_array_index_1079651_comb ^ p2_literal_1076353[p3_array_index_1079652_comb] ^ p2_literal_1076351[p3_array_index_1079637_comb] ^ p2_literal_1076349[p3_array_index_1079654_comb] ^ p2_literal_1076347[p3_array_index_1079639_comb] ^ p2_literal_1076345[p3_array_index_1079640_comb] ^ p3_array_index_1079641_comb;
  assign p3_res7__165_comb = p2_literal_1076345[p3_res7__164_comb] ^ p2_literal_1076347[p3_res7__163_comb] ^ p3_array_index_1079287_comb ^ p3_array_index_1079288_comb ^ p3_array_index_1079289_comb ^ p3_array_index_1079290_comb ^ p3_array_index_1079198_comb ^ p2_literal_1076358[p3_array_index_1079199_comb] ^ p3_array_index_1079200_comb ^ p3_array_index_1079235_comb ^ p2_literal_1076353[p3_array_index_1079202_comb] ^ p2_literal_1076351[p3_array_index_1079219_comb] ^ p2_literal_1076349[p3_array_index_1079204_comb] ^ p2_literal_1076347[p3_array_index_1079221_comb] ^ p2_literal_1076345[p3_array_index_1079206_comb] ^ p3_array_index_1079207_comb;
  assign p3_array_index_1079720_comb = p2_literal_1076349[p3_res7__562_comb];
  assign p3_array_index_1079721_comb = p2_literal_1076351[p3_res7__561_comb];
  assign p3_array_index_1079722_comb = p2_literal_1076353[p3_res7__560_comb];
  assign p3_array_index_1079723_comb = p2_literal_1076355[p3_array_index_1079630_comb];
  assign p3_array_index_1079301_comb = p2_literal_1076351[p3_res7__162_comb];
  assign p3_array_index_1079302_comb = p2_literal_1076353[p3_res7__161_comb];
  assign p3_array_index_1079303_comb = p2_literal_1076355[p3_res7__160_comb];
  assign p3_res7__565_comb = p2_literal_1076345[p3_res7__564_comb] ^ p2_literal_1076347[p3_res7__563_comb] ^ p3_array_index_1079720_comb ^ p3_array_index_1079721_comb ^ p3_array_index_1079722_comb ^ p3_array_index_1079723_comb ^ p3_array_index_1079631_comb ^ p2_literal_1076358[p3_array_index_1079632_comb] ^ p3_array_index_1079633_comb ^ p3_array_index_1079668_comb ^ p2_literal_1076353[p3_array_index_1079635_comb] ^ p2_literal_1076351[p3_array_index_1079652_comb] ^ p2_literal_1076349[p3_array_index_1079637_comb] ^ p2_literal_1076347[p3_array_index_1079654_comb] ^ p2_literal_1076345[p3_array_index_1079639_comb] ^ p3_array_index_1079640_comb;
  assign p3_res7__166_comb = p2_literal_1076345[p3_res7__165_comb] ^ p2_literal_1076347[p3_res7__164_comb] ^ p2_literal_1076349[p3_res7__163_comb] ^ p3_array_index_1079301_comb ^ p3_array_index_1079302_comb ^ p3_array_index_1079303_comb ^ p3_array_index_1079197_comb ^ p2_literal_1076358[p3_array_index_1079198_comb] ^ p3_array_index_1079199_comb ^ p3_array_index_1079249_comb ^ p3_array_index_1079217_comb ^ p2_literal_1076351[p3_array_index_1079202_comb] ^ p2_literal_1076349[p3_array_index_1079219_comb] ^ p2_literal_1076347[p3_array_index_1079204_comb] ^ p2_literal_1076345[p3_array_index_1079221_comb] ^ p3_array_index_1079206_comb;
  assign p3_array_index_1079734_comb = p2_literal_1076351[p3_res7__562_comb];
  assign p3_array_index_1079735_comb = p2_literal_1076353[p3_res7__561_comb];
  assign p3_array_index_1079736_comb = p2_literal_1076355[p3_res7__560_comb];
  assign p3_array_index_1079313_comb = p2_literal_1076351[p3_res7__163_comb];
  assign p3_array_index_1079314_comb = p2_literal_1076353[p3_res7__162_comb];
  assign p3_array_index_1079315_comb = p2_literal_1076355[p3_res7__161_comb];
  assign p3_res7__566_comb = p2_literal_1076345[p3_res7__565_comb] ^ p2_literal_1076347[p3_res7__564_comb] ^ p2_literal_1076349[p3_res7__563_comb] ^ p3_array_index_1079734_comb ^ p3_array_index_1079735_comb ^ p3_array_index_1079736_comb ^ p3_array_index_1079630_comb ^ p2_literal_1076358[p3_array_index_1079631_comb] ^ p3_array_index_1079632_comb ^ p3_array_index_1079682_comb ^ p3_array_index_1079650_comb ^ p2_literal_1076351[p3_array_index_1079635_comb] ^ p2_literal_1076349[p3_array_index_1079652_comb] ^ p2_literal_1076347[p3_array_index_1079637_comb] ^ p2_literal_1076345[p3_array_index_1079654_comb] ^ p3_array_index_1079639_comb;
  assign p3_res7__167_comb = p2_literal_1076345[p3_res7__166_comb] ^ p2_literal_1076347[p3_res7__165_comb] ^ p2_literal_1076349[p3_res7__164_comb] ^ p3_array_index_1079313_comb ^ p3_array_index_1079314_comb ^ p3_array_index_1079315_comb ^ p3_res7__160_comb ^ p2_literal_1076358[p3_array_index_1079197_comb] ^ p3_array_index_1079198_comb ^ p3_array_index_1079263_comb ^ p3_array_index_1079234_comb ^ p2_literal_1076351[p3_array_index_1079201_comb] ^ p2_literal_1076349[p3_array_index_1079202_comb] ^ p2_literal_1076347[p3_array_index_1079219_comb] ^ p2_literal_1076345[p3_array_index_1079204_comb] ^ p3_array_index_1079221_comb;
  assign p3_array_index_1079746_comb = p2_literal_1076351[p3_res7__563_comb];
  assign p3_array_index_1079747_comb = p2_literal_1076353[p3_res7__562_comb];
  assign p3_array_index_1079748_comb = p2_literal_1076355[p3_res7__561_comb];
  assign p3_array_index_1079326_comb = p2_literal_1076353[p3_res7__163_comb];
  assign p3_array_index_1079327_comb = p2_literal_1076355[p3_res7__162_comb];
  assign p3_res7__567_comb = p2_literal_1076345[p3_res7__566_comb] ^ p2_literal_1076347[p3_res7__565_comb] ^ p2_literal_1076349[p3_res7__564_comb] ^ p3_array_index_1079746_comb ^ p3_array_index_1079747_comb ^ p3_array_index_1079748_comb ^ p3_res7__560_comb ^ p2_literal_1076358[p3_array_index_1079630_comb] ^ p3_array_index_1079631_comb ^ p3_array_index_1079696_comb ^ p3_array_index_1079667_comb ^ p2_literal_1076351[p3_array_index_1079634_comb] ^ p2_literal_1076349[p3_array_index_1079635_comb] ^ p2_literal_1076347[p3_array_index_1079652_comb] ^ p2_literal_1076345[p3_array_index_1079637_comb] ^ p3_array_index_1079654_comb;
  assign p3_res7__168_comb = p2_literal_1076345[p3_res7__167_comb] ^ p2_literal_1076347[p3_res7__166_comb] ^ p2_literal_1076349[p3_res7__165_comb] ^ p2_literal_1076351[p3_res7__164_comb] ^ p3_array_index_1079326_comb ^ p3_array_index_1079327_comb ^ p3_res7__161_comb ^ p2_literal_1076358[p3_res7__160_comb] ^ p3_array_index_1079197_comb ^ p3_array_index_1079277_comb ^ p3_array_index_1079248_comb ^ p3_array_index_1079216_comb ^ p2_literal_1076349[p3_array_index_1079201_comb] ^ p2_literal_1076347[p3_array_index_1079202_comb] ^ p2_literal_1076345[p3_array_index_1079219_comb] ^ p3_array_index_1079204_comb;
  assign p3_array_index_1079759_comb = p2_literal_1076353[p3_res7__563_comb];
  assign p3_array_index_1079760_comb = p2_literal_1076355[p3_res7__562_comb];
  assign p3_array_index_1079337_comb = p2_literal_1076353[p3_res7__164_comb];
  assign p3_array_index_1079338_comb = p2_literal_1076355[p3_res7__163_comb];
  assign p3_res7__568_comb = p2_literal_1076345[p3_res7__567_comb] ^ p2_literal_1076347[p3_res7__566_comb] ^ p2_literal_1076349[p3_res7__565_comb] ^ p2_literal_1076351[p3_res7__564_comb] ^ p3_array_index_1079759_comb ^ p3_array_index_1079760_comb ^ p3_res7__561_comb ^ p2_literal_1076358[p3_res7__560_comb] ^ p3_array_index_1079630_comb ^ p3_array_index_1079710_comb ^ p3_array_index_1079681_comb ^ p3_array_index_1079649_comb ^ p2_literal_1076349[p3_array_index_1079634_comb] ^ p2_literal_1076347[p3_array_index_1079635_comb] ^ p2_literal_1076345[p3_array_index_1079652_comb] ^ p3_array_index_1079637_comb;
  assign p3_res7__169_comb = p2_literal_1076345[p3_res7__168_comb] ^ p2_literal_1076347[p3_res7__167_comb] ^ p2_literal_1076349[p3_res7__166_comb] ^ p2_literal_1076351[p3_res7__165_comb] ^ p3_array_index_1079337_comb ^ p3_array_index_1079338_comb ^ p3_res7__162_comb ^ p2_literal_1076358[p3_res7__161_comb] ^ p3_res7__160_comb ^ p3_array_index_1079290_comb ^ p3_array_index_1079262_comb ^ p3_array_index_1079233_comb ^ p2_literal_1076349[p3_array_index_1079200_comb] ^ p2_literal_1076347[p3_array_index_1079201_comb] ^ p2_literal_1076345[p3_array_index_1079202_comb] ^ p3_array_index_1079219_comb;
  assign p3_array_index_1079770_comb = p2_literal_1076353[p3_res7__564_comb];
  assign p3_array_index_1079771_comb = p2_literal_1076355[p3_res7__563_comb];
  assign p3_array_index_1079349_comb = p2_literal_1076355[p3_res7__164_comb];
  assign p3_res7__569_comb = p2_literal_1076345[p3_res7__568_comb] ^ p2_literal_1076347[p3_res7__567_comb] ^ p2_literal_1076349[p3_res7__566_comb] ^ p2_literal_1076351[p3_res7__565_comb] ^ p3_array_index_1079770_comb ^ p3_array_index_1079771_comb ^ p3_res7__562_comb ^ p2_literal_1076358[p3_res7__561_comb] ^ p3_res7__560_comb ^ p3_array_index_1079723_comb ^ p3_array_index_1079695_comb ^ p3_array_index_1079666_comb ^ p2_literal_1076349[p3_array_index_1079633_comb] ^ p2_literal_1076347[p3_array_index_1079634_comb] ^ p2_literal_1076345[p3_array_index_1079635_comb] ^ p3_array_index_1079652_comb;
  assign p3_res7__170_comb = p2_literal_1076345[p3_res7__169_comb] ^ p2_literal_1076347[p3_res7__168_comb] ^ p2_literal_1076349[p3_res7__167_comb] ^ p2_literal_1076351[p3_res7__166_comb] ^ p2_literal_1076353[p3_res7__165_comb] ^ p3_array_index_1079349_comb ^ p3_res7__163_comb ^ p2_literal_1076358[p3_res7__162_comb] ^ p3_res7__161_comb ^ p3_array_index_1079303_comb ^ p3_array_index_1079276_comb ^ p3_array_index_1079247_comb ^ p3_array_index_1079215_comb ^ p2_literal_1076347[p3_array_index_1079200_comb] ^ p2_literal_1076345[p3_array_index_1079201_comb] ^ p3_array_index_1079202_comb;
  assign p3_array_index_1079782_comb = p2_literal_1076355[p3_res7__564_comb];
  assign p3_array_index_1079359_comb = p2_literal_1076355[p3_res7__165_comb];
  assign p3_res7__570_comb = p2_literal_1076345[p3_res7__569_comb] ^ p2_literal_1076347[p3_res7__568_comb] ^ p2_literal_1076349[p3_res7__567_comb] ^ p2_literal_1076351[p3_res7__566_comb] ^ p2_literal_1076353[p3_res7__565_comb] ^ p3_array_index_1079782_comb ^ p3_res7__563_comb ^ p2_literal_1076358[p3_res7__562_comb] ^ p3_res7__561_comb ^ p3_array_index_1079736_comb ^ p3_array_index_1079709_comb ^ p3_array_index_1079680_comb ^ p3_array_index_1079648_comb ^ p2_literal_1076347[p3_array_index_1079633_comb] ^ p2_literal_1076345[p3_array_index_1079634_comb] ^ p3_array_index_1079635_comb;
  assign p3_res7__171_comb = p2_literal_1076345[p3_res7__170_comb] ^ p2_literal_1076347[p3_res7__169_comb] ^ p2_literal_1076349[p3_res7__168_comb] ^ p2_literal_1076351[p3_res7__167_comb] ^ p2_literal_1076353[p3_res7__166_comb] ^ p3_array_index_1079359_comb ^ p3_res7__164_comb ^ p2_literal_1076358[p3_res7__163_comb] ^ p3_res7__162_comb ^ p3_array_index_1079315_comb ^ p3_array_index_1079289_comb ^ p3_array_index_1079261_comb ^ p3_array_index_1079232_comb ^ p2_literal_1076347[p3_array_index_1079199_comb] ^ p2_literal_1076345[p3_array_index_1079200_comb] ^ p3_array_index_1079201_comb;
  assign p3_array_index_1079792_comb = p2_literal_1076355[p3_res7__565_comb];
  assign p3_res7__571_comb = p2_literal_1076345[p3_res7__570_comb] ^ p2_literal_1076347[p3_res7__569_comb] ^ p2_literal_1076349[p3_res7__568_comb] ^ p2_literal_1076351[p3_res7__567_comb] ^ p2_literal_1076353[p3_res7__566_comb] ^ p3_array_index_1079792_comb ^ p3_res7__564_comb ^ p2_literal_1076358[p3_res7__563_comb] ^ p3_res7__562_comb ^ p3_array_index_1079748_comb ^ p3_array_index_1079722_comb ^ p3_array_index_1079694_comb ^ p3_array_index_1079665_comb ^ p2_literal_1076347[p3_array_index_1079632_comb] ^ p2_literal_1076345[p3_array_index_1079633_comb] ^ p3_array_index_1079634_comb;
  assign p3_res7__172_comb = p2_literal_1076345[p3_res7__171_comb] ^ p2_literal_1076347[p3_res7__170_comb] ^ p2_literal_1076349[p3_res7__169_comb] ^ p2_literal_1076351[p3_res7__168_comb] ^ p2_literal_1076353[p3_res7__167_comb] ^ p2_literal_1076355[p3_res7__166_comb] ^ p3_res7__165_comb ^ p2_literal_1076358[p3_res7__164_comb] ^ p3_res7__163_comb ^ p3_array_index_1079327_comb ^ p3_array_index_1079302_comb ^ p3_array_index_1079275_comb ^ p3_array_index_1079246_comb ^ p3_array_index_1079214_comb ^ p2_literal_1076345[p3_array_index_1079199_comb] ^ p3_array_index_1079200_comb;
  assign p3_res7__572_comb = p2_literal_1076345[p3_res7__571_comb] ^ p2_literal_1076347[p3_res7__570_comb] ^ p2_literal_1076349[p3_res7__569_comb] ^ p2_literal_1076351[p3_res7__568_comb] ^ p2_literal_1076353[p3_res7__567_comb] ^ p2_literal_1076355[p3_res7__566_comb] ^ p3_res7__565_comb ^ p2_literal_1076358[p3_res7__564_comb] ^ p3_res7__563_comb ^ p3_array_index_1079760_comb ^ p3_array_index_1079735_comb ^ p3_array_index_1079708_comb ^ p3_array_index_1079679_comb ^ p3_array_index_1079647_comb ^ p2_literal_1076345[p3_array_index_1079632_comb] ^ p3_array_index_1079633_comb;
  assign p3_res7__173_comb = p2_literal_1076345[p3_res7__172_comb] ^ p2_literal_1076347[p3_res7__171_comb] ^ p2_literal_1076349[p3_res7__170_comb] ^ p2_literal_1076351[p3_res7__169_comb] ^ p2_literal_1076353[p3_res7__168_comb] ^ p2_literal_1076355[p3_res7__167_comb] ^ p3_res7__166_comb ^ p2_literal_1076358[p3_res7__165_comb] ^ p3_res7__164_comb ^ p3_array_index_1079338_comb ^ p3_array_index_1079314_comb ^ p3_array_index_1079288_comb ^ p3_array_index_1079260_comb ^ p3_array_index_1079231_comb ^ p2_literal_1076345[p3_array_index_1079198_comb] ^ p3_array_index_1079199_comb;
  assign p3_res7__573_comb = p2_literal_1076345[p3_res7__572_comb] ^ p2_literal_1076347[p3_res7__571_comb] ^ p2_literal_1076349[p3_res7__570_comb] ^ p2_literal_1076351[p3_res7__569_comb] ^ p2_literal_1076353[p3_res7__568_comb] ^ p2_literal_1076355[p3_res7__567_comb] ^ p3_res7__566_comb ^ p2_literal_1076358[p3_res7__565_comb] ^ p3_res7__564_comb ^ p3_array_index_1079771_comb ^ p3_array_index_1079747_comb ^ p3_array_index_1079721_comb ^ p3_array_index_1079693_comb ^ p3_array_index_1079664_comb ^ p2_literal_1076345[p3_array_index_1079631_comb] ^ p3_array_index_1079632_comb;
  assign p3_res7__174_comb = p2_literal_1076345[p3_res7__173_comb] ^ p2_literal_1076347[p3_res7__172_comb] ^ p2_literal_1076349[p3_res7__171_comb] ^ p2_literal_1076351[p3_res7__170_comb] ^ p2_literal_1076353[p3_res7__169_comb] ^ p2_literal_1076355[p3_res7__168_comb] ^ p3_res7__167_comb ^ p2_literal_1076358[p3_res7__166_comb] ^ p3_res7__165_comb ^ p3_array_index_1079349_comb ^ p3_array_index_1079326_comb ^ p3_array_index_1079301_comb ^ p3_array_index_1079274_comb ^ p3_array_index_1079245_comb ^ p3_array_index_1079213_comb ^ p3_array_index_1079198_comb;
  assign p3_res7__574_comb = p2_literal_1076345[p3_res7__573_comb] ^ p2_literal_1076347[p3_res7__572_comb] ^ p2_literal_1076349[p3_res7__571_comb] ^ p2_literal_1076351[p3_res7__570_comb] ^ p2_literal_1076353[p3_res7__569_comb] ^ p2_literal_1076355[p3_res7__568_comb] ^ p3_res7__567_comb ^ p2_literal_1076358[p3_res7__566_comb] ^ p3_res7__565_comb ^ p3_array_index_1079782_comb ^ p3_array_index_1079759_comb ^ p3_array_index_1079734_comb ^ p3_array_index_1079707_comb ^ p3_array_index_1079678_comb ^ p3_array_index_1079646_comb ^ p3_array_index_1079631_comb;
  assign p3_res7__175_comb = p2_literal_1076345[p3_res7__174_comb] ^ p2_literal_1076347[p3_res7__173_comb] ^ p2_literal_1076349[p3_res7__172_comb] ^ p2_literal_1076351[p3_res7__171_comb] ^ p2_literal_1076353[p3_res7__170_comb] ^ p2_literal_1076355[p3_res7__169_comb] ^ p3_res7__168_comb ^ p2_literal_1076358[p3_res7__167_comb] ^ p3_res7__166_comb ^ p3_array_index_1079359_comb ^ p3_array_index_1079337_comb ^ p3_array_index_1079313_comb ^ p3_array_index_1079287_comb ^ p3_array_index_1079259_comb ^ p3_array_index_1079230_comb ^ p3_array_index_1079197_comb;
  assign p3_res__10_comb = {p3_res7__175_comb, p3_res7__174_comb, p3_res7__173_comb, p3_res7__172_comb, p3_res7__171_comb, p3_res7__170_comb, p3_res7__169_comb, p3_res7__168_comb, p3_res7__167_comb, p3_res7__166_comb, p3_res7__165_comb, p3_res7__164_comb, p3_res7__163_comb, p3_res7__162_comb, p3_res7__161_comb, p3_res7__160_comb};
  assign p3_res7__575_comb = p2_literal_1076345[p3_res7__574_comb] ^ p2_literal_1076347[p3_res7__573_comb] ^ p2_literal_1076349[p3_res7__572_comb] ^ p2_literal_1076351[p3_res7__571_comb] ^ p2_literal_1076353[p3_res7__570_comb] ^ p2_literal_1076355[p3_res7__569_comb] ^ p3_res7__568_comb ^ p2_literal_1076358[p3_res7__567_comb] ^ p3_res7__566_comb ^ p3_array_index_1079792_comb ^ p3_array_index_1079770_comb ^ p3_array_index_1079746_comb ^ p3_array_index_1079720_comb ^ p3_array_index_1079692_comb ^ p3_array_index_1079663_comb ^ p3_array_index_1079630_comb;
  assign p3_xor_1079399_comb = p3_res__10_comb ^ p3_xor_1078963_comb;
  assign p3_res__35_comb = {p3_res7__575_comb, p3_res7__574_comb, p3_res7__573_comb, p3_res7__572_comb, p3_res7__571_comb, p3_res7__570_comb, p3_res7__569_comb, p3_res7__568_comb, p3_res7__567_comb, p3_res7__566_comb, p3_res7__565_comb, p3_res7__564_comb, p3_res7__563_comb, p3_res7__562_comb, p3_res7__561_comb, p3_res7__560_comb};

  // Registers for pipe stage 3:
  reg [127:0] p3_xor_1079181;
  reg [127:0] p3_xor_1079399;
  reg [127:0] p3_res__35;
  reg [7:0] p4_arr[256];
  reg [7:0] p4_literal_1076345[256];
  reg [7:0] p4_literal_1076347[256];
  reg [7:0] p4_literal_1076349[256];
  reg [7:0] p4_literal_1076351[256];
  reg [7:0] p4_literal_1076353[256];
  reg [7:0] p4_literal_1076355[256];
  reg [7:0] p4_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p3_xor_1079181 <= p3_xor_1079181_comb;
    p3_xor_1079399 <= p3_xor_1079399_comb;
    p3_res__35 <= p3_res__35_comb;
    p4_arr <= p3_arr;
    p4_literal_1076345 <= p3_literal_1076345;
    p4_literal_1076347 <= p3_literal_1076347;
    p4_literal_1076349 <= p3_literal_1076349;
    p4_literal_1076351 <= p3_literal_1076351;
    p4_literal_1076353 <= p3_literal_1076353;
    p4_literal_1076355 <= p3_literal_1076355;
    p4_literal_1076358 <= p3_literal_1076358;
  end

  // ===== Pipe stage 4:
  wire [127:0] p4_addedKey__52_comb;
  wire [7:0] p4_array_index_1079869_comb;
  wire [7:0] p4_array_index_1079870_comb;
  wire [7:0] p4_array_index_1079871_comb;
  wire [7:0] p4_array_index_1079872_comb;
  wire [7:0] p4_array_index_1079873_comb;
  wire [7:0] p4_array_index_1079874_comb;
  wire [7:0] p4_array_index_1079876_comb;
  wire [7:0] p4_array_index_1079878_comb;
  wire [7:0] p4_array_index_1079879_comb;
  wire [7:0] p4_array_index_1079880_comb;
  wire [7:0] p4_array_index_1079881_comb;
  wire [7:0] p4_array_index_1079882_comb;
  wire [7:0] p4_array_index_1079883_comb;
  wire [7:0] p4_array_index_1079885_comb;
  wire [7:0] p4_array_index_1079886_comb;
  wire [7:0] p4_array_index_1079887_comb;
  wire [7:0] p4_array_index_1079888_comb;
  wire [7:0] p4_array_index_1079889_comb;
  wire [7:0] p4_array_index_1079890_comb;
  wire [7:0] p4_array_index_1079891_comb;
  wire [7:0] p4_array_index_1079893_comb;
  wire [7:0] p4_res7__176_comb;
  wire [7:0] p4_array_index_1079902_comb;
  wire [7:0] p4_array_index_1079903_comb;
  wire [7:0] p4_array_index_1079904_comb;
  wire [7:0] p4_array_index_1079905_comb;
  wire [7:0] p4_array_index_1079906_comb;
  wire [7:0] p4_array_index_1079907_comb;
  wire [7:0] p4_res7__177_comb;
  wire [7:0] p4_array_index_1079917_comb;
  wire [7:0] p4_array_index_1079918_comb;
  wire [7:0] p4_array_index_1079919_comb;
  wire [7:0] p4_array_index_1079920_comb;
  wire [7:0] p4_array_index_1079921_comb;
  wire [7:0] p4_res7__178_comb;
  wire [7:0] p4_array_index_1079931_comb;
  wire [7:0] p4_array_index_1079932_comb;
  wire [7:0] p4_array_index_1079933_comb;
  wire [7:0] p4_array_index_1079934_comb;
  wire [7:0] p4_array_index_1079935_comb;
  wire [7:0] p4_res7__179_comb;
  wire [7:0] p4_array_index_1079946_comb;
  wire [7:0] p4_array_index_1079947_comb;
  wire [7:0] p4_array_index_1079948_comb;
  wire [7:0] p4_array_index_1079949_comb;
  wire [7:0] p4_res7__180_comb;
  wire [7:0] p4_array_index_1079959_comb;
  wire [7:0] p4_array_index_1079960_comb;
  wire [7:0] p4_array_index_1079961_comb;
  wire [7:0] p4_array_index_1079962_comb;
  wire [7:0] p4_res7__181_comb;
  wire [7:0] p4_array_index_1079973_comb;
  wire [7:0] p4_array_index_1079974_comb;
  wire [7:0] p4_array_index_1079975_comb;
  wire [7:0] p4_res7__182_comb;
  wire [7:0] p4_array_index_1079985_comb;
  wire [7:0] p4_array_index_1079986_comb;
  wire [7:0] p4_array_index_1079987_comb;
  wire [7:0] p4_res7__183_comb;
  wire [7:0] p4_array_index_1079998_comb;
  wire [7:0] p4_array_index_1079999_comb;
  wire [7:0] p4_res7__184_comb;
  wire [7:0] p4_array_index_1080009_comb;
  wire [7:0] p4_array_index_1080010_comb;
  wire [7:0] p4_res7__185_comb;
  wire [7:0] p4_array_index_1080021_comb;
  wire [7:0] p4_res7__186_comb;
  wire [7:0] p4_array_index_1080031_comb;
  wire [7:0] p4_res7__187_comb;
  wire [7:0] p4_res7__188_comb;
  wire [7:0] p4_res7__189_comb;
  wire [7:0] p4_res7__190_comb;
  wire [7:0] p4_res7__191_comb;
  wire [127:0] p4_res__11_comb;
  wire [127:0] p4_xor_1080071_comb;
  wire [127:0] p4_addedKey__53_comb;
  wire [7:0] p4_array_index_1080087_comb;
  wire [7:0] p4_array_index_1080088_comb;
  wire [7:0] p4_array_index_1080089_comb;
  wire [7:0] p4_array_index_1080090_comb;
  wire [7:0] p4_array_index_1080091_comb;
  wire [7:0] p4_array_index_1080092_comb;
  wire [7:0] p4_array_index_1080094_comb;
  wire [7:0] p4_array_index_1080096_comb;
  wire [7:0] p4_array_index_1080097_comb;
  wire [7:0] p4_array_index_1080098_comb;
  wire [7:0] p4_array_index_1080099_comb;
  wire [7:0] p4_array_index_1080100_comb;
  wire [7:0] p4_array_index_1080101_comb;
  wire [7:0] p4_array_index_1080103_comb;
  wire [7:0] p4_array_index_1080104_comb;
  wire [7:0] p4_array_index_1080105_comb;
  wire [7:0] p4_array_index_1080106_comb;
  wire [7:0] p4_array_index_1080107_comb;
  wire [7:0] p4_array_index_1080108_comb;
  wire [7:0] p4_array_index_1080109_comb;
  wire [7:0] p4_array_index_1080111_comb;
  wire [7:0] p4_res7__192_comb;
  wire [7:0] p4_array_index_1080120_comb;
  wire [7:0] p4_array_index_1080121_comb;
  wire [7:0] p4_array_index_1080122_comb;
  wire [7:0] p4_array_index_1080123_comb;
  wire [7:0] p4_array_index_1080124_comb;
  wire [7:0] p4_array_index_1080125_comb;
  wire [7:0] p4_res7__193_comb;
  wire [7:0] p4_array_index_1080135_comb;
  wire [7:0] p4_array_index_1080136_comb;
  wire [7:0] p4_array_index_1080137_comb;
  wire [7:0] p4_array_index_1080138_comb;
  wire [7:0] p4_array_index_1080139_comb;
  wire [7:0] p4_res7__194_comb;
  wire [7:0] p4_array_index_1080149_comb;
  wire [7:0] p4_array_index_1080150_comb;
  wire [7:0] p4_array_index_1080151_comb;
  wire [7:0] p4_array_index_1080152_comb;
  wire [7:0] p4_array_index_1080153_comb;
  wire [7:0] p4_res7__195_comb;
  wire [7:0] p4_array_index_1080164_comb;
  wire [7:0] p4_array_index_1080165_comb;
  wire [7:0] p4_array_index_1080166_comb;
  wire [7:0] p4_array_index_1080167_comb;
  wire [7:0] p4_res7__196_comb;
  wire [7:0] p4_array_index_1080177_comb;
  wire [7:0] p4_array_index_1080178_comb;
  wire [7:0] p4_array_index_1080179_comb;
  wire [7:0] p4_array_index_1080180_comb;
  wire [7:0] p4_res7__197_comb;
  wire [7:0] p4_array_index_1080191_comb;
  wire [7:0] p4_array_index_1080192_comb;
  wire [7:0] p4_array_index_1080193_comb;
  wire [7:0] p4_res7__198_comb;
  wire [7:0] p4_array_index_1080203_comb;
  wire [7:0] p4_array_index_1080204_comb;
  wire [7:0] p4_array_index_1080205_comb;
  wire [7:0] p4_res7__199_comb;
  wire [7:0] p4_array_index_1080216_comb;
  wire [7:0] p4_array_index_1080217_comb;
  wire [7:0] p4_res7__200_comb;
  wire [7:0] p4_array_index_1080227_comb;
  wire [7:0] p4_array_index_1080228_comb;
  wire [7:0] p4_res7__201_comb;
  wire [7:0] p4_array_index_1080239_comb;
  wire [7:0] p4_res7__202_comb;
  wire [7:0] p4_array_index_1080249_comb;
  wire [7:0] p4_res7__203_comb;
  wire [7:0] p4_res7__204_comb;
  wire [7:0] p4_res7__205_comb;
  wire [7:0] p4_res7__206_comb;
  wire [7:0] p4_res7__207_comb;
  wire [127:0] p4_res__12_comb;
  wire [127:0] p4_xor_1080289_comb;
  wire [127:0] p4_addedKey__54_comb;
  wire [7:0] p4_array_index_1080305_comb;
  wire [7:0] p4_array_index_1080306_comb;
  wire [7:0] p4_array_index_1080307_comb;
  wire [7:0] p4_array_index_1080308_comb;
  wire [7:0] p4_array_index_1080309_comb;
  wire [7:0] p4_array_index_1080310_comb;
  wire [7:0] p4_array_index_1080312_comb;
  wire [7:0] p4_array_index_1080314_comb;
  wire [7:0] p4_array_index_1080315_comb;
  wire [7:0] p4_array_index_1080316_comb;
  wire [7:0] p4_array_index_1080317_comb;
  wire [7:0] p4_array_index_1080318_comb;
  wire [7:0] p4_array_index_1080319_comb;
  wire [7:0] p4_array_index_1080321_comb;
  wire [7:0] p4_array_index_1080322_comb;
  wire [7:0] p4_array_index_1080323_comb;
  wire [7:0] p4_array_index_1080324_comb;
  wire [7:0] p4_array_index_1080325_comb;
  wire [7:0] p4_array_index_1080326_comb;
  wire [7:0] p4_array_index_1080327_comb;
  wire [7:0] p4_array_index_1080329_comb;
  wire [7:0] p4_res7__208_comb;
  wire [7:0] p4_array_index_1080338_comb;
  wire [7:0] p4_array_index_1080339_comb;
  wire [7:0] p4_array_index_1080340_comb;
  wire [7:0] p4_array_index_1080341_comb;
  wire [7:0] p4_array_index_1080342_comb;
  wire [7:0] p4_array_index_1080343_comb;
  wire [7:0] p4_res7__209_comb;
  wire [7:0] p4_array_index_1080353_comb;
  wire [7:0] p4_array_index_1080354_comb;
  wire [7:0] p4_array_index_1080355_comb;
  wire [7:0] p4_array_index_1080356_comb;
  wire [7:0] p4_array_index_1080357_comb;
  wire [7:0] p4_res7__210_comb;
  wire [7:0] p4_array_index_1080367_comb;
  wire [7:0] p4_array_index_1080368_comb;
  wire [7:0] p4_array_index_1080369_comb;
  wire [7:0] p4_array_index_1080370_comb;
  wire [7:0] p4_array_index_1080371_comb;
  wire [7:0] p4_res7__211_comb;
  wire [7:0] p4_array_index_1080382_comb;
  wire [7:0] p4_array_index_1080383_comb;
  wire [7:0] p4_array_index_1080384_comb;
  wire [7:0] p4_array_index_1080385_comb;
  wire [7:0] p4_res7__212_comb;
  wire [7:0] p4_array_index_1080395_comb;
  wire [7:0] p4_array_index_1080396_comb;
  wire [7:0] p4_array_index_1080397_comb;
  wire [7:0] p4_array_index_1080398_comb;
  wire [7:0] p4_res7__213_comb;
  wire [7:0] p4_array_index_1080409_comb;
  wire [7:0] p4_array_index_1080410_comb;
  wire [7:0] p4_array_index_1080411_comb;
  wire [7:0] p4_res7__214_comb;
  wire [7:0] p4_array_index_1080421_comb;
  wire [7:0] p4_array_index_1080422_comb;
  wire [7:0] p4_array_index_1080423_comb;
  wire [7:0] p4_res7__215_comb;
  wire [7:0] p4_array_index_1080434_comb;
  wire [7:0] p4_array_index_1080435_comb;
  wire [7:0] p4_res7__216_comb;
  wire [7:0] p4_array_index_1080445_comb;
  wire [7:0] p4_array_index_1080446_comb;
  wire [7:0] p4_res7__217_comb;
  wire [7:0] p4_array_index_1080457_comb;
  wire [7:0] p4_res7__218_comb;
  wire [7:0] p4_array_index_1080467_comb;
  wire [7:0] p4_res7__219_comb;
  wire [7:0] p4_res7__220_comb;
  wire [7:0] p4_res7__221_comb;
  wire [7:0] p4_res7__222_comb;
  wire [7:0] p4_res7__223_comb;
  wire [127:0] p4_res__13_comb;
  wire [127:0] p4_xor_1080507_comb;
  wire [127:0] p4_addedKey__55_comb;
  wire [7:0] p4_array_index_1080523_comb;
  wire [7:0] p4_array_index_1080524_comb;
  wire [7:0] p4_array_index_1080525_comb;
  wire [7:0] p4_array_index_1080526_comb;
  wire [7:0] p4_array_index_1080527_comb;
  wire [7:0] p4_array_index_1080528_comb;
  wire [7:0] p4_array_index_1080530_comb;
  wire [7:0] p4_array_index_1080532_comb;
  wire [7:0] p4_array_index_1080533_comb;
  wire [7:0] p4_array_index_1080534_comb;
  wire [7:0] p4_array_index_1080535_comb;
  wire [7:0] p4_array_index_1080536_comb;
  wire [7:0] p4_array_index_1080537_comb;
  wire [7:0] p4_array_index_1080539_comb;
  wire [7:0] p4_array_index_1080540_comb;
  wire [7:0] p4_array_index_1080541_comb;
  wire [7:0] p4_array_index_1080542_comb;
  wire [7:0] p4_array_index_1080543_comb;
  wire [7:0] p4_array_index_1080544_comb;
  wire [7:0] p4_array_index_1080545_comb;
  wire [7:0] p4_array_index_1080547_comb;
  wire [7:0] p4_res7__224_comb;
  wire [7:0] p4_array_index_1080556_comb;
  wire [7:0] p4_array_index_1080557_comb;
  wire [7:0] p4_array_index_1080558_comb;
  wire [7:0] p4_array_index_1080559_comb;
  wire [7:0] p4_array_index_1080560_comb;
  wire [7:0] p4_array_index_1080561_comb;
  wire [7:0] p4_res7__225_comb;
  wire [7:0] p4_array_index_1080571_comb;
  wire [7:0] p4_array_index_1080572_comb;
  wire [7:0] p4_array_index_1080573_comb;
  wire [7:0] p4_array_index_1080574_comb;
  wire [7:0] p4_array_index_1080575_comb;
  wire [7:0] p4_res7__226_comb;
  wire [7:0] p4_array_index_1080585_comb;
  wire [7:0] p4_array_index_1080586_comb;
  wire [7:0] p4_array_index_1080587_comb;
  wire [7:0] p4_array_index_1080588_comb;
  wire [7:0] p4_array_index_1080589_comb;
  wire [7:0] p4_res7__227_comb;
  wire [7:0] p4_array_index_1080600_comb;
  wire [7:0] p4_array_index_1080601_comb;
  wire [7:0] p4_array_index_1080602_comb;
  wire [7:0] p4_array_index_1080603_comb;
  wire [7:0] p4_res7__228_comb;
  wire [7:0] p4_array_index_1080613_comb;
  wire [7:0] p4_array_index_1080614_comb;
  wire [7:0] p4_array_index_1080615_comb;
  wire [7:0] p4_array_index_1080616_comb;
  wire [7:0] p4_res7__229_comb;
  wire [7:0] p4_array_index_1080627_comb;
  wire [7:0] p4_array_index_1080628_comb;
  wire [7:0] p4_array_index_1080629_comb;
  wire [7:0] p4_res7__230_comb;
  wire [7:0] p4_array_index_1080639_comb;
  wire [7:0] p4_array_index_1080640_comb;
  wire [7:0] p4_array_index_1080641_comb;
  wire [7:0] p4_res7__231_comb;
  wire [7:0] p4_array_index_1080652_comb;
  wire [7:0] p4_array_index_1080653_comb;
  wire [7:0] p4_res7__232_comb;
  wire [7:0] p4_array_index_1080663_comb;
  wire [7:0] p4_array_index_1080664_comb;
  wire [7:0] p4_res7__233_comb;
  wire [7:0] p4_array_index_1080670_comb;
  wire [7:0] p4_array_index_1080671_comb;
  wire [7:0] p4_array_index_1080672_comb;
  wire [7:0] p4_array_index_1080673_comb;
  wire [7:0] p4_array_index_1080674_comb;
  wire [7:0] p4_array_index_1080675_comb;
  wire [7:0] p4_array_index_1080676_comb;
  wire [7:0] p4_array_index_1080677_comb;
  wire [7:0] p4_array_index_1080678_comb;
  assign p4_addedKey__52_comb = p3_xor_1079399 ^ 128'h8d94_2d1d_95e6_7d2c_1a67_10c0_d5ff_3f0c;
  assign p4_array_index_1079869_comb = p3_arr[p4_addedKey__52_comb[127:120]];
  assign p4_array_index_1079870_comb = p3_arr[p4_addedKey__52_comb[119:112]];
  assign p4_array_index_1079871_comb = p3_arr[p4_addedKey__52_comb[111:104]];
  assign p4_array_index_1079872_comb = p3_arr[p4_addedKey__52_comb[103:96]];
  assign p4_array_index_1079873_comb = p3_arr[p4_addedKey__52_comb[95:88]];
  assign p4_array_index_1079874_comb = p3_arr[p4_addedKey__52_comb[87:80]];
  assign p4_array_index_1079876_comb = p3_arr[p4_addedKey__52_comb[71:64]];
  assign p4_array_index_1079878_comb = p3_arr[p4_addedKey__52_comb[55:48]];
  assign p4_array_index_1079879_comb = p3_arr[p4_addedKey__52_comb[47:40]];
  assign p4_array_index_1079880_comb = p3_arr[p4_addedKey__52_comb[39:32]];
  assign p4_array_index_1079881_comb = p3_arr[p4_addedKey__52_comb[31:24]];
  assign p4_array_index_1079882_comb = p3_arr[p4_addedKey__52_comb[23:16]];
  assign p4_array_index_1079883_comb = p3_arr[p4_addedKey__52_comb[15:8]];
  assign p4_array_index_1079885_comb = p3_literal_1076345[p4_array_index_1079869_comb];
  assign p4_array_index_1079886_comb = p3_literal_1076347[p4_array_index_1079870_comb];
  assign p4_array_index_1079887_comb = p3_literal_1076349[p4_array_index_1079871_comb];
  assign p4_array_index_1079888_comb = p3_literal_1076351[p4_array_index_1079872_comb];
  assign p4_array_index_1079889_comb = p3_literal_1076353[p4_array_index_1079873_comb];
  assign p4_array_index_1079890_comb = p3_literal_1076355[p4_array_index_1079874_comb];
  assign p4_array_index_1079891_comb = p3_arr[p4_addedKey__52_comb[79:72]];
  assign p4_array_index_1079893_comb = p3_arr[p4_addedKey__52_comb[63:56]];
  assign p4_res7__176_comb = p4_array_index_1079885_comb ^ p4_array_index_1079886_comb ^ p4_array_index_1079887_comb ^ p4_array_index_1079888_comb ^ p4_array_index_1079889_comb ^ p4_array_index_1079890_comb ^ p4_array_index_1079891_comb ^ p3_literal_1076358[p4_array_index_1079876_comb] ^ p4_array_index_1079893_comb ^ p3_literal_1076355[p4_array_index_1079878_comb] ^ p3_literal_1076353[p4_array_index_1079879_comb] ^ p3_literal_1076351[p4_array_index_1079880_comb] ^ p3_literal_1076349[p4_array_index_1079881_comb] ^ p3_literal_1076347[p4_array_index_1079882_comb] ^ p3_literal_1076345[p4_array_index_1079883_comb] ^ p3_arr[p4_addedKey__52_comb[7:0]];
  assign p4_array_index_1079902_comb = p3_literal_1076345[p4_res7__176_comb];
  assign p4_array_index_1079903_comb = p3_literal_1076347[p4_array_index_1079869_comb];
  assign p4_array_index_1079904_comb = p3_literal_1076349[p4_array_index_1079870_comb];
  assign p4_array_index_1079905_comb = p3_literal_1076351[p4_array_index_1079871_comb];
  assign p4_array_index_1079906_comb = p3_literal_1076353[p4_array_index_1079872_comb];
  assign p4_array_index_1079907_comb = p3_literal_1076355[p4_array_index_1079873_comb];
  assign p4_res7__177_comb = p4_array_index_1079902_comb ^ p4_array_index_1079903_comb ^ p4_array_index_1079904_comb ^ p4_array_index_1079905_comb ^ p4_array_index_1079906_comb ^ p4_array_index_1079907_comb ^ p4_array_index_1079874_comb ^ p3_literal_1076358[p4_array_index_1079891_comb] ^ p4_array_index_1079876_comb ^ p3_literal_1076355[p4_array_index_1079893_comb] ^ p3_literal_1076353[p4_array_index_1079878_comb] ^ p3_literal_1076351[p4_array_index_1079879_comb] ^ p3_literal_1076349[p4_array_index_1079880_comb] ^ p3_literal_1076347[p4_array_index_1079881_comb] ^ p3_literal_1076345[p4_array_index_1079882_comb] ^ p4_array_index_1079883_comb;
  assign p4_array_index_1079917_comb = p3_literal_1076347[p4_res7__176_comb];
  assign p4_array_index_1079918_comb = p3_literal_1076349[p4_array_index_1079869_comb];
  assign p4_array_index_1079919_comb = p3_literal_1076351[p4_array_index_1079870_comb];
  assign p4_array_index_1079920_comb = p3_literal_1076353[p4_array_index_1079871_comb];
  assign p4_array_index_1079921_comb = p3_literal_1076355[p4_array_index_1079872_comb];
  assign p4_res7__178_comb = p3_literal_1076345[p4_res7__177_comb] ^ p4_array_index_1079917_comb ^ p4_array_index_1079918_comb ^ p4_array_index_1079919_comb ^ p4_array_index_1079920_comb ^ p4_array_index_1079921_comb ^ p4_array_index_1079873_comb ^ p3_literal_1076358[p4_array_index_1079874_comb] ^ p4_array_index_1079891_comb ^ p3_literal_1076355[p4_array_index_1079876_comb] ^ p3_literal_1076353[p4_array_index_1079893_comb] ^ p3_literal_1076351[p4_array_index_1079878_comb] ^ p3_literal_1076349[p4_array_index_1079879_comb] ^ p3_literal_1076347[p4_array_index_1079880_comb] ^ p3_literal_1076345[p4_array_index_1079881_comb] ^ p4_array_index_1079882_comb;
  assign p4_array_index_1079931_comb = p3_literal_1076347[p4_res7__177_comb];
  assign p4_array_index_1079932_comb = p3_literal_1076349[p4_res7__176_comb];
  assign p4_array_index_1079933_comb = p3_literal_1076351[p4_array_index_1079869_comb];
  assign p4_array_index_1079934_comb = p3_literal_1076353[p4_array_index_1079870_comb];
  assign p4_array_index_1079935_comb = p3_literal_1076355[p4_array_index_1079871_comb];
  assign p4_res7__179_comb = p3_literal_1076345[p4_res7__178_comb] ^ p4_array_index_1079931_comb ^ p4_array_index_1079932_comb ^ p4_array_index_1079933_comb ^ p4_array_index_1079934_comb ^ p4_array_index_1079935_comb ^ p4_array_index_1079872_comb ^ p3_literal_1076358[p4_array_index_1079873_comb] ^ p4_array_index_1079874_comb ^ p3_literal_1076355[p4_array_index_1079891_comb] ^ p3_literal_1076353[p4_array_index_1079876_comb] ^ p3_literal_1076351[p4_array_index_1079893_comb] ^ p3_literal_1076349[p4_array_index_1079878_comb] ^ p3_literal_1076347[p4_array_index_1079879_comb] ^ p3_literal_1076345[p4_array_index_1079880_comb] ^ p4_array_index_1079881_comb;
  assign p4_array_index_1079946_comb = p3_literal_1076349[p4_res7__177_comb];
  assign p4_array_index_1079947_comb = p3_literal_1076351[p4_res7__176_comb];
  assign p4_array_index_1079948_comb = p3_literal_1076353[p4_array_index_1079869_comb];
  assign p4_array_index_1079949_comb = p3_literal_1076355[p4_array_index_1079870_comb];
  assign p4_res7__180_comb = p3_literal_1076345[p4_res7__179_comb] ^ p3_literal_1076347[p4_res7__178_comb] ^ p4_array_index_1079946_comb ^ p4_array_index_1079947_comb ^ p4_array_index_1079948_comb ^ p4_array_index_1079949_comb ^ p4_array_index_1079871_comb ^ p3_literal_1076358[p4_array_index_1079872_comb] ^ p4_array_index_1079873_comb ^ p4_array_index_1079890_comb ^ p3_literal_1076353[p4_array_index_1079891_comb] ^ p3_literal_1076351[p4_array_index_1079876_comb] ^ p3_literal_1076349[p4_array_index_1079893_comb] ^ p3_literal_1076347[p4_array_index_1079878_comb] ^ p3_literal_1076345[p4_array_index_1079879_comb] ^ p4_array_index_1079880_comb;
  assign p4_array_index_1079959_comb = p3_literal_1076349[p4_res7__178_comb];
  assign p4_array_index_1079960_comb = p3_literal_1076351[p4_res7__177_comb];
  assign p4_array_index_1079961_comb = p3_literal_1076353[p4_res7__176_comb];
  assign p4_array_index_1079962_comb = p3_literal_1076355[p4_array_index_1079869_comb];
  assign p4_res7__181_comb = p3_literal_1076345[p4_res7__180_comb] ^ p3_literal_1076347[p4_res7__179_comb] ^ p4_array_index_1079959_comb ^ p4_array_index_1079960_comb ^ p4_array_index_1079961_comb ^ p4_array_index_1079962_comb ^ p4_array_index_1079870_comb ^ p3_literal_1076358[p4_array_index_1079871_comb] ^ p4_array_index_1079872_comb ^ p4_array_index_1079907_comb ^ p3_literal_1076353[p4_array_index_1079874_comb] ^ p3_literal_1076351[p4_array_index_1079891_comb] ^ p3_literal_1076349[p4_array_index_1079876_comb] ^ p3_literal_1076347[p4_array_index_1079893_comb] ^ p3_literal_1076345[p4_array_index_1079878_comb] ^ p4_array_index_1079879_comb;
  assign p4_array_index_1079973_comb = p3_literal_1076351[p4_res7__178_comb];
  assign p4_array_index_1079974_comb = p3_literal_1076353[p4_res7__177_comb];
  assign p4_array_index_1079975_comb = p3_literal_1076355[p4_res7__176_comb];
  assign p4_res7__182_comb = p3_literal_1076345[p4_res7__181_comb] ^ p3_literal_1076347[p4_res7__180_comb] ^ p3_literal_1076349[p4_res7__179_comb] ^ p4_array_index_1079973_comb ^ p4_array_index_1079974_comb ^ p4_array_index_1079975_comb ^ p4_array_index_1079869_comb ^ p3_literal_1076358[p4_array_index_1079870_comb] ^ p4_array_index_1079871_comb ^ p4_array_index_1079921_comb ^ p4_array_index_1079889_comb ^ p3_literal_1076351[p4_array_index_1079874_comb] ^ p3_literal_1076349[p4_array_index_1079891_comb] ^ p3_literal_1076347[p4_array_index_1079876_comb] ^ p3_literal_1076345[p4_array_index_1079893_comb] ^ p4_array_index_1079878_comb;
  assign p4_array_index_1079985_comb = p3_literal_1076351[p4_res7__179_comb];
  assign p4_array_index_1079986_comb = p3_literal_1076353[p4_res7__178_comb];
  assign p4_array_index_1079987_comb = p3_literal_1076355[p4_res7__177_comb];
  assign p4_res7__183_comb = p3_literal_1076345[p4_res7__182_comb] ^ p3_literal_1076347[p4_res7__181_comb] ^ p3_literal_1076349[p4_res7__180_comb] ^ p4_array_index_1079985_comb ^ p4_array_index_1079986_comb ^ p4_array_index_1079987_comb ^ p4_res7__176_comb ^ p3_literal_1076358[p4_array_index_1079869_comb] ^ p4_array_index_1079870_comb ^ p4_array_index_1079935_comb ^ p4_array_index_1079906_comb ^ p3_literal_1076351[p4_array_index_1079873_comb] ^ p3_literal_1076349[p4_array_index_1079874_comb] ^ p3_literal_1076347[p4_array_index_1079891_comb] ^ p3_literal_1076345[p4_array_index_1079876_comb] ^ p4_array_index_1079893_comb;
  assign p4_array_index_1079998_comb = p3_literal_1076353[p4_res7__179_comb];
  assign p4_array_index_1079999_comb = p3_literal_1076355[p4_res7__178_comb];
  assign p4_res7__184_comb = p3_literal_1076345[p4_res7__183_comb] ^ p3_literal_1076347[p4_res7__182_comb] ^ p3_literal_1076349[p4_res7__181_comb] ^ p3_literal_1076351[p4_res7__180_comb] ^ p4_array_index_1079998_comb ^ p4_array_index_1079999_comb ^ p4_res7__177_comb ^ p3_literal_1076358[p4_res7__176_comb] ^ p4_array_index_1079869_comb ^ p4_array_index_1079949_comb ^ p4_array_index_1079920_comb ^ p4_array_index_1079888_comb ^ p3_literal_1076349[p4_array_index_1079873_comb] ^ p3_literal_1076347[p4_array_index_1079874_comb] ^ p3_literal_1076345[p4_array_index_1079891_comb] ^ p4_array_index_1079876_comb;
  assign p4_array_index_1080009_comb = p3_literal_1076353[p4_res7__180_comb];
  assign p4_array_index_1080010_comb = p3_literal_1076355[p4_res7__179_comb];
  assign p4_res7__185_comb = p3_literal_1076345[p4_res7__184_comb] ^ p3_literal_1076347[p4_res7__183_comb] ^ p3_literal_1076349[p4_res7__182_comb] ^ p3_literal_1076351[p4_res7__181_comb] ^ p4_array_index_1080009_comb ^ p4_array_index_1080010_comb ^ p4_res7__178_comb ^ p3_literal_1076358[p4_res7__177_comb] ^ p4_res7__176_comb ^ p4_array_index_1079962_comb ^ p4_array_index_1079934_comb ^ p4_array_index_1079905_comb ^ p3_literal_1076349[p4_array_index_1079872_comb] ^ p3_literal_1076347[p4_array_index_1079873_comb] ^ p3_literal_1076345[p4_array_index_1079874_comb] ^ p4_array_index_1079891_comb;
  assign p4_array_index_1080021_comb = p3_literal_1076355[p4_res7__180_comb];
  assign p4_res7__186_comb = p3_literal_1076345[p4_res7__185_comb] ^ p3_literal_1076347[p4_res7__184_comb] ^ p3_literal_1076349[p4_res7__183_comb] ^ p3_literal_1076351[p4_res7__182_comb] ^ p3_literal_1076353[p4_res7__181_comb] ^ p4_array_index_1080021_comb ^ p4_res7__179_comb ^ p3_literal_1076358[p4_res7__178_comb] ^ p4_res7__177_comb ^ p4_array_index_1079975_comb ^ p4_array_index_1079948_comb ^ p4_array_index_1079919_comb ^ p4_array_index_1079887_comb ^ p3_literal_1076347[p4_array_index_1079872_comb] ^ p3_literal_1076345[p4_array_index_1079873_comb] ^ p4_array_index_1079874_comb;
  assign p4_array_index_1080031_comb = p3_literal_1076355[p4_res7__181_comb];
  assign p4_res7__187_comb = p3_literal_1076345[p4_res7__186_comb] ^ p3_literal_1076347[p4_res7__185_comb] ^ p3_literal_1076349[p4_res7__184_comb] ^ p3_literal_1076351[p4_res7__183_comb] ^ p3_literal_1076353[p4_res7__182_comb] ^ p4_array_index_1080031_comb ^ p4_res7__180_comb ^ p3_literal_1076358[p4_res7__179_comb] ^ p4_res7__178_comb ^ p4_array_index_1079987_comb ^ p4_array_index_1079961_comb ^ p4_array_index_1079933_comb ^ p4_array_index_1079904_comb ^ p3_literal_1076347[p4_array_index_1079871_comb] ^ p3_literal_1076345[p4_array_index_1079872_comb] ^ p4_array_index_1079873_comb;
  assign p4_res7__188_comb = p3_literal_1076345[p4_res7__187_comb] ^ p3_literal_1076347[p4_res7__186_comb] ^ p3_literal_1076349[p4_res7__185_comb] ^ p3_literal_1076351[p4_res7__184_comb] ^ p3_literal_1076353[p4_res7__183_comb] ^ p3_literal_1076355[p4_res7__182_comb] ^ p4_res7__181_comb ^ p3_literal_1076358[p4_res7__180_comb] ^ p4_res7__179_comb ^ p4_array_index_1079999_comb ^ p4_array_index_1079974_comb ^ p4_array_index_1079947_comb ^ p4_array_index_1079918_comb ^ p4_array_index_1079886_comb ^ p3_literal_1076345[p4_array_index_1079871_comb] ^ p4_array_index_1079872_comb;
  assign p4_res7__189_comb = p3_literal_1076345[p4_res7__188_comb] ^ p3_literal_1076347[p4_res7__187_comb] ^ p3_literal_1076349[p4_res7__186_comb] ^ p3_literal_1076351[p4_res7__185_comb] ^ p3_literal_1076353[p4_res7__184_comb] ^ p3_literal_1076355[p4_res7__183_comb] ^ p4_res7__182_comb ^ p3_literal_1076358[p4_res7__181_comb] ^ p4_res7__180_comb ^ p4_array_index_1080010_comb ^ p4_array_index_1079986_comb ^ p4_array_index_1079960_comb ^ p4_array_index_1079932_comb ^ p4_array_index_1079903_comb ^ p3_literal_1076345[p4_array_index_1079870_comb] ^ p4_array_index_1079871_comb;
  assign p4_res7__190_comb = p3_literal_1076345[p4_res7__189_comb] ^ p3_literal_1076347[p4_res7__188_comb] ^ p3_literal_1076349[p4_res7__187_comb] ^ p3_literal_1076351[p4_res7__186_comb] ^ p3_literal_1076353[p4_res7__185_comb] ^ p3_literal_1076355[p4_res7__184_comb] ^ p4_res7__183_comb ^ p3_literal_1076358[p4_res7__182_comb] ^ p4_res7__181_comb ^ p4_array_index_1080021_comb ^ p4_array_index_1079998_comb ^ p4_array_index_1079973_comb ^ p4_array_index_1079946_comb ^ p4_array_index_1079917_comb ^ p4_array_index_1079885_comb ^ p4_array_index_1079870_comb;
  assign p4_res7__191_comb = p3_literal_1076345[p4_res7__190_comb] ^ p3_literal_1076347[p4_res7__189_comb] ^ p3_literal_1076349[p4_res7__188_comb] ^ p3_literal_1076351[p4_res7__187_comb] ^ p3_literal_1076353[p4_res7__186_comb] ^ p3_literal_1076355[p4_res7__185_comb] ^ p4_res7__184_comb ^ p3_literal_1076358[p4_res7__183_comb] ^ p4_res7__182_comb ^ p4_array_index_1080031_comb ^ p4_array_index_1080009_comb ^ p4_array_index_1079985_comb ^ p4_array_index_1079959_comb ^ p4_array_index_1079931_comb ^ p4_array_index_1079902_comb ^ p4_array_index_1079869_comb;
  assign p4_res__11_comb = {p4_res7__191_comb, p4_res7__190_comb, p4_res7__189_comb, p4_res7__188_comb, p4_res7__187_comb, p4_res7__186_comb, p4_res7__185_comb, p4_res7__184_comb, p4_res7__183_comb, p4_res7__182_comb, p4_res7__181_comb, p4_res7__180_comb, p4_res7__179_comb, p4_res7__178_comb, p4_res7__177_comb, p4_res7__176_comb};
  assign p4_xor_1080071_comb = p4_res__11_comb ^ p3_xor_1079181;
  assign p4_addedKey__53_comb = p4_xor_1080071_comb ^ 128'he336_5b6f_f9ae_0794_4740_add0_087b_ab0d;
  assign p4_array_index_1080087_comb = p3_arr[p4_addedKey__53_comb[127:120]];
  assign p4_array_index_1080088_comb = p3_arr[p4_addedKey__53_comb[119:112]];
  assign p4_array_index_1080089_comb = p3_arr[p4_addedKey__53_comb[111:104]];
  assign p4_array_index_1080090_comb = p3_arr[p4_addedKey__53_comb[103:96]];
  assign p4_array_index_1080091_comb = p3_arr[p4_addedKey__53_comb[95:88]];
  assign p4_array_index_1080092_comb = p3_arr[p4_addedKey__53_comb[87:80]];
  assign p4_array_index_1080094_comb = p3_arr[p4_addedKey__53_comb[71:64]];
  assign p4_array_index_1080096_comb = p3_arr[p4_addedKey__53_comb[55:48]];
  assign p4_array_index_1080097_comb = p3_arr[p4_addedKey__53_comb[47:40]];
  assign p4_array_index_1080098_comb = p3_arr[p4_addedKey__53_comb[39:32]];
  assign p4_array_index_1080099_comb = p3_arr[p4_addedKey__53_comb[31:24]];
  assign p4_array_index_1080100_comb = p3_arr[p4_addedKey__53_comb[23:16]];
  assign p4_array_index_1080101_comb = p3_arr[p4_addedKey__53_comb[15:8]];
  assign p4_array_index_1080103_comb = p3_literal_1076345[p4_array_index_1080087_comb];
  assign p4_array_index_1080104_comb = p3_literal_1076347[p4_array_index_1080088_comb];
  assign p4_array_index_1080105_comb = p3_literal_1076349[p4_array_index_1080089_comb];
  assign p4_array_index_1080106_comb = p3_literal_1076351[p4_array_index_1080090_comb];
  assign p4_array_index_1080107_comb = p3_literal_1076353[p4_array_index_1080091_comb];
  assign p4_array_index_1080108_comb = p3_literal_1076355[p4_array_index_1080092_comb];
  assign p4_array_index_1080109_comb = p3_arr[p4_addedKey__53_comb[79:72]];
  assign p4_array_index_1080111_comb = p3_arr[p4_addedKey__53_comb[63:56]];
  assign p4_res7__192_comb = p4_array_index_1080103_comb ^ p4_array_index_1080104_comb ^ p4_array_index_1080105_comb ^ p4_array_index_1080106_comb ^ p4_array_index_1080107_comb ^ p4_array_index_1080108_comb ^ p4_array_index_1080109_comb ^ p3_literal_1076358[p4_array_index_1080094_comb] ^ p4_array_index_1080111_comb ^ p3_literal_1076355[p4_array_index_1080096_comb] ^ p3_literal_1076353[p4_array_index_1080097_comb] ^ p3_literal_1076351[p4_array_index_1080098_comb] ^ p3_literal_1076349[p4_array_index_1080099_comb] ^ p3_literal_1076347[p4_array_index_1080100_comb] ^ p3_literal_1076345[p4_array_index_1080101_comb] ^ p3_arr[p4_addedKey__53_comb[7:0]];
  assign p4_array_index_1080120_comb = p3_literal_1076345[p4_res7__192_comb];
  assign p4_array_index_1080121_comb = p3_literal_1076347[p4_array_index_1080087_comb];
  assign p4_array_index_1080122_comb = p3_literal_1076349[p4_array_index_1080088_comb];
  assign p4_array_index_1080123_comb = p3_literal_1076351[p4_array_index_1080089_comb];
  assign p4_array_index_1080124_comb = p3_literal_1076353[p4_array_index_1080090_comb];
  assign p4_array_index_1080125_comb = p3_literal_1076355[p4_array_index_1080091_comb];
  assign p4_res7__193_comb = p4_array_index_1080120_comb ^ p4_array_index_1080121_comb ^ p4_array_index_1080122_comb ^ p4_array_index_1080123_comb ^ p4_array_index_1080124_comb ^ p4_array_index_1080125_comb ^ p4_array_index_1080092_comb ^ p3_literal_1076358[p4_array_index_1080109_comb] ^ p4_array_index_1080094_comb ^ p3_literal_1076355[p4_array_index_1080111_comb] ^ p3_literal_1076353[p4_array_index_1080096_comb] ^ p3_literal_1076351[p4_array_index_1080097_comb] ^ p3_literal_1076349[p4_array_index_1080098_comb] ^ p3_literal_1076347[p4_array_index_1080099_comb] ^ p3_literal_1076345[p4_array_index_1080100_comb] ^ p4_array_index_1080101_comb;
  assign p4_array_index_1080135_comb = p3_literal_1076347[p4_res7__192_comb];
  assign p4_array_index_1080136_comb = p3_literal_1076349[p4_array_index_1080087_comb];
  assign p4_array_index_1080137_comb = p3_literal_1076351[p4_array_index_1080088_comb];
  assign p4_array_index_1080138_comb = p3_literal_1076353[p4_array_index_1080089_comb];
  assign p4_array_index_1080139_comb = p3_literal_1076355[p4_array_index_1080090_comb];
  assign p4_res7__194_comb = p3_literal_1076345[p4_res7__193_comb] ^ p4_array_index_1080135_comb ^ p4_array_index_1080136_comb ^ p4_array_index_1080137_comb ^ p4_array_index_1080138_comb ^ p4_array_index_1080139_comb ^ p4_array_index_1080091_comb ^ p3_literal_1076358[p4_array_index_1080092_comb] ^ p4_array_index_1080109_comb ^ p3_literal_1076355[p4_array_index_1080094_comb] ^ p3_literal_1076353[p4_array_index_1080111_comb] ^ p3_literal_1076351[p4_array_index_1080096_comb] ^ p3_literal_1076349[p4_array_index_1080097_comb] ^ p3_literal_1076347[p4_array_index_1080098_comb] ^ p3_literal_1076345[p4_array_index_1080099_comb] ^ p4_array_index_1080100_comb;
  assign p4_array_index_1080149_comb = p3_literal_1076347[p4_res7__193_comb];
  assign p4_array_index_1080150_comb = p3_literal_1076349[p4_res7__192_comb];
  assign p4_array_index_1080151_comb = p3_literal_1076351[p4_array_index_1080087_comb];
  assign p4_array_index_1080152_comb = p3_literal_1076353[p4_array_index_1080088_comb];
  assign p4_array_index_1080153_comb = p3_literal_1076355[p4_array_index_1080089_comb];
  assign p4_res7__195_comb = p3_literal_1076345[p4_res7__194_comb] ^ p4_array_index_1080149_comb ^ p4_array_index_1080150_comb ^ p4_array_index_1080151_comb ^ p4_array_index_1080152_comb ^ p4_array_index_1080153_comb ^ p4_array_index_1080090_comb ^ p3_literal_1076358[p4_array_index_1080091_comb] ^ p4_array_index_1080092_comb ^ p3_literal_1076355[p4_array_index_1080109_comb] ^ p3_literal_1076353[p4_array_index_1080094_comb] ^ p3_literal_1076351[p4_array_index_1080111_comb] ^ p3_literal_1076349[p4_array_index_1080096_comb] ^ p3_literal_1076347[p4_array_index_1080097_comb] ^ p3_literal_1076345[p4_array_index_1080098_comb] ^ p4_array_index_1080099_comb;
  assign p4_array_index_1080164_comb = p3_literal_1076349[p4_res7__193_comb];
  assign p4_array_index_1080165_comb = p3_literal_1076351[p4_res7__192_comb];
  assign p4_array_index_1080166_comb = p3_literal_1076353[p4_array_index_1080087_comb];
  assign p4_array_index_1080167_comb = p3_literal_1076355[p4_array_index_1080088_comb];
  assign p4_res7__196_comb = p3_literal_1076345[p4_res7__195_comb] ^ p3_literal_1076347[p4_res7__194_comb] ^ p4_array_index_1080164_comb ^ p4_array_index_1080165_comb ^ p4_array_index_1080166_comb ^ p4_array_index_1080167_comb ^ p4_array_index_1080089_comb ^ p3_literal_1076358[p4_array_index_1080090_comb] ^ p4_array_index_1080091_comb ^ p4_array_index_1080108_comb ^ p3_literal_1076353[p4_array_index_1080109_comb] ^ p3_literal_1076351[p4_array_index_1080094_comb] ^ p3_literal_1076349[p4_array_index_1080111_comb] ^ p3_literal_1076347[p4_array_index_1080096_comb] ^ p3_literal_1076345[p4_array_index_1080097_comb] ^ p4_array_index_1080098_comb;
  assign p4_array_index_1080177_comb = p3_literal_1076349[p4_res7__194_comb];
  assign p4_array_index_1080178_comb = p3_literal_1076351[p4_res7__193_comb];
  assign p4_array_index_1080179_comb = p3_literal_1076353[p4_res7__192_comb];
  assign p4_array_index_1080180_comb = p3_literal_1076355[p4_array_index_1080087_comb];
  assign p4_res7__197_comb = p3_literal_1076345[p4_res7__196_comb] ^ p3_literal_1076347[p4_res7__195_comb] ^ p4_array_index_1080177_comb ^ p4_array_index_1080178_comb ^ p4_array_index_1080179_comb ^ p4_array_index_1080180_comb ^ p4_array_index_1080088_comb ^ p3_literal_1076358[p4_array_index_1080089_comb] ^ p4_array_index_1080090_comb ^ p4_array_index_1080125_comb ^ p3_literal_1076353[p4_array_index_1080092_comb] ^ p3_literal_1076351[p4_array_index_1080109_comb] ^ p3_literal_1076349[p4_array_index_1080094_comb] ^ p3_literal_1076347[p4_array_index_1080111_comb] ^ p3_literal_1076345[p4_array_index_1080096_comb] ^ p4_array_index_1080097_comb;
  assign p4_array_index_1080191_comb = p3_literal_1076351[p4_res7__194_comb];
  assign p4_array_index_1080192_comb = p3_literal_1076353[p4_res7__193_comb];
  assign p4_array_index_1080193_comb = p3_literal_1076355[p4_res7__192_comb];
  assign p4_res7__198_comb = p3_literal_1076345[p4_res7__197_comb] ^ p3_literal_1076347[p4_res7__196_comb] ^ p3_literal_1076349[p4_res7__195_comb] ^ p4_array_index_1080191_comb ^ p4_array_index_1080192_comb ^ p4_array_index_1080193_comb ^ p4_array_index_1080087_comb ^ p3_literal_1076358[p4_array_index_1080088_comb] ^ p4_array_index_1080089_comb ^ p4_array_index_1080139_comb ^ p4_array_index_1080107_comb ^ p3_literal_1076351[p4_array_index_1080092_comb] ^ p3_literal_1076349[p4_array_index_1080109_comb] ^ p3_literal_1076347[p4_array_index_1080094_comb] ^ p3_literal_1076345[p4_array_index_1080111_comb] ^ p4_array_index_1080096_comb;
  assign p4_array_index_1080203_comb = p3_literal_1076351[p4_res7__195_comb];
  assign p4_array_index_1080204_comb = p3_literal_1076353[p4_res7__194_comb];
  assign p4_array_index_1080205_comb = p3_literal_1076355[p4_res7__193_comb];
  assign p4_res7__199_comb = p3_literal_1076345[p4_res7__198_comb] ^ p3_literal_1076347[p4_res7__197_comb] ^ p3_literal_1076349[p4_res7__196_comb] ^ p4_array_index_1080203_comb ^ p4_array_index_1080204_comb ^ p4_array_index_1080205_comb ^ p4_res7__192_comb ^ p3_literal_1076358[p4_array_index_1080087_comb] ^ p4_array_index_1080088_comb ^ p4_array_index_1080153_comb ^ p4_array_index_1080124_comb ^ p3_literal_1076351[p4_array_index_1080091_comb] ^ p3_literal_1076349[p4_array_index_1080092_comb] ^ p3_literal_1076347[p4_array_index_1080109_comb] ^ p3_literal_1076345[p4_array_index_1080094_comb] ^ p4_array_index_1080111_comb;
  assign p4_array_index_1080216_comb = p3_literal_1076353[p4_res7__195_comb];
  assign p4_array_index_1080217_comb = p3_literal_1076355[p4_res7__194_comb];
  assign p4_res7__200_comb = p3_literal_1076345[p4_res7__199_comb] ^ p3_literal_1076347[p4_res7__198_comb] ^ p3_literal_1076349[p4_res7__197_comb] ^ p3_literal_1076351[p4_res7__196_comb] ^ p4_array_index_1080216_comb ^ p4_array_index_1080217_comb ^ p4_res7__193_comb ^ p3_literal_1076358[p4_res7__192_comb] ^ p4_array_index_1080087_comb ^ p4_array_index_1080167_comb ^ p4_array_index_1080138_comb ^ p4_array_index_1080106_comb ^ p3_literal_1076349[p4_array_index_1080091_comb] ^ p3_literal_1076347[p4_array_index_1080092_comb] ^ p3_literal_1076345[p4_array_index_1080109_comb] ^ p4_array_index_1080094_comb;
  assign p4_array_index_1080227_comb = p3_literal_1076353[p4_res7__196_comb];
  assign p4_array_index_1080228_comb = p3_literal_1076355[p4_res7__195_comb];
  assign p4_res7__201_comb = p3_literal_1076345[p4_res7__200_comb] ^ p3_literal_1076347[p4_res7__199_comb] ^ p3_literal_1076349[p4_res7__198_comb] ^ p3_literal_1076351[p4_res7__197_comb] ^ p4_array_index_1080227_comb ^ p4_array_index_1080228_comb ^ p4_res7__194_comb ^ p3_literal_1076358[p4_res7__193_comb] ^ p4_res7__192_comb ^ p4_array_index_1080180_comb ^ p4_array_index_1080152_comb ^ p4_array_index_1080123_comb ^ p3_literal_1076349[p4_array_index_1080090_comb] ^ p3_literal_1076347[p4_array_index_1080091_comb] ^ p3_literal_1076345[p4_array_index_1080092_comb] ^ p4_array_index_1080109_comb;
  assign p4_array_index_1080239_comb = p3_literal_1076355[p4_res7__196_comb];
  assign p4_res7__202_comb = p3_literal_1076345[p4_res7__201_comb] ^ p3_literal_1076347[p4_res7__200_comb] ^ p3_literal_1076349[p4_res7__199_comb] ^ p3_literal_1076351[p4_res7__198_comb] ^ p3_literal_1076353[p4_res7__197_comb] ^ p4_array_index_1080239_comb ^ p4_res7__195_comb ^ p3_literal_1076358[p4_res7__194_comb] ^ p4_res7__193_comb ^ p4_array_index_1080193_comb ^ p4_array_index_1080166_comb ^ p4_array_index_1080137_comb ^ p4_array_index_1080105_comb ^ p3_literal_1076347[p4_array_index_1080090_comb] ^ p3_literal_1076345[p4_array_index_1080091_comb] ^ p4_array_index_1080092_comb;
  assign p4_array_index_1080249_comb = p3_literal_1076355[p4_res7__197_comb];
  assign p4_res7__203_comb = p3_literal_1076345[p4_res7__202_comb] ^ p3_literal_1076347[p4_res7__201_comb] ^ p3_literal_1076349[p4_res7__200_comb] ^ p3_literal_1076351[p4_res7__199_comb] ^ p3_literal_1076353[p4_res7__198_comb] ^ p4_array_index_1080249_comb ^ p4_res7__196_comb ^ p3_literal_1076358[p4_res7__195_comb] ^ p4_res7__194_comb ^ p4_array_index_1080205_comb ^ p4_array_index_1080179_comb ^ p4_array_index_1080151_comb ^ p4_array_index_1080122_comb ^ p3_literal_1076347[p4_array_index_1080089_comb] ^ p3_literal_1076345[p4_array_index_1080090_comb] ^ p4_array_index_1080091_comb;
  assign p4_res7__204_comb = p3_literal_1076345[p4_res7__203_comb] ^ p3_literal_1076347[p4_res7__202_comb] ^ p3_literal_1076349[p4_res7__201_comb] ^ p3_literal_1076351[p4_res7__200_comb] ^ p3_literal_1076353[p4_res7__199_comb] ^ p3_literal_1076355[p4_res7__198_comb] ^ p4_res7__197_comb ^ p3_literal_1076358[p4_res7__196_comb] ^ p4_res7__195_comb ^ p4_array_index_1080217_comb ^ p4_array_index_1080192_comb ^ p4_array_index_1080165_comb ^ p4_array_index_1080136_comb ^ p4_array_index_1080104_comb ^ p3_literal_1076345[p4_array_index_1080089_comb] ^ p4_array_index_1080090_comb;
  assign p4_res7__205_comb = p3_literal_1076345[p4_res7__204_comb] ^ p3_literal_1076347[p4_res7__203_comb] ^ p3_literal_1076349[p4_res7__202_comb] ^ p3_literal_1076351[p4_res7__201_comb] ^ p3_literal_1076353[p4_res7__200_comb] ^ p3_literal_1076355[p4_res7__199_comb] ^ p4_res7__198_comb ^ p3_literal_1076358[p4_res7__197_comb] ^ p4_res7__196_comb ^ p4_array_index_1080228_comb ^ p4_array_index_1080204_comb ^ p4_array_index_1080178_comb ^ p4_array_index_1080150_comb ^ p4_array_index_1080121_comb ^ p3_literal_1076345[p4_array_index_1080088_comb] ^ p4_array_index_1080089_comb;
  assign p4_res7__206_comb = p3_literal_1076345[p4_res7__205_comb] ^ p3_literal_1076347[p4_res7__204_comb] ^ p3_literal_1076349[p4_res7__203_comb] ^ p3_literal_1076351[p4_res7__202_comb] ^ p3_literal_1076353[p4_res7__201_comb] ^ p3_literal_1076355[p4_res7__200_comb] ^ p4_res7__199_comb ^ p3_literal_1076358[p4_res7__198_comb] ^ p4_res7__197_comb ^ p4_array_index_1080239_comb ^ p4_array_index_1080216_comb ^ p4_array_index_1080191_comb ^ p4_array_index_1080164_comb ^ p4_array_index_1080135_comb ^ p4_array_index_1080103_comb ^ p4_array_index_1080088_comb;
  assign p4_res7__207_comb = p3_literal_1076345[p4_res7__206_comb] ^ p3_literal_1076347[p4_res7__205_comb] ^ p3_literal_1076349[p4_res7__204_comb] ^ p3_literal_1076351[p4_res7__203_comb] ^ p3_literal_1076353[p4_res7__202_comb] ^ p3_literal_1076355[p4_res7__201_comb] ^ p4_res7__200_comb ^ p3_literal_1076358[p4_res7__199_comb] ^ p4_res7__198_comb ^ p4_array_index_1080249_comb ^ p4_array_index_1080227_comb ^ p4_array_index_1080203_comb ^ p4_array_index_1080177_comb ^ p4_array_index_1080149_comb ^ p4_array_index_1080120_comb ^ p4_array_index_1080087_comb;
  assign p4_res__12_comb = {p4_res7__207_comb, p4_res7__206_comb, p4_res7__205_comb, p4_res7__204_comb, p4_res7__203_comb, p4_res7__202_comb, p4_res7__201_comb, p4_res7__200_comb, p4_res7__199_comb, p4_res7__198_comb, p4_res7__197_comb, p4_res7__196_comb, p4_res7__195_comb, p4_res7__194_comb, p4_res7__193_comb, p4_res7__192_comb};
  assign p4_xor_1080289_comb = p4_res__12_comb ^ p3_xor_1079399;
  assign p4_addedKey__54_comb = p4_xor_1080289_comb ^ 128'h5113_c1f9_4d76_899f_a029_a9e0_ac34_d40e;
  assign p4_array_index_1080305_comb = p3_arr[p4_addedKey__54_comb[127:120]];
  assign p4_array_index_1080306_comb = p3_arr[p4_addedKey__54_comb[119:112]];
  assign p4_array_index_1080307_comb = p3_arr[p4_addedKey__54_comb[111:104]];
  assign p4_array_index_1080308_comb = p3_arr[p4_addedKey__54_comb[103:96]];
  assign p4_array_index_1080309_comb = p3_arr[p4_addedKey__54_comb[95:88]];
  assign p4_array_index_1080310_comb = p3_arr[p4_addedKey__54_comb[87:80]];
  assign p4_array_index_1080312_comb = p3_arr[p4_addedKey__54_comb[71:64]];
  assign p4_array_index_1080314_comb = p3_arr[p4_addedKey__54_comb[55:48]];
  assign p4_array_index_1080315_comb = p3_arr[p4_addedKey__54_comb[47:40]];
  assign p4_array_index_1080316_comb = p3_arr[p4_addedKey__54_comb[39:32]];
  assign p4_array_index_1080317_comb = p3_arr[p4_addedKey__54_comb[31:24]];
  assign p4_array_index_1080318_comb = p3_arr[p4_addedKey__54_comb[23:16]];
  assign p4_array_index_1080319_comb = p3_arr[p4_addedKey__54_comb[15:8]];
  assign p4_array_index_1080321_comb = p3_literal_1076345[p4_array_index_1080305_comb];
  assign p4_array_index_1080322_comb = p3_literal_1076347[p4_array_index_1080306_comb];
  assign p4_array_index_1080323_comb = p3_literal_1076349[p4_array_index_1080307_comb];
  assign p4_array_index_1080324_comb = p3_literal_1076351[p4_array_index_1080308_comb];
  assign p4_array_index_1080325_comb = p3_literal_1076353[p4_array_index_1080309_comb];
  assign p4_array_index_1080326_comb = p3_literal_1076355[p4_array_index_1080310_comb];
  assign p4_array_index_1080327_comb = p3_arr[p4_addedKey__54_comb[79:72]];
  assign p4_array_index_1080329_comb = p3_arr[p4_addedKey__54_comb[63:56]];
  assign p4_res7__208_comb = p4_array_index_1080321_comb ^ p4_array_index_1080322_comb ^ p4_array_index_1080323_comb ^ p4_array_index_1080324_comb ^ p4_array_index_1080325_comb ^ p4_array_index_1080326_comb ^ p4_array_index_1080327_comb ^ p3_literal_1076358[p4_array_index_1080312_comb] ^ p4_array_index_1080329_comb ^ p3_literal_1076355[p4_array_index_1080314_comb] ^ p3_literal_1076353[p4_array_index_1080315_comb] ^ p3_literal_1076351[p4_array_index_1080316_comb] ^ p3_literal_1076349[p4_array_index_1080317_comb] ^ p3_literal_1076347[p4_array_index_1080318_comb] ^ p3_literal_1076345[p4_array_index_1080319_comb] ^ p3_arr[p4_addedKey__54_comb[7:0]];
  assign p4_array_index_1080338_comb = p3_literal_1076345[p4_res7__208_comb];
  assign p4_array_index_1080339_comb = p3_literal_1076347[p4_array_index_1080305_comb];
  assign p4_array_index_1080340_comb = p3_literal_1076349[p4_array_index_1080306_comb];
  assign p4_array_index_1080341_comb = p3_literal_1076351[p4_array_index_1080307_comb];
  assign p4_array_index_1080342_comb = p3_literal_1076353[p4_array_index_1080308_comb];
  assign p4_array_index_1080343_comb = p3_literal_1076355[p4_array_index_1080309_comb];
  assign p4_res7__209_comb = p4_array_index_1080338_comb ^ p4_array_index_1080339_comb ^ p4_array_index_1080340_comb ^ p4_array_index_1080341_comb ^ p4_array_index_1080342_comb ^ p4_array_index_1080343_comb ^ p4_array_index_1080310_comb ^ p3_literal_1076358[p4_array_index_1080327_comb] ^ p4_array_index_1080312_comb ^ p3_literal_1076355[p4_array_index_1080329_comb] ^ p3_literal_1076353[p4_array_index_1080314_comb] ^ p3_literal_1076351[p4_array_index_1080315_comb] ^ p3_literal_1076349[p4_array_index_1080316_comb] ^ p3_literal_1076347[p4_array_index_1080317_comb] ^ p3_literal_1076345[p4_array_index_1080318_comb] ^ p4_array_index_1080319_comb;
  assign p4_array_index_1080353_comb = p3_literal_1076347[p4_res7__208_comb];
  assign p4_array_index_1080354_comb = p3_literal_1076349[p4_array_index_1080305_comb];
  assign p4_array_index_1080355_comb = p3_literal_1076351[p4_array_index_1080306_comb];
  assign p4_array_index_1080356_comb = p3_literal_1076353[p4_array_index_1080307_comb];
  assign p4_array_index_1080357_comb = p3_literal_1076355[p4_array_index_1080308_comb];
  assign p4_res7__210_comb = p3_literal_1076345[p4_res7__209_comb] ^ p4_array_index_1080353_comb ^ p4_array_index_1080354_comb ^ p4_array_index_1080355_comb ^ p4_array_index_1080356_comb ^ p4_array_index_1080357_comb ^ p4_array_index_1080309_comb ^ p3_literal_1076358[p4_array_index_1080310_comb] ^ p4_array_index_1080327_comb ^ p3_literal_1076355[p4_array_index_1080312_comb] ^ p3_literal_1076353[p4_array_index_1080329_comb] ^ p3_literal_1076351[p4_array_index_1080314_comb] ^ p3_literal_1076349[p4_array_index_1080315_comb] ^ p3_literal_1076347[p4_array_index_1080316_comb] ^ p3_literal_1076345[p4_array_index_1080317_comb] ^ p4_array_index_1080318_comb;
  assign p4_array_index_1080367_comb = p3_literal_1076347[p4_res7__209_comb];
  assign p4_array_index_1080368_comb = p3_literal_1076349[p4_res7__208_comb];
  assign p4_array_index_1080369_comb = p3_literal_1076351[p4_array_index_1080305_comb];
  assign p4_array_index_1080370_comb = p3_literal_1076353[p4_array_index_1080306_comb];
  assign p4_array_index_1080371_comb = p3_literal_1076355[p4_array_index_1080307_comb];
  assign p4_res7__211_comb = p3_literal_1076345[p4_res7__210_comb] ^ p4_array_index_1080367_comb ^ p4_array_index_1080368_comb ^ p4_array_index_1080369_comb ^ p4_array_index_1080370_comb ^ p4_array_index_1080371_comb ^ p4_array_index_1080308_comb ^ p3_literal_1076358[p4_array_index_1080309_comb] ^ p4_array_index_1080310_comb ^ p3_literal_1076355[p4_array_index_1080327_comb] ^ p3_literal_1076353[p4_array_index_1080312_comb] ^ p3_literal_1076351[p4_array_index_1080329_comb] ^ p3_literal_1076349[p4_array_index_1080314_comb] ^ p3_literal_1076347[p4_array_index_1080315_comb] ^ p3_literal_1076345[p4_array_index_1080316_comb] ^ p4_array_index_1080317_comb;
  assign p4_array_index_1080382_comb = p3_literal_1076349[p4_res7__209_comb];
  assign p4_array_index_1080383_comb = p3_literal_1076351[p4_res7__208_comb];
  assign p4_array_index_1080384_comb = p3_literal_1076353[p4_array_index_1080305_comb];
  assign p4_array_index_1080385_comb = p3_literal_1076355[p4_array_index_1080306_comb];
  assign p4_res7__212_comb = p3_literal_1076345[p4_res7__211_comb] ^ p3_literal_1076347[p4_res7__210_comb] ^ p4_array_index_1080382_comb ^ p4_array_index_1080383_comb ^ p4_array_index_1080384_comb ^ p4_array_index_1080385_comb ^ p4_array_index_1080307_comb ^ p3_literal_1076358[p4_array_index_1080308_comb] ^ p4_array_index_1080309_comb ^ p4_array_index_1080326_comb ^ p3_literal_1076353[p4_array_index_1080327_comb] ^ p3_literal_1076351[p4_array_index_1080312_comb] ^ p3_literal_1076349[p4_array_index_1080329_comb] ^ p3_literal_1076347[p4_array_index_1080314_comb] ^ p3_literal_1076345[p4_array_index_1080315_comb] ^ p4_array_index_1080316_comb;
  assign p4_array_index_1080395_comb = p3_literal_1076349[p4_res7__210_comb];
  assign p4_array_index_1080396_comb = p3_literal_1076351[p4_res7__209_comb];
  assign p4_array_index_1080397_comb = p3_literal_1076353[p4_res7__208_comb];
  assign p4_array_index_1080398_comb = p3_literal_1076355[p4_array_index_1080305_comb];
  assign p4_res7__213_comb = p3_literal_1076345[p4_res7__212_comb] ^ p3_literal_1076347[p4_res7__211_comb] ^ p4_array_index_1080395_comb ^ p4_array_index_1080396_comb ^ p4_array_index_1080397_comb ^ p4_array_index_1080398_comb ^ p4_array_index_1080306_comb ^ p3_literal_1076358[p4_array_index_1080307_comb] ^ p4_array_index_1080308_comb ^ p4_array_index_1080343_comb ^ p3_literal_1076353[p4_array_index_1080310_comb] ^ p3_literal_1076351[p4_array_index_1080327_comb] ^ p3_literal_1076349[p4_array_index_1080312_comb] ^ p3_literal_1076347[p4_array_index_1080329_comb] ^ p3_literal_1076345[p4_array_index_1080314_comb] ^ p4_array_index_1080315_comb;
  assign p4_array_index_1080409_comb = p3_literal_1076351[p4_res7__210_comb];
  assign p4_array_index_1080410_comb = p3_literal_1076353[p4_res7__209_comb];
  assign p4_array_index_1080411_comb = p3_literal_1076355[p4_res7__208_comb];
  assign p4_res7__214_comb = p3_literal_1076345[p4_res7__213_comb] ^ p3_literal_1076347[p4_res7__212_comb] ^ p3_literal_1076349[p4_res7__211_comb] ^ p4_array_index_1080409_comb ^ p4_array_index_1080410_comb ^ p4_array_index_1080411_comb ^ p4_array_index_1080305_comb ^ p3_literal_1076358[p4_array_index_1080306_comb] ^ p4_array_index_1080307_comb ^ p4_array_index_1080357_comb ^ p4_array_index_1080325_comb ^ p3_literal_1076351[p4_array_index_1080310_comb] ^ p3_literal_1076349[p4_array_index_1080327_comb] ^ p3_literal_1076347[p4_array_index_1080312_comb] ^ p3_literal_1076345[p4_array_index_1080329_comb] ^ p4_array_index_1080314_comb;
  assign p4_array_index_1080421_comb = p3_literal_1076351[p4_res7__211_comb];
  assign p4_array_index_1080422_comb = p3_literal_1076353[p4_res7__210_comb];
  assign p4_array_index_1080423_comb = p3_literal_1076355[p4_res7__209_comb];
  assign p4_res7__215_comb = p3_literal_1076345[p4_res7__214_comb] ^ p3_literal_1076347[p4_res7__213_comb] ^ p3_literal_1076349[p4_res7__212_comb] ^ p4_array_index_1080421_comb ^ p4_array_index_1080422_comb ^ p4_array_index_1080423_comb ^ p4_res7__208_comb ^ p3_literal_1076358[p4_array_index_1080305_comb] ^ p4_array_index_1080306_comb ^ p4_array_index_1080371_comb ^ p4_array_index_1080342_comb ^ p3_literal_1076351[p4_array_index_1080309_comb] ^ p3_literal_1076349[p4_array_index_1080310_comb] ^ p3_literal_1076347[p4_array_index_1080327_comb] ^ p3_literal_1076345[p4_array_index_1080312_comb] ^ p4_array_index_1080329_comb;
  assign p4_array_index_1080434_comb = p3_literal_1076353[p4_res7__211_comb];
  assign p4_array_index_1080435_comb = p3_literal_1076355[p4_res7__210_comb];
  assign p4_res7__216_comb = p3_literal_1076345[p4_res7__215_comb] ^ p3_literal_1076347[p4_res7__214_comb] ^ p3_literal_1076349[p4_res7__213_comb] ^ p3_literal_1076351[p4_res7__212_comb] ^ p4_array_index_1080434_comb ^ p4_array_index_1080435_comb ^ p4_res7__209_comb ^ p3_literal_1076358[p4_res7__208_comb] ^ p4_array_index_1080305_comb ^ p4_array_index_1080385_comb ^ p4_array_index_1080356_comb ^ p4_array_index_1080324_comb ^ p3_literal_1076349[p4_array_index_1080309_comb] ^ p3_literal_1076347[p4_array_index_1080310_comb] ^ p3_literal_1076345[p4_array_index_1080327_comb] ^ p4_array_index_1080312_comb;
  assign p4_array_index_1080445_comb = p3_literal_1076353[p4_res7__212_comb];
  assign p4_array_index_1080446_comb = p3_literal_1076355[p4_res7__211_comb];
  assign p4_res7__217_comb = p3_literal_1076345[p4_res7__216_comb] ^ p3_literal_1076347[p4_res7__215_comb] ^ p3_literal_1076349[p4_res7__214_comb] ^ p3_literal_1076351[p4_res7__213_comb] ^ p4_array_index_1080445_comb ^ p4_array_index_1080446_comb ^ p4_res7__210_comb ^ p3_literal_1076358[p4_res7__209_comb] ^ p4_res7__208_comb ^ p4_array_index_1080398_comb ^ p4_array_index_1080370_comb ^ p4_array_index_1080341_comb ^ p3_literal_1076349[p4_array_index_1080308_comb] ^ p3_literal_1076347[p4_array_index_1080309_comb] ^ p3_literal_1076345[p4_array_index_1080310_comb] ^ p4_array_index_1080327_comb;
  assign p4_array_index_1080457_comb = p3_literal_1076355[p4_res7__212_comb];
  assign p4_res7__218_comb = p3_literal_1076345[p4_res7__217_comb] ^ p3_literal_1076347[p4_res7__216_comb] ^ p3_literal_1076349[p4_res7__215_comb] ^ p3_literal_1076351[p4_res7__214_comb] ^ p3_literal_1076353[p4_res7__213_comb] ^ p4_array_index_1080457_comb ^ p4_res7__211_comb ^ p3_literal_1076358[p4_res7__210_comb] ^ p4_res7__209_comb ^ p4_array_index_1080411_comb ^ p4_array_index_1080384_comb ^ p4_array_index_1080355_comb ^ p4_array_index_1080323_comb ^ p3_literal_1076347[p4_array_index_1080308_comb] ^ p3_literal_1076345[p4_array_index_1080309_comb] ^ p4_array_index_1080310_comb;
  assign p4_array_index_1080467_comb = p3_literal_1076355[p4_res7__213_comb];
  assign p4_res7__219_comb = p3_literal_1076345[p4_res7__218_comb] ^ p3_literal_1076347[p4_res7__217_comb] ^ p3_literal_1076349[p4_res7__216_comb] ^ p3_literal_1076351[p4_res7__215_comb] ^ p3_literal_1076353[p4_res7__214_comb] ^ p4_array_index_1080467_comb ^ p4_res7__212_comb ^ p3_literal_1076358[p4_res7__211_comb] ^ p4_res7__210_comb ^ p4_array_index_1080423_comb ^ p4_array_index_1080397_comb ^ p4_array_index_1080369_comb ^ p4_array_index_1080340_comb ^ p3_literal_1076347[p4_array_index_1080307_comb] ^ p3_literal_1076345[p4_array_index_1080308_comb] ^ p4_array_index_1080309_comb;
  assign p4_res7__220_comb = p3_literal_1076345[p4_res7__219_comb] ^ p3_literal_1076347[p4_res7__218_comb] ^ p3_literal_1076349[p4_res7__217_comb] ^ p3_literal_1076351[p4_res7__216_comb] ^ p3_literal_1076353[p4_res7__215_comb] ^ p3_literal_1076355[p4_res7__214_comb] ^ p4_res7__213_comb ^ p3_literal_1076358[p4_res7__212_comb] ^ p4_res7__211_comb ^ p4_array_index_1080435_comb ^ p4_array_index_1080410_comb ^ p4_array_index_1080383_comb ^ p4_array_index_1080354_comb ^ p4_array_index_1080322_comb ^ p3_literal_1076345[p4_array_index_1080307_comb] ^ p4_array_index_1080308_comb;
  assign p4_res7__221_comb = p3_literal_1076345[p4_res7__220_comb] ^ p3_literal_1076347[p4_res7__219_comb] ^ p3_literal_1076349[p4_res7__218_comb] ^ p3_literal_1076351[p4_res7__217_comb] ^ p3_literal_1076353[p4_res7__216_comb] ^ p3_literal_1076355[p4_res7__215_comb] ^ p4_res7__214_comb ^ p3_literal_1076358[p4_res7__213_comb] ^ p4_res7__212_comb ^ p4_array_index_1080446_comb ^ p4_array_index_1080422_comb ^ p4_array_index_1080396_comb ^ p4_array_index_1080368_comb ^ p4_array_index_1080339_comb ^ p3_literal_1076345[p4_array_index_1080306_comb] ^ p4_array_index_1080307_comb;
  assign p4_res7__222_comb = p3_literal_1076345[p4_res7__221_comb] ^ p3_literal_1076347[p4_res7__220_comb] ^ p3_literal_1076349[p4_res7__219_comb] ^ p3_literal_1076351[p4_res7__218_comb] ^ p3_literal_1076353[p4_res7__217_comb] ^ p3_literal_1076355[p4_res7__216_comb] ^ p4_res7__215_comb ^ p3_literal_1076358[p4_res7__214_comb] ^ p4_res7__213_comb ^ p4_array_index_1080457_comb ^ p4_array_index_1080434_comb ^ p4_array_index_1080409_comb ^ p4_array_index_1080382_comb ^ p4_array_index_1080353_comb ^ p4_array_index_1080321_comb ^ p4_array_index_1080306_comb;
  assign p4_res7__223_comb = p3_literal_1076345[p4_res7__222_comb] ^ p3_literal_1076347[p4_res7__221_comb] ^ p3_literal_1076349[p4_res7__220_comb] ^ p3_literal_1076351[p4_res7__219_comb] ^ p3_literal_1076353[p4_res7__218_comb] ^ p3_literal_1076355[p4_res7__217_comb] ^ p4_res7__216_comb ^ p3_literal_1076358[p4_res7__215_comb] ^ p4_res7__214_comb ^ p4_array_index_1080467_comb ^ p4_array_index_1080445_comb ^ p4_array_index_1080421_comb ^ p4_array_index_1080395_comb ^ p4_array_index_1080367_comb ^ p4_array_index_1080338_comb ^ p4_array_index_1080305_comb;
  assign p4_res__13_comb = {p4_res7__223_comb, p4_res7__222_comb, p4_res7__221_comb, p4_res7__220_comb, p4_res7__219_comb, p4_res7__218_comb, p4_res7__217_comb, p4_res7__216_comb, p4_res7__215_comb, p4_res7__214_comb, p4_res7__213_comb, p4_res7__212_comb, p4_res7__211_comb, p4_res7__210_comb, p4_res7__209_comb, p4_res7__208_comb};
  assign p4_xor_1080507_comb = p4_res__13_comb ^ p4_xor_1080071_comb;
  assign p4_addedKey__55_comb = p4_xor_1080507_comb ^ 128'h3fb1_b78b_213e_f327_fd0e_14f0_71b0_400f;
  assign p4_array_index_1080523_comb = p3_arr[p4_addedKey__55_comb[127:120]];
  assign p4_array_index_1080524_comb = p3_arr[p4_addedKey__55_comb[119:112]];
  assign p4_array_index_1080525_comb = p3_arr[p4_addedKey__55_comb[111:104]];
  assign p4_array_index_1080526_comb = p3_arr[p4_addedKey__55_comb[103:96]];
  assign p4_array_index_1080527_comb = p3_arr[p4_addedKey__55_comb[95:88]];
  assign p4_array_index_1080528_comb = p3_arr[p4_addedKey__55_comb[87:80]];
  assign p4_array_index_1080530_comb = p3_arr[p4_addedKey__55_comb[71:64]];
  assign p4_array_index_1080532_comb = p3_arr[p4_addedKey__55_comb[55:48]];
  assign p4_array_index_1080533_comb = p3_arr[p4_addedKey__55_comb[47:40]];
  assign p4_array_index_1080534_comb = p3_arr[p4_addedKey__55_comb[39:32]];
  assign p4_array_index_1080535_comb = p3_arr[p4_addedKey__55_comb[31:24]];
  assign p4_array_index_1080536_comb = p3_arr[p4_addedKey__55_comb[23:16]];
  assign p4_array_index_1080537_comb = p3_arr[p4_addedKey__55_comb[15:8]];
  assign p4_array_index_1080539_comb = p3_literal_1076345[p4_array_index_1080523_comb];
  assign p4_array_index_1080540_comb = p3_literal_1076347[p4_array_index_1080524_comb];
  assign p4_array_index_1080541_comb = p3_literal_1076349[p4_array_index_1080525_comb];
  assign p4_array_index_1080542_comb = p3_literal_1076351[p4_array_index_1080526_comb];
  assign p4_array_index_1080543_comb = p3_literal_1076353[p4_array_index_1080527_comb];
  assign p4_array_index_1080544_comb = p3_literal_1076355[p4_array_index_1080528_comb];
  assign p4_array_index_1080545_comb = p3_arr[p4_addedKey__55_comb[79:72]];
  assign p4_array_index_1080547_comb = p3_arr[p4_addedKey__55_comb[63:56]];
  assign p4_res7__224_comb = p4_array_index_1080539_comb ^ p4_array_index_1080540_comb ^ p4_array_index_1080541_comb ^ p4_array_index_1080542_comb ^ p4_array_index_1080543_comb ^ p4_array_index_1080544_comb ^ p4_array_index_1080545_comb ^ p3_literal_1076358[p4_array_index_1080530_comb] ^ p4_array_index_1080547_comb ^ p3_literal_1076355[p4_array_index_1080532_comb] ^ p3_literal_1076353[p4_array_index_1080533_comb] ^ p3_literal_1076351[p4_array_index_1080534_comb] ^ p3_literal_1076349[p4_array_index_1080535_comb] ^ p3_literal_1076347[p4_array_index_1080536_comb] ^ p3_literal_1076345[p4_array_index_1080537_comb] ^ p3_arr[p4_addedKey__55_comb[7:0]];
  assign p4_array_index_1080556_comb = p3_literal_1076345[p4_res7__224_comb];
  assign p4_array_index_1080557_comb = p3_literal_1076347[p4_array_index_1080523_comb];
  assign p4_array_index_1080558_comb = p3_literal_1076349[p4_array_index_1080524_comb];
  assign p4_array_index_1080559_comb = p3_literal_1076351[p4_array_index_1080525_comb];
  assign p4_array_index_1080560_comb = p3_literal_1076353[p4_array_index_1080526_comb];
  assign p4_array_index_1080561_comb = p3_literal_1076355[p4_array_index_1080527_comb];
  assign p4_res7__225_comb = p4_array_index_1080556_comb ^ p4_array_index_1080557_comb ^ p4_array_index_1080558_comb ^ p4_array_index_1080559_comb ^ p4_array_index_1080560_comb ^ p4_array_index_1080561_comb ^ p4_array_index_1080528_comb ^ p3_literal_1076358[p4_array_index_1080545_comb] ^ p4_array_index_1080530_comb ^ p3_literal_1076355[p4_array_index_1080547_comb] ^ p3_literal_1076353[p4_array_index_1080532_comb] ^ p3_literal_1076351[p4_array_index_1080533_comb] ^ p3_literal_1076349[p4_array_index_1080534_comb] ^ p3_literal_1076347[p4_array_index_1080535_comb] ^ p3_literal_1076345[p4_array_index_1080536_comb] ^ p4_array_index_1080537_comb;
  assign p4_array_index_1080571_comb = p3_literal_1076347[p4_res7__224_comb];
  assign p4_array_index_1080572_comb = p3_literal_1076349[p4_array_index_1080523_comb];
  assign p4_array_index_1080573_comb = p3_literal_1076351[p4_array_index_1080524_comb];
  assign p4_array_index_1080574_comb = p3_literal_1076353[p4_array_index_1080525_comb];
  assign p4_array_index_1080575_comb = p3_literal_1076355[p4_array_index_1080526_comb];
  assign p4_res7__226_comb = p3_literal_1076345[p4_res7__225_comb] ^ p4_array_index_1080571_comb ^ p4_array_index_1080572_comb ^ p4_array_index_1080573_comb ^ p4_array_index_1080574_comb ^ p4_array_index_1080575_comb ^ p4_array_index_1080527_comb ^ p3_literal_1076358[p4_array_index_1080528_comb] ^ p4_array_index_1080545_comb ^ p3_literal_1076355[p4_array_index_1080530_comb] ^ p3_literal_1076353[p4_array_index_1080547_comb] ^ p3_literal_1076351[p4_array_index_1080532_comb] ^ p3_literal_1076349[p4_array_index_1080533_comb] ^ p3_literal_1076347[p4_array_index_1080534_comb] ^ p3_literal_1076345[p4_array_index_1080535_comb] ^ p4_array_index_1080536_comb;
  assign p4_array_index_1080585_comb = p3_literal_1076347[p4_res7__225_comb];
  assign p4_array_index_1080586_comb = p3_literal_1076349[p4_res7__224_comb];
  assign p4_array_index_1080587_comb = p3_literal_1076351[p4_array_index_1080523_comb];
  assign p4_array_index_1080588_comb = p3_literal_1076353[p4_array_index_1080524_comb];
  assign p4_array_index_1080589_comb = p3_literal_1076355[p4_array_index_1080525_comb];
  assign p4_res7__227_comb = p3_literal_1076345[p4_res7__226_comb] ^ p4_array_index_1080585_comb ^ p4_array_index_1080586_comb ^ p4_array_index_1080587_comb ^ p4_array_index_1080588_comb ^ p4_array_index_1080589_comb ^ p4_array_index_1080526_comb ^ p3_literal_1076358[p4_array_index_1080527_comb] ^ p4_array_index_1080528_comb ^ p3_literal_1076355[p4_array_index_1080545_comb] ^ p3_literal_1076353[p4_array_index_1080530_comb] ^ p3_literal_1076351[p4_array_index_1080547_comb] ^ p3_literal_1076349[p4_array_index_1080532_comb] ^ p3_literal_1076347[p4_array_index_1080533_comb] ^ p3_literal_1076345[p4_array_index_1080534_comb] ^ p4_array_index_1080535_comb;
  assign p4_array_index_1080600_comb = p3_literal_1076349[p4_res7__225_comb];
  assign p4_array_index_1080601_comb = p3_literal_1076351[p4_res7__224_comb];
  assign p4_array_index_1080602_comb = p3_literal_1076353[p4_array_index_1080523_comb];
  assign p4_array_index_1080603_comb = p3_literal_1076355[p4_array_index_1080524_comb];
  assign p4_res7__228_comb = p3_literal_1076345[p4_res7__227_comb] ^ p3_literal_1076347[p4_res7__226_comb] ^ p4_array_index_1080600_comb ^ p4_array_index_1080601_comb ^ p4_array_index_1080602_comb ^ p4_array_index_1080603_comb ^ p4_array_index_1080525_comb ^ p3_literal_1076358[p4_array_index_1080526_comb] ^ p4_array_index_1080527_comb ^ p4_array_index_1080544_comb ^ p3_literal_1076353[p4_array_index_1080545_comb] ^ p3_literal_1076351[p4_array_index_1080530_comb] ^ p3_literal_1076349[p4_array_index_1080547_comb] ^ p3_literal_1076347[p4_array_index_1080532_comb] ^ p3_literal_1076345[p4_array_index_1080533_comb] ^ p4_array_index_1080534_comb;
  assign p4_array_index_1080613_comb = p3_literal_1076349[p4_res7__226_comb];
  assign p4_array_index_1080614_comb = p3_literal_1076351[p4_res7__225_comb];
  assign p4_array_index_1080615_comb = p3_literal_1076353[p4_res7__224_comb];
  assign p4_array_index_1080616_comb = p3_literal_1076355[p4_array_index_1080523_comb];
  assign p4_res7__229_comb = p3_literal_1076345[p4_res7__228_comb] ^ p3_literal_1076347[p4_res7__227_comb] ^ p4_array_index_1080613_comb ^ p4_array_index_1080614_comb ^ p4_array_index_1080615_comb ^ p4_array_index_1080616_comb ^ p4_array_index_1080524_comb ^ p3_literal_1076358[p4_array_index_1080525_comb] ^ p4_array_index_1080526_comb ^ p4_array_index_1080561_comb ^ p3_literal_1076353[p4_array_index_1080528_comb] ^ p3_literal_1076351[p4_array_index_1080545_comb] ^ p3_literal_1076349[p4_array_index_1080530_comb] ^ p3_literal_1076347[p4_array_index_1080547_comb] ^ p3_literal_1076345[p4_array_index_1080532_comb] ^ p4_array_index_1080533_comb;
  assign p4_array_index_1080627_comb = p3_literal_1076351[p4_res7__226_comb];
  assign p4_array_index_1080628_comb = p3_literal_1076353[p4_res7__225_comb];
  assign p4_array_index_1080629_comb = p3_literal_1076355[p4_res7__224_comb];
  assign p4_res7__230_comb = p3_literal_1076345[p4_res7__229_comb] ^ p3_literal_1076347[p4_res7__228_comb] ^ p3_literal_1076349[p4_res7__227_comb] ^ p4_array_index_1080627_comb ^ p4_array_index_1080628_comb ^ p4_array_index_1080629_comb ^ p4_array_index_1080523_comb ^ p3_literal_1076358[p4_array_index_1080524_comb] ^ p4_array_index_1080525_comb ^ p4_array_index_1080575_comb ^ p4_array_index_1080543_comb ^ p3_literal_1076351[p4_array_index_1080528_comb] ^ p3_literal_1076349[p4_array_index_1080545_comb] ^ p3_literal_1076347[p4_array_index_1080530_comb] ^ p3_literal_1076345[p4_array_index_1080547_comb] ^ p4_array_index_1080532_comb;
  assign p4_array_index_1080639_comb = p3_literal_1076351[p4_res7__227_comb];
  assign p4_array_index_1080640_comb = p3_literal_1076353[p4_res7__226_comb];
  assign p4_array_index_1080641_comb = p3_literal_1076355[p4_res7__225_comb];
  assign p4_res7__231_comb = p3_literal_1076345[p4_res7__230_comb] ^ p3_literal_1076347[p4_res7__229_comb] ^ p3_literal_1076349[p4_res7__228_comb] ^ p4_array_index_1080639_comb ^ p4_array_index_1080640_comb ^ p4_array_index_1080641_comb ^ p4_res7__224_comb ^ p3_literal_1076358[p4_array_index_1080523_comb] ^ p4_array_index_1080524_comb ^ p4_array_index_1080589_comb ^ p4_array_index_1080560_comb ^ p3_literal_1076351[p4_array_index_1080527_comb] ^ p3_literal_1076349[p4_array_index_1080528_comb] ^ p3_literal_1076347[p4_array_index_1080545_comb] ^ p3_literal_1076345[p4_array_index_1080530_comb] ^ p4_array_index_1080547_comb;
  assign p4_array_index_1080652_comb = p3_literal_1076353[p4_res7__227_comb];
  assign p4_array_index_1080653_comb = p3_literal_1076355[p4_res7__226_comb];
  assign p4_res7__232_comb = p3_literal_1076345[p4_res7__231_comb] ^ p3_literal_1076347[p4_res7__230_comb] ^ p3_literal_1076349[p4_res7__229_comb] ^ p3_literal_1076351[p4_res7__228_comb] ^ p4_array_index_1080652_comb ^ p4_array_index_1080653_comb ^ p4_res7__225_comb ^ p3_literal_1076358[p4_res7__224_comb] ^ p4_array_index_1080523_comb ^ p4_array_index_1080603_comb ^ p4_array_index_1080574_comb ^ p4_array_index_1080542_comb ^ p3_literal_1076349[p4_array_index_1080527_comb] ^ p3_literal_1076347[p4_array_index_1080528_comb] ^ p3_literal_1076345[p4_array_index_1080545_comb] ^ p4_array_index_1080530_comb;
  assign p4_array_index_1080663_comb = p3_literal_1076353[p4_res7__228_comb];
  assign p4_array_index_1080664_comb = p3_literal_1076355[p4_res7__227_comb];
  assign p4_res7__233_comb = p3_literal_1076345[p4_res7__232_comb] ^ p3_literal_1076347[p4_res7__231_comb] ^ p3_literal_1076349[p4_res7__230_comb] ^ p3_literal_1076351[p4_res7__229_comb] ^ p4_array_index_1080663_comb ^ p4_array_index_1080664_comb ^ p4_res7__226_comb ^ p3_literal_1076358[p4_res7__225_comb] ^ p4_res7__224_comb ^ p4_array_index_1080616_comb ^ p4_array_index_1080588_comb ^ p4_array_index_1080559_comb ^ p3_literal_1076349[p4_array_index_1080526_comb] ^ p3_literal_1076347[p4_array_index_1080527_comb] ^ p3_literal_1076345[p4_array_index_1080528_comb] ^ p4_array_index_1080545_comb;
  assign p4_array_index_1080670_comb = p3_literal_1076345[p4_res7__233_comb];
  assign p4_array_index_1080671_comb = p3_literal_1076347[p4_res7__232_comb];
  assign p4_array_index_1080672_comb = p3_literal_1076349[p4_res7__231_comb];
  assign p4_array_index_1080673_comb = p3_literal_1076351[p4_res7__230_comb];
  assign p4_array_index_1080674_comb = p3_literal_1076353[p4_res7__229_comb];
  assign p4_array_index_1080675_comb = p3_literal_1076355[p4_res7__228_comb];
  assign p4_array_index_1080676_comb = p3_literal_1076358[p4_res7__226_comb];
  assign p4_array_index_1080677_comb = p3_literal_1076347[p4_array_index_1080526_comb];
  assign p4_array_index_1080678_comb = p3_literal_1076345[p4_array_index_1080527_comb];

  // Registers for pipe stage 4:
  reg [127:0] p4_xor_1080289;
  reg [127:0] p4_xor_1080507;
  reg [7:0] p4_array_index_1080523;
  reg [7:0] p4_array_index_1080524;
  reg [7:0] p4_array_index_1080525;
  reg [7:0] p4_array_index_1080526;
  reg [7:0] p4_array_index_1080527;
  reg [7:0] p4_array_index_1080528;
  reg [7:0] p4_array_index_1080539;
  reg [7:0] p4_array_index_1080540;
  reg [7:0] p4_array_index_1080541;
  reg [7:0] p4_res7__224;
  reg [7:0] p4_array_index_1080556;
  reg [7:0] p4_array_index_1080557;
  reg [7:0] p4_array_index_1080558;
  reg [7:0] p4_res7__225;
  reg [7:0] p4_array_index_1080571;
  reg [7:0] p4_array_index_1080572;
  reg [7:0] p4_array_index_1080573;
  reg [7:0] p4_res7__226;
  reg [7:0] p4_array_index_1080585;
  reg [7:0] p4_array_index_1080586;
  reg [7:0] p4_array_index_1080587;
  reg [7:0] p4_res7__227;
  reg [7:0] p4_array_index_1080600;
  reg [7:0] p4_array_index_1080601;
  reg [7:0] p4_array_index_1080602;
  reg [7:0] p4_res7__228;
  reg [7:0] p4_array_index_1080613;
  reg [7:0] p4_array_index_1080614;
  reg [7:0] p4_array_index_1080615;
  reg [7:0] p4_res7__229;
  reg [7:0] p4_array_index_1080627;
  reg [7:0] p4_array_index_1080628;
  reg [7:0] p4_array_index_1080629;
  reg [7:0] p4_res7__230;
  reg [7:0] p4_array_index_1080639;
  reg [7:0] p4_array_index_1080640;
  reg [7:0] p4_array_index_1080641;
  reg [7:0] p4_res7__231;
  reg [7:0] p4_array_index_1080652;
  reg [7:0] p4_array_index_1080653;
  reg [7:0] p4_res7__232;
  reg [7:0] p4_array_index_1080663;
  reg [7:0] p4_array_index_1080664;
  reg [7:0] p4_res7__233;
  reg [7:0] p4_array_index_1080670;
  reg [7:0] p4_array_index_1080671;
  reg [7:0] p4_array_index_1080672;
  reg [7:0] p4_array_index_1080673;
  reg [7:0] p4_array_index_1080674;
  reg [7:0] p4_array_index_1080675;
  reg [7:0] p4_array_index_1080676;
  reg [7:0] p4_array_index_1080677;
  reg [7:0] p4_array_index_1080678;
  reg [127:0] p4_res__35;
  reg [7:0] p5_arr[256];
  reg [7:0] p5_literal_1076345[256];
  reg [7:0] p5_literal_1076347[256];
  reg [7:0] p5_literal_1076349[256];
  reg [7:0] p5_literal_1076351[256];
  reg [7:0] p5_literal_1076353[256];
  reg [7:0] p5_literal_1076355[256];
  reg [7:0] p5_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p4_xor_1080289 <= p4_xor_1080289_comb;
    p4_xor_1080507 <= p4_xor_1080507_comb;
    p4_array_index_1080523 <= p4_array_index_1080523_comb;
    p4_array_index_1080524 <= p4_array_index_1080524_comb;
    p4_array_index_1080525 <= p4_array_index_1080525_comb;
    p4_array_index_1080526 <= p4_array_index_1080526_comb;
    p4_array_index_1080527 <= p4_array_index_1080527_comb;
    p4_array_index_1080528 <= p4_array_index_1080528_comb;
    p4_array_index_1080539 <= p4_array_index_1080539_comb;
    p4_array_index_1080540 <= p4_array_index_1080540_comb;
    p4_array_index_1080541 <= p4_array_index_1080541_comb;
    p4_res7__224 <= p4_res7__224_comb;
    p4_array_index_1080556 <= p4_array_index_1080556_comb;
    p4_array_index_1080557 <= p4_array_index_1080557_comb;
    p4_array_index_1080558 <= p4_array_index_1080558_comb;
    p4_res7__225 <= p4_res7__225_comb;
    p4_array_index_1080571 <= p4_array_index_1080571_comb;
    p4_array_index_1080572 <= p4_array_index_1080572_comb;
    p4_array_index_1080573 <= p4_array_index_1080573_comb;
    p4_res7__226 <= p4_res7__226_comb;
    p4_array_index_1080585 <= p4_array_index_1080585_comb;
    p4_array_index_1080586 <= p4_array_index_1080586_comb;
    p4_array_index_1080587 <= p4_array_index_1080587_comb;
    p4_res7__227 <= p4_res7__227_comb;
    p4_array_index_1080600 <= p4_array_index_1080600_comb;
    p4_array_index_1080601 <= p4_array_index_1080601_comb;
    p4_array_index_1080602 <= p4_array_index_1080602_comb;
    p4_res7__228 <= p4_res7__228_comb;
    p4_array_index_1080613 <= p4_array_index_1080613_comb;
    p4_array_index_1080614 <= p4_array_index_1080614_comb;
    p4_array_index_1080615 <= p4_array_index_1080615_comb;
    p4_res7__229 <= p4_res7__229_comb;
    p4_array_index_1080627 <= p4_array_index_1080627_comb;
    p4_array_index_1080628 <= p4_array_index_1080628_comb;
    p4_array_index_1080629 <= p4_array_index_1080629_comb;
    p4_res7__230 <= p4_res7__230_comb;
    p4_array_index_1080639 <= p4_array_index_1080639_comb;
    p4_array_index_1080640 <= p4_array_index_1080640_comb;
    p4_array_index_1080641 <= p4_array_index_1080641_comb;
    p4_res7__231 <= p4_res7__231_comb;
    p4_array_index_1080652 <= p4_array_index_1080652_comb;
    p4_array_index_1080653 <= p4_array_index_1080653_comb;
    p4_res7__232 <= p4_res7__232_comb;
    p4_array_index_1080663 <= p4_array_index_1080663_comb;
    p4_array_index_1080664 <= p4_array_index_1080664_comb;
    p4_res7__233 <= p4_res7__233_comb;
    p4_array_index_1080670 <= p4_array_index_1080670_comb;
    p4_array_index_1080671 <= p4_array_index_1080671_comb;
    p4_array_index_1080672 <= p4_array_index_1080672_comb;
    p4_array_index_1080673 <= p4_array_index_1080673_comb;
    p4_array_index_1080674 <= p4_array_index_1080674_comb;
    p4_array_index_1080675 <= p4_array_index_1080675_comb;
    p4_array_index_1080676 <= p4_array_index_1080676_comb;
    p4_array_index_1080677 <= p4_array_index_1080677_comb;
    p4_array_index_1080678 <= p4_array_index_1080678_comb;
    p4_res__35 <= p3_res__35;
    p5_arr <= p4_arr;
    p5_literal_1076345 <= p4_literal_1076345;
    p5_literal_1076347 <= p4_literal_1076347;
    p5_literal_1076349 <= p4_literal_1076349;
    p5_literal_1076351 <= p4_literal_1076351;
    p5_literal_1076353 <= p4_literal_1076353;
    p5_literal_1076355 <= p4_literal_1076355;
    p5_literal_1076358 <= p4_literal_1076358;
  end

  // ===== Pipe stage 5:
  wire [7:0] p5_res7__234_comb;
  wire [7:0] p5_array_index_1080813_comb;
  wire [7:0] p5_res7__235_comb;
  wire [7:0] p5_res7__236_comb;
  wire [7:0] p5_res7__237_comb;
  wire [7:0] p5_res7__238_comb;
  wire [7:0] p5_res7__239_comb;
  wire [127:0] p5_res__14_comb;
  wire [127:0] p5_k5_comb;
  wire [127:0] p5_addedKey__56_comb;
  wire [7:0] p5_array_index_1080869_comb;
  wire [7:0] p5_array_index_1080870_comb;
  wire [7:0] p5_array_index_1080871_comb;
  wire [7:0] p5_array_index_1080872_comb;
  wire [7:0] p5_array_index_1080873_comb;
  wire [7:0] p5_array_index_1080874_comb;
  wire [7:0] p5_array_index_1080876_comb;
  wire [7:0] p5_array_index_1080878_comb;
  wire [7:0] p5_array_index_1080879_comb;
  wire [7:0] p5_array_index_1080880_comb;
  wire [7:0] p5_array_index_1080881_comb;
  wire [7:0] p5_array_index_1080882_comb;
  wire [7:0] p5_array_index_1080883_comb;
  wire [7:0] p5_array_index_1080885_comb;
  wire [7:0] p5_array_index_1080886_comb;
  wire [7:0] p5_array_index_1080887_comb;
  wire [7:0] p5_array_index_1080888_comb;
  wire [7:0] p5_array_index_1080889_comb;
  wire [7:0] p5_array_index_1080890_comb;
  wire [7:0] p5_array_index_1080891_comb;
  wire [7:0] p5_array_index_1080893_comb;
  wire [7:0] p5_res7__240_comb;
  wire [7:0] p5_array_index_1080902_comb;
  wire [7:0] p5_array_index_1080903_comb;
  wire [7:0] p5_array_index_1080904_comb;
  wire [7:0] p5_array_index_1080905_comb;
  wire [7:0] p5_array_index_1080906_comb;
  wire [7:0] p5_array_index_1080907_comb;
  wire [7:0] p5_res7__241_comb;
  wire [7:0] p5_array_index_1080917_comb;
  wire [7:0] p5_array_index_1080918_comb;
  wire [7:0] p5_array_index_1080919_comb;
  wire [7:0] p5_array_index_1080920_comb;
  wire [7:0] p5_array_index_1080921_comb;
  wire [7:0] p5_res7__242_comb;
  wire [7:0] p5_array_index_1080931_comb;
  wire [7:0] p5_array_index_1080932_comb;
  wire [7:0] p5_array_index_1080933_comb;
  wire [7:0] p5_array_index_1080934_comb;
  wire [7:0] p5_array_index_1080935_comb;
  wire [7:0] p5_res7__243_comb;
  wire [7:0] p5_array_index_1080946_comb;
  wire [7:0] p5_array_index_1080947_comb;
  wire [7:0] p5_array_index_1080948_comb;
  wire [7:0] p5_array_index_1080949_comb;
  wire [7:0] p5_res7__244_comb;
  wire [7:0] p5_array_index_1080959_comb;
  wire [7:0] p5_array_index_1080960_comb;
  wire [7:0] p5_array_index_1080961_comb;
  wire [7:0] p5_array_index_1080962_comb;
  wire [7:0] p5_res7__245_comb;
  wire [7:0] p5_array_index_1080973_comb;
  wire [7:0] p5_array_index_1080974_comb;
  wire [7:0] p5_array_index_1080975_comb;
  wire [7:0] p5_res7__246_comb;
  wire [7:0] p5_array_index_1080985_comb;
  wire [7:0] p5_array_index_1080986_comb;
  wire [7:0] p5_array_index_1080987_comb;
  wire [7:0] p5_res7__247_comb;
  wire [7:0] p5_array_index_1080998_comb;
  wire [7:0] p5_array_index_1080999_comb;
  wire [7:0] p5_res7__248_comb;
  wire [7:0] p5_array_index_1081009_comb;
  wire [7:0] p5_array_index_1081010_comb;
  wire [7:0] p5_res7__249_comb;
  wire [7:0] p5_array_index_1081021_comb;
  wire [7:0] p5_res7__250_comb;
  wire [7:0] p5_array_index_1081031_comb;
  wire [7:0] p5_res7__251_comb;
  wire [7:0] p5_res7__252_comb;
  wire [7:0] p5_res7__253_comb;
  wire [7:0] p5_res7__254_comb;
  wire [7:0] p5_res7__255_comb;
  wire [127:0] p5_res__15_comb;
  wire [127:0] p5_k4_comb;
  wire [127:0] p5_addedKey__57_comb;
  wire [7:0] p5_array_index_1081087_comb;
  wire [7:0] p5_array_index_1081088_comb;
  wire [7:0] p5_array_index_1081089_comb;
  wire [7:0] p5_array_index_1081090_comb;
  wire [7:0] p5_array_index_1081091_comb;
  wire [7:0] p5_array_index_1081092_comb;
  wire [7:0] p5_array_index_1081094_comb;
  wire [7:0] p5_array_index_1081096_comb;
  wire [7:0] p5_array_index_1081097_comb;
  wire [7:0] p5_array_index_1081098_comb;
  wire [7:0] p5_array_index_1081099_comb;
  wire [7:0] p5_array_index_1081100_comb;
  wire [7:0] p5_array_index_1081101_comb;
  wire [7:0] p5_array_index_1081103_comb;
  wire [7:0] p5_array_index_1081104_comb;
  wire [7:0] p5_array_index_1081105_comb;
  wire [7:0] p5_array_index_1081106_comb;
  wire [7:0] p5_array_index_1081107_comb;
  wire [7:0] p5_array_index_1081108_comb;
  wire [7:0] p5_array_index_1081109_comb;
  wire [7:0] p5_array_index_1081111_comb;
  wire [7:0] p5_res7__256_comb;
  wire [7:0] p5_array_index_1081120_comb;
  wire [7:0] p5_array_index_1081121_comb;
  wire [7:0] p5_array_index_1081122_comb;
  wire [7:0] p5_array_index_1081123_comb;
  wire [7:0] p5_array_index_1081124_comb;
  wire [7:0] p5_array_index_1081125_comb;
  wire [7:0] p5_res7__257_comb;
  wire [7:0] p5_array_index_1081135_comb;
  wire [7:0] p5_array_index_1081136_comb;
  wire [7:0] p5_array_index_1081137_comb;
  wire [7:0] p5_array_index_1081138_comb;
  wire [7:0] p5_array_index_1081139_comb;
  wire [7:0] p5_res7__258_comb;
  wire [7:0] p5_array_index_1081149_comb;
  wire [7:0] p5_array_index_1081150_comb;
  wire [7:0] p5_array_index_1081151_comb;
  wire [7:0] p5_array_index_1081152_comb;
  wire [7:0] p5_array_index_1081153_comb;
  wire [7:0] p5_res7__259_comb;
  wire [7:0] p5_array_index_1081164_comb;
  wire [7:0] p5_array_index_1081165_comb;
  wire [7:0] p5_array_index_1081166_comb;
  wire [7:0] p5_array_index_1081167_comb;
  wire [7:0] p5_res7__260_comb;
  wire [7:0] p5_array_index_1081177_comb;
  wire [7:0] p5_array_index_1081178_comb;
  wire [7:0] p5_array_index_1081179_comb;
  wire [7:0] p5_array_index_1081180_comb;
  wire [7:0] p5_res7__261_comb;
  wire [7:0] p5_array_index_1081191_comb;
  wire [7:0] p5_array_index_1081192_comb;
  wire [7:0] p5_array_index_1081193_comb;
  wire [127:0] p5_addedKey__36_comb;
  wire [7:0] p5_res7__262_comb;
  wire [7:0] p5_array_index_1081203_comb;
  wire [7:0] p5_array_index_1081204_comb;
  wire [7:0] p5_array_index_1081205_comb;
  wire [7:0] p5_array_index_1081625_comb;
  wire [7:0] p5_array_index_1081626_comb;
  wire [7:0] p5_array_index_1081627_comb;
  wire [7:0] p5_array_index_1081628_comb;
  wire [7:0] p5_array_index_1081629_comb;
  wire [7:0] p5_array_index_1081630_comb;
  wire [7:0] p5_array_index_1081632_comb;
  wire [7:0] p5_array_index_1081634_comb;
  wire [7:0] p5_array_index_1081635_comb;
  wire [7:0] p5_array_index_1081636_comb;
  wire [7:0] p5_array_index_1081637_comb;
  wire [7:0] p5_array_index_1081638_comb;
  wire [7:0] p5_array_index_1081639_comb;
  wire [7:0] p5_res7__263_comb;
  wire [7:0] p5_array_index_1081641_comb;
  wire [7:0] p5_array_index_1081642_comb;
  wire [7:0] p5_array_index_1081643_comb;
  wire [7:0] p5_array_index_1081644_comb;
  wire [7:0] p5_array_index_1081645_comb;
  wire [7:0] p5_array_index_1081646_comb;
  wire [7:0] p5_array_index_1081647_comb;
  wire [7:0] p5_array_index_1081649_comb;
  wire [7:0] p5_array_index_1081216_comb;
  wire [7:0] p5_array_index_1081217_comb;
  wire [7:0] p5_res7__576_comb;
  wire [7:0] p5_res7__264_comb;
  wire [7:0] p5_array_index_1081658_comb;
  wire [7:0] p5_array_index_1081659_comb;
  wire [7:0] p5_array_index_1081660_comb;
  wire [7:0] p5_array_index_1081661_comb;
  wire [7:0] p5_array_index_1081662_comb;
  wire [7:0] p5_array_index_1081663_comb;
  wire [7:0] p5_array_index_1081227_comb;
  wire [7:0] p5_array_index_1081228_comb;
  wire [7:0] p5_res7__577_comb;
  wire [7:0] p5_res7__265_comb;
  wire [7:0] p5_array_index_1081673_comb;
  wire [7:0] p5_array_index_1081674_comb;
  wire [7:0] p5_array_index_1081675_comb;
  wire [7:0] p5_array_index_1081676_comb;
  wire [7:0] p5_array_index_1081677_comb;
  wire [7:0] p5_array_index_1081239_comb;
  wire [7:0] p5_res7__578_comb;
  wire [7:0] p5_res7__266_comb;
  wire [7:0] p5_array_index_1081687_comb;
  wire [7:0] p5_array_index_1081688_comb;
  wire [7:0] p5_array_index_1081689_comb;
  wire [7:0] p5_array_index_1081690_comb;
  wire [7:0] p5_array_index_1081691_comb;
  wire [7:0] p5_array_index_1081249_comb;
  wire [7:0] p5_res7__579_comb;
  wire [7:0] p5_res7__267_comb;
  wire [7:0] p5_array_index_1081702_comb;
  wire [7:0] p5_array_index_1081703_comb;
  wire [7:0] p5_array_index_1081704_comb;
  wire [7:0] p5_array_index_1081705_comb;
  wire [7:0] p5_res7__580_comb;
  wire [7:0] p5_res7__268_comb;
  wire [7:0] p5_array_index_1081715_comb;
  wire [7:0] p5_array_index_1081716_comb;
  wire [7:0] p5_array_index_1081717_comb;
  wire [7:0] p5_array_index_1081718_comb;
  wire [7:0] p5_res7__581_comb;
  wire [7:0] p5_res7__269_comb;
  wire [7:0] p5_array_index_1081729_comb;
  wire [7:0] p5_array_index_1081730_comb;
  wire [7:0] p5_array_index_1081731_comb;
  wire [7:0] p5_res7__582_comb;
  wire [7:0] p5_res7__270_comb;
  wire [7:0] p5_array_index_1081741_comb;
  wire [7:0] p5_array_index_1081742_comb;
  wire [7:0] p5_array_index_1081743_comb;
  wire [7:0] p5_res7__583_comb;
  wire [7:0] p5_res7__271_comb;
  wire [7:0] p5_array_index_1081754_comb;
  wire [7:0] p5_array_index_1081755_comb;
  wire [127:0] p5_res__16_comb;
  wire [7:0] p5_res7__584_comb;
  wire [127:0] p5_xor_1081289_comb;
  wire [7:0] p5_array_index_1081765_comb;
  wire [7:0] p5_array_index_1081766_comb;
  wire [127:0] p5_addedKey__58_comb;
  wire [7:0] p5_res7__585_comb;
  wire [7:0] p5_array_index_1081777_comb;
  wire [7:0] p5_array_index_1081305_comb;
  wire [7:0] p5_array_index_1081306_comb;
  wire [7:0] p5_array_index_1081307_comb;
  wire [7:0] p5_array_index_1081308_comb;
  wire [7:0] p5_array_index_1081309_comb;
  wire [7:0] p5_array_index_1081310_comb;
  wire [7:0] p5_array_index_1081312_comb;
  wire [7:0] p5_array_index_1081314_comb;
  wire [7:0] p5_array_index_1081315_comb;
  wire [7:0] p5_array_index_1081316_comb;
  wire [7:0] p5_array_index_1081317_comb;
  wire [7:0] p5_array_index_1081318_comb;
  wire [7:0] p5_array_index_1081319_comb;
  wire [7:0] p5_res7__586_comb;
  wire [7:0] p5_array_index_1081321_comb;
  wire [7:0] p5_array_index_1081322_comb;
  wire [7:0] p5_array_index_1081323_comb;
  wire [7:0] p5_array_index_1081324_comb;
  wire [7:0] p5_array_index_1081325_comb;
  wire [7:0] p5_array_index_1081326_comb;
  wire [7:0] p5_array_index_1081327_comb;
  wire [7:0] p5_array_index_1081329_comb;
  wire [7:0] p5_array_index_1081787_comb;
  wire [7:0] p5_res7__272_comb;
  wire [7:0] p5_res7__587_comb;
  wire [7:0] p5_array_index_1081338_comb;
  wire [7:0] p5_array_index_1081339_comb;
  wire [7:0] p5_array_index_1081340_comb;
  wire [7:0] p5_array_index_1081341_comb;
  wire [7:0] p5_array_index_1081342_comb;
  wire [7:0] p5_array_index_1081343_comb;
  wire [7:0] p5_res7__273_comb;
  wire [7:0] p5_res7__588_comb;
  wire [7:0] p5_array_index_1081353_comb;
  wire [7:0] p5_array_index_1081354_comb;
  wire [7:0] p5_array_index_1081355_comb;
  wire [7:0] p5_array_index_1081356_comb;
  wire [7:0] p5_array_index_1081357_comb;
  wire [7:0] p5_res7__274_comb;
  wire [7:0] p5_res7__589_comb;
  wire [7:0] p5_array_index_1081367_comb;
  wire [7:0] p5_array_index_1081368_comb;
  wire [7:0] p5_array_index_1081369_comb;
  wire [7:0] p5_array_index_1081370_comb;
  wire [7:0] p5_array_index_1081371_comb;
  wire [7:0] p5_res7__275_comb;
  wire [7:0] p5_res7__590_comb;
  wire [7:0] p5_array_index_1081382_comb;
  wire [7:0] p5_array_index_1081383_comb;
  wire [7:0] p5_array_index_1081384_comb;
  wire [7:0] p5_array_index_1081385_comb;
  wire [7:0] p5_res7__276_comb;
  wire [7:0] p5_res7__591_comb;
  wire [7:0] p5_array_index_1081395_comb;
  wire [7:0] p5_array_index_1081396_comb;
  wire [7:0] p5_array_index_1081397_comb;
  wire [7:0] p5_array_index_1081398_comb;
  wire [127:0] p5_res__36_comb;
  wire [7:0] p5_res7__277_comb;
  wire [127:0] p5_addedKey__37_comb;
  wire [7:0] p5_array_index_1081409_comb;
  wire [7:0] p5_array_index_1081410_comb;
  wire [7:0] p5_array_index_1081411_comb;
  wire [7:0] p5_res7__278_comb;
  wire [7:0] p5_array_index_1081841_comb;
  wire [7:0] p5_array_index_1081842_comb;
  wire [7:0] p5_array_index_1081843_comb;
  wire [7:0] p5_array_index_1081844_comb;
  wire [7:0] p5_array_index_1081845_comb;
  wire [7:0] p5_array_index_1081846_comb;
  wire [7:0] p5_array_index_1081848_comb;
  wire [7:0] p5_array_index_1081850_comb;
  wire [7:0] p5_array_index_1081851_comb;
  wire [7:0] p5_array_index_1081852_comb;
  wire [7:0] p5_array_index_1081853_comb;
  wire [7:0] p5_array_index_1081854_comb;
  wire [7:0] p5_array_index_1081855_comb;
  wire [7:0] p5_array_index_1081421_comb;
  wire [7:0] p5_array_index_1081422_comb;
  wire [7:0] p5_array_index_1081423_comb;
  wire [7:0] p5_array_index_1081857_comb;
  wire [7:0] p5_array_index_1081858_comb;
  wire [7:0] p5_array_index_1081859_comb;
  wire [7:0] p5_array_index_1081860_comb;
  wire [7:0] p5_array_index_1081861_comb;
  wire [7:0] p5_array_index_1081862_comb;
  wire [7:0] p5_array_index_1081863_comb;
  wire [7:0] p5_array_index_1081865_comb;
  wire [7:0] p5_res7__279_comb;
  wire [7:0] p5_res7__592_comb;
  wire [7:0] p5_array_index_1081434_comb;
  wire [7:0] p5_array_index_1081435_comb;
  wire [7:0] p5_array_index_1081874_comb;
  wire [7:0] p5_array_index_1081875_comb;
  wire [7:0] p5_array_index_1081876_comb;
  wire [7:0] p5_array_index_1081877_comb;
  wire [7:0] p5_array_index_1081878_comb;
  wire [7:0] p5_array_index_1081879_comb;
  wire [7:0] p5_res7__280_comb;
  wire [7:0] p5_res7__593_comb;
  wire [7:0] p5_array_index_1081445_comb;
  wire [7:0] p5_array_index_1081446_comb;
  wire [7:0] p5_array_index_1081889_comb;
  wire [7:0] p5_array_index_1081890_comb;
  wire [7:0] p5_array_index_1081891_comb;
  wire [7:0] p5_array_index_1081892_comb;
  wire [7:0] p5_array_index_1081893_comb;
  wire [7:0] p5_res7__281_comb;
  wire [7:0] p5_res7__594_comb;
  wire [7:0] p5_array_index_1081457_comb;
  wire [7:0] p5_array_index_1081903_comb;
  wire [7:0] p5_array_index_1081904_comb;
  wire [7:0] p5_array_index_1081905_comb;
  wire [7:0] p5_array_index_1081906_comb;
  wire [7:0] p5_array_index_1081907_comb;
  wire [7:0] p5_res7__282_comb;
  wire [7:0] p5_res7__595_comb;
  wire [7:0] p5_array_index_1081467_comb;
  wire [7:0] p5_array_index_1081918_comb;
  wire [7:0] p5_array_index_1081919_comb;
  wire [7:0] p5_array_index_1081920_comb;
  wire [7:0] p5_array_index_1081921_comb;
  wire [7:0] p5_res7__283_comb;
  wire [7:0] p5_res7__596_comb;
  wire [7:0] p5_array_index_1081931_comb;
  wire [7:0] p5_array_index_1081932_comb;
  wire [7:0] p5_array_index_1081933_comb;
  wire [7:0] p5_array_index_1081934_comb;
  wire [7:0] p5_res7__284_comb;
  wire [7:0] p5_res7__597_comb;
  wire [7:0] p5_array_index_1081945_comb;
  wire [7:0] p5_array_index_1081946_comb;
  wire [7:0] p5_array_index_1081947_comb;
  wire [7:0] p5_res7__285_comb;
  wire [7:0] p5_res7__598_comb;
  wire [7:0] p5_array_index_1081957_comb;
  wire [7:0] p5_array_index_1081958_comb;
  wire [7:0] p5_array_index_1081959_comb;
  wire [7:0] p5_res7__286_comb;
  wire [7:0] p5_res7__599_comb;
  wire [7:0] p5_array_index_1081970_comb;
  wire [7:0] p5_array_index_1081971_comb;
  wire [7:0] p5_res7__287_comb;
  wire [7:0] p5_res7__600_comb;
  wire [127:0] p5_res__17_comb;
  wire [7:0] p5_array_index_1081981_comb;
  wire [7:0] p5_array_index_1081982_comb;
  wire [127:0] p5_xor_1081507_comb;
  wire [7:0] p5_res7__601_comb;
  wire [127:0] p5_addedKey__59_comb;
  wire [7:0] p5_array_index_1081993_comb;
  wire [7:0] p5_res7__602_comb;
  wire [7:0] p5_array_index_1081523_comb;
  wire [7:0] p5_array_index_1081524_comb;
  wire [7:0] p5_array_index_1081525_comb;
  wire [7:0] p5_array_index_1081526_comb;
  wire [7:0] p5_array_index_1081527_comb;
  wire [7:0] p5_array_index_1081528_comb;
  wire [7:0] p5_array_index_1081530_comb;
  wire [7:0] p5_array_index_1081532_comb;
  wire [7:0] p5_array_index_1081533_comb;
  wire [7:0] p5_array_index_1081534_comb;
  wire [7:0] p5_array_index_1081535_comb;
  wire [7:0] p5_array_index_1081536_comb;
  wire [7:0] p5_array_index_1081537_comb;
  wire [7:0] p5_array_index_1082003_comb;
  wire [7:0] p5_array_index_1081539_comb;
  wire [7:0] p5_array_index_1081540_comb;
  wire [7:0] p5_array_index_1081541_comb;
  wire [7:0] p5_array_index_1081542_comb;
  wire [7:0] p5_array_index_1081543_comb;
  wire [7:0] p5_array_index_1081544_comb;
  wire [7:0] p5_array_index_1081545_comb;
  wire [7:0] p5_array_index_1081547_comb;
  wire [7:0] p5_res7__603_comb;
  wire [7:0] p5_res7__288_comb;
  wire [7:0] p5_array_index_1081556_comb;
  wire [7:0] p5_array_index_1081557_comb;
  wire [7:0] p5_array_index_1081558_comb;
  wire [7:0] p5_array_index_1081559_comb;
  wire [7:0] p5_array_index_1081560_comb;
  wire [7:0] p5_array_index_1081561_comb;
  wire [7:0] p5_res7__604_comb;
  wire [7:0] p5_res7__289_comb;
  wire [7:0] p5_array_index_1081571_comb;
  wire [7:0] p5_array_index_1081572_comb;
  wire [7:0] p5_array_index_1081573_comb;
  wire [7:0] p5_array_index_1081574_comb;
  wire [7:0] p5_array_index_1081575_comb;
  wire [7:0] p5_res7__605_comb;
  wire [7:0] p5_res7__290_comb;
  wire [7:0] p5_array_index_1081585_comb;
  wire [7:0] p5_array_index_1081586_comb;
  wire [7:0] p5_array_index_1081587_comb;
  wire [7:0] p5_array_index_1081588_comb;
  wire [7:0] p5_array_index_1081589_comb;
  wire [7:0] p5_res7__606_comb;
  wire [7:0] p5_res7__291_comb;
  wire [7:0] p5_array_index_1081600_comb;
  wire [7:0] p5_array_index_1081601_comb;
  wire [7:0] p5_array_index_1081602_comb;
  wire [7:0] p5_array_index_1081603_comb;
  wire [7:0] p5_res7__607_comb;
  wire [7:0] p5_res7__292_comb;
  wire [127:0] p5_res__37_comb;
  assign p5_res7__234_comb = p4_array_index_1080670 ^ p4_array_index_1080671 ^ p4_array_index_1080672 ^ p4_array_index_1080673 ^ p4_array_index_1080674 ^ p4_array_index_1080675 ^ p4_res7__227 ^ p4_array_index_1080676 ^ p4_res7__225 ^ p4_array_index_1080629 ^ p4_array_index_1080602 ^ p4_array_index_1080573 ^ p4_array_index_1080541 ^ p4_array_index_1080677 ^ p4_array_index_1080678 ^ p4_array_index_1080528;
  assign p5_array_index_1080813_comb = p4_literal_1076355[p4_res7__229];
  assign p5_res7__235_comb = p4_literal_1076345[p5_res7__234_comb] ^ p4_literal_1076347[p4_res7__233] ^ p4_literal_1076349[p4_res7__232] ^ p4_literal_1076351[p4_res7__231] ^ p4_literal_1076353[p4_res7__230] ^ p5_array_index_1080813_comb ^ p4_res7__228 ^ p4_literal_1076358[p4_res7__227] ^ p4_res7__226 ^ p4_array_index_1080641 ^ p4_array_index_1080615 ^ p4_array_index_1080587 ^ p4_array_index_1080558 ^ p4_literal_1076347[p4_array_index_1080525] ^ p4_literal_1076345[p4_array_index_1080526] ^ p4_array_index_1080527;
  assign p5_res7__236_comb = p4_literal_1076345[p5_res7__235_comb] ^ p4_literal_1076347[p5_res7__234_comb] ^ p4_literal_1076349[p4_res7__233] ^ p4_literal_1076351[p4_res7__232] ^ p4_literal_1076353[p4_res7__231] ^ p4_literal_1076355[p4_res7__230] ^ p4_res7__229 ^ p4_literal_1076358[p4_res7__228] ^ p4_res7__227 ^ p4_array_index_1080653 ^ p4_array_index_1080628 ^ p4_array_index_1080601 ^ p4_array_index_1080572 ^ p4_array_index_1080540 ^ p4_literal_1076345[p4_array_index_1080525] ^ p4_array_index_1080526;
  assign p5_res7__237_comb = p4_literal_1076345[p5_res7__236_comb] ^ p4_literal_1076347[p5_res7__235_comb] ^ p4_literal_1076349[p5_res7__234_comb] ^ p4_literal_1076351[p4_res7__233] ^ p4_literal_1076353[p4_res7__232] ^ p4_literal_1076355[p4_res7__231] ^ p4_res7__230 ^ p4_literal_1076358[p4_res7__229] ^ p4_res7__228 ^ p4_array_index_1080664 ^ p4_array_index_1080640 ^ p4_array_index_1080614 ^ p4_array_index_1080586 ^ p4_array_index_1080557 ^ p4_literal_1076345[p4_array_index_1080524] ^ p4_array_index_1080525;
  assign p5_res7__238_comb = p4_literal_1076345[p5_res7__237_comb] ^ p4_literal_1076347[p5_res7__236_comb] ^ p4_literal_1076349[p5_res7__235_comb] ^ p4_literal_1076351[p5_res7__234_comb] ^ p4_literal_1076353[p4_res7__233] ^ p4_literal_1076355[p4_res7__232] ^ p4_res7__231 ^ p4_literal_1076358[p4_res7__230] ^ p4_res7__229 ^ p4_array_index_1080675 ^ p4_array_index_1080652 ^ p4_array_index_1080627 ^ p4_array_index_1080600 ^ p4_array_index_1080571 ^ p4_array_index_1080539 ^ p4_array_index_1080524;
  assign p5_res7__239_comb = p4_literal_1076345[p5_res7__238_comb] ^ p4_literal_1076347[p5_res7__237_comb] ^ p4_literal_1076349[p5_res7__236_comb] ^ p4_literal_1076351[p5_res7__235_comb] ^ p4_literal_1076353[p5_res7__234_comb] ^ p4_literal_1076355[p4_res7__233] ^ p4_res7__232 ^ p4_literal_1076358[p4_res7__231] ^ p4_res7__230 ^ p5_array_index_1080813_comb ^ p4_array_index_1080663 ^ p4_array_index_1080639 ^ p4_array_index_1080613 ^ p4_array_index_1080585 ^ p4_array_index_1080556 ^ p4_array_index_1080523;
  assign p5_res__14_comb = {p5_res7__239_comb, p5_res7__238_comb, p5_res7__237_comb, p5_res7__236_comb, p5_res7__235_comb, p5_res7__234_comb, p4_res7__233, p4_res7__232, p4_res7__231, p4_res7__230, p4_res7__229, p4_res7__228, p4_res7__227, p4_res7__226, p4_res7__225, p4_res7__224};
  assign p5_k5_comb = p5_res__14_comb ^ p4_xor_1080289;
  assign p5_addedKey__56_comb = p5_k5_comb ^ 128'h2fb2_6c2c_0f0a_acd1_9935_81c3_4e97_5410;
  assign p5_array_index_1080869_comb = p4_arr[p5_addedKey__56_comb[127:120]];
  assign p5_array_index_1080870_comb = p4_arr[p5_addedKey__56_comb[119:112]];
  assign p5_array_index_1080871_comb = p4_arr[p5_addedKey__56_comb[111:104]];
  assign p5_array_index_1080872_comb = p4_arr[p5_addedKey__56_comb[103:96]];
  assign p5_array_index_1080873_comb = p4_arr[p5_addedKey__56_comb[95:88]];
  assign p5_array_index_1080874_comb = p4_arr[p5_addedKey__56_comb[87:80]];
  assign p5_array_index_1080876_comb = p4_arr[p5_addedKey__56_comb[71:64]];
  assign p5_array_index_1080878_comb = p4_arr[p5_addedKey__56_comb[55:48]];
  assign p5_array_index_1080879_comb = p4_arr[p5_addedKey__56_comb[47:40]];
  assign p5_array_index_1080880_comb = p4_arr[p5_addedKey__56_comb[39:32]];
  assign p5_array_index_1080881_comb = p4_arr[p5_addedKey__56_comb[31:24]];
  assign p5_array_index_1080882_comb = p4_arr[p5_addedKey__56_comb[23:16]];
  assign p5_array_index_1080883_comb = p4_arr[p5_addedKey__56_comb[15:8]];
  assign p5_array_index_1080885_comb = p4_literal_1076345[p5_array_index_1080869_comb];
  assign p5_array_index_1080886_comb = p4_literal_1076347[p5_array_index_1080870_comb];
  assign p5_array_index_1080887_comb = p4_literal_1076349[p5_array_index_1080871_comb];
  assign p5_array_index_1080888_comb = p4_literal_1076351[p5_array_index_1080872_comb];
  assign p5_array_index_1080889_comb = p4_literal_1076353[p5_array_index_1080873_comb];
  assign p5_array_index_1080890_comb = p4_literal_1076355[p5_array_index_1080874_comb];
  assign p5_array_index_1080891_comb = p4_arr[p5_addedKey__56_comb[79:72]];
  assign p5_array_index_1080893_comb = p4_arr[p5_addedKey__56_comb[63:56]];
  assign p5_res7__240_comb = p5_array_index_1080885_comb ^ p5_array_index_1080886_comb ^ p5_array_index_1080887_comb ^ p5_array_index_1080888_comb ^ p5_array_index_1080889_comb ^ p5_array_index_1080890_comb ^ p5_array_index_1080891_comb ^ p4_literal_1076358[p5_array_index_1080876_comb] ^ p5_array_index_1080893_comb ^ p4_literal_1076355[p5_array_index_1080878_comb] ^ p4_literal_1076353[p5_array_index_1080879_comb] ^ p4_literal_1076351[p5_array_index_1080880_comb] ^ p4_literal_1076349[p5_array_index_1080881_comb] ^ p4_literal_1076347[p5_array_index_1080882_comb] ^ p4_literal_1076345[p5_array_index_1080883_comb] ^ p4_arr[p5_addedKey__56_comb[7:0]];
  assign p5_array_index_1080902_comb = p4_literal_1076345[p5_res7__240_comb];
  assign p5_array_index_1080903_comb = p4_literal_1076347[p5_array_index_1080869_comb];
  assign p5_array_index_1080904_comb = p4_literal_1076349[p5_array_index_1080870_comb];
  assign p5_array_index_1080905_comb = p4_literal_1076351[p5_array_index_1080871_comb];
  assign p5_array_index_1080906_comb = p4_literal_1076353[p5_array_index_1080872_comb];
  assign p5_array_index_1080907_comb = p4_literal_1076355[p5_array_index_1080873_comb];
  assign p5_res7__241_comb = p5_array_index_1080902_comb ^ p5_array_index_1080903_comb ^ p5_array_index_1080904_comb ^ p5_array_index_1080905_comb ^ p5_array_index_1080906_comb ^ p5_array_index_1080907_comb ^ p5_array_index_1080874_comb ^ p4_literal_1076358[p5_array_index_1080891_comb] ^ p5_array_index_1080876_comb ^ p4_literal_1076355[p5_array_index_1080893_comb] ^ p4_literal_1076353[p5_array_index_1080878_comb] ^ p4_literal_1076351[p5_array_index_1080879_comb] ^ p4_literal_1076349[p5_array_index_1080880_comb] ^ p4_literal_1076347[p5_array_index_1080881_comb] ^ p4_literal_1076345[p5_array_index_1080882_comb] ^ p5_array_index_1080883_comb;
  assign p5_array_index_1080917_comb = p4_literal_1076347[p5_res7__240_comb];
  assign p5_array_index_1080918_comb = p4_literal_1076349[p5_array_index_1080869_comb];
  assign p5_array_index_1080919_comb = p4_literal_1076351[p5_array_index_1080870_comb];
  assign p5_array_index_1080920_comb = p4_literal_1076353[p5_array_index_1080871_comb];
  assign p5_array_index_1080921_comb = p4_literal_1076355[p5_array_index_1080872_comb];
  assign p5_res7__242_comb = p4_literal_1076345[p5_res7__241_comb] ^ p5_array_index_1080917_comb ^ p5_array_index_1080918_comb ^ p5_array_index_1080919_comb ^ p5_array_index_1080920_comb ^ p5_array_index_1080921_comb ^ p5_array_index_1080873_comb ^ p4_literal_1076358[p5_array_index_1080874_comb] ^ p5_array_index_1080891_comb ^ p4_literal_1076355[p5_array_index_1080876_comb] ^ p4_literal_1076353[p5_array_index_1080893_comb] ^ p4_literal_1076351[p5_array_index_1080878_comb] ^ p4_literal_1076349[p5_array_index_1080879_comb] ^ p4_literal_1076347[p5_array_index_1080880_comb] ^ p4_literal_1076345[p5_array_index_1080881_comb] ^ p5_array_index_1080882_comb;
  assign p5_array_index_1080931_comb = p4_literal_1076347[p5_res7__241_comb];
  assign p5_array_index_1080932_comb = p4_literal_1076349[p5_res7__240_comb];
  assign p5_array_index_1080933_comb = p4_literal_1076351[p5_array_index_1080869_comb];
  assign p5_array_index_1080934_comb = p4_literal_1076353[p5_array_index_1080870_comb];
  assign p5_array_index_1080935_comb = p4_literal_1076355[p5_array_index_1080871_comb];
  assign p5_res7__243_comb = p4_literal_1076345[p5_res7__242_comb] ^ p5_array_index_1080931_comb ^ p5_array_index_1080932_comb ^ p5_array_index_1080933_comb ^ p5_array_index_1080934_comb ^ p5_array_index_1080935_comb ^ p5_array_index_1080872_comb ^ p4_literal_1076358[p5_array_index_1080873_comb] ^ p5_array_index_1080874_comb ^ p4_literal_1076355[p5_array_index_1080891_comb] ^ p4_literal_1076353[p5_array_index_1080876_comb] ^ p4_literal_1076351[p5_array_index_1080893_comb] ^ p4_literal_1076349[p5_array_index_1080878_comb] ^ p4_literal_1076347[p5_array_index_1080879_comb] ^ p4_literal_1076345[p5_array_index_1080880_comb] ^ p5_array_index_1080881_comb;
  assign p5_array_index_1080946_comb = p4_literal_1076349[p5_res7__241_comb];
  assign p5_array_index_1080947_comb = p4_literal_1076351[p5_res7__240_comb];
  assign p5_array_index_1080948_comb = p4_literal_1076353[p5_array_index_1080869_comb];
  assign p5_array_index_1080949_comb = p4_literal_1076355[p5_array_index_1080870_comb];
  assign p5_res7__244_comb = p4_literal_1076345[p5_res7__243_comb] ^ p4_literal_1076347[p5_res7__242_comb] ^ p5_array_index_1080946_comb ^ p5_array_index_1080947_comb ^ p5_array_index_1080948_comb ^ p5_array_index_1080949_comb ^ p5_array_index_1080871_comb ^ p4_literal_1076358[p5_array_index_1080872_comb] ^ p5_array_index_1080873_comb ^ p5_array_index_1080890_comb ^ p4_literal_1076353[p5_array_index_1080891_comb] ^ p4_literal_1076351[p5_array_index_1080876_comb] ^ p4_literal_1076349[p5_array_index_1080893_comb] ^ p4_literal_1076347[p5_array_index_1080878_comb] ^ p4_literal_1076345[p5_array_index_1080879_comb] ^ p5_array_index_1080880_comb;
  assign p5_array_index_1080959_comb = p4_literal_1076349[p5_res7__242_comb];
  assign p5_array_index_1080960_comb = p4_literal_1076351[p5_res7__241_comb];
  assign p5_array_index_1080961_comb = p4_literal_1076353[p5_res7__240_comb];
  assign p5_array_index_1080962_comb = p4_literal_1076355[p5_array_index_1080869_comb];
  assign p5_res7__245_comb = p4_literal_1076345[p5_res7__244_comb] ^ p4_literal_1076347[p5_res7__243_comb] ^ p5_array_index_1080959_comb ^ p5_array_index_1080960_comb ^ p5_array_index_1080961_comb ^ p5_array_index_1080962_comb ^ p5_array_index_1080870_comb ^ p4_literal_1076358[p5_array_index_1080871_comb] ^ p5_array_index_1080872_comb ^ p5_array_index_1080907_comb ^ p4_literal_1076353[p5_array_index_1080874_comb] ^ p4_literal_1076351[p5_array_index_1080891_comb] ^ p4_literal_1076349[p5_array_index_1080876_comb] ^ p4_literal_1076347[p5_array_index_1080893_comb] ^ p4_literal_1076345[p5_array_index_1080878_comb] ^ p5_array_index_1080879_comb;
  assign p5_array_index_1080973_comb = p4_literal_1076351[p5_res7__242_comb];
  assign p5_array_index_1080974_comb = p4_literal_1076353[p5_res7__241_comb];
  assign p5_array_index_1080975_comb = p4_literal_1076355[p5_res7__240_comb];
  assign p5_res7__246_comb = p4_literal_1076345[p5_res7__245_comb] ^ p4_literal_1076347[p5_res7__244_comb] ^ p4_literal_1076349[p5_res7__243_comb] ^ p5_array_index_1080973_comb ^ p5_array_index_1080974_comb ^ p5_array_index_1080975_comb ^ p5_array_index_1080869_comb ^ p4_literal_1076358[p5_array_index_1080870_comb] ^ p5_array_index_1080871_comb ^ p5_array_index_1080921_comb ^ p5_array_index_1080889_comb ^ p4_literal_1076351[p5_array_index_1080874_comb] ^ p4_literal_1076349[p5_array_index_1080891_comb] ^ p4_literal_1076347[p5_array_index_1080876_comb] ^ p4_literal_1076345[p5_array_index_1080893_comb] ^ p5_array_index_1080878_comb;
  assign p5_array_index_1080985_comb = p4_literal_1076351[p5_res7__243_comb];
  assign p5_array_index_1080986_comb = p4_literal_1076353[p5_res7__242_comb];
  assign p5_array_index_1080987_comb = p4_literal_1076355[p5_res7__241_comb];
  assign p5_res7__247_comb = p4_literal_1076345[p5_res7__246_comb] ^ p4_literal_1076347[p5_res7__245_comb] ^ p4_literal_1076349[p5_res7__244_comb] ^ p5_array_index_1080985_comb ^ p5_array_index_1080986_comb ^ p5_array_index_1080987_comb ^ p5_res7__240_comb ^ p4_literal_1076358[p5_array_index_1080869_comb] ^ p5_array_index_1080870_comb ^ p5_array_index_1080935_comb ^ p5_array_index_1080906_comb ^ p4_literal_1076351[p5_array_index_1080873_comb] ^ p4_literal_1076349[p5_array_index_1080874_comb] ^ p4_literal_1076347[p5_array_index_1080891_comb] ^ p4_literal_1076345[p5_array_index_1080876_comb] ^ p5_array_index_1080893_comb;
  assign p5_array_index_1080998_comb = p4_literal_1076353[p5_res7__243_comb];
  assign p5_array_index_1080999_comb = p4_literal_1076355[p5_res7__242_comb];
  assign p5_res7__248_comb = p4_literal_1076345[p5_res7__247_comb] ^ p4_literal_1076347[p5_res7__246_comb] ^ p4_literal_1076349[p5_res7__245_comb] ^ p4_literal_1076351[p5_res7__244_comb] ^ p5_array_index_1080998_comb ^ p5_array_index_1080999_comb ^ p5_res7__241_comb ^ p4_literal_1076358[p5_res7__240_comb] ^ p5_array_index_1080869_comb ^ p5_array_index_1080949_comb ^ p5_array_index_1080920_comb ^ p5_array_index_1080888_comb ^ p4_literal_1076349[p5_array_index_1080873_comb] ^ p4_literal_1076347[p5_array_index_1080874_comb] ^ p4_literal_1076345[p5_array_index_1080891_comb] ^ p5_array_index_1080876_comb;
  assign p5_array_index_1081009_comb = p4_literal_1076353[p5_res7__244_comb];
  assign p5_array_index_1081010_comb = p4_literal_1076355[p5_res7__243_comb];
  assign p5_res7__249_comb = p4_literal_1076345[p5_res7__248_comb] ^ p4_literal_1076347[p5_res7__247_comb] ^ p4_literal_1076349[p5_res7__246_comb] ^ p4_literal_1076351[p5_res7__245_comb] ^ p5_array_index_1081009_comb ^ p5_array_index_1081010_comb ^ p5_res7__242_comb ^ p4_literal_1076358[p5_res7__241_comb] ^ p5_res7__240_comb ^ p5_array_index_1080962_comb ^ p5_array_index_1080934_comb ^ p5_array_index_1080905_comb ^ p4_literal_1076349[p5_array_index_1080872_comb] ^ p4_literal_1076347[p5_array_index_1080873_comb] ^ p4_literal_1076345[p5_array_index_1080874_comb] ^ p5_array_index_1080891_comb;
  assign p5_array_index_1081021_comb = p4_literal_1076355[p5_res7__244_comb];
  assign p5_res7__250_comb = p4_literal_1076345[p5_res7__249_comb] ^ p4_literal_1076347[p5_res7__248_comb] ^ p4_literal_1076349[p5_res7__247_comb] ^ p4_literal_1076351[p5_res7__246_comb] ^ p4_literal_1076353[p5_res7__245_comb] ^ p5_array_index_1081021_comb ^ p5_res7__243_comb ^ p4_literal_1076358[p5_res7__242_comb] ^ p5_res7__241_comb ^ p5_array_index_1080975_comb ^ p5_array_index_1080948_comb ^ p5_array_index_1080919_comb ^ p5_array_index_1080887_comb ^ p4_literal_1076347[p5_array_index_1080872_comb] ^ p4_literal_1076345[p5_array_index_1080873_comb] ^ p5_array_index_1080874_comb;
  assign p5_array_index_1081031_comb = p4_literal_1076355[p5_res7__245_comb];
  assign p5_res7__251_comb = p4_literal_1076345[p5_res7__250_comb] ^ p4_literal_1076347[p5_res7__249_comb] ^ p4_literal_1076349[p5_res7__248_comb] ^ p4_literal_1076351[p5_res7__247_comb] ^ p4_literal_1076353[p5_res7__246_comb] ^ p5_array_index_1081031_comb ^ p5_res7__244_comb ^ p4_literal_1076358[p5_res7__243_comb] ^ p5_res7__242_comb ^ p5_array_index_1080987_comb ^ p5_array_index_1080961_comb ^ p5_array_index_1080933_comb ^ p5_array_index_1080904_comb ^ p4_literal_1076347[p5_array_index_1080871_comb] ^ p4_literal_1076345[p5_array_index_1080872_comb] ^ p5_array_index_1080873_comb;
  assign p5_res7__252_comb = p4_literal_1076345[p5_res7__251_comb] ^ p4_literal_1076347[p5_res7__250_comb] ^ p4_literal_1076349[p5_res7__249_comb] ^ p4_literal_1076351[p5_res7__248_comb] ^ p4_literal_1076353[p5_res7__247_comb] ^ p4_literal_1076355[p5_res7__246_comb] ^ p5_res7__245_comb ^ p4_literal_1076358[p5_res7__244_comb] ^ p5_res7__243_comb ^ p5_array_index_1080999_comb ^ p5_array_index_1080974_comb ^ p5_array_index_1080947_comb ^ p5_array_index_1080918_comb ^ p5_array_index_1080886_comb ^ p4_literal_1076345[p5_array_index_1080871_comb] ^ p5_array_index_1080872_comb;
  assign p5_res7__253_comb = p4_literal_1076345[p5_res7__252_comb] ^ p4_literal_1076347[p5_res7__251_comb] ^ p4_literal_1076349[p5_res7__250_comb] ^ p4_literal_1076351[p5_res7__249_comb] ^ p4_literal_1076353[p5_res7__248_comb] ^ p4_literal_1076355[p5_res7__247_comb] ^ p5_res7__246_comb ^ p4_literal_1076358[p5_res7__245_comb] ^ p5_res7__244_comb ^ p5_array_index_1081010_comb ^ p5_array_index_1080986_comb ^ p5_array_index_1080960_comb ^ p5_array_index_1080932_comb ^ p5_array_index_1080903_comb ^ p4_literal_1076345[p5_array_index_1080870_comb] ^ p5_array_index_1080871_comb;
  assign p5_res7__254_comb = p4_literal_1076345[p5_res7__253_comb] ^ p4_literal_1076347[p5_res7__252_comb] ^ p4_literal_1076349[p5_res7__251_comb] ^ p4_literal_1076351[p5_res7__250_comb] ^ p4_literal_1076353[p5_res7__249_comb] ^ p4_literal_1076355[p5_res7__248_comb] ^ p5_res7__247_comb ^ p4_literal_1076358[p5_res7__246_comb] ^ p5_res7__245_comb ^ p5_array_index_1081021_comb ^ p5_array_index_1080998_comb ^ p5_array_index_1080973_comb ^ p5_array_index_1080946_comb ^ p5_array_index_1080917_comb ^ p5_array_index_1080885_comb ^ p5_array_index_1080870_comb;
  assign p5_res7__255_comb = p4_literal_1076345[p5_res7__254_comb] ^ p4_literal_1076347[p5_res7__253_comb] ^ p4_literal_1076349[p5_res7__252_comb] ^ p4_literal_1076351[p5_res7__251_comb] ^ p4_literal_1076353[p5_res7__250_comb] ^ p4_literal_1076355[p5_res7__249_comb] ^ p5_res7__248_comb ^ p4_literal_1076358[p5_res7__247_comb] ^ p5_res7__246_comb ^ p5_array_index_1081031_comb ^ p5_array_index_1081009_comb ^ p5_array_index_1080985_comb ^ p5_array_index_1080959_comb ^ p5_array_index_1080931_comb ^ p5_array_index_1080902_comb ^ p5_array_index_1080869_comb;
  assign p5_res__15_comb = {p5_res7__255_comb, p5_res7__254_comb, p5_res7__253_comb, p5_res7__252_comb, p5_res7__251_comb, p5_res7__250_comb, p5_res7__249_comb, p5_res7__248_comb, p5_res7__247_comb, p5_res7__246_comb, p5_res7__245_comb, p5_res7__244_comb, p5_res7__243_comb, p5_res7__242_comb, p5_res7__241_comb, p5_res7__240_comb};
  assign p5_k4_comb = p5_res__15_comb ^ p4_xor_1080507;
  assign p5_addedKey__57_comb = p5_k4_comb ^ 128'h4110_1a5e_6342_d669_c412_3cd3_9313_c011;
  assign p5_array_index_1081087_comb = p4_arr[p5_addedKey__57_comb[127:120]];
  assign p5_array_index_1081088_comb = p4_arr[p5_addedKey__57_comb[119:112]];
  assign p5_array_index_1081089_comb = p4_arr[p5_addedKey__57_comb[111:104]];
  assign p5_array_index_1081090_comb = p4_arr[p5_addedKey__57_comb[103:96]];
  assign p5_array_index_1081091_comb = p4_arr[p5_addedKey__57_comb[95:88]];
  assign p5_array_index_1081092_comb = p4_arr[p5_addedKey__57_comb[87:80]];
  assign p5_array_index_1081094_comb = p4_arr[p5_addedKey__57_comb[71:64]];
  assign p5_array_index_1081096_comb = p4_arr[p5_addedKey__57_comb[55:48]];
  assign p5_array_index_1081097_comb = p4_arr[p5_addedKey__57_comb[47:40]];
  assign p5_array_index_1081098_comb = p4_arr[p5_addedKey__57_comb[39:32]];
  assign p5_array_index_1081099_comb = p4_arr[p5_addedKey__57_comb[31:24]];
  assign p5_array_index_1081100_comb = p4_arr[p5_addedKey__57_comb[23:16]];
  assign p5_array_index_1081101_comb = p4_arr[p5_addedKey__57_comb[15:8]];
  assign p5_array_index_1081103_comb = p4_literal_1076345[p5_array_index_1081087_comb];
  assign p5_array_index_1081104_comb = p4_literal_1076347[p5_array_index_1081088_comb];
  assign p5_array_index_1081105_comb = p4_literal_1076349[p5_array_index_1081089_comb];
  assign p5_array_index_1081106_comb = p4_literal_1076351[p5_array_index_1081090_comb];
  assign p5_array_index_1081107_comb = p4_literal_1076353[p5_array_index_1081091_comb];
  assign p5_array_index_1081108_comb = p4_literal_1076355[p5_array_index_1081092_comb];
  assign p5_array_index_1081109_comb = p4_arr[p5_addedKey__57_comb[79:72]];
  assign p5_array_index_1081111_comb = p4_arr[p5_addedKey__57_comb[63:56]];
  assign p5_res7__256_comb = p5_array_index_1081103_comb ^ p5_array_index_1081104_comb ^ p5_array_index_1081105_comb ^ p5_array_index_1081106_comb ^ p5_array_index_1081107_comb ^ p5_array_index_1081108_comb ^ p5_array_index_1081109_comb ^ p4_literal_1076358[p5_array_index_1081094_comb] ^ p5_array_index_1081111_comb ^ p4_literal_1076355[p5_array_index_1081096_comb] ^ p4_literal_1076353[p5_array_index_1081097_comb] ^ p4_literal_1076351[p5_array_index_1081098_comb] ^ p4_literal_1076349[p5_array_index_1081099_comb] ^ p4_literal_1076347[p5_array_index_1081100_comb] ^ p4_literal_1076345[p5_array_index_1081101_comb] ^ p4_arr[p5_addedKey__57_comb[7:0]];
  assign p5_array_index_1081120_comb = p4_literal_1076345[p5_res7__256_comb];
  assign p5_array_index_1081121_comb = p4_literal_1076347[p5_array_index_1081087_comb];
  assign p5_array_index_1081122_comb = p4_literal_1076349[p5_array_index_1081088_comb];
  assign p5_array_index_1081123_comb = p4_literal_1076351[p5_array_index_1081089_comb];
  assign p5_array_index_1081124_comb = p4_literal_1076353[p5_array_index_1081090_comb];
  assign p5_array_index_1081125_comb = p4_literal_1076355[p5_array_index_1081091_comb];
  assign p5_res7__257_comb = p5_array_index_1081120_comb ^ p5_array_index_1081121_comb ^ p5_array_index_1081122_comb ^ p5_array_index_1081123_comb ^ p5_array_index_1081124_comb ^ p5_array_index_1081125_comb ^ p5_array_index_1081092_comb ^ p4_literal_1076358[p5_array_index_1081109_comb] ^ p5_array_index_1081094_comb ^ p4_literal_1076355[p5_array_index_1081111_comb] ^ p4_literal_1076353[p5_array_index_1081096_comb] ^ p4_literal_1076351[p5_array_index_1081097_comb] ^ p4_literal_1076349[p5_array_index_1081098_comb] ^ p4_literal_1076347[p5_array_index_1081099_comb] ^ p4_literal_1076345[p5_array_index_1081100_comb] ^ p5_array_index_1081101_comb;
  assign p5_array_index_1081135_comb = p4_literal_1076347[p5_res7__256_comb];
  assign p5_array_index_1081136_comb = p4_literal_1076349[p5_array_index_1081087_comb];
  assign p5_array_index_1081137_comb = p4_literal_1076351[p5_array_index_1081088_comb];
  assign p5_array_index_1081138_comb = p4_literal_1076353[p5_array_index_1081089_comb];
  assign p5_array_index_1081139_comb = p4_literal_1076355[p5_array_index_1081090_comb];
  assign p5_res7__258_comb = p4_literal_1076345[p5_res7__257_comb] ^ p5_array_index_1081135_comb ^ p5_array_index_1081136_comb ^ p5_array_index_1081137_comb ^ p5_array_index_1081138_comb ^ p5_array_index_1081139_comb ^ p5_array_index_1081091_comb ^ p4_literal_1076358[p5_array_index_1081092_comb] ^ p5_array_index_1081109_comb ^ p4_literal_1076355[p5_array_index_1081094_comb] ^ p4_literal_1076353[p5_array_index_1081111_comb] ^ p4_literal_1076351[p5_array_index_1081096_comb] ^ p4_literal_1076349[p5_array_index_1081097_comb] ^ p4_literal_1076347[p5_array_index_1081098_comb] ^ p4_literal_1076345[p5_array_index_1081099_comb] ^ p5_array_index_1081100_comb;
  assign p5_array_index_1081149_comb = p4_literal_1076347[p5_res7__257_comb];
  assign p5_array_index_1081150_comb = p4_literal_1076349[p5_res7__256_comb];
  assign p5_array_index_1081151_comb = p4_literal_1076351[p5_array_index_1081087_comb];
  assign p5_array_index_1081152_comb = p4_literal_1076353[p5_array_index_1081088_comb];
  assign p5_array_index_1081153_comb = p4_literal_1076355[p5_array_index_1081089_comb];
  assign p5_res7__259_comb = p4_literal_1076345[p5_res7__258_comb] ^ p5_array_index_1081149_comb ^ p5_array_index_1081150_comb ^ p5_array_index_1081151_comb ^ p5_array_index_1081152_comb ^ p5_array_index_1081153_comb ^ p5_array_index_1081090_comb ^ p4_literal_1076358[p5_array_index_1081091_comb] ^ p5_array_index_1081092_comb ^ p4_literal_1076355[p5_array_index_1081109_comb] ^ p4_literal_1076353[p5_array_index_1081094_comb] ^ p4_literal_1076351[p5_array_index_1081111_comb] ^ p4_literal_1076349[p5_array_index_1081096_comb] ^ p4_literal_1076347[p5_array_index_1081097_comb] ^ p4_literal_1076345[p5_array_index_1081098_comb] ^ p5_array_index_1081099_comb;
  assign p5_array_index_1081164_comb = p4_literal_1076349[p5_res7__257_comb];
  assign p5_array_index_1081165_comb = p4_literal_1076351[p5_res7__256_comb];
  assign p5_array_index_1081166_comb = p4_literal_1076353[p5_array_index_1081087_comb];
  assign p5_array_index_1081167_comb = p4_literal_1076355[p5_array_index_1081088_comb];
  assign p5_res7__260_comb = p4_literal_1076345[p5_res7__259_comb] ^ p4_literal_1076347[p5_res7__258_comb] ^ p5_array_index_1081164_comb ^ p5_array_index_1081165_comb ^ p5_array_index_1081166_comb ^ p5_array_index_1081167_comb ^ p5_array_index_1081089_comb ^ p4_literal_1076358[p5_array_index_1081090_comb] ^ p5_array_index_1081091_comb ^ p5_array_index_1081108_comb ^ p4_literal_1076353[p5_array_index_1081109_comb] ^ p4_literal_1076351[p5_array_index_1081094_comb] ^ p4_literal_1076349[p5_array_index_1081111_comb] ^ p4_literal_1076347[p5_array_index_1081096_comb] ^ p4_literal_1076345[p5_array_index_1081097_comb] ^ p5_array_index_1081098_comb;
  assign p5_array_index_1081177_comb = p4_literal_1076349[p5_res7__258_comb];
  assign p5_array_index_1081178_comb = p4_literal_1076351[p5_res7__257_comb];
  assign p5_array_index_1081179_comb = p4_literal_1076353[p5_res7__256_comb];
  assign p5_array_index_1081180_comb = p4_literal_1076355[p5_array_index_1081087_comb];
  assign p5_res7__261_comb = p4_literal_1076345[p5_res7__260_comb] ^ p4_literal_1076347[p5_res7__259_comb] ^ p5_array_index_1081177_comb ^ p5_array_index_1081178_comb ^ p5_array_index_1081179_comb ^ p5_array_index_1081180_comb ^ p5_array_index_1081088_comb ^ p4_literal_1076358[p5_array_index_1081089_comb] ^ p5_array_index_1081090_comb ^ p5_array_index_1081125_comb ^ p4_literal_1076353[p5_array_index_1081092_comb] ^ p4_literal_1076351[p5_array_index_1081109_comb] ^ p4_literal_1076349[p5_array_index_1081094_comb] ^ p4_literal_1076347[p5_array_index_1081111_comb] ^ p4_literal_1076345[p5_array_index_1081096_comb] ^ p5_array_index_1081097_comb;
  assign p5_array_index_1081191_comb = p4_literal_1076351[p5_res7__258_comb];
  assign p5_array_index_1081192_comb = p4_literal_1076353[p5_res7__257_comb];
  assign p5_array_index_1081193_comb = p4_literal_1076355[p5_res7__256_comb];
  assign p5_addedKey__36_comb = p5_k4_comb ^ p4_res__35;
  assign p5_res7__262_comb = p4_literal_1076345[p5_res7__261_comb] ^ p4_literal_1076347[p5_res7__260_comb] ^ p4_literal_1076349[p5_res7__259_comb] ^ p5_array_index_1081191_comb ^ p5_array_index_1081192_comb ^ p5_array_index_1081193_comb ^ p5_array_index_1081087_comb ^ p4_literal_1076358[p5_array_index_1081088_comb] ^ p5_array_index_1081089_comb ^ p5_array_index_1081139_comb ^ p5_array_index_1081107_comb ^ p4_literal_1076351[p5_array_index_1081092_comb] ^ p4_literal_1076349[p5_array_index_1081109_comb] ^ p4_literal_1076347[p5_array_index_1081094_comb] ^ p4_literal_1076345[p5_array_index_1081111_comb] ^ p5_array_index_1081096_comb;
  assign p5_array_index_1081203_comb = p4_literal_1076351[p5_res7__259_comb];
  assign p5_array_index_1081204_comb = p4_literal_1076353[p5_res7__258_comb];
  assign p5_array_index_1081205_comb = p4_literal_1076355[p5_res7__257_comb];
  assign p5_array_index_1081625_comb = p4_arr[p5_addedKey__36_comb[127:120]];
  assign p5_array_index_1081626_comb = p4_arr[p5_addedKey__36_comb[119:112]];
  assign p5_array_index_1081627_comb = p4_arr[p5_addedKey__36_comb[111:104]];
  assign p5_array_index_1081628_comb = p4_arr[p5_addedKey__36_comb[103:96]];
  assign p5_array_index_1081629_comb = p4_arr[p5_addedKey__36_comb[95:88]];
  assign p5_array_index_1081630_comb = p4_arr[p5_addedKey__36_comb[87:80]];
  assign p5_array_index_1081632_comb = p4_arr[p5_addedKey__36_comb[71:64]];
  assign p5_array_index_1081634_comb = p4_arr[p5_addedKey__36_comb[55:48]];
  assign p5_array_index_1081635_comb = p4_arr[p5_addedKey__36_comb[47:40]];
  assign p5_array_index_1081636_comb = p4_arr[p5_addedKey__36_comb[39:32]];
  assign p5_array_index_1081637_comb = p4_arr[p5_addedKey__36_comb[31:24]];
  assign p5_array_index_1081638_comb = p4_arr[p5_addedKey__36_comb[23:16]];
  assign p5_array_index_1081639_comb = p4_arr[p5_addedKey__36_comb[15:8]];
  assign p5_res7__263_comb = p4_literal_1076345[p5_res7__262_comb] ^ p4_literal_1076347[p5_res7__261_comb] ^ p4_literal_1076349[p5_res7__260_comb] ^ p5_array_index_1081203_comb ^ p5_array_index_1081204_comb ^ p5_array_index_1081205_comb ^ p5_res7__256_comb ^ p4_literal_1076358[p5_array_index_1081087_comb] ^ p5_array_index_1081088_comb ^ p5_array_index_1081153_comb ^ p5_array_index_1081124_comb ^ p4_literal_1076351[p5_array_index_1081091_comb] ^ p4_literal_1076349[p5_array_index_1081092_comb] ^ p4_literal_1076347[p5_array_index_1081109_comb] ^ p4_literal_1076345[p5_array_index_1081094_comb] ^ p5_array_index_1081111_comb;
  assign p5_array_index_1081641_comb = p4_literal_1076345[p5_array_index_1081625_comb];
  assign p5_array_index_1081642_comb = p4_literal_1076347[p5_array_index_1081626_comb];
  assign p5_array_index_1081643_comb = p4_literal_1076349[p5_array_index_1081627_comb];
  assign p5_array_index_1081644_comb = p4_literal_1076351[p5_array_index_1081628_comb];
  assign p5_array_index_1081645_comb = p4_literal_1076353[p5_array_index_1081629_comb];
  assign p5_array_index_1081646_comb = p4_literal_1076355[p5_array_index_1081630_comb];
  assign p5_array_index_1081647_comb = p4_arr[p5_addedKey__36_comb[79:72]];
  assign p5_array_index_1081649_comb = p4_arr[p5_addedKey__36_comb[63:56]];
  assign p5_array_index_1081216_comb = p4_literal_1076353[p5_res7__259_comb];
  assign p5_array_index_1081217_comb = p4_literal_1076355[p5_res7__258_comb];
  assign p5_res7__576_comb = p5_array_index_1081641_comb ^ p5_array_index_1081642_comb ^ p5_array_index_1081643_comb ^ p5_array_index_1081644_comb ^ p5_array_index_1081645_comb ^ p5_array_index_1081646_comb ^ p5_array_index_1081647_comb ^ p4_literal_1076358[p5_array_index_1081632_comb] ^ p5_array_index_1081649_comb ^ p4_literal_1076355[p5_array_index_1081634_comb] ^ p4_literal_1076353[p5_array_index_1081635_comb] ^ p4_literal_1076351[p5_array_index_1081636_comb] ^ p4_literal_1076349[p5_array_index_1081637_comb] ^ p4_literal_1076347[p5_array_index_1081638_comb] ^ p4_literal_1076345[p5_array_index_1081639_comb] ^ p4_arr[p5_addedKey__36_comb[7:0]];
  assign p5_res7__264_comb = p4_literal_1076345[p5_res7__263_comb] ^ p4_literal_1076347[p5_res7__262_comb] ^ p4_literal_1076349[p5_res7__261_comb] ^ p4_literal_1076351[p5_res7__260_comb] ^ p5_array_index_1081216_comb ^ p5_array_index_1081217_comb ^ p5_res7__257_comb ^ p4_literal_1076358[p5_res7__256_comb] ^ p5_array_index_1081087_comb ^ p5_array_index_1081167_comb ^ p5_array_index_1081138_comb ^ p5_array_index_1081106_comb ^ p4_literal_1076349[p5_array_index_1081091_comb] ^ p4_literal_1076347[p5_array_index_1081092_comb] ^ p4_literal_1076345[p5_array_index_1081109_comb] ^ p5_array_index_1081094_comb;
  assign p5_array_index_1081658_comb = p4_literal_1076345[p5_res7__576_comb];
  assign p5_array_index_1081659_comb = p4_literal_1076347[p5_array_index_1081625_comb];
  assign p5_array_index_1081660_comb = p4_literal_1076349[p5_array_index_1081626_comb];
  assign p5_array_index_1081661_comb = p4_literal_1076351[p5_array_index_1081627_comb];
  assign p5_array_index_1081662_comb = p4_literal_1076353[p5_array_index_1081628_comb];
  assign p5_array_index_1081663_comb = p4_literal_1076355[p5_array_index_1081629_comb];
  assign p5_array_index_1081227_comb = p4_literal_1076353[p5_res7__260_comb];
  assign p5_array_index_1081228_comb = p4_literal_1076355[p5_res7__259_comb];
  assign p5_res7__577_comb = p5_array_index_1081658_comb ^ p5_array_index_1081659_comb ^ p5_array_index_1081660_comb ^ p5_array_index_1081661_comb ^ p5_array_index_1081662_comb ^ p5_array_index_1081663_comb ^ p5_array_index_1081630_comb ^ p4_literal_1076358[p5_array_index_1081647_comb] ^ p5_array_index_1081632_comb ^ p4_literal_1076355[p5_array_index_1081649_comb] ^ p4_literal_1076353[p5_array_index_1081634_comb] ^ p4_literal_1076351[p5_array_index_1081635_comb] ^ p4_literal_1076349[p5_array_index_1081636_comb] ^ p4_literal_1076347[p5_array_index_1081637_comb] ^ p4_literal_1076345[p5_array_index_1081638_comb] ^ p5_array_index_1081639_comb;
  assign p5_res7__265_comb = p4_literal_1076345[p5_res7__264_comb] ^ p4_literal_1076347[p5_res7__263_comb] ^ p4_literal_1076349[p5_res7__262_comb] ^ p4_literal_1076351[p5_res7__261_comb] ^ p5_array_index_1081227_comb ^ p5_array_index_1081228_comb ^ p5_res7__258_comb ^ p4_literal_1076358[p5_res7__257_comb] ^ p5_res7__256_comb ^ p5_array_index_1081180_comb ^ p5_array_index_1081152_comb ^ p5_array_index_1081123_comb ^ p4_literal_1076349[p5_array_index_1081090_comb] ^ p4_literal_1076347[p5_array_index_1081091_comb] ^ p4_literal_1076345[p5_array_index_1081092_comb] ^ p5_array_index_1081109_comb;
  assign p5_array_index_1081673_comb = p4_literal_1076347[p5_res7__576_comb];
  assign p5_array_index_1081674_comb = p4_literal_1076349[p5_array_index_1081625_comb];
  assign p5_array_index_1081675_comb = p4_literal_1076351[p5_array_index_1081626_comb];
  assign p5_array_index_1081676_comb = p4_literal_1076353[p5_array_index_1081627_comb];
  assign p5_array_index_1081677_comb = p4_literal_1076355[p5_array_index_1081628_comb];
  assign p5_array_index_1081239_comb = p4_literal_1076355[p5_res7__260_comb];
  assign p5_res7__578_comb = p4_literal_1076345[p5_res7__577_comb] ^ p5_array_index_1081673_comb ^ p5_array_index_1081674_comb ^ p5_array_index_1081675_comb ^ p5_array_index_1081676_comb ^ p5_array_index_1081677_comb ^ p5_array_index_1081629_comb ^ p4_literal_1076358[p5_array_index_1081630_comb] ^ p5_array_index_1081647_comb ^ p4_literal_1076355[p5_array_index_1081632_comb] ^ p4_literal_1076353[p5_array_index_1081649_comb] ^ p4_literal_1076351[p5_array_index_1081634_comb] ^ p4_literal_1076349[p5_array_index_1081635_comb] ^ p4_literal_1076347[p5_array_index_1081636_comb] ^ p4_literal_1076345[p5_array_index_1081637_comb] ^ p5_array_index_1081638_comb;
  assign p5_res7__266_comb = p4_literal_1076345[p5_res7__265_comb] ^ p4_literal_1076347[p5_res7__264_comb] ^ p4_literal_1076349[p5_res7__263_comb] ^ p4_literal_1076351[p5_res7__262_comb] ^ p4_literal_1076353[p5_res7__261_comb] ^ p5_array_index_1081239_comb ^ p5_res7__259_comb ^ p4_literal_1076358[p5_res7__258_comb] ^ p5_res7__257_comb ^ p5_array_index_1081193_comb ^ p5_array_index_1081166_comb ^ p5_array_index_1081137_comb ^ p5_array_index_1081105_comb ^ p4_literal_1076347[p5_array_index_1081090_comb] ^ p4_literal_1076345[p5_array_index_1081091_comb] ^ p5_array_index_1081092_comb;
  assign p5_array_index_1081687_comb = p4_literal_1076347[p5_res7__577_comb];
  assign p5_array_index_1081688_comb = p4_literal_1076349[p5_res7__576_comb];
  assign p5_array_index_1081689_comb = p4_literal_1076351[p5_array_index_1081625_comb];
  assign p5_array_index_1081690_comb = p4_literal_1076353[p5_array_index_1081626_comb];
  assign p5_array_index_1081691_comb = p4_literal_1076355[p5_array_index_1081627_comb];
  assign p5_array_index_1081249_comb = p4_literal_1076355[p5_res7__261_comb];
  assign p5_res7__579_comb = p4_literal_1076345[p5_res7__578_comb] ^ p5_array_index_1081687_comb ^ p5_array_index_1081688_comb ^ p5_array_index_1081689_comb ^ p5_array_index_1081690_comb ^ p5_array_index_1081691_comb ^ p5_array_index_1081628_comb ^ p4_literal_1076358[p5_array_index_1081629_comb] ^ p5_array_index_1081630_comb ^ p4_literal_1076355[p5_array_index_1081647_comb] ^ p4_literal_1076353[p5_array_index_1081632_comb] ^ p4_literal_1076351[p5_array_index_1081649_comb] ^ p4_literal_1076349[p5_array_index_1081634_comb] ^ p4_literal_1076347[p5_array_index_1081635_comb] ^ p4_literal_1076345[p5_array_index_1081636_comb] ^ p5_array_index_1081637_comb;
  assign p5_res7__267_comb = p4_literal_1076345[p5_res7__266_comb] ^ p4_literal_1076347[p5_res7__265_comb] ^ p4_literal_1076349[p5_res7__264_comb] ^ p4_literal_1076351[p5_res7__263_comb] ^ p4_literal_1076353[p5_res7__262_comb] ^ p5_array_index_1081249_comb ^ p5_res7__260_comb ^ p4_literal_1076358[p5_res7__259_comb] ^ p5_res7__258_comb ^ p5_array_index_1081205_comb ^ p5_array_index_1081179_comb ^ p5_array_index_1081151_comb ^ p5_array_index_1081122_comb ^ p4_literal_1076347[p5_array_index_1081089_comb] ^ p4_literal_1076345[p5_array_index_1081090_comb] ^ p5_array_index_1081091_comb;
  assign p5_array_index_1081702_comb = p4_literal_1076349[p5_res7__577_comb];
  assign p5_array_index_1081703_comb = p4_literal_1076351[p5_res7__576_comb];
  assign p5_array_index_1081704_comb = p4_literal_1076353[p5_array_index_1081625_comb];
  assign p5_array_index_1081705_comb = p4_literal_1076355[p5_array_index_1081626_comb];
  assign p5_res7__580_comb = p4_literal_1076345[p5_res7__579_comb] ^ p4_literal_1076347[p5_res7__578_comb] ^ p5_array_index_1081702_comb ^ p5_array_index_1081703_comb ^ p5_array_index_1081704_comb ^ p5_array_index_1081705_comb ^ p5_array_index_1081627_comb ^ p4_literal_1076358[p5_array_index_1081628_comb] ^ p5_array_index_1081629_comb ^ p5_array_index_1081646_comb ^ p4_literal_1076353[p5_array_index_1081647_comb] ^ p4_literal_1076351[p5_array_index_1081632_comb] ^ p4_literal_1076349[p5_array_index_1081649_comb] ^ p4_literal_1076347[p5_array_index_1081634_comb] ^ p4_literal_1076345[p5_array_index_1081635_comb] ^ p5_array_index_1081636_comb;
  assign p5_res7__268_comb = p4_literal_1076345[p5_res7__267_comb] ^ p4_literal_1076347[p5_res7__266_comb] ^ p4_literal_1076349[p5_res7__265_comb] ^ p4_literal_1076351[p5_res7__264_comb] ^ p4_literal_1076353[p5_res7__263_comb] ^ p4_literal_1076355[p5_res7__262_comb] ^ p5_res7__261_comb ^ p4_literal_1076358[p5_res7__260_comb] ^ p5_res7__259_comb ^ p5_array_index_1081217_comb ^ p5_array_index_1081192_comb ^ p5_array_index_1081165_comb ^ p5_array_index_1081136_comb ^ p5_array_index_1081104_comb ^ p4_literal_1076345[p5_array_index_1081089_comb] ^ p5_array_index_1081090_comb;
  assign p5_array_index_1081715_comb = p4_literal_1076349[p5_res7__578_comb];
  assign p5_array_index_1081716_comb = p4_literal_1076351[p5_res7__577_comb];
  assign p5_array_index_1081717_comb = p4_literal_1076353[p5_res7__576_comb];
  assign p5_array_index_1081718_comb = p4_literal_1076355[p5_array_index_1081625_comb];
  assign p5_res7__581_comb = p4_literal_1076345[p5_res7__580_comb] ^ p4_literal_1076347[p5_res7__579_comb] ^ p5_array_index_1081715_comb ^ p5_array_index_1081716_comb ^ p5_array_index_1081717_comb ^ p5_array_index_1081718_comb ^ p5_array_index_1081626_comb ^ p4_literal_1076358[p5_array_index_1081627_comb] ^ p5_array_index_1081628_comb ^ p5_array_index_1081663_comb ^ p4_literal_1076353[p5_array_index_1081630_comb] ^ p4_literal_1076351[p5_array_index_1081647_comb] ^ p4_literal_1076349[p5_array_index_1081632_comb] ^ p4_literal_1076347[p5_array_index_1081649_comb] ^ p4_literal_1076345[p5_array_index_1081634_comb] ^ p5_array_index_1081635_comb;
  assign p5_res7__269_comb = p4_literal_1076345[p5_res7__268_comb] ^ p4_literal_1076347[p5_res7__267_comb] ^ p4_literal_1076349[p5_res7__266_comb] ^ p4_literal_1076351[p5_res7__265_comb] ^ p4_literal_1076353[p5_res7__264_comb] ^ p4_literal_1076355[p5_res7__263_comb] ^ p5_res7__262_comb ^ p4_literal_1076358[p5_res7__261_comb] ^ p5_res7__260_comb ^ p5_array_index_1081228_comb ^ p5_array_index_1081204_comb ^ p5_array_index_1081178_comb ^ p5_array_index_1081150_comb ^ p5_array_index_1081121_comb ^ p4_literal_1076345[p5_array_index_1081088_comb] ^ p5_array_index_1081089_comb;
  assign p5_array_index_1081729_comb = p4_literal_1076351[p5_res7__578_comb];
  assign p5_array_index_1081730_comb = p4_literal_1076353[p5_res7__577_comb];
  assign p5_array_index_1081731_comb = p4_literal_1076355[p5_res7__576_comb];
  assign p5_res7__582_comb = p4_literal_1076345[p5_res7__581_comb] ^ p4_literal_1076347[p5_res7__580_comb] ^ p4_literal_1076349[p5_res7__579_comb] ^ p5_array_index_1081729_comb ^ p5_array_index_1081730_comb ^ p5_array_index_1081731_comb ^ p5_array_index_1081625_comb ^ p4_literal_1076358[p5_array_index_1081626_comb] ^ p5_array_index_1081627_comb ^ p5_array_index_1081677_comb ^ p5_array_index_1081645_comb ^ p4_literal_1076351[p5_array_index_1081630_comb] ^ p4_literal_1076349[p5_array_index_1081647_comb] ^ p4_literal_1076347[p5_array_index_1081632_comb] ^ p4_literal_1076345[p5_array_index_1081649_comb] ^ p5_array_index_1081634_comb;
  assign p5_res7__270_comb = p4_literal_1076345[p5_res7__269_comb] ^ p4_literal_1076347[p5_res7__268_comb] ^ p4_literal_1076349[p5_res7__267_comb] ^ p4_literal_1076351[p5_res7__266_comb] ^ p4_literal_1076353[p5_res7__265_comb] ^ p4_literal_1076355[p5_res7__264_comb] ^ p5_res7__263_comb ^ p4_literal_1076358[p5_res7__262_comb] ^ p5_res7__261_comb ^ p5_array_index_1081239_comb ^ p5_array_index_1081216_comb ^ p5_array_index_1081191_comb ^ p5_array_index_1081164_comb ^ p5_array_index_1081135_comb ^ p5_array_index_1081103_comb ^ p5_array_index_1081088_comb;
  assign p5_array_index_1081741_comb = p4_literal_1076351[p5_res7__579_comb];
  assign p5_array_index_1081742_comb = p4_literal_1076353[p5_res7__578_comb];
  assign p5_array_index_1081743_comb = p4_literal_1076355[p5_res7__577_comb];
  assign p5_res7__583_comb = p4_literal_1076345[p5_res7__582_comb] ^ p4_literal_1076347[p5_res7__581_comb] ^ p4_literal_1076349[p5_res7__580_comb] ^ p5_array_index_1081741_comb ^ p5_array_index_1081742_comb ^ p5_array_index_1081743_comb ^ p5_res7__576_comb ^ p4_literal_1076358[p5_array_index_1081625_comb] ^ p5_array_index_1081626_comb ^ p5_array_index_1081691_comb ^ p5_array_index_1081662_comb ^ p4_literal_1076351[p5_array_index_1081629_comb] ^ p4_literal_1076349[p5_array_index_1081630_comb] ^ p4_literal_1076347[p5_array_index_1081647_comb] ^ p4_literal_1076345[p5_array_index_1081632_comb] ^ p5_array_index_1081649_comb;
  assign p5_res7__271_comb = p4_literal_1076345[p5_res7__270_comb] ^ p4_literal_1076347[p5_res7__269_comb] ^ p4_literal_1076349[p5_res7__268_comb] ^ p4_literal_1076351[p5_res7__267_comb] ^ p4_literal_1076353[p5_res7__266_comb] ^ p4_literal_1076355[p5_res7__265_comb] ^ p5_res7__264_comb ^ p4_literal_1076358[p5_res7__263_comb] ^ p5_res7__262_comb ^ p5_array_index_1081249_comb ^ p5_array_index_1081227_comb ^ p5_array_index_1081203_comb ^ p5_array_index_1081177_comb ^ p5_array_index_1081149_comb ^ p5_array_index_1081120_comb ^ p5_array_index_1081087_comb;
  assign p5_array_index_1081754_comb = p4_literal_1076353[p5_res7__579_comb];
  assign p5_array_index_1081755_comb = p4_literal_1076355[p5_res7__578_comb];
  assign p5_res__16_comb = {p5_res7__271_comb, p5_res7__270_comb, p5_res7__269_comb, p5_res7__268_comb, p5_res7__267_comb, p5_res7__266_comb, p5_res7__265_comb, p5_res7__264_comb, p5_res7__263_comb, p5_res7__262_comb, p5_res7__261_comb, p5_res7__260_comb, p5_res7__259_comb, p5_res7__258_comb, p5_res7__257_comb, p5_res7__256_comb};
  assign p5_res7__584_comb = p4_literal_1076345[p5_res7__583_comb] ^ p4_literal_1076347[p5_res7__582_comb] ^ p4_literal_1076349[p5_res7__581_comb] ^ p4_literal_1076351[p5_res7__580_comb] ^ p5_array_index_1081754_comb ^ p5_array_index_1081755_comb ^ p5_res7__577_comb ^ p4_literal_1076358[p5_res7__576_comb] ^ p5_array_index_1081625_comb ^ p5_array_index_1081705_comb ^ p5_array_index_1081676_comb ^ p5_array_index_1081644_comb ^ p4_literal_1076349[p5_array_index_1081629_comb] ^ p4_literal_1076347[p5_array_index_1081630_comb] ^ p4_literal_1076345[p5_array_index_1081647_comb] ^ p5_array_index_1081632_comb;
  assign p5_xor_1081289_comb = p5_res__16_comb ^ p5_k5_comb;
  assign p5_array_index_1081765_comb = p4_literal_1076353[p5_res7__580_comb];
  assign p5_array_index_1081766_comb = p4_literal_1076355[p5_res7__579_comb];
  assign p5_addedKey__58_comb = p5_xor_1081289_comb ^ 128'hf335_80c8_d79a_5862_237b_38e3_375c_bf12;
  assign p5_res7__585_comb = p4_literal_1076345[p5_res7__584_comb] ^ p4_literal_1076347[p5_res7__583_comb] ^ p4_literal_1076349[p5_res7__582_comb] ^ p4_literal_1076351[p5_res7__581_comb] ^ p5_array_index_1081765_comb ^ p5_array_index_1081766_comb ^ p5_res7__578_comb ^ p4_literal_1076358[p5_res7__577_comb] ^ p5_res7__576_comb ^ p5_array_index_1081718_comb ^ p5_array_index_1081690_comb ^ p5_array_index_1081661_comb ^ p4_literal_1076349[p5_array_index_1081628_comb] ^ p4_literal_1076347[p5_array_index_1081629_comb] ^ p4_literal_1076345[p5_array_index_1081630_comb] ^ p5_array_index_1081647_comb;
  assign p5_array_index_1081777_comb = p4_literal_1076355[p5_res7__580_comb];
  assign p5_array_index_1081305_comb = p4_arr[p5_addedKey__58_comb[127:120]];
  assign p5_array_index_1081306_comb = p4_arr[p5_addedKey__58_comb[119:112]];
  assign p5_array_index_1081307_comb = p4_arr[p5_addedKey__58_comb[111:104]];
  assign p5_array_index_1081308_comb = p4_arr[p5_addedKey__58_comb[103:96]];
  assign p5_array_index_1081309_comb = p4_arr[p5_addedKey__58_comb[95:88]];
  assign p5_array_index_1081310_comb = p4_arr[p5_addedKey__58_comb[87:80]];
  assign p5_array_index_1081312_comb = p4_arr[p5_addedKey__58_comb[71:64]];
  assign p5_array_index_1081314_comb = p4_arr[p5_addedKey__58_comb[55:48]];
  assign p5_array_index_1081315_comb = p4_arr[p5_addedKey__58_comb[47:40]];
  assign p5_array_index_1081316_comb = p4_arr[p5_addedKey__58_comb[39:32]];
  assign p5_array_index_1081317_comb = p4_arr[p5_addedKey__58_comb[31:24]];
  assign p5_array_index_1081318_comb = p4_arr[p5_addedKey__58_comb[23:16]];
  assign p5_array_index_1081319_comb = p4_arr[p5_addedKey__58_comb[15:8]];
  assign p5_res7__586_comb = p4_literal_1076345[p5_res7__585_comb] ^ p4_literal_1076347[p5_res7__584_comb] ^ p4_literal_1076349[p5_res7__583_comb] ^ p4_literal_1076351[p5_res7__582_comb] ^ p4_literal_1076353[p5_res7__581_comb] ^ p5_array_index_1081777_comb ^ p5_res7__579_comb ^ p4_literal_1076358[p5_res7__578_comb] ^ p5_res7__577_comb ^ p5_array_index_1081731_comb ^ p5_array_index_1081704_comb ^ p5_array_index_1081675_comb ^ p5_array_index_1081643_comb ^ p4_literal_1076347[p5_array_index_1081628_comb] ^ p4_literal_1076345[p5_array_index_1081629_comb] ^ p5_array_index_1081630_comb;
  assign p5_array_index_1081321_comb = p4_literal_1076345[p5_array_index_1081305_comb];
  assign p5_array_index_1081322_comb = p4_literal_1076347[p5_array_index_1081306_comb];
  assign p5_array_index_1081323_comb = p4_literal_1076349[p5_array_index_1081307_comb];
  assign p5_array_index_1081324_comb = p4_literal_1076351[p5_array_index_1081308_comb];
  assign p5_array_index_1081325_comb = p4_literal_1076353[p5_array_index_1081309_comb];
  assign p5_array_index_1081326_comb = p4_literal_1076355[p5_array_index_1081310_comb];
  assign p5_array_index_1081327_comb = p4_arr[p5_addedKey__58_comb[79:72]];
  assign p5_array_index_1081329_comb = p4_arr[p5_addedKey__58_comb[63:56]];
  assign p5_array_index_1081787_comb = p4_literal_1076355[p5_res7__581_comb];
  assign p5_res7__272_comb = p5_array_index_1081321_comb ^ p5_array_index_1081322_comb ^ p5_array_index_1081323_comb ^ p5_array_index_1081324_comb ^ p5_array_index_1081325_comb ^ p5_array_index_1081326_comb ^ p5_array_index_1081327_comb ^ p4_literal_1076358[p5_array_index_1081312_comb] ^ p5_array_index_1081329_comb ^ p4_literal_1076355[p5_array_index_1081314_comb] ^ p4_literal_1076353[p5_array_index_1081315_comb] ^ p4_literal_1076351[p5_array_index_1081316_comb] ^ p4_literal_1076349[p5_array_index_1081317_comb] ^ p4_literal_1076347[p5_array_index_1081318_comb] ^ p4_literal_1076345[p5_array_index_1081319_comb] ^ p4_arr[p5_addedKey__58_comb[7:0]];
  assign p5_res7__587_comb = p4_literal_1076345[p5_res7__586_comb] ^ p4_literal_1076347[p5_res7__585_comb] ^ p4_literal_1076349[p5_res7__584_comb] ^ p4_literal_1076351[p5_res7__583_comb] ^ p4_literal_1076353[p5_res7__582_comb] ^ p5_array_index_1081787_comb ^ p5_res7__580_comb ^ p4_literal_1076358[p5_res7__579_comb] ^ p5_res7__578_comb ^ p5_array_index_1081743_comb ^ p5_array_index_1081717_comb ^ p5_array_index_1081689_comb ^ p5_array_index_1081660_comb ^ p4_literal_1076347[p5_array_index_1081627_comb] ^ p4_literal_1076345[p5_array_index_1081628_comb] ^ p5_array_index_1081629_comb;
  assign p5_array_index_1081338_comb = p4_literal_1076345[p5_res7__272_comb];
  assign p5_array_index_1081339_comb = p4_literal_1076347[p5_array_index_1081305_comb];
  assign p5_array_index_1081340_comb = p4_literal_1076349[p5_array_index_1081306_comb];
  assign p5_array_index_1081341_comb = p4_literal_1076351[p5_array_index_1081307_comb];
  assign p5_array_index_1081342_comb = p4_literal_1076353[p5_array_index_1081308_comb];
  assign p5_array_index_1081343_comb = p4_literal_1076355[p5_array_index_1081309_comb];
  assign p5_res7__273_comb = p5_array_index_1081338_comb ^ p5_array_index_1081339_comb ^ p5_array_index_1081340_comb ^ p5_array_index_1081341_comb ^ p5_array_index_1081342_comb ^ p5_array_index_1081343_comb ^ p5_array_index_1081310_comb ^ p4_literal_1076358[p5_array_index_1081327_comb] ^ p5_array_index_1081312_comb ^ p4_literal_1076355[p5_array_index_1081329_comb] ^ p4_literal_1076353[p5_array_index_1081314_comb] ^ p4_literal_1076351[p5_array_index_1081315_comb] ^ p4_literal_1076349[p5_array_index_1081316_comb] ^ p4_literal_1076347[p5_array_index_1081317_comb] ^ p4_literal_1076345[p5_array_index_1081318_comb] ^ p5_array_index_1081319_comb;
  assign p5_res7__588_comb = p4_literal_1076345[p5_res7__587_comb] ^ p4_literal_1076347[p5_res7__586_comb] ^ p4_literal_1076349[p5_res7__585_comb] ^ p4_literal_1076351[p5_res7__584_comb] ^ p4_literal_1076353[p5_res7__583_comb] ^ p4_literal_1076355[p5_res7__582_comb] ^ p5_res7__581_comb ^ p4_literal_1076358[p5_res7__580_comb] ^ p5_res7__579_comb ^ p5_array_index_1081755_comb ^ p5_array_index_1081730_comb ^ p5_array_index_1081703_comb ^ p5_array_index_1081674_comb ^ p5_array_index_1081642_comb ^ p4_literal_1076345[p5_array_index_1081627_comb] ^ p5_array_index_1081628_comb;
  assign p5_array_index_1081353_comb = p4_literal_1076347[p5_res7__272_comb];
  assign p5_array_index_1081354_comb = p4_literal_1076349[p5_array_index_1081305_comb];
  assign p5_array_index_1081355_comb = p4_literal_1076351[p5_array_index_1081306_comb];
  assign p5_array_index_1081356_comb = p4_literal_1076353[p5_array_index_1081307_comb];
  assign p5_array_index_1081357_comb = p4_literal_1076355[p5_array_index_1081308_comb];
  assign p5_res7__274_comb = p4_literal_1076345[p5_res7__273_comb] ^ p5_array_index_1081353_comb ^ p5_array_index_1081354_comb ^ p5_array_index_1081355_comb ^ p5_array_index_1081356_comb ^ p5_array_index_1081357_comb ^ p5_array_index_1081309_comb ^ p4_literal_1076358[p5_array_index_1081310_comb] ^ p5_array_index_1081327_comb ^ p4_literal_1076355[p5_array_index_1081312_comb] ^ p4_literal_1076353[p5_array_index_1081329_comb] ^ p4_literal_1076351[p5_array_index_1081314_comb] ^ p4_literal_1076349[p5_array_index_1081315_comb] ^ p4_literal_1076347[p5_array_index_1081316_comb] ^ p4_literal_1076345[p5_array_index_1081317_comb] ^ p5_array_index_1081318_comb;
  assign p5_res7__589_comb = p4_literal_1076345[p5_res7__588_comb] ^ p4_literal_1076347[p5_res7__587_comb] ^ p4_literal_1076349[p5_res7__586_comb] ^ p4_literal_1076351[p5_res7__585_comb] ^ p4_literal_1076353[p5_res7__584_comb] ^ p4_literal_1076355[p5_res7__583_comb] ^ p5_res7__582_comb ^ p4_literal_1076358[p5_res7__581_comb] ^ p5_res7__580_comb ^ p5_array_index_1081766_comb ^ p5_array_index_1081742_comb ^ p5_array_index_1081716_comb ^ p5_array_index_1081688_comb ^ p5_array_index_1081659_comb ^ p4_literal_1076345[p5_array_index_1081626_comb] ^ p5_array_index_1081627_comb;
  assign p5_array_index_1081367_comb = p4_literal_1076347[p5_res7__273_comb];
  assign p5_array_index_1081368_comb = p4_literal_1076349[p5_res7__272_comb];
  assign p5_array_index_1081369_comb = p4_literal_1076351[p5_array_index_1081305_comb];
  assign p5_array_index_1081370_comb = p4_literal_1076353[p5_array_index_1081306_comb];
  assign p5_array_index_1081371_comb = p4_literal_1076355[p5_array_index_1081307_comb];
  assign p5_res7__275_comb = p4_literal_1076345[p5_res7__274_comb] ^ p5_array_index_1081367_comb ^ p5_array_index_1081368_comb ^ p5_array_index_1081369_comb ^ p5_array_index_1081370_comb ^ p5_array_index_1081371_comb ^ p5_array_index_1081308_comb ^ p4_literal_1076358[p5_array_index_1081309_comb] ^ p5_array_index_1081310_comb ^ p4_literal_1076355[p5_array_index_1081327_comb] ^ p4_literal_1076353[p5_array_index_1081312_comb] ^ p4_literal_1076351[p5_array_index_1081329_comb] ^ p4_literal_1076349[p5_array_index_1081314_comb] ^ p4_literal_1076347[p5_array_index_1081315_comb] ^ p4_literal_1076345[p5_array_index_1081316_comb] ^ p5_array_index_1081317_comb;
  assign p5_res7__590_comb = p4_literal_1076345[p5_res7__589_comb] ^ p4_literal_1076347[p5_res7__588_comb] ^ p4_literal_1076349[p5_res7__587_comb] ^ p4_literal_1076351[p5_res7__586_comb] ^ p4_literal_1076353[p5_res7__585_comb] ^ p4_literal_1076355[p5_res7__584_comb] ^ p5_res7__583_comb ^ p4_literal_1076358[p5_res7__582_comb] ^ p5_res7__581_comb ^ p5_array_index_1081777_comb ^ p5_array_index_1081754_comb ^ p5_array_index_1081729_comb ^ p5_array_index_1081702_comb ^ p5_array_index_1081673_comb ^ p5_array_index_1081641_comb ^ p5_array_index_1081626_comb;
  assign p5_array_index_1081382_comb = p4_literal_1076349[p5_res7__273_comb];
  assign p5_array_index_1081383_comb = p4_literal_1076351[p5_res7__272_comb];
  assign p5_array_index_1081384_comb = p4_literal_1076353[p5_array_index_1081305_comb];
  assign p5_array_index_1081385_comb = p4_literal_1076355[p5_array_index_1081306_comb];
  assign p5_res7__276_comb = p4_literal_1076345[p5_res7__275_comb] ^ p4_literal_1076347[p5_res7__274_comb] ^ p5_array_index_1081382_comb ^ p5_array_index_1081383_comb ^ p5_array_index_1081384_comb ^ p5_array_index_1081385_comb ^ p5_array_index_1081307_comb ^ p4_literal_1076358[p5_array_index_1081308_comb] ^ p5_array_index_1081309_comb ^ p5_array_index_1081326_comb ^ p4_literal_1076353[p5_array_index_1081327_comb] ^ p4_literal_1076351[p5_array_index_1081312_comb] ^ p4_literal_1076349[p5_array_index_1081329_comb] ^ p4_literal_1076347[p5_array_index_1081314_comb] ^ p4_literal_1076345[p5_array_index_1081315_comb] ^ p5_array_index_1081316_comb;
  assign p5_res7__591_comb = p4_literal_1076345[p5_res7__590_comb] ^ p4_literal_1076347[p5_res7__589_comb] ^ p4_literal_1076349[p5_res7__588_comb] ^ p4_literal_1076351[p5_res7__587_comb] ^ p4_literal_1076353[p5_res7__586_comb] ^ p4_literal_1076355[p5_res7__585_comb] ^ p5_res7__584_comb ^ p4_literal_1076358[p5_res7__583_comb] ^ p5_res7__582_comb ^ p5_array_index_1081787_comb ^ p5_array_index_1081765_comb ^ p5_array_index_1081741_comb ^ p5_array_index_1081715_comb ^ p5_array_index_1081687_comb ^ p5_array_index_1081658_comb ^ p5_array_index_1081625_comb;
  assign p5_array_index_1081395_comb = p4_literal_1076349[p5_res7__274_comb];
  assign p5_array_index_1081396_comb = p4_literal_1076351[p5_res7__273_comb];
  assign p5_array_index_1081397_comb = p4_literal_1076353[p5_res7__272_comb];
  assign p5_array_index_1081398_comb = p4_literal_1076355[p5_array_index_1081305_comb];
  assign p5_res__36_comb = {p5_res7__591_comb, p5_res7__590_comb, p5_res7__589_comb, p5_res7__588_comb, p5_res7__587_comb, p5_res7__586_comb, p5_res7__585_comb, p5_res7__584_comb, p5_res7__583_comb, p5_res7__582_comb, p5_res7__581_comb, p5_res7__580_comb, p5_res7__579_comb, p5_res7__578_comb, p5_res7__577_comb, p5_res7__576_comb};
  assign p5_res7__277_comb = p4_literal_1076345[p5_res7__276_comb] ^ p4_literal_1076347[p5_res7__275_comb] ^ p5_array_index_1081395_comb ^ p5_array_index_1081396_comb ^ p5_array_index_1081397_comb ^ p5_array_index_1081398_comb ^ p5_array_index_1081306_comb ^ p4_literal_1076358[p5_array_index_1081307_comb] ^ p5_array_index_1081308_comb ^ p5_array_index_1081343_comb ^ p4_literal_1076353[p5_array_index_1081310_comb] ^ p4_literal_1076351[p5_array_index_1081327_comb] ^ p4_literal_1076349[p5_array_index_1081312_comb] ^ p4_literal_1076347[p5_array_index_1081329_comb] ^ p4_literal_1076345[p5_array_index_1081314_comb] ^ p5_array_index_1081315_comb;
  assign p5_addedKey__37_comb = p5_k5_comb ^ p5_res__36_comb;
  assign p5_array_index_1081409_comb = p4_literal_1076351[p5_res7__274_comb];
  assign p5_array_index_1081410_comb = p4_literal_1076353[p5_res7__273_comb];
  assign p5_array_index_1081411_comb = p4_literal_1076355[p5_res7__272_comb];
  assign p5_res7__278_comb = p4_literal_1076345[p5_res7__277_comb] ^ p4_literal_1076347[p5_res7__276_comb] ^ p4_literal_1076349[p5_res7__275_comb] ^ p5_array_index_1081409_comb ^ p5_array_index_1081410_comb ^ p5_array_index_1081411_comb ^ p5_array_index_1081305_comb ^ p4_literal_1076358[p5_array_index_1081306_comb] ^ p5_array_index_1081307_comb ^ p5_array_index_1081357_comb ^ p5_array_index_1081325_comb ^ p4_literal_1076351[p5_array_index_1081310_comb] ^ p4_literal_1076349[p5_array_index_1081327_comb] ^ p4_literal_1076347[p5_array_index_1081312_comb] ^ p4_literal_1076345[p5_array_index_1081329_comb] ^ p5_array_index_1081314_comb;
  assign p5_array_index_1081841_comb = p4_arr[p5_addedKey__37_comb[127:120]];
  assign p5_array_index_1081842_comb = p4_arr[p5_addedKey__37_comb[119:112]];
  assign p5_array_index_1081843_comb = p4_arr[p5_addedKey__37_comb[111:104]];
  assign p5_array_index_1081844_comb = p4_arr[p5_addedKey__37_comb[103:96]];
  assign p5_array_index_1081845_comb = p4_arr[p5_addedKey__37_comb[95:88]];
  assign p5_array_index_1081846_comb = p4_arr[p5_addedKey__37_comb[87:80]];
  assign p5_array_index_1081848_comb = p4_arr[p5_addedKey__37_comb[71:64]];
  assign p5_array_index_1081850_comb = p4_arr[p5_addedKey__37_comb[55:48]];
  assign p5_array_index_1081851_comb = p4_arr[p5_addedKey__37_comb[47:40]];
  assign p5_array_index_1081852_comb = p4_arr[p5_addedKey__37_comb[39:32]];
  assign p5_array_index_1081853_comb = p4_arr[p5_addedKey__37_comb[31:24]];
  assign p5_array_index_1081854_comb = p4_arr[p5_addedKey__37_comb[23:16]];
  assign p5_array_index_1081855_comb = p4_arr[p5_addedKey__37_comb[15:8]];
  assign p5_array_index_1081421_comb = p4_literal_1076351[p5_res7__275_comb];
  assign p5_array_index_1081422_comb = p4_literal_1076353[p5_res7__274_comb];
  assign p5_array_index_1081423_comb = p4_literal_1076355[p5_res7__273_comb];
  assign p5_array_index_1081857_comb = p4_literal_1076345[p5_array_index_1081841_comb];
  assign p5_array_index_1081858_comb = p4_literal_1076347[p5_array_index_1081842_comb];
  assign p5_array_index_1081859_comb = p4_literal_1076349[p5_array_index_1081843_comb];
  assign p5_array_index_1081860_comb = p4_literal_1076351[p5_array_index_1081844_comb];
  assign p5_array_index_1081861_comb = p4_literal_1076353[p5_array_index_1081845_comb];
  assign p5_array_index_1081862_comb = p4_literal_1076355[p5_array_index_1081846_comb];
  assign p5_array_index_1081863_comb = p4_arr[p5_addedKey__37_comb[79:72]];
  assign p5_array_index_1081865_comb = p4_arr[p5_addedKey__37_comb[63:56]];
  assign p5_res7__279_comb = p4_literal_1076345[p5_res7__278_comb] ^ p4_literal_1076347[p5_res7__277_comb] ^ p4_literal_1076349[p5_res7__276_comb] ^ p5_array_index_1081421_comb ^ p5_array_index_1081422_comb ^ p5_array_index_1081423_comb ^ p5_res7__272_comb ^ p4_literal_1076358[p5_array_index_1081305_comb] ^ p5_array_index_1081306_comb ^ p5_array_index_1081371_comb ^ p5_array_index_1081342_comb ^ p4_literal_1076351[p5_array_index_1081309_comb] ^ p4_literal_1076349[p5_array_index_1081310_comb] ^ p4_literal_1076347[p5_array_index_1081327_comb] ^ p4_literal_1076345[p5_array_index_1081312_comb] ^ p5_array_index_1081329_comb;
  assign p5_res7__592_comb = p5_array_index_1081857_comb ^ p5_array_index_1081858_comb ^ p5_array_index_1081859_comb ^ p5_array_index_1081860_comb ^ p5_array_index_1081861_comb ^ p5_array_index_1081862_comb ^ p5_array_index_1081863_comb ^ p4_literal_1076358[p5_array_index_1081848_comb] ^ p5_array_index_1081865_comb ^ p4_literal_1076355[p5_array_index_1081850_comb] ^ p4_literal_1076353[p5_array_index_1081851_comb] ^ p4_literal_1076351[p5_array_index_1081852_comb] ^ p4_literal_1076349[p5_array_index_1081853_comb] ^ p4_literal_1076347[p5_array_index_1081854_comb] ^ p4_literal_1076345[p5_array_index_1081855_comb] ^ p4_arr[p5_addedKey__37_comb[7:0]];
  assign p5_array_index_1081434_comb = p4_literal_1076353[p5_res7__275_comb];
  assign p5_array_index_1081435_comb = p4_literal_1076355[p5_res7__274_comb];
  assign p5_array_index_1081874_comb = p4_literal_1076345[p5_res7__592_comb];
  assign p5_array_index_1081875_comb = p4_literal_1076347[p5_array_index_1081841_comb];
  assign p5_array_index_1081876_comb = p4_literal_1076349[p5_array_index_1081842_comb];
  assign p5_array_index_1081877_comb = p4_literal_1076351[p5_array_index_1081843_comb];
  assign p5_array_index_1081878_comb = p4_literal_1076353[p5_array_index_1081844_comb];
  assign p5_array_index_1081879_comb = p4_literal_1076355[p5_array_index_1081845_comb];
  assign p5_res7__280_comb = p4_literal_1076345[p5_res7__279_comb] ^ p4_literal_1076347[p5_res7__278_comb] ^ p4_literal_1076349[p5_res7__277_comb] ^ p4_literal_1076351[p5_res7__276_comb] ^ p5_array_index_1081434_comb ^ p5_array_index_1081435_comb ^ p5_res7__273_comb ^ p4_literal_1076358[p5_res7__272_comb] ^ p5_array_index_1081305_comb ^ p5_array_index_1081385_comb ^ p5_array_index_1081356_comb ^ p5_array_index_1081324_comb ^ p4_literal_1076349[p5_array_index_1081309_comb] ^ p4_literal_1076347[p5_array_index_1081310_comb] ^ p4_literal_1076345[p5_array_index_1081327_comb] ^ p5_array_index_1081312_comb;
  assign p5_res7__593_comb = p5_array_index_1081874_comb ^ p5_array_index_1081875_comb ^ p5_array_index_1081876_comb ^ p5_array_index_1081877_comb ^ p5_array_index_1081878_comb ^ p5_array_index_1081879_comb ^ p5_array_index_1081846_comb ^ p4_literal_1076358[p5_array_index_1081863_comb] ^ p5_array_index_1081848_comb ^ p4_literal_1076355[p5_array_index_1081865_comb] ^ p4_literal_1076353[p5_array_index_1081850_comb] ^ p4_literal_1076351[p5_array_index_1081851_comb] ^ p4_literal_1076349[p5_array_index_1081852_comb] ^ p4_literal_1076347[p5_array_index_1081853_comb] ^ p4_literal_1076345[p5_array_index_1081854_comb] ^ p5_array_index_1081855_comb;
  assign p5_array_index_1081445_comb = p4_literal_1076353[p5_res7__276_comb];
  assign p5_array_index_1081446_comb = p4_literal_1076355[p5_res7__275_comb];
  assign p5_array_index_1081889_comb = p4_literal_1076347[p5_res7__592_comb];
  assign p5_array_index_1081890_comb = p4_literal_1076349[p5_array_index_1081841_comb];
  assign p5_array_index_1081891_comb = p4_literal_1076351[p5_array_index_1081842_comb];
  assign p5_array_index_1081892_comb = p4_literal_1076353[p5_array_index_1081843_comb];
  assign p5_array_index_1081893_comb = p4_literal_1076355[p5_array_index_1081844_comb];
  assign p5_res7__281_comb = p4_literal_1076345[p5_res7__280_comb] ^ p4_literal_1076347[p5_res7__279_comb] ^ p4_literal_1076349[p5_res7__278_comb] ^ p4_literal_1076351[p5_res7__277_comb] ^ p5_array_index_1081445_comb ^ p5_array_index_1081446_comb ^ p5_res7__274_comb ^ p4_literal_1076358[p5_res7__273_comb] ^ p5_res7__272_comb ^ p5_array_index_1081398_comb ^ p5_array_index_1081370_comb ^ p5_array_index_1081341_comb ^ p4_literal_1076349[p5_array_index_1081308_comb] ^ p4_literal_1076347[p5_array_index_1081309_comb] ^ p4_literal_1076345[p5_array_index_1081310_comb] ^ p5_array_index_1081327_comb;
  assign p5_res7__594_comb = p4_literal_1076345[p5_res7__593_comb] ^ p5_array_index_1081889_comb ^ p5_array_index_1081890_comb ^ p5_array_index_1081891_comb ^ p5_array_index_1081892_comb ^ p5_array_index_1081893_comb ^ p5_array_index_1081845_comb ^ p4_literal_1076358[p5_array_index_1081846_comb] ^ p5_array_index_1081863_comb ^ p4_literal_1076355[p5_array_index_1081848_comb] ^ p4_literal_1076353[p5_array_index_1081865_comb] ^ p4_literal_1076351[p5_array_index_1081850_comb] ^ p4_literal_1076349[p5_array_index_1081851_comb] ^ p4_literal_1076347[p5_array_index_1081852_comb] ^ p4_literal_1076345[p5_array_index_1081853_comb] ^ p5_array_index_1081854_comb;
  assign p5_array_index_1081457_comb = p4_literal_1076355[p5_res7__276_comb];
  assign p5_array_index_1081903_comb = p4_literal_1076347[p5_res7__593_comb];
  assign p5_array_index_1081904_comb = p4_literal_1076349[p5_res7__592_comb];
  assign p5_array_index_1081905_comb = p4_literal_1076351[p5_array_index_1081841_comb];
  assign p5_array_index_1081906_comb = p4_literal_1076353[p5_array_index_1081842_comb];
  assign p5_array_index_1081907_comb = p4_literal_1076355[p5_array_index_1081843_comb];
  assign p5_res7__282_comb = p4_literal_1076345[p5_res7__281_comb] ^ p4_literal_1076347[p5_res7__280_comb] ^ p4_literal_1076349[p5_res7__279_comb] ^ p4_literal_1076351[p5_res7__278_comb] ^ p4_literal_1076353[p5_res7__277_comb] ^ p5_array_index_1081457_comb ^ p5_res7__275_comb ^ p4_literal_1076358[p5_res7__274_comb] ^ p5_res7__273_comb ^ p5_array_index_1081411_comb ^ p5_array_index_1081384_comb ^ p5_array_index_1081355_comb ^ p5_array_index_1081323_comb ^ p4_literal_1076347[p5_array_index_1081308_comb] ^ p4_literal_1076345[p5_array_index_1081309_comb] ^ p5_array_index_1081310_comb;
  assign p5_res7__595_comb = p4_literal_1076345[p5_res7__594_comb] ^ p5_array_index_1081903_comb ^ p5_array_index_1081904_comb ^ p5_array_index_1081905_comb ^ p5_array_index_1081906_comb ^ p5_array_index_1081907_comb ^ p5_array_index_1081844_comb ^ p4_literal_1076358[p5_array_index_1081845_comb] ^ p5_array_index_1081846_comb ^ p4_literal_1076355[p5_array_index_1081863_comb] ^ p4_literal_1076353[p5_array_index_1081848_comb] ^ p4_literal_1076351[p5_array_index_1081865_comb] ^ p4_literal_1076349[p5_array_index_1081850_comb] ^ p4_literal_1076347[p5_array_index_1081851_comb] ^ p4_literal_1076345[p5_array_index_1081852_comb] ^ p5_array_index_1081853_comb;
  assign p5_array_index_1081467_comb = p4_literal_1076355[p5_res7__277_comb];
  assign p5_array_index_1081918_comb = p4_literal_1076349[p5_res7__593_comb];
  assign p5_array_index_1081919_comb = p4_literal_1076351[p5_res7__592_comb];
  assign p5_array_index_1081920_comb = p4_literal_1076353[p5_array_index_1081841_comb];
  assign p5_array_index_1081921_comb = p4_literal_1076355[p5_array_index_1081842_comb];
  assign p5_res7__283_comb = p4_literal_1076345[p5_res7__282_comb] ^ p4_literal_1076347[p5_res7__281_comb] ^ p4_literal_1076349[p5_res7__280_comb] ^ p4_literal_1076351[p5_res7__279_comb] ^ p4_literal_1076353[p5_res7__278_comb] ^ p5_array_index_1081467_comb ^ p5_res7__276_comb ^ p4_literal_1076358[p5_res7__275_comb] ^ p5_res7__274_comb ^ p5_array_index_1081423_comb ^ p5_array_index_1081397_comb ^ p5_array_index_1081369_comb ^ p5_array_index_1081340_comb ^ p4_literal_1076347[p5_array_index_1081307_comb] ^ p4_literal_1076345[p5_array_index_1081308_comb] ^ p5_array_index_1081309_comb;
  assign p5_res7__596_comb = p4_literal_1076345[p5_res7__595_comb] ^ p4_literal_1076347[p5_res7__594_comb] ^ p5_array_index_1081918_comb ^ p5_array_index_1081919_comb ^ p5_array_index_1081920_comb ^ p5_array_index_1081921_comb ^ p5_array_index_1081843_comb ^ p4_literal_1076358[p5_array_index_1081844_comb] ^ p5_array_index_1081845_comb ^ p5_array_index_1081862_comb ^ p4_literal_1076353[p5_array_index_1081863_comb] ^ p4_literal_1076351[p5_array_index_1081848_comb] ^ p4_literal_1076349[p5_array_index_1081865_comb] ^ p4_literal_1076347[p5_array_index_1081850_comb] ^ p4_literal_1076345[p5_array_index_1081851_comb] ^ p5_array_index_1081852_comb;
  assign p5_array_index_1081931_comb = p4_literal_1076349[p5_res7__594_comb];
  assign p5_array_index_1081932_comb = p4_literal_1076351[p5_res7__593_comb];
  assign p5_array_index_1081933_comb = p4_literal_1076353[p5_res7__592_comb];
  assign p5_array_index_1081934_comb = p4_literal_1076355[p5_array_index_1081841_comb];
  assign p5_res7__284_comb = p4_literal_1076345[p5_res7__283_comb] ^ p4_literal_1076347[p5_res7__282_comb] ^ p4_literal_1076349[p5_res7__281_comb] ^ p4_literal_1076351[p5_res7__280_comb] ^ p4_literal_1076353[p5_res7__279_comb] ^ p4_literal_1076355[p5_res7__278_comb] ^ p5_res7__277_comb ^ p4_literal_1076358[p5_res7__276_comb] ^ p5_res7__275_comb ^ p5_array_index_1081435_comb ^ p5_array_index_1081410_comb ^ p5_array_index_1081383_comb ^ p5_array_index_1081354_comb ^ p5_array_index_1081322_comb ^ p4_literal_1076345[p5_array_index_1081307_comb] ^ p5_array_index_1081308_comb;
  assign p5_res7__597_comb = p4_literal_1076345[p5_res7__596_comb] ^ p4_literal_1076347[p5_res7__595_comb] ^ p5_array_index_1081931_comb ^ p5_array_index_1081932_comb ^ p5_array_index_1081933_comb ^ p5_array_index_1081934_comb ^ p5_array_index_1081842_comb ^ p4_literal_1076358[p5_array_index_1081843_comb] ^ p5_array_index_1081844_comb ^ p5_array_index_1081879_comb ^ p4_literal_1076353[p5_array_index_1081846_comb] ^ p4_literal_1076351[p5_array_index_1081863_comb] ^ p4_literal_1076349[p5_array_index_1081848_comb] ^ p4_literal_1076347[p5_array_index_1081865_comb] ^ p4_literal_1076345[p5_array_index_1081850_comb] ^ p5_array_index_1081851_comb;
  assign p5_array_index_1081945_comb = p4_literal_1076351[p5_res7__594_comb];
  assign p5_array_index_1081946_comb = p4_literal_1076353[p5_res7__593_comb];
  assign p5_array_index_1081947_comb = p4_literal_1076355[p5_res7__592_comb];
  assign p5_res7__285_comb = p4_literal_1076345[p5_res7__284_comb] ^ p4_literal_1076347[p5_res7__283_comb] ^ p4_literal_1076349[p5_res7__282_comb] ^ p4_literal_1076351[p5_res7__281_comb] ^ p4_literal_1076353[p5_res7__280_comb] ^ p4_literal_1076355[p5_res7__279_comb] ^ p5_res7__278_comb ^ p4_literal_1076358[p5_res7__277_comb] ^ p5_res7__276_comb ^ p5_array_index_1081446_comb ^ p5_array_index_1081422_comb ^ p5_array_index_1081396_comb ^ p5_array_index_1081368_comb ^ p5_array_index_1081339_comb ^ p4_literal_1076345[p5_array_index_1081306_comb] ^ p5_array_index_1081307_comb;
  assign p5_res7__598_comb = p4_literal_1076345[p5_res7__597_comb] ^ p4_literal_1076347[p5_res7__596_comb] ^ p4_literal_1076349[p5_res7__595_comb] ^ p5_array_index_1081945_comb ^ p5_array_index_1081946_comb ^ p5_array_index_1081947_comb ^ p5_array_index_1081841_comb ^ p4_literal_1076358[p5_array_index_1081842_comb] ^ p5_array_index_1081843_comb ^ p5_array_index_1081893_comb ^ p5_array_index_1081861_comb ^ p4_literal_1076351[p5_array_index_1081846_comb] ^ p4_literal_1076349[p5_array_index_1081863_comb] ^ p4_literal_1076347[p5_array_index_1081848_comb] ^ p4_literal_1076345[p5_array_index_1081865_comb] ^ p5_array_index_1081850_comb;
  assign p5_array_index_1081957_comb = p4_literal_1076351[p5_res7__595_comb];
  assign p5_array_index_1081958_comb = p4_literal_1076353[p5_res7__594_comb];
  assign p5_array_index_1081959_comb = p4_literal_1076355[p5_res7__593_comb];
  assign p5_res7__286_comb = p4_literal_1076345[p5_res7__285_comb] ^ p4_literal_1076347[p5_res7__284_comb] ^ p4_literal_1076349[p5_res7__283_comb] ^ p4_literal_1076351[p5_res7__282_comb] ^ p4_literal_1076353[p5_res7__281_comb] ^ p4_literal_1076355[p5_res7__280_comb] ^ p5_res7__279_comb ^ p4_literal_1076358[p5_res7__278_comb] ^ p5_res7__277_comb ^ p5_array_index_1081457_comb ^ p5_array_index_1081434_comb ^ p5_array_index_1081409_comb ^ p5_array_index_1081382_comb ^ p5_array_index_1081353_comb ^ p5_array_index_1081321_comb ^ p5_array_index_1081306_comb;
  assign p5_res7__599_comb = p4_literal_1076345[p5_res7__598_comb] ^ p4_literal_1076347[p5_res7__597_comb] ^ p4_literal_1076349[p5_res7__596_comb] ^ p5_array_index_1081957_comb ^ p5_array_index_1081958_comb ^ p5_array_index_1081959_comb ^ p5_res7__592_comb ^ p4_literal_1076358[p5_array_index_1081841_comb] ^ p5_array_index_1081842_comb ^ p5_array_index_1081907_comb ^ p5_array_index_1081878_comb ^ p4_literal_1076351[p5_array_index_1081845_comb] ^ p4_literal_1076349[p5_array_index_1081846_comb] ^ p4_literal_1076347[p5_array_index_1081863_comb] ^ p4_literal_1076345[p5_array_index_1081848_comb] ^ p5_array_index_1081865_comb;
  assign p5_array_index_1081970_comb = p4_literal_1076353[p5_res7__595_comb];
  assign p5_array_index_1081971_comb = p4_literal_1076355[p5_res7__594_comb];
  assign p5_res7__287_comb = p4_literal_1076345[p5_res7__286_comb] ^ p4_literal_1076347[p5_res7__285_comb] ^ p4_literal_1076349[p5_res7__284_comb] ^ p4_literal_1076351[p5_res7__283_comb] ^ p4_literal_1076353[p5_res7__282_comb] ^ p4_literal_1076355[p5_res7__281_comb] ^ p5_res7__280_comb ^ p4_literal_1076358[p5_res7__279_comb] ^ p5_res7__278_comb ^ p5_array_index_1081467_comb ^ p5_array_index_1081445_comb ^ p5_array_index_1081421_comb ^ p5_array_index_1081395_comb ^ p5_array_index_1081367_comb ^ p5_array_index_1081338_comb ^ p5_array_index_1081305_comb;
  assign p5_res7__600_comb = p4_literal_1076345[p5_res7__599_comb] ^ p4_literal_1076347[p5_res7__598_comb] ^ p4_literal_1076349[p5_res7__597_comb] ^ p4_literal_1076351[p5_res7__596_comb] ^ p5_array_index_1081970_comb ^ p5_array_index_1081971_comb ^ p5_res7__593_comb ^ p4_literal_1076358[p5_res7__592_comb] ^ p5_array_index_1081841_comb ^ p5_array_index_1081921_comb ^ p5_array_index_1081892_comb ^ p5_array_index_1081860_comb ^ p4_literal_1076349[p5_array_index_1081845_comb] ^ p4_literal_1076347[p5_array_index_1081846_comb] ^ p4_literal_1076345[p5_array_index_1081863_comb] ^ p5_array_index_1081848_comb;
  assign p5_res__17_comb = {p5_res7__287_comb, p5_res7__286_comb, p5_res7__285_comb, p5_res7__284_comb, p5_res7__283_comb, p5_res7__282_comb, p5_res7__281_comb, p5_res7__280_comb, p5_res7__279_comb, p5_res7__278_comb, p5_res7__277_comb, p5_res7__276_comb, p5_res7__275_comb, p5_res7__274_comb, p5_res7__273_comb, p5_res7__272_comb};
  assign p5_array_index_1081981_comb = p4_literal_1076353[p5_res7__596_comb];
  assign p5_array_index_1081982_comb = p4_literal_1076355[p5_res7__595_comb];
  assign p5_xor_1081507_comb = p5_res__17_comb ^ p5_k4_comb;
  assign p5_res7__601_comb = p4_literal_1076345[p5_res7__600_comb] ^ p4_literal_1076347[p5_res7__599_comb] ^ p4_literal_1076349[p5_res7__598_comb] ^ p4_literal_1076351[p5_res7__597_comb] ^ p5_array_index_1081981_comb ^ p5_array_index_1081982_comb ^ p5_res7__594_comb ^ p4_literal_1076358[p5_res7__593_comb] ^ p5_res7__592_comb ^ p5_array_index_1081934_comb ^ p5_array_index_1081906_comb ^ p5_array_index_1081877_comb ^ p4_literal_1076349[p5_array_index_1081844_comb] ^ p4_literal_1076347[p5_array_index_1081845_comb] ^ p4_literal_1076345[p5_array_index_1081846_comb] ^ p5_array_index_1081863_comb;
  assign p5_addedKey__59_comb = p5_xor_1081507_comb ^ 128'h9d97_f6ba_bbd2_22da_7e5c_85f3_ead8_2b13;
  assign p5_array_index_1081993_comb = p4_literal_1076355[p5_res7__596_comb];
  assign p5_res7__602_comb = p4_literal_1076345[p5_res7__601_comb] ^ p4_literal_1076347[p5_res7__600_comb] ^ p4_literal_1076349[p5_res7__599_comb] ^ p4_literal_1076351[p5_res7__598_comb] ^ p4_literal_1076353[p5_res7__597_comb] ^ p5_array_index_1081993_comb ^ p5_res7__595_comb ^ p4_literal_1076358[p5_res7__594_comb] ^ p5_res7__593_comb ^ p5_array_index_1081947_comb ^ p5_array_index_1081920_comb ^ p5_array_index_1081891_comb ^ p5_array_index_1081859_comb ^ p4_literal_1076347[p5_array_index_1081844_comb] ^ p4_literal_1076345[p5_array_index_1081845_comb] ^ p5_array_index_1081846_comb;
  assign p5_array_index_1081523_comb = p4_arr[p5_addedKey__59_comb[127:120]];
  assign p5_array_index_1081524_comb = p4_arr[p5_addedKey__59_comb[119:112]];
  assign p5_array_index_1081525_comb = p4_arr[p5_addedKey__59_comb[111:104]];
  assign p5_array_index_1081526_comb = p4_arr[p5_addedKey__59_comb[103:96]];
  assign p5_array_index_1081527_comb = p4_arr[p5_addedKey__59_comb[95:88]];
  assign p5_array_index_1081528_comb = p4_arr[p5_addedKey__59_comb[87:80]];
  assign p5_array_index_1081530_comb = p4_arr[p5_addedKey__59_comb[71:64]];
  assign p5_array_index_1081532_comb = p4_arr[p5_addedKey__59_comb[55:48]];
  assign p5_array_index_1081533_comb = p4_arr[p5_addedKey__59_comb[47:40]];
  assign p5_array_index_1081534_comb = p4_arr[p5_addedKey__59_comb[39:32]];
  assign p5_array_index_1081535_comb = p4_arr[p5_addedKey__59_comb[31:24]];
  assign p5_array_index_1081536_comb = p4_arr[p5_addedKey__59_comb[23:16]];
  assign p5_array_index_1081537_comb = p4_arr[p5_addedKey__59_comb[15:8]];
  assign p5_array_index_1082003_comb = p4_literal_1076355[p5_res7__597_comb];
  assign p5_array_index_1081539_comb = p4_literal_1076345[p5_array_index_1081523_comb];
  assign p5_array_index_1081540_comb = p4_literal_1076347[p5_array_index_1081524_comb];
  assign p5_array_index_1081541_comb = p4_literal_1076349[p5_array_index_1081525_comb];
  assign p5_array_index_1081542_comb = p4_literal_1076351[p5_array_index_1081526_comb];
  assign p5_array_index_1081543_comb = p4_literal_1076353[p5_array_index_1081527_comb];
  assign p5_array_index_1081544_comb = p4_literal_1076355[p5_array_index_1081528_comb];
  assign p5_array_index_1081545_comb = p4_arr[p5_addedKey__59_comb[79:72]];
  assign p5_array_index_1081547_comb = p4_arr[p5_addedKey__59_comb[63:56]];
  assign p5_res7__603_comb = p4_literal_1076345[p5_res7__602_comb] ^ p4_literal_1076347[p5_res7__601_comb] ^ p4_literal_1076349[p5_res7__600_comb] ^ p4_literal_1076351[p5_res7__599_comb] ^ p4_literal_1076353[p5_res7__598_comb] ^ p5_array_index_1082003_comb ^ p5_res7__596_comb ^ p4_literal_1076358[p5_res7__595_comb] ^ p5_res7__594_comb ^ p5_array_index_1081959_comb ^ p5_array_index_1081933_comb ^ p5_array_index_1081905_comb ^ p5_array_index_1081876_comb ^ p4_literal_1076347[p5_array_index_1081843_comb] ^ p4_literal_1076345[p5_array_index_1081844_comb] ^ p5_array_index_1081845_comb;
  assign p5_res7__288_comb = p5_array_index_1081539_comb ^ p5_array_index_1081540_comb ^ p5_array_index_1081541_comb ^ p5_array_index_1081542_comb ^ p5_array_index_1081543_comb ^ p5_array_index_1081544_comb ^ p5_array_index_1081545_comb ^ p4_literal_1076358[p5_array_index_1081530_comb] ^ p5_array_index_1081547_comb ^ p4_literal_1076355[p5_array_index_1081532_comb] ^ p4_literal_1076353[p5_array_index_1081533_comb] ^ p4_literal_1076351[p5_array_index_1081534_comb] ^ p4_literal_1076349[p5_array_index_1081535_comb] ^ p4_literal_1076347[p5_array_index_1081536_comb] ^ p4_literal_1076345[p5_array_index_1081537_comb] ^ p4_arr[p5_addedKey__59_comb[7:0]];
  assign p5_array_index_1081556_comb = p4_literal_1076345[p5_res7__288_comb];
  assign p5_array_index_1081557_comb = p4_literal_1076347[p5_array_index_1081523_comb];
  assign p5_array_index_1081558_comb = p4_literal_1076349[p5_array_index_1081524_comb];
  assign p5_array_index_1081559_comb = p4_literal_1076351[p5_array_index_1081525_comb];
  assign p5_array_index_1081560_comb = p4_literal_1076353[p5_array_index_1081526_comb];
  assign p5_array_index_1081561_comb = p4_literal_1076355[p5_array_index_1081527_comb];
  assign p5_res7__604_comb = p4_literal_1076345[p5_res7__603_comb] ^ p4_literal_1076347[p5_res7__602_comb] ^ p4_literal_1076349[p5_res7__601_comb] ^ p4_literal_1076351[p5_res7__600_comb] ^ p4_literal_1076353[p5_res7__599_comb] ^ p4_literal_1076355[p5_res7__598_comb] ^ p5_res7__597_comb ^ p4_literal_1076358[p5_res7__596_comb] ^ p5_res7__595_comb ^ p5_array_index_1081971_comb ^ p5_array_index_1081946_comb ^ p5_array_index_1081919_comb ^ p5_array_index_1081890_comb ^ p5_array_index_1081858_comb ^ p4_literal_1076345[p5_array_index_1081843_comb] ^ p5_array_index_1081844_comb;
  assign p5_res7__289_comb = p5_array_index_1081556_comb ^ p5_array_index_1081557_comb ^ p5_array_index_1081558_comb ^ p5_array_index_1081559_comb ^ p5_array_index_1081560_comb ^ p5_array_index_1081561_comb ^ p5_array_index_1081528_comb ^ p4_literal_1076358[p5_array_index_1081545_comb] ^ p5_array_index_1081530_comb ^ p4_literal_1076355[p5_array_index_1081547_comb] ^ p4_literal_1076353[p5_array_index_1081532_comb] ^ p4_literal_1076351[p5_array_index_1081533_comb] ^ p4_literal_1076349[p5_array_index_1081534_comb] ^ p4_literal_1076347[p5_array_index_1081535_comb] ^ p4_literal_1076345[p5_array_index_1081536_comb] ^ p5_array_index_1081537_comb;
  assign p5_array_index_1081571_comb = p4_literal_1076347[p5_res7__288_comb];
  assign p5_array_index_1081572_comb = p4_literal_1076349[p5_array_index_1081523_comb];
  assign p5_array_index_1081573_comb = p4_literal_1076351[p5_array_index_1081524_comb];
  assign p5_array_index_1081574_comb = p4_literal_1076353[p5_array_index_1081525_comb];
  assign p5_array_index_1081575_comb = p4_literal_1076355[p5_array_index_1081526_comb];
  assign p5_res7__605_comb = p4_literal_1076345[p5_res7__604_comb] ^ p4_literal_1076347[p5_res7__603_comb] ^ p4_literal_1076349[p5_res7__602_comb] ^ p4_literal_1076351[p5_res7__601_comb] ^ p4_literal_1076353[p5_res7__600_comb] ^ p4_literal_1076355[p5_res7__599_comb] ^ p5_res7__598_comb ^ p4_literal_1076358[p5_res7__597_comb] ^ p5_res7__596_comb ^ p5_array_index_1081982_comb ^ p5_array_index_1081958_comb ^ p5_array_index_1081932_comb ^ p5_array_index_1081904_comb ^ p5_array_index_1081875_comb ^ p4_literal_1076345[p5_array_index_1081842_comb] ^ p5_array_index_1081843_comb;
  assign p5_res7__290_comb = p4_literal_1076345[p5_res7__289_comb] ^ p5_array_index_1081571_comb ^ p5_array_index_1081572_comb ^ p5_array_index_1081573_comb ^ p5_array_index_1081574_comb ^ p5_array_index_1081575_comb ^ p5_array_index_1081527_comb ^ p4_literal_1076358[p5_array_index_1081528_comb] ^ p5_array_index_1081545_comb ^ p4_literal_1076355[p5_array_index_1081530_comb] ^ p4_literal_1076353[p5_array_index_1081547_comb] ^ p4_literal_1076351[p5_array_index_1081532_comb] ^ p4_literal_1076349[p5_array_index_1081533_comb] ^ p4_literal_1076347[p5_array_index_1081534_comb] ^ p4_literal_1076345[p5_array_index_1081535_comb] ^ p5_array_index_1081536_comb;
  assign p5_array_index_1081585_comb = p4_literal_1076347[p5_res7__289_comb];
  assign p5_array_index_1081586_comb = p4_literal_1076349[p5_res7__288_comb];
  assign p5_array_index_1081587_comb = p4_literal_1076351[p5_array_index_1081523_comb];
  assign p5_array_index_1081588_comb = p4_literal_1076353[p5_array_index_1081524_comb];
  assign p5_array_index_1081589_comb = p4_literal_1076355[p5_array_index_1081525_comb];
  assign p5_res7__606_comb = p4_literal_1076345[p5_res7__605_comb] ^ p4_literal_1076347[p5_res7__604_comb] ^ p4_literal_1076349[p5_res7__603_comb] ^ p4_literal_1076351[p5_res7__602_comb] ^ p4_literal_1076353[p5_res7__601_comb] ^ p4_literal_1076355[p5_res7__600_comb] ^ p5_res7__599_comb ^ p4_literal_1076358[p5_res7__598_comb] ^ p5_res7__597_comb ^ p5_array_index_1081993_comb ^ p5_array_index_1081970_comb ^ p5_array_index_1081945_comb ^ p5_array_index_1081918_comb ^ p5_array_index_1081889_comb ^ p5_array_index_1081857_comb ^ p5_array_index_1081842_comb;
  assign p5_res7__291_comb = p4_literal_1076345[p5_res7__290_comb] ^ p5_array_index_1081585_comb ^ p5_array_index_1081586_comb ^ p5_array_index_1081587_comb ^ p5_array_index_1081588_comb ^ p5_array_index_1081589_comb ^ p5_array_index_1081526_comb ^ p4_literal_1076358[p5_array_index_1081527_comb] ^ p5_array_index_1081528_comb ^ p4_literal_1076355[p5_array_index_1081545_comb] ^ p4_literal_1076353[p5_array_index_1081530_comb] ^ p4_literal_1076351[p5_array_index_1081547_comb] ^ p4_literal_1076349[p5_array_index_1081532_comb] ^ p4_literal_1076347[p5_array_index_1081533_comb] ^ p4_literal_1076345[p5_array_index_1081534_comb] ^ p5_array_index_1081535_comb;
  assign p5_array_index_1081600_comb = p4_literal_1076349[p5_res7__289_comb];
  assign p5_array_index_1081601_comb = p4_literal_1076351[p5_res7__288_comb];
  assign p5_array_index_1081602_comb = p4_literal_1076353[p5_array_index_1081523_comb];
  assign p5_array_index_1081603_comb = p4_literal_1076355[p5_array_index_1081524_comb];
  assign p5_res7__607_comb = p4_literal_1076345[p5_res7__606_comb] ^ p4_literal_1076347[p5_res7__605_comb] ^ p4_literal_1076349[p5_res7__604_comb] ^ p4_literal_1076351[p5_res7__603_comb] ^ p4_literal_1076353[p5_res7__602_comb] ^ p4_literal_1076355[p5_res7__601_comb] ^ p5_res7__600_comb ^ p4_literal_1076358[p5_res7__599_comb] ^ p5_res7__598_comb ^ p5_array_index_1082003_comb ^ p5_array_index_1081981_comb ^ p5_array_index_1081957_comb ^ p5_array_index_1081931_comb ^ p5_array_index_1081903_comb ^ p5_array_index_1081874_comb ^ p5_array_index_1081841_comb;
  assign p5_res7__292_comb = p4_literal_1076345[p5_res7__291_comb] ^ p4_literal_1076347[p5_res7__290_comb] ^ p5_array_index_1081600_comb ^ p5_array_index_1081601_comb ^ p5_array_index_1081602_comb ^ p5_array_index_1081603_comb ^ p5_array_index_1081525_comb ^ p4_literal_1076358[p5_array_index_1081526_comb] ^ p5_array_index_1081527_comb ^ p5_array_index_1081544_comb ^ p4_literal_1076353[p5_array_index_1081545_comb] ^ p4_literal_1076351[p5_array_index_1081530_comb] ^ p4_literal_1076349[p5_array_index_1081547_comb] ^ p4_literal_1076347[p5_array_index_1081532_comb] ^ p4_literal_1076345[p5_array_index_1081533_comb] ^ p5_array_index_1081534_comb;
  assign p5_res__37_comb = {p5_res7__607_comb, p5_res7__606_comb, p5_res7__605_comb, p5_res7__604_comb, p5_res7__603_comb, p5_res7__602_comb, p5_res7__601_comb, p5_res7__600_comb, p5_res7__599_comb, p5_res7__598_comb, p5_res7__597_comb, p5_res7__596_comb, p5_res7__595_comb, p5_res7__594_comb, p5_res7__593_comb, p5_res7__592_comb};

  // Registers for pipe stage 5:
  reg [127:0] p5_xor_1081289;
  reg [127:0] p5_xor_1081507;
  reg [7:0] p5_array_index_1081523;
  reg [7:0] p5_array_index_1081524;
  reg [7:0] p5_array_index_1081525;
  reg [7:0] p5_array_index_1081526;
  reg [7:0] p5_array_index_1081527;
  reg [7:0] p5_array_index_1081528;
  reg [7:0] p5_array_index_1081530;
  reg [7:0] p5_array_index_1081532;
  reg [7:0] p5_array_index_1081533;
  reg [7:0] p5_array_index_1081539;
  reg [7:0] p5_array_index_1081540;
  reg [7:0] p5_array_index_1081541;
  reg [7:0] p5_array_index_1081542;
  reg [7:0] p5_array_index_1081543;
  reg [7:0] p5_array_index_1081545;
  reg [7:0] p5_array_index_1081547;
  reg [7:0] p5_res7__288;
  reg [7:0] p5_array_index_1081556;
  reg [7:0] p5_array_index_1081557;
  reg [7:0] p5_array_index_1081558;
  reg [7:0] p5_array_index_1081559;
  reg [7:0] p5_array_index_1081560;
  reg [7:0] p5_array_index_1081561;
  reg [7:0] p5_res7__289;
  reg [7:0] p5_array_index_1081571;
  reg [7:0] p5_array_index_1081572;
  reg [7:0] p5_array_index_1081573;
  reg [7:0] p5_array_index_1081574;
  reg [7:0] p5_array_index_1081575;
  reg [7:0] p5_res7__290;
  reg [7:0] p5_array_index_1081585;
  reg [7:0] p5_array_index_1081586;
  reg [7:0] p5_array_index_1081587;
  reg [7:0] p5_array_index_1081588;
  reg [7:0] p5_array_index_1081589;
  reg [7:0] p5_res7__291;
  reg [7:0] p5_array_index_1081600;
  reg [7:0] p5_array_index_1081601;
  reg [7:0] p5_array_index_1081602;
  reg [7:0] p5_array_index_1081603;
  reg [7:0] p5_res7__292;
  reg [127:0] p5_res__37;
  reg [7:0] p6_arr[256];
  reg [7:0] p6_literal_1076345[256];
  reg [7:0] p6_literal_1076347[256];
  reg [7:0] p6_literal_1076349[256];
  reg [7:0] p6_literal_1076351[256];
  reg [7:0] p6_literal_1076353[256];
  reg [7:0] p6_literal_1076355[256];
  reg [7:0] p6_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p5_xor_1081289 <= p5_xor_1081289_comb;
    p5_xor_1081507 <= p5_xor_1081507_comb;
    p5_array_index_1081523 <= p5_array_index_1081523_comb;
    p5_array_index_1081524 <= p5_array_index_1081524_comb;
    p5_array_index_1081525 <= p5_array_index_1081525_comb;
    p5_array_index_1081526 <= p5_array_index_1081526_comb;
    p5_array_index_1081527 <= p5_array_index_1081527_comb;
    p5_array_index_1081528 <= p5_array_index_1081528_comb;
    p5_array_index_1081530 <= p5_array_index_1081530_comb;
    p5_array_index_1081532 <= p5_array_index_1081532_comb;
    p5_array_index_1081533 <= p5_array_index_1081533_comb;
    p5_array_index_1081539 <= p5_array_index_1081539_comb;
    p5_array_index_1081540 <= p5_array_index_1081540_comb;
    p5_array_index_1081541 <= p5_array_index_1081541_comb;
    p5_array_index_1081542 <= p5_array_index_1081542_comb;
    p5_array_index_1081543 <= p5_array_index_1081543_comb;
    p5_array_index_1081545 <= p5_array_index_1081545_comb;
    p5_array_index_1081547 <= p5_array_index_1081547_comb;
    p5_res7__288 <= p5_res7__288_comb;
    p5_array_index_1081556 <= p5_array_index_1081556_comb;
    p5_array_index_1081557 <= p5_array_index_1081557_comb;
    p5_array_index_1081558 <= p5_array_index_1081558_comb;
    p5_array_index_1081559 <= p5_array_index_1081559_comb;
    p5_array_index_1081560 <= p5_array_index_1081560_comb;
    p5_array_index_1081561 <= p5_array_index_1081561_comb;
    p5_res7__289 <= p5_res7__289_comb;
    p5_array_index_1081571 <= p5_array_index_1081571_comb;
    p5_array_index_1081572 <= p5_array_index_1081572_comb;
    p5_array_index_1081573 <= p5_array_index_1081573_comb;
    p5_array_index_1081574 <= p5_array_index_1081574_comb;
    p5_array_index_1081575 <= p5_array_index_1081575_comb;
    p5_res7__290 <= p5_res7__290_comb;
    p5_array_index_1081585 <= p5_array_index_1081585_comb;
    p5_array_index_1081586 <= p5_array_index_1081586_comb;
    p5_array_index_1081587 <= p5_array_index_1081587_comb;
    p5_array_index_1081588 <= p5_array_index_1081588_comb;
    p5_array_index_1081589 <= p5_array_index_1081589_comb;
    p5_res7__291 <= p5_res7__291_comb;
    p5_array_index_1081600 <= p5_array_index_1081600_comb;
    p5_array_index_1081601 <= p5_array_index_1081601_comb;
    p5_array_index_1081602 <= p5_array_index_1081602_comb;
    p5_array_index_1081603 <= p5_array_index_1081603_comb;
    p5_res7__292 <= p5_res7__292_comb;
    p5_res__37 <= p5_res__37_comb;
    p6_arr <= p5_arr;
    p6_literal_1076345 <= p5_literal_1076345;
    p6_literal_1076347 <= p5_literal_1076347;
    p6_literal_1076349 <= p5_literal_1076349;
    p6_literal_1076351 <= p5_literal_1076351;
    p6_literal_1076353 <= p5_literal_1076353;
    p6_literal_1076355 <= p5_literal_1076355;
    p6_literal_1076358 <= p5_literal_1076358;
  end

  // ===== Pipe stage 6:
  wire [7:0] p6_array_index_1082149_comb;
  wire [7:0] p6_array_index_1082150_comb;
  wire [7:0] p6_array_index_1082151_comb;
  wire [7:0] p6_array_index_1082152_comb;
  wire [7:0] p6_res7__293_comb;
  wire [7:0] p6_array_index_1082163_comb;
  wire [7:0] p6_array_index_1082164_comb;
  wire [7:0] p6_array_index_1082165_comb;
  wire [7:0] p6_res7__294_comb;
  wire [7:0] p6_array_index_1082175_comb;
  wire [7:0] p6_array_index_1082176_comb;
  wire [7:0] p6_array_index_1082177_comb;
  wire [7:0] p6_res7__295_comb;
  wire [7:0] p6_array_index_1082188_comb;
  wire [7:0] p6_array_index_1082189_comb;
  wire [7:0] p6_res7__296_comb;
  wire [7:0] p6_array_index_1082199_comb;
  wire [7:0] p6_array_index_1082200_comb;
  wire [7:0] p6_res7__297_comb;
  wire [7:0] p6_array_index_1082211_comb;
  wire [7:0] p6_res7__298_comb;
  wire [7:0] p6_array_index_1082221_comb;
  wire [7:0] p6_res7__299_comb;
  wire [7:0] p6_res7__300_comb;
  wire [7:0] p6_res7__301_comb;
  wire [7:0] p6_res7__302_comb;
  wire [7:0] p6_res7__303_comb;
  wire [127:0] p6_res__18_comb;
  wire [127:0] p6_xor_1082261_comb;
  wire [127:0] p6_addedKey__60_comb;
  wire [7:0] p6_array_index_1082277_comb;
  wire [7:0] p6_array_index_1082278_comb;
  wire [7:0] p6_array_index_1082279_comb;
  wire [7:0] p6_array_index_1082280_comb;
  wire [7:0] p6_array_index_1082281_comb;
  wire [7:0] p6_array_index_1082282_comb;
  wire [7:0] p6_array_index_1082284_comb;
  wire [7:0] p6_array_index_1082286_comb;
  wire [7:0] p6_array_index_1082287_comb;
  wire [7:0] p6_array_index_1082288_comb;
  wire [7:0] p6_array_index_1082289_comb;
  wire [7:0] p6_array_index_1082290_comb;
  wire [7:0] p6_array_index_1082291_comb;
  wire [7:0] p6_array_index_1082293_comb;
  wire [7:0] p6_array_index_1082294_comb;
  wire [7:0] p6_array_index_1082295_comb;
  wire [7:0] p6_array_index_1082296_comb;
  wire [7:0] p6_array_index_1082297_comb;
  wire [7:0] p6_array_index_1082298_comb;
  wire [7:0] p6_array_index_1082299_comb;
  wire [7:0] p6_array_index_1082301_comb;
  wire [7:0] p6_res7__304_comb;
  wire [7:0] p6_array_index_1082310_comb;
  wire [7:0] p6_array_index_1082311_comb;
  wire [7:0] p6_array_index_1082312_comb;
  wire [7:0] p6_array_index_1082313_comb;
  wire [7:0] p6_array_index_1082314_comb;
  wire [7:0] p6_array_index_1082315_comb;
  wire [7:0] p6_res7__305_comb;
  wire [7:0] p6_array_index_1082325_comb;
  wire [7:0] p6_array_index_1082326_comb;
  wire [7:0] p6_array_index_1082327_comb;
  wire [7:0] p6_array_index_1082328_comb;
  wire [7:0] p6_array_index_1082329_comb;
  wire [7:0] p6_res7__306_comb;
  wire [7:0] p6_array_index_1082339_comb;
  wire [7:0] p6_array_index_1082340_comb;
  wire [7:0] p6_array_index_1082341_comb;
  wire [7:0] p6_array_index_1082342_comb;
  wire [7:0] p6_array_index_1082343_comb;
  wire [7:0] p6_res7__307_comb;
  wire [7:0] p6_array_index_1082354_comb;
  wire [7:0] p6_array_index_1082355_comb;
  wire [7:0] p6_array_index_1082356_comb;
  wire [7:0] p6_array_index_1082357_comb;
  wire [7:0] p6_res7__308_comb;
  wire [7:0] p6_array_index_1082367_comb;
  wire [7:0] p6_array_index_1082368_comb;
  wire [7:0] p6_array_index_1082369_comb;
  wire [7:0] p6_array_index_1082370_comb;
  wire [7:0] p6_res7__309_comb;
  wire [7:0] p6_array_index_1082381_comb;
  wire [7:0] p6_array_index_1082382_comb;
  wire [7:0] p6_array_index_1082383_comb;
  wire [7:0] p6_res7__310_comb;
  wire [7:0] p6_array_index_1082393_comb;
  wire [7:0] p6_array_index_1082394_comb;
  wire [7:0] p6_array_index_1082395_comb;
  wire [7:0] p6_res7__311_comb;
  wire [7:0] p6_array_index_1082406_comb;
  wire [7:0] p6_array_index_1082407_comb;
  wire [7:0] p6_res7__312_comb;
  wire [7:0] p6_array_index_1082417_comb;
  wire [7:0] p6_array_index_1082418_comb;
  wire [7:0] p6_res7__313_comb;
  wire [7:0] p6_array_index_1082429_comb;
  wire [7:0] p6_res7__314_comb;
  wire [7:0] p6_array_index_1082439_comb;
  wire [7:0] p6_res7__315_comb;
  wire [7:0] p6_res7__316_comb;
  wire [7:0] p6_res7__317_comb;
  wire [7:0] p6_res7__318_comb;
  wire [7:0] p6_res7__319_comb;
  wire [127:0] p6_res__19_comb;
  wire [127:0] p6_xor_1082479_comb;
  wire [127:0] p6_addedKey__61_comb;
  wire [7:0] p6_array_index_1082495_comb;
  wire [7:0] p6_array_index_1082496_comb;
  wire [7:0] p6_array_index_1082497_comb;
  wire [7:0] p6_array_index_1082498_comb;
  wire [7:0] p6_array_index_1082499_comb;
  wire [7:0] p6_array_index_1082500_comb;
  wire [7:0] p6_array_index_1082502_comb;
  wire [7:0] p6_array_index_1082504_comb;
  wire [7:0] p6_array_index_1082505_comb;
  wire [7:0] p6_array_index_1082506_comb;
  wire [7:0] p6_array_index_1082507_comb;
  wire [7:0] p6_array_index_1082508_comb;
  wire [7:0] p6_array_index_1082509_comb;
  wire [7:0] p6_array_index_1082511_comb;
  wire [7:0] p6_array_index_1082512_comb;
  wire [7:0] p6_array_index_1082513_comb;
  wire [7:0] p6_array_index_1082514_comb;
  wire [7:0] p6_array_index_1082515_comb;
  wire [7:0] p6_array_index_1082516_comb;
  wire [7:0] p6_array_index_1082517_comb;
  wire [7:0] p6_array_index_1082519_comb;
  wire [7:0] p6_res7__320_comb;
  wire [7:0] p6_array_index_1082528_comb;
  wire [7:0] p6_array_index_1082529_comb;
  wire [7:0] p6_array_index_1082530_comb;
  wire [7:0] p6_array_index_1082531_comb;
  wire [7:0] p6_array_index_1082532_comb;
  wire [7:0] p6_array_index_1082533_comb;
  wire [7:0] p6_res7__321_comb;
  wire [7:0] p6_array_index_1082543_comb;
  wire [7:0] p6_array_index_1082544_comb;
  wire [7:0] p6_array_index_1082545_comb;
  wire [7:0] p6_array_index_1082546_comb;
  wire [7:0] p6_array_index_1082547_comb;
  wire [7:0] p6_res7__322_comb;
  wire [7:0] p6_array_index_1082557_comb;
  wire [7:0] p6_array_index_1082558_comb;
  wire [7:0] p6_array_index_1082559_comb;
  wire [7:0] p6_array_index_1082560_comb;
  wire [7:0] p6_array_index_1082561_comb;
  wire [7:0] p6_res7__323_comb;
  wire [7:0] p6_array_index_1082572_comb;
  wire [7:0] p6_array_index_1082573_comb;
  wire [7:0] p6_array_index_1082574_comb;
  wire [7:0] p6_array_index_1082575_comb;
  wire [7:0] p6_res7__324_comb;
  wire [7:0] p6_array_index_1082585_comb;
  wire [7:0] p6_array_index_1082586_comb;
  wire [7:0] p6_array_index_1082587_comb;
  wire [7:0] p6_array_index_1082588_comb;
  wire [7:0] p6_res7__325_comb;
  wire [7:0] p6_array_index_1082599_comb;
  wire [7:0] p6_array_index_1082600_comb;
  wire [7:0] p6_array_index_1082601_comb;
  wire [7:0] p6_res7__326_comb;
  wire [7:0] p6_array_index_1082611_comb;
  wire [7:0] p6_array_index_1082612_comb;
  wire [7:0] p6_array_index_1082613_comb;
  wire [7:0] p6_res7__327_comb;
  wire [7:0] p6_array_index_1082624_comb;
  wire [7:0] p6_array_index_1082625_comb;
  wire [7:0] p6_res7__328_comb;
  wire [7:0] p6_array_index_1082635_comb;
  wire [7:0] p6_array_index_1082636_comb;
  wire [7:0] p6_res7__329_comb;
  wire [7:0] p6_array_index_1082647_comb;
  wire [7:0] p6_res7__330_comb;
  wire [7:0] p6_array_index_1082657_comb;
  wire [7:0] p6_res7__331_comb;
  wire [7:0] p6_res7__332_comb;
  wire [7:0] p6_res7__333_comb;
  wire [7:0] p6_res7__334_comb;
  wire [7:0] p6_res7__335_comb;
  wire [127:0] p6_res__20_comb;
  wire [127:0] p6_xor_1082697_comb;
  wire [127:0] p6_addedKey__62_comb;
  wire [7:0] p6_array_index_1082713_comb;
  wire [7:0] p6_array_index_1082714_comb;
  wire [7:0] p6_array_index_1082715_comb;
  wire [7:0] p6_array_index_1082716_comb;
  wire [7:0] p6_array_index_1082717_comb;
  wire [7:0] p6_array_index_1082718_comb;
  wire [7:0] p6_array_index_1082720_comb;
  wire [7:0] p6_array_index_1082722_comb;
  wire [7:0] p6_array_index_1082723_comb;
  wire [7:0] p6_array_index_1082724_comb;
  wire [7:0] p6_array_index_1082725_comb;
  wire [7:0] p6_array_index_1082726_comb;
  wire [7:0] p6_array_index_1082727_comb;
  wire [7:0] p6_array_index_1082729_comb;
  wire [7:0] p6_array_index_1082730_comb;
  wire [7:0] p6_array_index_1082731_comb;
  wire [7:0] p6_array_index_1082732_comb;
  wire [7:0] p6_array_index_1082733_comb;
  wire [7:0] p6_array_index_1082734_comb;
  wire [7:0] p6_array_index_1082735_comb;
  wire [7:0] p6_array_index_1082737_comb;
  wire [7:0] p6_res7__336_comb;
  wire [7:0] p6_array_index_1082746_comb;
  wire [7:0] p6_array_index_1082747_comb;
  wire [7:0] p6_array_index_1082748_comb;
  wire [7:0] p6_array_index_1082749_comb;
  wire [7:0] p6_array_index_1082750_comb;
  wire [7:0] p6_array_index_1082751_comb;
  wire [7:0] p6_res7__337_comb;
  wire [7:0] p6_array_index_1082761_comb;
  wire [7:0] p6_array_index_1082762_comb;
  wire [7:0] p6_array_index_1082763_comb;
  wire [7:0] p6_array_index_1082764_comb;
  wire [7:0] p6_array_index_1082765_comb;
  wire [7:0] p6_res7__338_comb;
  wire [7:0] p6_array_index_1082775_comb;
  wire [7:0] p6_array_index_1082776_comb;
  wire [7:0] p6_array_index_1082777_comb;
  wire [7:0] p6_array_index_1082778_comb;
  wire [7:0] p6_array_index_1082779_comb;
  wire [7:0] p6_res7__339_comb;
  wire [7:0] p6_array_index_1082790_comb;
  wire [7:0] p6_array_index_1082791_comb;
  wire [7:0] p6_array_index_1082792_comb;
  wire [7:0] p6_array_index_1082793_comb;
  wire [7:0] p6_res7__340_comb;
  wire [7:0] p6_array_index_1082803_comb;
  wire [7:0] p6_array_index_1082804_comb;
  wire [7:0] p6_array_index_1082805_comb;
  wire [7:0] p6_array_index_1082806_comb;
  wire [7:0] p6_res7__341_comb;
  wire [7:0] p6_array_index_1082817_comb;
  wire [7:0] p6_array_index_1082818_comb;
  wire [7:0] p6_array_index_1082819_comb;
  wire [7:0] p6_res7__342_comb;
  wire [7:0] p6_array_index_1082829_comb;
  wire [7:0] p6_array_index_1082830_comb;
  wire [7:0] p6_array_index_1082831_comb;
  wire [7:0] p6_res7__343_comb;
  wire [7:0] p6_array_index_1082842_comb;
  wire [7:0] p6_array_index_1082843_comb;
  wire [7:0] p6_res7__344_comb;
  wire [7:0] p6_array_index_1082853_comb;
  wire [7:0] p6_array_index_1082854_comb;
  wire [7:0] p6_res7__345_comb;
  wire [7:0] p6_array_index_1082865_comb;
  wire [7:0] p6_res7__346_comb;
  wire [7:0] p6_array_index_1082875_comb;
  wire [7:0] p6_res7__347_comb;
  wire [7:0] p6_res7__348_comb;
  wire [7:0] p6_res7__349_comb;
  wire [7:0] p6_res7__350_comb;
  wire [7:0] p6_res7__351_comb;
  wire [127:0] p6_res__21_comb;
  wire [127:0] p6_xor_1082915_comb;
  assign p6_array_index_1082149_comb = p5_literal_1076349[p5_res7__290];
  assign p6_array_index_1082150_comb = p5_literal_1076351[p5_res7__289];
  assign p6_array_index_1082151_comb = p5_literal_1076353[p5_res7__288];
  assign p6_array_index_1082152_comb = p5_literal_1076355[p5_array_index_1081523];
  assign p6_res7__293_comb = p5_literal_1076345[p5_res7__292] ^ p5_literal_1076347[p5_res7__291] ^ p6_array_index_1082149_comb ^ p6_array_index_1082150_comb ^ p6_array_index_1082151_comb ^ p6_array_index_1082152_comb ^ p5_array_index_1081524 ^ p5_literal_1076358[p5_array_index_1081525] ^ p5_array_index_1081526 ^ p5_array_index_1081561 ^ p5_literal_1076353[p5_array_index_1081528] ^ p5_literal_1076351[p5_array_index_1081545] ^ p5_literal_1076349[p5_array_index_1081530] ^ p5_literal_1076347[p5_array_index_1081547] ^ p5_literal_1076345[p5_array_index_1081532] ^ p5_array_index_1081533;
  assign p6_array_index_1082163_comb = p5_literal_1076351[p5_res7__290];
  assign p6_array_index_1082164_comb = p5_literal_1076353[p5_res7__289];
  assign p6_array_index_1082165_comb = p5_literal_1076355[p5_res7__288];
  assign p6_res7__294_comb = p5_literal_1076345[p6_res7__293_comb] ^ p5_literal_1076347[p5_res7__292] ^ p5_literal_1076349[p5_res7__291] ^ p6_array_index_1082163_comb ^ p6_array_index_1082164_comb ^ p6_array_index_1082165_comb ^ p5_array_index_1081523 ^ p5_literal_1076358[p5_array_index_1081524] ^ p5_array_index_1081525 ^ p5_array_index_1081575 ^ p5_array_index_1081543 ^ p5_literal_1076351[p5_array_index_1081528] ^ p5_literal_1076349[p5_array_index_1081545] ^ p5_literal_1076347[p5_array_index_1081530] ^ p5_literal_1076345[p5_array_index_1081547] ^ p5_array_index_1081532;
  assign p6_array_index_1082175_comb = p5_literal_1076351[p5_res7__291];
  assign p6_array_index_1082176_comb = p5_literal_1076353[p5_res7__290];
  assign p6_array_index_1082177_comb = p5_literal_1076355[p5_res7__289];
  assign p6_res7__295_comb = p5_literal_1076345[p6_res7__294_comb] ^ p5_literal_1076347[p6_res7__293_comb] ^ p5_literal_1076349[p5_res7__292] ^ p6_array_index_1082175_comb ^ p6_array_index_1082176_comb ^ p6_array_index_1082177_comb ^ p5_res7__288 ^ p5_literal_1076358[p5_array_index_1081523] ^ p5_array_index_1081524 ^ p5_array_index_1081589 ^ p5_array_index_1081560 ^ p5_literal_1076351[p5_array_index_1081527] ^ p5_literal_1076349[p5_array_index_1081528] ^ p5_literal_1076347[p5_array_index_1081545] ^ p5_literal_1076345[p5_array_index_1081530] ^ p5_array_index_1081547;
  assign p6_array_index_1082188_comb = p5_literal_1076353[p5_res7__291];
  assign p6_array_index_1082189_comb = p5_literal_1076355[p5_res7__290];
  assign p6_res7__296_comb = p5_literal_1076345[p6_res7__295_comb] ^ p5_literal_1076347[p6_res7__294_comb] ^ p5_literal_1076349[p6_res7__293_comb] ^ p5_literal_1076351[p5_res7__292] ^ p6_array_index_1082188_comb ^ p6_array_index_1082189_comb ^ p5_res7__289 ^ p5_literal_1076358[p5_res7__288] ^ p5_array_index_1081523 ^ p5_array_index_1081603 ^ p5_array_index_1081574 ^ p5_array_index_1081542 ^ p5_literal_1076349[p5_array_index_1081527] ^ p5_literal_1076347[p5_array_index_1081528] ^ p5_literal_1076345[p5_array_index_1081545] ^ p5_array_index_1081530;
  assign p6_array_index_1082199_comb = p5_literal_1076353[p5_res7__292];
  assign p6_array_index_1082200_comb = p5_literal_1076355[p5_res7__291];
  assign p6_res7__297_comb = p5_literal_1076345[p6_res7__296_comb] ^ p5_literal_1076347[p6_res7__295_comb] ^ p5_literal_1076349[p6_res7__294_comb] ^ p5_literal_1076351[p6_res7__293_comb] ^ p6_array_index_1082199_comb ^ p6_array_index_1082200_comb ^ p5_res7__290 ^ p5_literal_1076358[p5_res7__289] ^ p5_res7__288 ^ p6_array_index_1082152_comb ^ p5_array_index_1081588 ^ p5_array_index_1081559 ^ p5_literal_1076349[p5_array_index_1081526] ^ p5_literal_1076347[p5_array_index_1081527] ^ p5_literal_1076345[p5_array_index_1081528] ^ p5_array_index_1081545;
  assign p6_array_index_1082211_comb = p5_literal_1076355[p5_res7__292];
  assign p6_res7__298_comb = p5_literal_1076345[p6_res7__297_comb] ^ p5_literal_1076347[p6_res7__296_comb] ^ p5_literal_1076349[p6_res7__295_comb] ^ p5_literal_1076351[p6_res7__294_comb] ^ p5_literal_1076353[p6_res7__293_comb] ^ p6_array_index_1082211_comb ^ p5_res7__291 ^ p5_literal_1076358[p5_res7__290] ^ p5_res7__289 ^ p6_array_index_1082165_comb ^ p5_array_index_1081602 ^ p5_array_index_1081573 ^ p5_array_index_1081541 ^ p5_literal_1076347[p5_array_index_1081526] ^ p5_literal_1076345[p5_array_index_1081527] ^ p5_array_index_1081528;
  assign p6_array_index_1082221_comb = p5_literal_1076355[p6_res7__293_comb];
  assign p6_res7__299_comb = p5_literal_1076345[p6_res7__298_comb] ^ p5_literal_1076347[p6_res7__297_comb] ^ p5_literal_1076349[p6_res7__296_comb] ^ p5_literal_1076351[p6_res7__295_comb] ^ p5_literal_1076353[p6_res7__294_comb] ^ p6_array_index_1082221_comb ^ p5_res7__292 ^ p5_literal_1076358[p5_res7__291] ^ p5_res7__290 ^ p6_array_index_1082177_comb ^ p6_array_index_1082151_comb ^ p5_array_index_1081587 ^ p5_array_index_1081558 ^ p5_literal_1076347[p5_array_index_1081525] ^ p5_literal_1076345[p5_array_index_1081526] ^ p5_array_index_1081527;
  assign p6_res7__300_comb = p5_literal_1076345[p6_res7__299_comb] ^ p5_literal_1076347[p6_res7__298_comb] ^ p5_literal_1076349[p6_res7__297_comb] ^ p5_literal_1076351[p6_res7__296_comb] ^ p5_literal_1076353[p6_res7__295_comb] ^ p5_literal_1076355[p6_res7__294_comb] ^ p6_res7__293_comb ^ p5_literal_1076358[p5_res7__292] ^ p5_res7__291 ^ p6_array_index_1082189_comb ^ p6_array_index_1082164_comb ^ p5_array_index_1081601 ^ p5_array_index_1081572 ^ p5_array_index_1081540 ^ p5_literal_1076345[p5_array_index_1081525] ^ p5_array_index_1081526;
  assign p6_res7__301_comb = p5_literal_1076345[p6_res7__300_comb] ^ p5_literal_1076347[p6_res7__299_comb] ^ p5_literal_1076349[p6_res7__298_comb] ^ p5_literal_1076351[p6_res7__297_comb] ^ p5_literal_1076353[p6_res7__296_comb] ^ p5_literal_1076355[p6_res7__295_comb] ^ p6_res7__294_comb ^ p5_literal_1076358[p6_res7__293_comb] ^ p5_res7__292 ^ p6_array_index_1082200_comb ^ p6_array_index_1082176_comb ^ p6_array_index_1082150_comb ^ p5_array_index_1081586 ^ p5_array_index_1081557 ^ p5_literal_1076345[p5_array_index_1081524] ^ p5_array_index_1081525;
  assign p6_res7__302_comb = p5_literal_1076345[p6_res7__301_comb] ^ p5_literal_1076347[p6_res7__300_comb] ^ p5_literal_1076349[p6_res7__299_comb] ^ p5_literal_1076351[p6_res7__298_comb] ^ p5_literal_1076353[p6_res7__297_comb] ^ p5_literal_1076355[p6_res7__296_comb] ^ p6_res7__295_comb ^ p5_literal_1076358[p6_res7__294_comb] ^ p6_res7__293_comb ^ p6_array_index_1082211_comb ^ p6_array_index_1082188_comb ^ p6_array_index_1082163_comb ^ p5_array_index_1081600 ^ p5_array_index_1081571 ^ p5_array_index_1081539 ^ p5_array_index_1081524;
  assign p6_res7__303_comb = p5_literal_1076345[p6_res7__302_comb] ^ p5_literal_1076347[p6_res7__301_comb] ^ p5_literal_1076349[p6_res7__300_comb] ^ p5_literal_1076351[p6_res7__299_comb] ^ p5_literal_1076353[p6_res7__298_comb] ^ p5_literal_1076355[p6_res7__297_comb] ^ p6_res7__296_comb ^ p5_literal_1076358[p6_res7__295_comb] ^ p6_res7__294_comb ^ p6_array_index_1082221_comb ^ p6_array_index_1082199_comb ^ p6_array_index_1082175_comb ^ p6_array_index_1082149_comb ^ p5_array_index_1081585 ^ p5_array_index_1081556 ^ p5_array_index_1081523;
  assign p6_res__18_comb = {p6_res7__303_comb, p6_res7__302_comb, p6_res7__301_comb, p6_res7__300_comb, p6_res7__299_comb, p6_res7__298_comb, p6_res7__297_comb, p6_res7__296_comb, p6_res7__295_comb, p6_res7__294_comb, p6_res7__293_comb, p5_res7__292, p5_res7__291, p5_res7__290, p5_res7__289, p5_res7__288};
  assign p6_xor_1082261_comb = p6_res__18_comb ^ p5_xor_1081289;
  assign p6_addedKey__60_comb = p6_xor_1082261_comb ^ 128'h547f_7727_7ce9_8774_2ea9_3083_bcc2_4114;
  assign p6_array_index_1082277_comb = p5_arr[p6_addedKey__60_comb[127:120]];
  assign p6_array_index_1082278_comb = p5_arr[p6_addedKey__60_comb[119:112]];
  assign p6_array_index_1082279_comb = p5_arr[p6_addedKey__60_comb[111:104]];
  assign p6_array_index_1082280_comb = p5_arr[p6_addedKey__60_comb[103:96]];
  assign p6_array_index_1082281_comb = p5_arr[p6_addedKey__60_comb[95:88]];
  assign p6_array_index_1082282_comb = p5_arr[p6_addedKey__60_comb[87:80]];
  assign p6_array_index_1082284_comb = p5_arr[p6_addedKey__60_comb[71:64]];
  assign p6_array_index_1082286_comb = p5_arr[p6_addedKey__60_comb[55:48]];
  assign p6_array_index_1082287_comb = p5_arr[p6_addedKey__60_comb[47:40]];
  assign p6_array_index_1082288_comb = p5_arr[p6_addedKey__60_comb[39:32]];
  assign p6_array_index_1082289_comb = p5_arr[p6_addedKey__60_comb[31:24]];
  assign p6_array_index_1082290_comb = p5_arr[p6_addedKey__60_comb[23:16]];
  assign p6_array_index_1082291_comb = p5_arr[p6_addedKey__60_comb[15:8]];
  assign p6_array_index_1082293_comb = p5_literal_1076345[p6_array_index_1082277_comb];
  assign p6_array_index_1082294_comb = p5_literal_1076347[p6_array_index_1082278_comb];
  assign p6_array_index_1082295_comb = p5_literal_1076349[p6_array_index_1082279_comb];
  assign p6_array_index_1082296_comb = p5_literal_1076351[p6_array_index_1082280_comb];
  assign p6_array_index_1082297_comb = p5_literal_1076353[p6_array_index_1082281_comb];
  assign p6_array_index_1082298_comb = p5_literal_1076355[p6_array_index_1082282_comb];
  assign p6_array_index_1082299_comb = p5_arr[p6_addedKey__60_comb[79:72]];
  assign p6_array_index_1082301_comb = p5_arr[p6_addedKey__60_comb[63:56]];
  assign p6_res7__304_comb = p6_array_index_1082293_comb ^ p6_array_index_1082294_comb ^ p6_array_index_1082295_comb ^ p6_array_index_1082296_comb ^ p6_array_index_1082297_comb ^ p6_array_index_1082298_comb ^ p6_array_index_1082299_comb ^ p5_literal_1076358[p6_array_index_1082284_comb] ^ p6_array_index_1082301_comb ^ p5_literal_1076355[p6_array_index_1082286_comb] ^ p5_literal_1076353[p6_array_index_1082287_comb] ^ p5_literal_1076351[p6_array_index_1082288_comb] ^ p5_literal_1076349[p6_array_index_1082289_comb] ^ p5_literal_1076347[p6_array_index_1082290_comb] ^ p5_literal_1076345[p6_array_index_1082291_comb] ^ p5_arr[p6_addedKey__60_comb[7:0]];
  assign p6_array_index_1082310_comb = p5_literal_1076345[p6_res7__304_comb];
  assign p6_array_index_1082311_comb = p5_literal_1076347[p6_array_index_1082277_comb];
  assign p6_array_index_1082312_comb = p5_literal_1076349[p6_array_index_1082278_comb];
  assign p6_array_index_1082313_comb = p5_literal_1076351[p6_array_index_1082279_comb];
  assign p6_array_index_1082314_comb = p5_literal_1076353[p6_array_index_1082280_comb];
  assign p6_array_index_1082315_comb = p5_literal_1076355[p6_array_index_1082281_comb];
  assign p6_res7__305_comb = p6_array_index_1082310_comb ^ p6_array_index_1082311_comb ^ p6_array_index_1082312_comb ^ p6_array_index_1082313_comb ^ p6_array_index_1082314_comb ^ p6_array_index_1082315_comb ^ p6_array_index_1082282_comb ^ p5_literal_1076358[p6_array_index_1082299_comb] ^ p6_array_index_1082284_comb ^ p5_literal_1076355[p6_array_index_1082301_comb] ^ p5_literal_1076353[p6_array_index_1082286_comb] ^ p5_literal_1076351[p6_array_index_1082287_comb] ^ p5_literal_1076349[p6_array_index_1082288_comb] ^ p5_literal_1076347[p6_array_index_1082289_comb] ^ p5_literal_1076345[p6_array_index_1082290_comb] ^ p6_array_index_1082291_comb;
  assign p6_array_index_1082325_comb = p5_literal_1076347[p6_res7__304_comb];
  assign p6_array_index_1082326_comb = p5_literal_1076349[p6_array_index_1082277_comb];
  assign p6_array_index_1082327_comb = p5_literal_1076351[p6_array_index_1082278_comb];
  assign p6_array_index_1082328_comb = p5_literal_1076353[p6_array_index_1082279_comb];
  assign p6_array_index_1082329_comb = p5_literal_1076355[p6_array_index_1082280_comb];
  assign p6_res7__306_comb = p5_literal_1076345[p6_res7__305_comb] ^ p6_array_index_1082325_comb ^ p6_array_index_1082326_comb ^ p6_array_index_1082327_comb ^ p6_array_index_1082328_comb ^ p6_array_index_1082329_comb ^ p6_array_index_1082281_comb ^ p5_literal_1076358[p6_array_index_1082282_comb] ^ p6_array_index_1082299_comb ^ p5_literal_1076355[p6_array_index_1082284_comb] ^ p5_literal_1076353[p6_array_index_1082301_comb] ^ p5_literal_1076351[p6_array_index_1082286_comb] ^ p5_literal_1076349[p6_array_index_1082287_comb] ^ p5_literal_1076347[p6_array_index_1082288_comb] ^ p5_literal_1076345[p6_array_index_1082289_comb] ^ p6_array_index_1082290_comb;
  assign p6_array_index_1082339_comb = p5_literal_1076347[p6_res7__305_comb];
  assign p6_array_index_1082340_comb = p5_literal_1076349[p6_res7__304_comb];
  assign p6_array_index_1082341_comb = p5_literal_1076351[p6_array_index_1082277_comb];
  assign p6_array_index_1082342_comb = p5_literal_1076353[p6_array_index_1082278_comb];
  assign p6_array_index_1082343_comb = p5_literal_1076355[p6_array_index_1082279_comb];
  assign p6_res7__307_comb = p5_literal_1076345[p6_res7__306_comb] ^ p6_array_index_1082339_comb ^ p6_array_index_1082340_comb ^ p6_array_index_1082341_comb ^ p6_array_index_1082342_comb ^ p6_array_index_1082343_comb ^ p6_array_index_1082280_comb ^ p5_literal_1076358[p6_array_index_1082281_comb] ^ p6_array_index_1082282_comb ^ p5_literal_1076355[p6_array_index_1082299_comb] ^ p5_literal_1076353[p6_array_index_1082284_comb] ^ p5_literal_1076351[p6_array_index_1082301_comb] ^ p5_literal_1076349[p6_array_index_1082286_comb] ^ p5_literal_1076347[p6_array_index_1082287_comb] ^ p5_literal_1076345[p6_array_index_1082288_comb] ^ p6_array_index_1082289_comb;
  assign p6_array_index_1082354_comb = p5_literal_1076349[p6_res7__305_comb];
  assign p6_array_index_1082355_comb = p5_literal_1076351[p6_res7__304_comb];
  assign p6_array_index_1082356_comb = p5_literal_1076353[p6_array_index_1082277_comb];
  assign p6_array_index_1082357_comb = p5_literal_1076355[p6_array_index_1082278_comb];
  assign p6_res7__308_comb = p5_literal_1076345[p6_res7__307_comb] ^ p5_literal_1076347[p6_res7__306_comb] ^ p6_array_index_1082354_comb ^ p6_array_index_1082355_comb ^ p6_array_index_1082356_comb ^ p6_array_index_1082357_comb ^ p6_array_index_1082279_comb ^ p5_literal_1076358[p6_array_index_1082280_comb] ^ p6_array_index_1082281_comb ^ p6_array_index_1082298_comb ^ p5_literal_1076353[p6_array_index_1082299_comb] ^ p5_literal_1076351[p6_array_index_1082284_comb] ^ p5_literal_1076349[p6_array_index_1082301_comb] ^ p5_literal_1076347[p6_array_index_1082286_comb] ^ p5_literal_1076345[p6_array_index_1082287_comb] ^ p6_array_index_1082288_comb;
  assign p6_array_index_1082367_comb = p5_literal_1076349[p6_res7__306_comb];
  assign p6_array_index_1082368_comb = p5_literal_1076351[p6_res7__305_comb];
  assign p6_array_index_1082369_comb = p5_literal_1076353[p6_res7__304_comb];
  assign p6_array_index_1082370_comb = p5_literal_1076355[p6_array_index_1082277_comb];
  assign p6_res7__309_comb = p5_literal_1076345[p6_res7__308_comb] ^ p5_literal_1076347[p6_res7__307_comb] ^ p6_array_index_1082367_comb ^ p6_array_index_1082368_comb ^ p6_array_index_1082369_comb ^ p6_array_index_1082370_comb ^ p6_array_index_1082278_comb ^ p5_literal_1076358[p6_array_index_1082279_comb] ^ p6_array_index_1082280_comb ^ p6_array_index_1082315_comb ^ p5_literal_1076353[p6_array_index_1082282_comb] ^ p5_literal_1076351[p6_array_index_1082299_comb] ^ p5_literal_1076349[p6_array_index_1082284_comb] ^ p5_literal_1076347[p6_array_index_1082301_comb] ^ p5_literal_1076345[p6_array_index_1082286_comb] ^ p6_array_index_1082287_comb;
  assign p6_array_index_1082381_comb = p5_literal_1076351[p6_res7__306_comb];
  assign p6_array_index_1082382_comb = p5_literal_1076353[p6_res7__305_comb];
  assign p6_array_index_1082383_comb = p5_literal_1076355[p6_res7__304_comb];
  assign p6_res7__310_comb = p5_literal_1076345[p6_res7__309_comb] ^ p5_literal_1076347[p6_res7__308_comb] ^ p5_literal_1076349[p6_res7__307_comb] ^ p6_array_index_1082381_comb ^ p6_array_index_1082382_comb ^ p6_array_index_1082383_comb ^ p6_array_index_1082277_comb ^ p5_literal_1076358[p6_array_index_1082278_comb] ^ p6_array_index_1082279_comb ^ p6_array_index_1082329_comb ^ p6_array_index_1082297_comb ^ p5_literal_1076351[p6_array_index_1082282_comb] ^ p5_literal_1076349[p6_array_index_1082299_comb] ^ p5_literal_1076347[p6_array_index_1082284_comb] ^ p5_literal_1076345[p6_array_index_1082301_comb] ^ p6_array_index_1082286_comb;
  assign p6_array_index_1082393_comb = p5_literal_1076351[p6_res7__307_comb];
  assign p6_array_index_1082394_comb = p5_literal_1076353[p6_res7__306_comb];
  assign p6_array_index_1082395_comb = p5_literal_1076355[p6_res7__305_comb];
  assign p6_res7__311_comb = p5_literal_1076345[p6_res7__310_comb] ^ p5_literal_1076347[p6_res7__309_comb] ^ p5_literal_1076349[p6_res7__308_comb] ^ p6_array_index_1082393_comb ^ p6_array_index_1082394_comb ^ p6_array_index_1082395_comb ^ p6_res7__304_comb ^ p5_literal_1076358[p6_array_index_1082277_comb] ^ p6_array_index_1082278_comb ^ p6_array_index_1082343_comb ^ p6_array_index_1082314_comb ^ p5_literal_1076351[p6_array_index_1082281_comb] ^ p5_literal_1076349[p6_array_index_1082282_comb] ^ p5_literal_1076347[p6_array_index_1082299_comb] ^ p5_literal_1076345[p6_array_index_1082284_comb] ^ p6_array_index_1082301_comb;
  assign p6_array_index_1082406_comb = p5_literal_1076353[p6_res7__307_comb];
  assign p6_array_index_1082407_comb = p5_literal_1076355[p6_res7__306_comb];
  assign p6_res7__312_comb = p5_literal_1076345[p6_res7__311_comb] ^ p5_literal_1076347[p6_res7__310_comb] ^ p5_literal_1076349[p6_res7__309_comb] ^ p5_literal_1076351[p6_res7__308_comb] ^ p6_array_index_1082406_comb ^ p6_array_index_1082407_comb ^ p6_res7__305_comb ^ p5_literal_1076358[p6_res7__304_comb] ^ p6_array_index_1082277_comb ^ p6_array_index_1082357_comb ^ p6_array_index_1082328_comb ^ p6_array_index_1082296_comb ^ p5_literal_1076349[p6_array_index_1082281_comb] ^ p5_literal_1076347[p6_array_index_1082282_comb] ^ p5_literal_1076345[p6_array_index_1082299_comb] ^ p6_array_index_1082284_comb;
  assign p6_array_index_1082417_comb = p5_literal_1076353[p6_res7__308_comb];
  assign p6_array_index_1082418_comb = p5_literal_1076355[p6_res7__307_comb];
  assign p6_res7__313_comb = p5_literal_1076345[p6_res7__312_comb] ^ p5_literal_1076347[p6_res7__311_comb] ^ p5_literal_1076349[p6_res7__310_comb] ^ p5_literal_1076351[p6_res7__309_comb] ^ p6_array_index_1082417_comb ^ p6_array_index_1082418_comb ^ p6_res7__306_comb ^ p5_literal_1076358[p6_res7__305_comb] ^ p6_res7__304_comb ^ p6_array_index_1082370_comb ^ p6_array_index_1082342_comb ^ p6_array_index_1082313_comb ^ p5_literal_1076349[p6_array_index_1082280_comb] ^ p5_literal_1076347[p6_array_index_1082281_comb] ^ p5_literal_1076345[p6_array_index_1082282_comb] ^ p6_array_index_1082299_comb;
  assign p6_array_index_1082429_comb = p5_literal_1076355[p6_res7__308_comb];
  assign p6_res7__314_comb = p5_literal_1076345[p6_res7__313_comb] ^ p5_literal_1076347[p6_res7__312_comb] ^ p5_literal_1076349[p6_res7__311_comb] ^ p5_literal_1076351[p6_res7__310_comb] ^ p5_literal_1076353[p6_res7__309_comb] ^ p6_array_index_1082429_comb ^ p6_res7__307_comb ^ p5_literal_1076358[p6_res7__306_comb] ^ p6_res7__305_comb ^ p6_array_index_1082383_comb ^ p6_array_index_1082356_comb ^ p6_array_index_1082327_comb ^ p6_array_index_1082295_comb ^ p5_literal_1076347[p6_array_index_1082280_comb] ^ p5_literal_1076345[p6_array_index_1082281_comb] ^ p6_array_index_1082282_comb;
  assign p6_array_index_1082439_comb = p5_literal_1076355[p6_res7__309_comb];
  assign p6_res7__315_comb = p5_literal_1076345[p6_res7__314_comb] ^ p5_literal_1076347[p6_res7__313_comb] ^ p5_literal_1076349[p6_res7__312_comb] ^ p5_literal_1076351[p6_res7__311_comb] ^ p5_literal_1076353[p6_res7__310_comb] ^ p6_array_index_1082439_comb ^ p6_res7__308_comb ^ p5_literal_1076358[p6_res7__307_comb] ^ p6_res7__306_comb ^ p6_array_index_1082395_comb ^ p6_array_index_1082369_comb ^ p6_array_index_1082341_comb ^ p6_array_index_1082312_comb ^ p5_literal_1076347[p6_array_index_1082279_comb] ^ p5_literal_1076345[p6_array_index_1082280_comb] ^ p6_array_index_1082281_comb;
  assign p6_res7__316_comb = p5_literal_1076345[p6_res7__315_comb] ^ p5_literal_1076347[p6_res7__314_comb] ^ p5_literal_1076349[p6_res7__313_comb] ^ p5_literal_1076351[p6_res7__312_comb] ^ p5_literal_1076353[p6_res7__311_comb] ^ p5_literal_1076355[p6_res7__310_comb] ^ p6_res7__309_comb ^ p5_literal_1076358[p6_res7__308_comb] ^ p6_res7__307_comb ^ p6_array_index_1082407_comb ^ p6_array_index_1082382_comb ^ p6_array_index_1082355_comb ^ p6_array_index_1082326_comb ^ p6_array_index_1082294_comb ^ p5_literal_1076345[p6_array_index_1082279_comb] ^ p6_array_index_1082280_comb;
  assign p6_res7__317_comb = p5_literal_1076345[p6_res7__316_comb] ^ p5_literal_1076347[p6_res7__315_comb] ^ p5_literal_1076349[p6_res7__314_comb] ^ p5_literal_1076351[p6_res7__313_comb] ^ p5_literal_1076353[p6_res7__312_comb] ^ p5_literal_1076355[p6_res7__311_comb] ^ p6_res7__310_comb ^ p5_literal_1076358[p6_res7__309_comb] ^ p6_res7__308_comb ^ p6_array_index_1082418_comb ^ p6_array_index_1082394_comb ^ p6_array_index_1082368_comb ^ p6_array_index_1082340_comb ^ p6_array_index_1082311_comb ^ p5_literal_1076345[p6_array_index_1082278_comb] ^ p6_array_index_1082279_comb;
  assign p6_res7__318_comb = p5_literal_1076345[p6_res7__317_comb] ^ p5_literal_1076347[p6_res7__316_comb] ^ p5_literal_1076349[p6_res7__315_comb] ^ p5_literal_1076351[p6_res7__314_comb] ^ p5_literal_1076353[p6_res7__313_comb] ^ p5_literal_1076355[p6_res7__312_comb] ^ p6_res7__311_comb ^ p5_literal_1076358[p6_res7__310_comb] ^ p6_res7__309_comb ^ p6_array_index_1082429_comb ^ p6_array_index_1082406_comb ^ p6_array_index_1082381_comb ^ p6_array_index_1082354_comb ^ p6_array_index_1082325_comb ^ p6_array_index_1082293_comb ^ p6_array_index_1082278_comb;
  assign p6_res7__319_comb = p5_literal_1076345[p6_res7__318_comb] ^ p5_literal_1076347[p6_res7__317_comb] ^ p5_literal_1076349[p6_res7__316_comb] ^ p5_literal_1076351[p6_res7__315_comb] ^ p5_literal_1076353[p6_res7__314_comb] ^ p5_literal_1076355[p6_res7__313_comb] ^ p6_res7__312_comb ^ p5_literal_1076358[p6_res7__311_comb] ^ p6_res7__310_comb ^ p6_array_index_1082439_comb ^ p6_array_index_1082417_comb ^ p6_array_index_1082393_comb ^ p6_array_index_1082367_comb ^ p6_array_index_1082339_comb ^ p6_array_index_1082310_comb ^ p6_array_index_1082277_comb;
  assign p6_res__19_comb = {p6_res7__319_comb, p6_res7__318_comb, p6_res7__317_comb, p6_res7__316_comb, p6_res7__315_comb, p6_res7__314_comb, p6_res7__313_comb, p6_res7__312_comb, p6_res7__311_comb, p6_res7__310_comb, p6_res7__309_comb, p6_res7__308_comb, p6_res7__307_comb, p6_res7__306_comb, p6_res7__305_comb, p6_res7__304_comb};
  assign p6_xor_1082479_comb = p6_res__19_comb ^ p5_xor_1081507;
  assign p6_addedKey__61_comb = p6_xor_1082479_comb ^ 128'h3add_0155_10a1_fdcc_738e_8d93_6146_d515;
  assign p6_array_index_1082495_comb = p5_arr[p6_addedKey__61_comb[127:120]];
  assign p6_array_index_1082496_comb = p5_arr[p6_addedKey__61_comb[119:112]];
  assign p6_array_index_1082497_comb = p5_arr[p6_addedKey__61_comb[111:104]];
  assign p6_array_index_1082498_comb = p5_arr[p6_addedKey__61_comb[103:96]];
  assign p6_array_index_1082499_comb = p5_arr[p6_addedKey__61_comb[95:88]];
  assign p6_array_index_1082500_comb = p5_arr[p6_addedKey__61_comb[87:80]];
  assign p6_array_index_1082502_comb = p5_arr[p6_addedKey__61_comb[71:64]];
  assign p6_array_index_1082504_comb = p5_arr[p6_addedKey__61_comb[55:48]];
  assign p6_array_index_1082505_comb = p5_arr[p6_addedKey__61_comb[47:40]];
  assign p6_array_index_1082506_comb = p5_arr[p6_addedKey__61_comb[39:32]];
  assign p6_array_index_1082507_comb = p5_arr[p6_addedKey__61_comb[31:24]];
  assign p6_array_index_1082508_comb = p5_arr[p6_addedKey__61_comb[23:16]];
  assign p6_array_index_1082509_comb = p5_arr[p6_addedKey__61_comb[15:8]];
  assign p6_array_index_1082511_comb = p5_literal_1076345[p6_array_index_1082495_comb];
  assign p6_array_index_1082512_comb = p5_literal_1076347[p6_array_index_1082496_comb];
  assign p6_array_index_1082513_comb = p5_literal_1076349[p6_array_index_1082497_comb];
  assign p6_array_index_1082514_comb = p5_literal_1076351[p6_array_index_1082498_comb];
  assign p6_array_index_1082515_comb = p5_literal_1076353[p6_array_index_1082499_comb];
  assign p6_array_index_1082516_comb = p5_literal_1076355[p6_array_index_1082500_comb];
  assign p6_array_index_1082517_comb = p5_arr[p6_addedKey__61_comb[79:72]];
  assign p6_array_index_1082519_comb = p5_arr[p6_addedKey__61_comb[63:56]];
  assign p6_res7__320_comb = p6_array_index_1082511_comb ^ p6_array_index_1082512_comb ^ p6_array_index_1082513_comb ^ p6_array_index_1082514_comb ^ p6_array_index_1082515_comb ^ p6_array_index_1082516_comb ^ p6_array_index_1082517_comb ^ p5_literal_1076358[p6_array_index_1082502_comb] ^ p6_array_index_1082519_comb ^ p5_literal_1076355[p6_array_index_1082504_comb] ^ p5_literal_1076353[p6_array_index_1082505_comb] ^ p5_literal_1076351[p6_array_index_1082506_comb] ^ p5_literal_1076349[p6_array_index_1082507_comb] ^ p5_literal_1076347[p6_array_index_1082508_comb] ^ p5_literal_1076345[p6_array_index_1082509_comb] ^ p5_arr[p6_addedKey__61_comb[7:0]];
  assign p6_array_index_1082528_comb = p5_literal_1076345[p6_res7__320_comb];
  assign p6_array_index_1082529_comb = p5_literal_1076347[p6_array_index_1082495_comb];
  assign p6_array_index_1082530_comb = p5_literal_1076349[p6_array_index_1082496_comb];
  assign p6_array_index_1082531_comb = p5_literal_1076351[p6_array_index_1082497_comb];
  assign p6_array_index_1082532_comb = p5_literal_1076353[p6_array_index_1082498_comb];
  assign p6_array_index_1082533_comb = p5_literal_1076355[p6_array_index_1082499_comb];
  assign p6_res7__321_comb = p6_array_index_1082528_comb ^ p6_array_index_1082529_comb ^ p6_array_index_1082530_comb ^ p6_array_index_1082531_comb ^ p6_array_index_1082532_comb ^ p6_array_index_1082533_comb ^ p6_array_index_1082500_comb ^ p5_literal_1076358[p6_array_index_1082517_comb] ^ p6_array_index_1082502_comb ^ p5_literal_1076355[p6_array_index_1082519_comb] ^ p5_literal_1076353[p6_array_index_1082504_comb] ^ p5_literal_1076351[p6_array_index_1082505_comb] ^ p5_literal_1076349[p6_array_index_1082506_comb] ^ p5_literal_1076347[p6_array_index_1082507_comb] ^ p5_literal_1076345[p6_array_index_1082508_comb] ^ p6_array_index_1082509_comb;
  assign p6_array_index_1082543_comb = p5_literal_1076347[p6_res7__320_comb];
  assign p6_array_index_1082544_comb = p5_literal_1076349[p6_array_index_1082495_comb];
  assign p6_array_index_1082545_comb = p5_literal_1076351[p6_array_index_1082496_comb];
  assign p6_array_index_1082546_comb = p5_literal_1076353[p6_array_index_1082497_comb];
  assign p6_array_index_1082547_comb = p5_literal_1076355[p6_array_index_1082498_comb];
  assign p6_res7__322_comb = p5_literal_1076345[p6_res7__321_comb] ^ p6_array_index_1082543_comb ^ p6_array_index_1082544_comb ^ p6_array_index_1082545_comb ^ p6_array_index_1082546_comb ^ p6_array_index_1082547_comb ^ p6_array_index_1082499_comb ^ p5_literal_1076358[p6_array_index_1082500_comb] ^ p6_array_index_1082517_comb ^ p5_literal_1076355[p6_array_index_1082502_comb] ^ p5_literal_1076353[p6_array_index_1082519_comb] ^ p5_literal_1076351[p6_array_index_1082504_comb] ^ p5_literal_1076349[p6_array_index_1082505_comb] ^ p5_literal_1076347[p6_array_index_1082506_comb] ^ p5_literal_1076345[p6_array_index_1082507_comb] ^ p6_array_index_1082508_comb;
  assign p6_array_index_1082557_comb = p5_literal_1076347[p6_res7__321_comb];
  assign p6_array_index_1082558_comb = p5_literal_1076349[p6_res7__320_comb];
  assign p6_array_index_1082559_comb = p5_literal_1076351[p6_array_index_1082495_comb];
  assign p6_array_index_1082560_comb = p5_literal_1076353[p6_array_index_1082496_comb];
  assign p6_array_index_1082561_comb = p5_literal_1076355[p6_array_index_1082497_comb];
  assign p6_res7__323_comb = p5_literal_1076345[p6_res7__322_comb] ^ p6_array_index_1082557_comb ^ p6_array_index_1082558_comb ^ p6_array_index_1082559_comb ^ p6_array_index_1082560_comb ^ p6_array_index_1082561_comb ^ p6_array_index_1082498_comb ^ p5_literal_1076358[p6_array_index_1082499_comb] ^ p6_array_index_1082500_comb ^ p5_literal_1076355[p6_array_index_1082517_comb] ^ p5_literal_1076353[p6_array_index_1082502_comb] ^ p5_literal_1076351[p6_array_index_1082519_comb] ^ p5_literal_1076349[p6_array_index_1082504_comb] ^ p5_literal_1076347[p6_array_index_1082505_comb] ^ p5_literal_1076345[p6_array_index_1082506_comb] ^ p6_array_index_1082507_comb;
  assign p6_array_index_1082572_comb = p5_literal_1076349[p6_res7__321_comb];
  assign p6_array_index_1082573_comb = p5_literal_1076351[p6_res7__320_comb];
  assign p6_array_index_1082574_comb = p5_literal_1076353[p6_array_index_1082495_comb];
  assign p6_array_index_1082575_comb = p5_literal_1076355[p6_array_index_1082496_comb];
  assign p6_res7__324_comb = p5_literal_1076345[p6_res7__323_comb] ^ p5_literal_1076347[p6_res7__322_comb] ^ p6_array_index_1082572_comb ^ p6_array_index_1082573_comb ^ p6_array_index_1082574_comb ^ p6_array_index_1082575_comb ^ p6_array_index_1082497_comb ^ p5_literal_1076358[p6_array_index_1082498_comb] ^ p6_array_index_1082499_comb ^ p6_array_index_1082516_comb ^ p5_literal_1076353[p6_array_index_1082517_comb] ^ p5_literal_1076351[p6_array_index_1082502_comb] ^ p5_literal_1076349[p6_array_index_1082519_comb] ^ p5_literal_1076347[p6_array_index_1082504_comb] ^ p5_literal_1076345[p6_array_index_1082505_comb] ^ p6_array_index_1082506_comb;
  assign p6_array_index_1082585_comb = p5_literal_1076349[p6_res7__322_comb];
  assign p6_array_index_1082586_comb = p5_literal_1076351[p6_res7__321_comb];
  assign p6_array_index_1082587_comb = p5_literal_1076353[p6_res7__320_comb];
  assign p6_array_index_1082588_comb = p5_literal_1076355[p6_array_index_1082495_comb];
  assign p6_res7__325_comb = p5_literal_1076345[p6_res7__324_comb] ^ p5_literal_1076347[p6_res7__323_comb] ^ p6_array_index_1082585_comb ^ p6_array_index_1082586_comb ^ p6_array_index_1082587_comb ^ p6_array_index_1082588_comb ^ p6_array_index_1082496_comb ^ p5_literal_1076358[p6_array_index_1082497_comb] ^ p6_array_index_1082498_comb ^ p6_array_index_1082533_comb ^ p5_literal_1076353[p6_array_index_1082500_comb] ^ p5_literal_1076351[p6_array_index_1082517_comb] ^ p5_literal_1076349[p6_array_index_1082502_comb] ^ p5_literal_1076347[p6_array_index_1082519_comb] ^ p5_literal_1076345[p6_array_index_1082504_comb] ^ p6_array_index_1082505_comb;
  assign p6_array_index_1082599_comb = p5_literal_1076351[p6_res7__322_comb];
  assign p6_array_index_1082600_comb = p5_literal_1076353[p6_res7__321_comb];
  assign p6_array_index_1082601_comb = p5_literal_1076355[p6_res7__320_comb];
  assign p6_res7__326_comb = p5_literal_1076345[p6_res7__325_comb] ^ p5_literal_1076347[p6_res7__324_comb] ^ p5_literal_1076349[p6_res7__323_comb] ^ p6_array_index_1082599_comb ^ p6_array_index_1082600_comb ^ p6_array_index_1082601_comb ^ p6_array_index_1082495_comb ^ p5_literal_1076358[p6_array_index_1082496_comb] ^ p6_array_index_1082497_comb ^ p6_array_index_1082547_comb ^ p6_array_index_1082515_comb ^ p5_literal_1076351[p6_array_index_1082500_comb] ^ p5_literal_1076349[p6_array_index_1082517_comb] ^ p5_literal_1076347[p6_array_index_1082502_comb] ^ p5_literal_1076345[p6_array_index_1082519_comb] ^ p6_array_index_1082504_comb;
  assign p6_array_index_1082611_comb = p5_literal_1076351[p6_res7__323_comb];
  assign p6_array_index_1082612_comb = p5_literal_1076353[p6_res7__322_comb];
  assign p6_array_index_1082613_comb = p5_literal_1076355[p6_res7__321_comb];
  assign p6_res7__327_comb = p5_literal_1076345[p6_res7__326_comb] ^ p5_literal_1076347[p6_res7__325_comb] ^ p5_literal_1076349[p6_res7__324_comb] ^ p6_array_index_1082611_comb ^ p6_array_index_1082612_comb ^ p6_array_index_1082613_comb ^ p6_res7__320_comb ^ p5_literal_1076358[p6_array_index_1082495_comb] ^ p6_array_index_1082496_comb ^ p6_array_index_1082561_comb ^ p6_array_index_1082532_comb ^ p5_literal_1076351[p6_array_index_1082499_comb] ^ p5_literal_1076349[p6_array_index_1082500_comb] ^ p5_literal_1076347[p6_array_index_1082517_comb] ^ p5_literal_1076345[p6_array_index_1082502_comb] ^ p6_array_index_1082519_comb;
  assign p6_array_index_1082624_comb = p5_literal_1076353[p6_res7__323_comb];
  assign p6_array_index_1082625_comb = p5_literal_1076355[p6_res7__322_comb];
  assign p6_res7__328_comb = p5_literal_1076345[p6_res7__327_comb] ^ p5_literal_1076347[p6_res7__326_comb] ^ p5_literal_1076349[p6_res7__325_comb] ^ p5_literal_1076351[p6_res7__324_comb] ^ p6_array_index_1082624_comb ^ p6_array_index_1082625_comb ^ p6_res7__321_comb ^ p5_literal_1076358[p6_res7__320_comb] ^ p6_array_index_1082495_comb ^ p6_array_index_1082575_comb ^ p6_array_index_1082546_comb ^ p6_array_index_1082514_comb ^ p5_literal_1076349[p6_array_index_1082499_comb] ^ p5_literal_1076347[p6_array_index_1082500_comb] ^ p5_literal_1076345[p6_array_index_1082517_comb] ^ p6_array_index_1082502_comb;
  assign p6_array_index_1082635_comb = p5_literal_1076353[p6_res7__324_comb];
  assign p6_array_index_1082636_comb = p5_literal_1076355[p6_res7__323_comb];
  assign p6_res7__329_comb = p5_literal_1076345[p6_res7__328_comb] ^ p5_literal_1076347[p6_res7__327_comb] ^ p5_literal_1076349[p6_res7__326_comb] ^ p5_literal_1076351[p6_res7__325_comb] ^ p6_array_index_1082635_comb ^ p6_array_index_1082636_comb ^ p6_res7__322_comb ^ p5_literal_1076358[p6_res7__321_comb] ^ p6_res7__320_comb ^ p6_array_index_1082588_comb ^ p6_array_index_1082560_comb ^ p6_array_index_1082531_comb ^ p5_literal_1076349[p6_array_index_1082498_comb] ^ p5_literal_1076347[p6_array_index_1082499_comb] ^ p5_literal_1076345[p6_array_index_1082500_comb] ^ p6_array_index_1082517_comb;
  assign p6_array_index_1082647_comb = p5_literal_1076355[p6_res7__324_comb];
  assign p6_res7__330_comb = p5_literal_1076345[p6_res7__329_comb] ^ p5_literal_1076347[p6_res7__328_comb] ^ p5_literal_1076349[p6_res7__327_comb] ^ p5_literal_1076351[p6_res7__326_comb] ^ p5_literal_1076353[p6_res7__325_comb] ^ p6_array_index_1082647_comb ^ p6_res7__323_comb ^ p5_literal_1076358[p6_res7__322_comb] ^ p6_res7__321_comb ^ p6_array_index_1082601_comb ^ p6_array_index_1082574_comb ^ p6_array_index_1082545_comb ^ p6_array_index_1082513_comb ^ p5_literal_1076347[p6_array_index_1082498_comb] ^ p5_literal_1076345[p6_array_index_1082499_comb] ^ p6_array_index_1082500_comb;
  assign p6_array_index_1082657_comb = p5_literal_1076355[p6_res7__325_comb];
  assign p6_res7__331_comb = p5_literal_1076345[p6_res7__330_comb] ^ p5_literal_1076347[p6_res7__329_comb] ^ p5_literal_1076349[p6_res7__328_comb] ^ p5_literal_1076351[p6_res7__327_comb] ^ p5_literal_1076353[p6_res7__326_comb] ^ p6_array_index_1082657_comb ^ p6_res7__324_comb ^ p5_literal_1076358[p6_res7__323_comb] ^ p6_res7__322_comb ^ p6_array_index_1082613_comb ^ p6_array_index_1082587_comb ^ p6_array_index_1082559_comb ^ p6_array_index_1082530_comb ^ p5_literal_1076347[p6_array_index_1082497_comb] ^ p5_literal_1076345[p6_array_index_1082498_comb] ^ p6_array_index_1082499_comb;
  assign p6_res7__332_comb = p5_literal_1076345[p6_res7__331_comb] ^ p5_literal_1076347[p6_res7__330_comb] ^ p5_literal_1076349[p6_res7__329_comb] ^ p5_literal_1076351[p6_res7__328_comb] ^ p5_literal_1076353[p6_res7__327_comb] ^ p5_literal_1076355[p6_res7__326_comb] ^ p6_res7__325_comb ^ p5_literal_1076358[p6_res7__324_comb] ^ p6_res7__323_comb ^ p6_array_index_1082625_comb ^ p6_array_index_1082600_comb ^ p6_array_index_1082573_comb ^ p6_array_index_1082544_comb ^ p6_array_index_1082512_comb ^ p5_literal_1076345[p6_array_index_1082497_comb] ^ p6_array_index_1082498_comb;
  assign p6_res7__333_comb = p5_literal_1076345[p6_res7__332_comb] ^ p5_literal_1076347[p6_res7__331_comb] ^ p5_literal_1076349[p6_res7__330_comb] ^ p5_literal_1076351[p6_res7__329_comb] ^ p5_literal_1076353[p6_res7__328_comb] ^ p5_literal_1076355[p6_res7__327_comb] ^ p6_res7__326_comb ^ p5_literal_1076358[p6_res7__325_comb] ^ p6_res7__324_comb ^ p6_array_index_1082636_comb ^ p6_array_index_1082612_comb ^ p6_array_index_1082586_comb ^ p6_array_index_1082558_comb ^ p6_array_index_1082529_comb ^ p5_literal_1076345[p6_array_index_1082496_comb] ^ p6_array_index_1082497_comb;
  assign p6_res7__334_comb = p5_literal_1076345[p6_res7__333_comb] ^ p5_literal_1076347[p6_res7__332_comb] ^ p5_literal_1076349[p6_res7__331_comb] ^ p5_literal_1076351[p6_res7__330_comb] ^ p5_literal_1076353[p6_res7__329_comb] ^ p5_literal_1076355[p6_res7__328_comb] ^ p6_res7__327_comb ^ p5_literal_1076358[p6_res7__326_comb] ^ p6_res7__325_comb ^ p6_array_index_1082647_comb ^ p6_array_index_1082624_comb ^ p6_array_index_1082599_comb ^ p6_array_index_1082572_comb ^ p6_array_index_1082543_comb ^ p6_array_index_1082511_comb ^ p6_array_index_1082496_comb;
  assign p6_res7__335_comb = p5_literal_1076345[p6_res7__334_comb] ^ p5_literal_1076347[p6_res7__333_comb] ^ p5_literal_1076349[p6_res7__332_comb] ^ p5_literal_1076351[p6_res7__331_comb] ^ p5_literal_1076353[p6_res7__330_comb] ^ p5_literal_1076355[p6_res7__329_comb] ^ p6_res7__328_comb ^ p5_literal_1076358[p6_res7__327_comb] ^ p6_res7__326_comb ^ p6_array_index_1082657_comb ^ p6_array_index_1082635_comb ^ p6_array_index_1082611_comb ^ p6_array_index_1082585_comb ^ p6_array_index_1082557_comb ^ p6_array_index_1082528_comb ^ p6_array_index_1082495_comb;
  assign p6_res__20_comb = {p6_res7__335_comb, p6_res7__334_comb, p6_res7__333_comb, p6_res7__332_comb, p6_res7__331_comb, p6_res7__330_comb, p6_res7__329_comb, p6_res7__328_comb, p6_res7__327_comb, p6_res7__326_comb, p6_res7__325_comb, p6_res7__324_comb, p6_res7__323_comb, p6_res7__322_comb, p6_res7__321_comb, p6_res7__320_comb};
  assign p6_xor_1082697_comb = p6_res__20_comb ^ p6_xor_1082261_comb;
  assign p6_addedKey__62_comb = p6_xor_1082697_comb ^ 128'h88f8_9bc3_a479_73c7_94e7_89a3_c509_aa16;
  assign p6_array_index_1082713_comb = p5_arr[p6_addedKey__62_comb[127:120]];
  assign p6_array_index_1082714_comb = p5_arr[p6_addedKey__62_comb[119:112]];
  assign p6_array_index_1082715_comb = p5_arr[p6_addedKey__62_comb[111:104]];
  assign p6_array_index_1082716_comb = p5_arr[p6_addedKey__62_comb[103:96]];
  assign p6_array_index_1082717_comb = p5_arr[p6_addedKey__62_comb[95:88]];
  assign p6_array_index_1082718_comb = p5_arr[p6_addedKey__62_comb[87:80]];
  assign p6_array_index_1082720_comb = p5_arr[p6_addedKey__62_comb[71:64]];
  assign p6_array_index_1082722_comb = p5_arr[p6_addedKey__62_comb[55:48]];
  assign p6_array_index_1082723_comb = p5_arr[p6_addedKey__62_comb[47:40]];
  assign p6_array_index_1082724_comb = p5_arr[p6_addedKey__62_comb[39:32]];
  assign p6_array_index_1082725_comb = p5_arr[p6_addedKey__62_comb[31:24]];
  assign p6_array_index_1082726_comb = p5_arr[p6_addedKey__62_comb[23:16]];
  assign p6_array_index_1082727_comb = p5_arr[p6_addedKey__62_comb[15:8]];
  assign p6_array_index_1082729_comb = p5_literal_1076345[p6_array_index_1082713_comb];
  assign p6_array_index_1082730_comb = p5_literal_1076347[p6_array_index_1082714_comb];
  assign p6_array_index_1082731_comb = p5_literal_1076349[p6_array_index_1082715_comb];
  assign p6_array_index_1082732_comb = p5_literal_1076351[p6_array_index_1082716_comb];
  assign p6_array_index_1082733_comb = p5_literal_1076353[p6_array_index_1082717_comb];
  assign p6_array_index_1082734_comb = p5_literal_1076355[p6_array_index_1082718_comb];
  assign p6_array_index_1082735_comb = p5_arr[p6_addedKey__62_comb[79:72]];
  assign p6_array_index_1082737_comb = p5_arr[p6_addedKey__62_comb[63:56]];
  assign p6_res7__336_comb = p6_array_index_1082729_comb ^ p6_array_index_1082730_comb ^ p6_array_index_1082731_comb ^ p6_array_index_1082732_comb ^ p6_array_index_1082733_comb ^ p6_array_index_1082734_comb ^ p6_array_index_1082735_comb ^ p5_literal_1076358[p6_array_index_1082720_comb] ^ p6_array_index_1082737_comb ^ p5_literal_1076355[p6_array_index_1082722_comb] ^ p5_literal_1076353[p6_array_index_1082723_comb] ^ p5_literal_1076351[p6_array_index_1082724_comb] ^ p5_literal_1076349[p6_array_index_1082725_comb] ^ p5_literal_1076347[p6_array_index_1082726_comb] ^ p5_literal_1076345[p6_array_index_1082727_comb] ^ p5_arr[p6_addedKey__62_comb[7:0]];
  assign p6_array_index_1082746_comb = p5_literal_1076345[p6_res7__336_comb];
  assign p6_array_index_1082747_comb = p5_literal_1076347[p6_array_index_1082713_comb];
  assign p6_array_index_1082748_comb = p5_literal_1076349[p6_array_index_1082714_comb];
  assign p6_array_index_1082749_comb = p5_literal_1076351[p6_array_index_1082715_comb];
  assign p6_array_index_1082750_comb = p5_literal_1076353[p6_array_index_1082716_comb];
  assign p6_array_index_1082751_comb = p5_literal_1076355[p6_array_index_1082717_comb];
  assign p6_res7__337_comb = p6_array_index_1082746_comb ^ p6_array_index_1082747_comb ^ p6_array_index_1082748_comb ^ p6_array_index_1082749_comb ^ p6_array_index_1082750_comb ^ p6_array_index_1082751_comb ^ p6_array_index_1082718_comb ^ p5_literal_1076358[p6_array_index_1082735_comb] ^ p6_array_index_1082720_comb ^ p5_literal_1076355[p6_array_index_1082737_comb] ^ p5_literal_1076353[p6_array_index_1082722_comb] ^ p5_literal_1076351[p6_array_index_1082723_comb] ^ p5_literal_1076349[p6_array_index_1082724_comb] ^ p5_literal_1076347[p6_array_index_1082725_comb] ^ p5_literal_1076345[p6_array_index_1082726_comb] ^ p6_array_index_1082727_comb;
  assign p6_array_index_1082761_comb = p5_literal_1076347[p6_res7__336_comb];
  assign p6_array_index_1082762_comb = p5_literal_1076349[p6_array_index_1082713_comb];
  assign p6_array_index_1082763_comb = p5_literal_1076351[p6_array_index_1082714_comb];
  assign p6_array_index_1082764_comb = p5_literal_1076353[p6_array_index_1082715_comb];
  assign p6_array_index_1082765_comb = p5_literal_1076355[p6_array_index_1082716_comb];
  assign p6_res7__338_comb = p5_literal_1076345[p6_res7__337_comb] ^ p6_array_index_1082761_comb ^ p6_array_index_1082762_comb ^ p6_array_index_1082763_comb ^ p6_array_index_1082764_comb ^ p6_array_index_1082765_comb ^ p6_array_index_1082717_comb ^ p5_literal_1076358[p6_array_index_1082718_comb] ^ p6_array_index_1082735_comb ^ p5_literal_1076355[p6_array_index_1082720_comb] ^ p5_literal_1076353[p6_array_index_1082737_comb] ^ p5_literal_1076351[p6_array_index_1082722_comb] ^ p5_literal_1076349[p6_array_index_1082723_comb] ^ p5_literal_1076347[p6_array_index_1082724_comb] ^ p5_literal_1076345[p6_array_index_1082725_comb] ^ p6_array_index_1082726_comb;
  assign p6_array_index_1082775_comb = p5_literal_1076347[p6_res7__337_comb];
  assign p6_array_index_1082776_comb = p5_literal_1076349[p6_res7__336_comb];
  assign p6_array_index_1082777_comb = p5_literal_1076351[p6_array_index_1082713_comb];
  assign p6_array_index_1082778_comb = p5_literal_1076353[p6_array_index_1082714_comb];
  assign p6_array_index_1082779_comb = p5_literal_1076355[p6_array_index_1082715_comb];
  assign p6_res7__339_comb = p5_literal_1076345[p6_res7__338_comb] ^ p6_array_index_1082775_comb ^ p6_array_index_1082776_comb ^ p6_array_index_1082777_comb ^ p6_array_index_1082778_comb ^ p6_array_index_1082779_comb ^ p6_array_index_1082716_comb ^ p5_literal_1076358[p6_array_index_1082717_comb] ^ p6_array_index_1082718_comb ^ p5_literal_1076355[p6_array_index_1082735_comb] ^ p5_literal_1076353[p6_array_index_1082720_comb] ^ p5_literal_1076351[p6_array_index_1082737_comb] ^ p5_literal_1076349[p6_array_index_1082722_comb] ^ p5_literal_1076347[p6_array_index_1082723_comb] ^ p5_literal_1076345[p6_array_index_1082724_comb] ^ p6_array_index_1082725_comb;
  assign p6_array_index_1082790_comb = p5_literal_1076349[p6_res7__337_comb];
  assign p6_array_index_1082791_comb = p5_literal_1076351[p6_res7__336_comb];
  assign p6_array_index_1082792_comb = p5_literal_1076353[p6_array_index_1082713_comb];
  assign p6_array_index_1082793_comb = p5_literal_1076355[p6_array_index_1082714_comb];
  assign p6_res7__340_comb = p5_literal_1076345[p6_res7__339_comb] ^ p5_literal_1076347[p6_res7__338_comb] ^ p6_array_index_1082790_comb ^ p6_array_index_1082791_comb ^ p6_array_index_1082792_comb ^ p6_array_index_1082793_comb ^ p6_array_index_1082715_comb ^ p5_literal_1076358[p6_array_index_1082716_comb] ^ p6_array_index_1082717_comb ^ p6_array_index_1082734_comb ^ p5_literal_1076353[p6_array_index_1082735_comb] ^ p5_literal_1076351[p6_array_index_1082720_comb] ^ p5_literal_1076349[p6_array_index_1082737_comb] ^ p5_literal_1076347[p6_array_index_1082722_comb] ^ p5_literal_1076345[p6_array_index_1082723_comb] ^ p6_array_index_1082724_comb;
  assign p6_array_index_1082803_comb = p5_literal_1076349[p6_res7__338_comb];
  assign p6_array_index_1082804_comb = p5_literal_1076351[p6_res7__337_comb];
  assign p6_array_index_1082805_comb = p5_literal_1076353[p6_res7__336_comb];
  assign p6_array_index_1082806_comb = p5_literal_1076355[p6_array_index_1082713_comb];
  assign p6_res7__341_comb = p5_literal_1076345[p6_res7__340_comb] ^ p5_literal_1076347[p6_res7__339_comb] ^ p6_array_index_1082803_comb ^ p6_array_index_1082804_comb ^ p6_array_index_1082805_comb ^ p6_array_index_1082806_comb ^ p6_array_index_1082714_comb ^ p5_literal_1076358[p6_array_index_1082715_comb] ^ p6_array_index_1082716_comb ^ p6_array_index_1082751_comb ^ p5_literal_1076353[p6_array_index_1082718_comb] ^ p5_literal_1076351[p6_array_index_1082735_comb] ^ p5_literal_1076349[p6_array_index_1082720_comb] ^ p5_literal_1076347[p6_array_index_1082737_comb] ^ p5_literal_1076345[p6_array_index_1082722_comb] ^ p6_array_index_1082723_comb;
  assign p6_array_index_1082817_comb = p5_literal_1076351[p6_res7__338_comb];
  assign p6_array_index_1082818_comb = p5_literal_1076353[p6_res7__337_comb];
  assign p6_array_index_1082819_comb = p5_literal_1076355[p6_res7__336_comb];
  assign p6_res7__342_comb = p5_literal_1076345[p6_res7__341_comb] ^ p5_literal_1076347[p6_res7__340_comb] ^ p5_literal_1076349[p6_res7__339_comb] ^ p6_array_index_1082817_comb ^ p6_array_index_1082818_comb ^ p6_array_index_1082819_comb ^ p6_array_index_1082713_comb ^ p5_literal_1076358[p6_array_index_1082714_comb] ^ p6_array_index_1082715_comb ^ p6_array_index_1082765_comb ^ p6_array_index_1082733_comb ^ p5_literal_1076351[p6_array_index_1082718_comb] ^ p5_literal_1076349[p6_array_index_1082735_comb] ^ p5_literal_1076347[p6_array_index_1082720_comb] ^ p5_literal_1076345[p6_array_index_1082737_comb] ^ p6_array_index_1082722_comb;
  assign p6_array_index_1082829_comb = p5_literal_1076351[p6_res7__339_comb];
  assign p6_array_index_1082830_comb = p5_literal_1076353[p6_res7__338_comb];
  assign p6_array_index_1082831_comb = p5_literal_1076355[p6_res7__337_comb];
  assign p6_res7__343_comb = p5_literal_1076345[p6_res7__342_comb] ^ p5_literal_1076347[p6_res7__341_comb] ^ p5_literal_1076349[p6_res7__340_comb] ^ p6_array_index_1082829_comb ^ p6_array_index_1082830_comb ^ p6_array_index_1082831_comb ^ p6_res7__336_comb ^ p5_literal_1076358[p6_array_index_1082713_comb] ^ p6_array_index_1082714_comb ^ p6_array_index_1082779_comb ^ p6_array_index_1082750_comb ^ p5_literal_1076351[p6_array_index_1082717_comb] ^ p5_literal_1076349[p6_array_index_1082718_comb] ^ p5_literal_1076347[p6_array_index_1082735_comb] ^ p5_literal_1076345[p6_array_index_1082720_comb] ^ p6_array_index_1082737_comb;
  assign p6_array_index_1082842_comb = p5_literal_1076353[p6_res7__339_comb];
  assign p6_array_index_1082843_comb = p5_literal_1076355[p6_res7__338_comb];
  assign p6_res7__344_comb = p5_literal_1076345[p6_res7__343_comb] ^ p5_literal_1076347[p6_res7__342_comb] ^ p5_literal_1076349[p6_res7__341_comb] ^ p5_literal_1076351[p6_res7__340_comb] ^ p6_array_index_1082842_comb ^ p6_array_index_1082843_comb ^ p6_res7__337_comb ^ p5_literal_1076358[p6_res7__336_comb] ^ p6_array_index_1082713_comb ^ p6_array_index_1082793_comb ^ p6_array_index_1082764_comb ^ p6_array_index_1082732_comb ^ p5_literal_1076349[p6_array_index_1082717_comb] ^ p5_literal_1076347[p6_array_index_1082718_comb] ^ p5_literal_1076345[p6_array_index_1082735_comb] ^ p6_array_index_1082720_comb;
  assign p6_array_index_1082853_comb = p5_literal_1076353[p6_res7__340_comb];
  assign p6_array_index_1082854_comb = p5_literal_1076355[p6_res7__339_comb];
  assign p6_res7__345_comb = p5_literal_1076345[p6_res7__344_comb] ^ p5_literal_1076347[p6_res7__343_comb] ^ p5_literal_1076349[p6_res7__342_comb] ^ p5_literal_1076351[p6_res7__341_comb] ^ p6_array_index_1082853_comb ^ p6_array_index_1082854_comb ^ p6_res7__338_comb ^ p5_literal_1076358[p6_res7__337_comb] ^ p6_res7__336_comb ^ p6_array_index_1082806_comb ^ p6_array_index_1082778_comb ^ p6_array_index_1082749_comb ^ p5_literal_1076349[p6_array_index_1082716_comb] ^ p5_literal_1076347[p6_array_index_1082717_comb] ^ p5_literal_1076345[p6_array_index_1082718_comb] ^ p6_array_index_1082735_comb;
  assign p6_array_index_1082865_comb = p5_literal_1076355[p6_res7__340_comb];
  assign p6_res7__346_comb = p5_literal_1076345[p6_res7__345_comb] ^ p5_literal_1076347[p6_res7__344_comb] ^ p5_literal_1076349[p6_res7__343_comb] ^ p5_literal_1076351[p6_res7__342_comb] ^ p5_literal_1076353[p6_res7__341_comb] ^ p6_array_index_1082865_comb ^ p6_res7__339_comb ^ p5_literal_1076358[p6_res7__338_comb] ^ p6_res7__337_comb ^ p6_array_index_1082819_comb ^ p6_array_index_1082792_comb ^ p6_array_index_1082763_comb ^ p6_array_index_1082731_comb ^ p5_literal_1076347[p6_array_index_1082716_comb] ^ p5_literal_1076345[p6_array_index_1082717_comb] ^ p6_array_index_1082718_comb;
  assign p6_array_index_1082875_comb = p5_literal_1076355[p6_res7__341_comb];
  assign p6_res7__347_comb = p5_literal_1076345[p6_res7__346_comb] ^ p5_literal_1076347[p6_res7__345_comb] ^ p5_literal_1076349[p6_res7__344_comb] ^ p5_literal_1076351[p6_res7__343_comb] ^ p5_literal_1076353[p6_res7__342_comb] ^ p6_array_index_1082875_comb ^ p6_res7__340_comb ^ p5_literal_1076358[p6_res7__339_comb] ^ p6_res7__338_comb ^ p6_array_index_1082831_comb ^ p6_array_index_1082805_comb ^ p6_array_index_1082777_comb ^ p6_array_index_1082748_comb ^ p5_literal_1076347[p6_array_index_1082715_comb] ^ p5_literal_1076345[p6_array_index_1082716_comb] ^ p6_array_index_1082717_comb;
  assign p6_res7__348_comb = p5_literal_1076345[p6_res7__347_comb] ^ p5_literal_1076347[p6_res7__346_comb] ^ p5_literal_1076349[p6_res7__345_comb] ^ p5_literal_1076351[p6_res7__344_comb] ^ p5_literal_1076353[p6_res7__343_comb] ^ p5_literal_1076355[p6_res7__342_comb] ^ p6_res7__341_comb ^ p5_literal_1076358[p6_res7__340_comb] ^ p6_res7__339_comb ^ p6_array_index_1082843_comb ^ p6_array_index_1082818_comb ^ p6_array_index_1082791_comb ^ p6_array_index_1082762_comb ^ p6_array_index_1082730_comb ^ p5_literal_1076345[p6_array_index_1082715_comb] ^ p6_array_index_1082716_comb;
  assign p6_res7__349_comb = p5_literal_1076345[p6_res7__348_comb] ^ p5_literal_1076347[p6_res7__347_comb] ^ p5_literal_1076349[p6_res7__346_comb] ^ p5_literal_1076351[p6_res7__345_comb] ^ p5_literal_1076353[p6_res7__344_comb] ^ p5_literal_1076355[p6_res7__343_comb] ^ p6_res7__342_comb ^ p5_literal_1076358[p6_res7__341_comb] ^ p6_res7__340_comb ^ p6_array_index_1082854_comb ^ p6_array_index_1082830_comb ^ p6_array_index_1082804_comb ^ p6_array_index_1082776_comb ^ p6_array_index_1082747_comb ^ p5_literal_1076345[p6_array_index_1082714_comb] ^ p6_array_index_1082715_comb;
  assign p6_res7__350_comb = p5_literal_1076345[p6_res7__349_comb] ^ p5_literal_1076347[p6_res7__348_comb] ^ p5_literal_1076349[p6_res7__347_comb] ^ p5_literal_1076351[p6_res7__346_comb] ^ p5_literal_1076353[p6_res7__345_comb] ^ p5_literal_1076355[p6_res7__344_comb] ^ p6_res7__343_comb ^ p5_literal_1076358[p6_res7__342_comb] ^ p6_res7__341_comb ^ p6_array_index_1082865_comb ^ p6_array_index_1082842_comb ^ p6_array_index_1082817_comb ^ p6_array_index_1082790_comb ^ p6_array_index_1082761_comb ^ p6_array_index_1082729_comb ^ p6_array_index_1082714_comb;
  assign p6_res7__351_comb = p5_literal_1076345[p6_res7__350_comb] ^ p5_literal_1076347[p6_res7__349_comb] ^ p5_literal_1076349[p6_res7__348_comb] ^ p5_literal_1076351[p6_res7__347_comb] ^ p5_literal_1076353[p6_res7__346_comb] ^ p5_literal_1076355[p6_res7__345_comb] ^ p6_res7__344_comb ^ p5_literal_1076358[p6_res7__343_comb] ^ p6_res7__342_comb ^ p6_array_index_1082875_comb ^ p6_array_index_1082853_comb ^ p6_array_index_1082829_comb ^ p6_array_index_1082803_comb ^ p6_array_index_1082775_comb ^ p6_array_index_1082746_comb ^ p6_array_index_1082713_comb;
  assign p6_res__21_comb = {p6_res7__351_comb, p6_res7__350_comb, p6_res7__349_comb, p6_res7__348_comb, p6_res7__347_comb, p6_res7__346_comb, p6_res7__345_comb, p6_res7__344_comb, p6_res7__343_comb, p6_res7__342_comb, p6_res7__341_comb, p6_res7__340_comb, p6_res7__339_comb, p6_res7__338_comb, p6_res7__337_comb, p6_res7__336_comb};
  assign p6_xor_1082915_comb = p6_res__21_comb ^ p6_xor_1082479_comb;

  // Registers for pipe stage 6:
  reg [127:0] p6_xor_1082697;
  reg [127:0] p6_xor_1082915;
  reg [127:0] p6_res__37;
  reg [7:0] p7_arr[256];
  reg [7:0] p7_literal_1076345[256];
  reg [7:0] p7_literal_1076347[256];
  reg [7:0] p7_literal_1076349[256];
  reg [7:0] p7_literal_1076351[256];
  reg [7:0] p7_literal_1076353[256];
  reg [7:0] p7_literal_1076355[256];
  reg [7:0] p7_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p6_xor_1082697 <= p6_xor_1082697_comb;
    p6_xor_1082915 <= p6_xor_1082915_comb;
    p6_res__37 <= p5_res__37;
    p7_arr <= p6_arr;
    p7_literal_1076345 <= p6_literal_1076345;
    p7_literal_1076347 <= p6_literal_1076347;
    p7_literal_1076349 <= p6_literal_1076349;
    p7_literal_1076351 <= p6_literal_1076351;
    p7_literal_1076353 <= p6_literal_1076353;
    p7_literal_1076355 <= p6_literal_1076355;
    p7_literal_1076358 <= p6_literal_1076358;
  end

  // ===== Pipe stage 7:
  wire [127:0] p7_addedKey__63_comb;
  wire [7:0] p7_array_index_1082953_comb;
  wire [7:0] p7_array_index_1082954_comb;
  wire [7:0] p7_array_index_1082955_comb;
  wire [7:0] p7_array_index_1082956_comb;
  wire [7:0] p7_array_index_1082957_comb;
  wire [7:0] p7_array_index_1082958_comb;
  wire [7:0] p7_array_index_1082960_comb;
  wire [7:0] p7_array_index_1082962_comb;
  wire [7:0] p7_array_index_1082963_comb;
  wire [7:0] p7_array_index_1082964_comb;
  wire [7:0] p7_array_index_1082965_comb;
  wire [7:0] p7_array_index_1082966_comb;
  wire [7:0] p7_array_index_1082967_comb;
  wire [7:0] p7_array_index_1082969_comb;
  wire [7:0] p7_array_index_1082970_comb;
  wire [7:0] p7_array_index_1082971_comb;
  wire [7:0] p7_array_index_1082972_comb;
  wire [7:0] p7_array_index_1082973_comb;
  wire [7:0] p7_array_index_1082974_comb;
  wire [7:0] p7_array_index_1082975_comb;
  wire [7:0] p7_array_index_1082977_comb;
  wire [7:0] p7_res7__352_comb;
  wire [7:0] p7_array_index_1082986_comb;
  wire [7:0] p7_array_index_1082987_comb;
  wire [7:0] p7_array_index_1082988_comb;
  wire [7:0] p7_array_index_1082989_comb;
  wire [7:0] p7_array_index_1082990_comb;
  wire [7:0] p7_array_index_1082991_comb;
  wire [7:0] p7_res7__353_comb;
  wire [7:0] p7_array_index_1083001_comb;
  wire [7:0] p7_array_index_1083002_comb;
  wire [7:0] p7_array_index_1083003_comb;
  wire [7:0] p7_array_index_1083004_comb;
  wire [7:0] p7_array_index_1083005_comb;
  wire [7:0] p7_res7__354_comb;
  wire [7:0] p7_array_index_1083015_comb;
  wire [7:0] p7_array_index_1083016_comb;
  wire [7:0] p7_array_index_1083017_comb;
  wire [7:0] p7_array_index_1083018_comb;
  wire [7:0] p7_array_index_1083019_comb;
  wire [7:0] p7_res7__355_comb;
  wire [7:0] p7_array_index_1083030_comb;
  wire [7:0] p7_array_index_1083031_comb;
  wire [7:0] p7_array_index_1083032_comb;
  wire [7:0] p7_array_index_1083033_comb;
  wire [7:0] p7_res7__356_comb;
  wire [7:0] p7_array_index_1083043_comb;
  wire [7:0] p7_array_index_1083044_comb;
  wire [7:0] p7_array_index_1083045_comb;
  wire [7:0] p7_array_index_1083046_comb;
  wire [7:0] p7_res7__357_comb;
  wire [7:0] p7_array_index_1083057_comb;
  wire [7:0] p7_array_index_1083058_comb;
  wire [7:0] p7_array_index_1083059_comb;
  wire [7:0] p7_res7__358_comb;
  wire [7:0] p7_array_index_1083069_comb;
  wire [7:0] p7_array_index_1083070_comb;
  wire [7:0] p7_array_index_1083071_comb;
  wire [7:0] p7_res7__359_comb;
  wire [7:0] p7_array_index_1083082_comb;
  wire [7:0] p7_array_index_1083083_comb;
  wire [7:0] p7_res7__360_comb;
  wire [7:0] p7_array_index_1083093_comb;
  wire [7:0] p7_array_index_1083094_comb;
  wire [7:0] p7_res7__361_comb;
  wire [7:0] p7_array_index_1083105_comb;
  wire [7:0] p7_res7__362_comb;
  wire [7:0] p7_array_index_1083115_comb;
  wire [7:0] p7_res7__363_comb;
  wire [7:0] p7_res7__364_comb;
  wire [7:0] p7_res7__365_comb;
  wire [7:0] p7_res7__366_comb;
  wire [7:0] p7_res7__367_comb;
  wire [127:0] p7_res__22_comb;
  wire [127:0] p7_k7_comb;
  wire [127:0] p7_addedKey__64_comb;
  wire [7:0] p7_array_index_1083171_comb;
  wire [7:0] p7_array_index_1083172_comb;
  wire [7:0] p7_array_index_1083173_comb;
  wire [7:0] p7_array_index_1083174_comb;
  wire [7:0] p7_array_index_1083175_comb;
  wire [7:0] p7_array_index_1083176_comb;
  wire [7:0] p7_array_index_1083178_comb;
  wire [7:0] p7_array_index_1083180_comb;
  wire [7:0] p7_array_index_1083181_comb;
  wire [7:0] p7_array_index_1083182_comb;
  wire [7:0] p7_array_index_1083183_comb;
  wire [7:0] p7_array_index_1083184_comb;
  wire [7:0] p7_array_index_1083185_comb;
  wire [7:0] p7_array_index_1083187_comb;
  wire [7:0] p7_array_index_1083188_comb;
  wire [7:0] p7_array_index_1083189_comb;
  wire [7:0] p7_array_index_1083190_comb;
  wire [7:0] p7_array_index_1083191_comb;
  wire [7:0] p7_array_index_1083192_comb;
  wire [7:0] p7_array_index_1083193_comb;
  wire [7:0] p7_array_index_1083195_comb;
  wire [7:0] p7_res7__368_comb;
  wire [7:0] p7_array_index_1083204_comb;
  wire [7:0] p7_array_index_1083205_comb;
  wire [7:0] p7_array_index_1083206_comb;
  wire [7:0] p7_array_index_1083207_comb;
  wire [7:0] p7_array_index_1083208_comb;
  wire [7:0] p7_array_index_1083209_comb;
  wire [7:0] p7_res7__369_comb;
  wire [7:0] p7_array_index_1083219_comb;
  wire [7:0] p7_array_index_1083220_comb;
  wire [7:0] p7_array_index_1083221_comb;
  wire [7:0] p7_array_index_1083222_comb;
  wire [7:0] p7_array_index_1083223_comb;
  wire [7:0] p7_res7__370_comb;
  wire [7:0] p7_array_index_1083233_comb;
  wire [7:0] p7_array_index_1083234_comb;
  wire [7:0] p7_array_index_1083235_comb;
  wire [7:0] p7_array_index_1083236_comb;
  wire [7:0] p7_array_index_1083237_comb;
  wire [7:0] p7_res7__371_comb;
  wire [7:0] p7_array_index_1083248_comb;
  wire [7:0] p7_array_index_1083249_comb;
  wire [7:0] p7_array_index_1083250_comb;
  wire [7:0] p7_array_index_1083251_comb;
  wire [7:0] p7_res7__372_comb;
  wire [7:0] p7_array_index_1083261_comb;
  wire [7:0] p7_array_index_1083262_comb;
  wire [7:0] p7_array_index_1083263_comb;
  wire [7:0] p7_array_index_1083264_comb;
  wire [7:0] p7_res7__373_comb;
  wire [7:0] p7_array_index_1083275_comb;
  wire [7:0] p7_array_index_1083276_comb;
  wire [7:0] p7_array_index_1083277_comb;
  wire [7:0] p7_res7__374_comb;
  wire [7:0] p7_array_index_1083287_comb;
  wire [7:0] p7_array_index_1083288_comb;
  wire [7:0] p7_array_index_1083289_comb;
  wire [7:0] p7_res7__375_comb;
  wire [7:0] p7_array_index_1083300_comb;
  wire [7:0] p7_array_index_1083301_comb;
  wire [7:0] p7_res7__376_comb;
  wire [7:0] p7_array_index_1083311_comb;
  wire [7:0] p7_array_index_1083312_comb;
  wire [7:0] p7_res7__377_comb;
  wire [7:0] p7_array_index_1083323_comb;
  wire [7:0] p7_res7__378_comb;
  wire [7:0] p7_array_index_1083333_comb;
  wire [7:0] p7_res7__379_comb;
  wire [7:0] p7_res7__380_comb;
  wire [7:0] p7_res7__381_comb;
  wire [7:0] p7_res7__382_comb;
  wire [7:0] p7_res7__383_comb;
  wire [127:0] p7_res__23_comb;
  wire [127:0] p7_k6_comb;
  wire [127:0] p7_addedKey__65_comb;
  wire [7:0] p7_array_index_1083389_comb;
  wire [7:0] p7_array_index_1083390_comb;
  wire [7:0] p7_array_index_1083391_comb;
  wire [7:0] p7_array_index_1083392_comb;
  wire [7:0] p7_array_index_1083393_comb;
  wire [7:0] p7_array_index_1083394_comb;
  wire [7:0] p7_array_index_1083396_comb;
  wire [7:0] p7_array_index_1083398_comb;
  wire [7:0] p7_array_index_1083399_comb;
  wire [7:0] p7_array_index_1083400_comb;
  wire [7:0] p7_array_index_1083401_comb;
  wire [7:0] p7_array_index_1083402_comb;
  wire [7:0] p7_array_index_1083403_comb;
  wire [7:0] p7_array_index_1083405_comb;
  wire [7:0] p7_array_index_1083406_comb;
  wire [7:0] p7_array_index_1083407_comb;
  wire [7:0] p7_array_index_1083408_comb;
  wire [7:0] p7_array_index_1083409_comb;
  wire [7:0] p7_array_index_1083410_comb;
  wire [7:0] p7_array_index_1083411_comb;
  wire [7:0] p7_array_index_1083413_comb;
  wire [7:0] p7_res7__384_comb;
  wire [7:0] p7_array_index_1083422_comb;
  wire [7:0] p7_array_index_1083423_comb;
  wire [7:0] p7_array_index_1083424_comb;
  wire [7:0] p7_array_index_1083425_comb;
  wire [7:0] p7_array_index_1083426_comb;
  wire [7:0] p7_array_index_1083427_comb;
  wire [7:0] p7_res7__385_comb;
  wire [7:0] p7_array_index_1083437_comb;
  wire [7:0] p7_array_index_1083438_comb;
  wire [7:0] p7_array_index_1083439_comb;
  wire [7:0] p7_array_index_1083440_comb;
  wire [7:0] p7_array_index_1083441_comb;
  wire [7:0] p7_res7__386_comb;
  wire [7:0] p7_array_index_1083451_comb;
  wire [7:0] p7_array_index_1083452_comb;
  wire [7:0] p7_array_index_1083453_comb;
  wire [7:0] p7_array_index_1083454_comb;
  wire [7:0] p7_array_index_1083455_comb;
  wire [7:0] p7_res7__387_comb;
  wire [7:0] p7_array_index_1083466_comb;
  wire [7:0] p7_array_index_1083467_comb;
  wire [7:0] p7_array_index_1083468_comb;
  wire [7:0] p7_array_index_1083469_comb;
  wire [7:0] p7_res7__388_comb;
  wire [7:0] p7_array_index_1083479_comb;
  wire [7:0] p7_array_index_1083480_comb;
  wire [7:0] p7_array_index_1083481_comb;
  wire [7:0] p7_array_index_1083482_comb;
  wire [7:0] p7_res7__389_comb;
  wire [7:0] p7_array_index_1083493_comb;
  wire [7:0] p7_array_index_1083494_comb;
  wire [7:0] p7_array_index_1083495_comb;
  wire [7:0] p7_res7__390_comb;
  wire [7:0] p7_array_index_1083505_comb;
  wire [7:0] p7_array_index_1083506_comb;
  wire [7:0] p7_array_index_1083507_comb;
  wire [7:0] p7_res7__391_comb;
  wire [7:0] p7_array_index_1083518_comb;
  wire [7:0] p7_array_index_1083519_comb;
  wire [7:0] p7_res7__392_comb;
  wire [7:0] p7_array_index_1083529_comb;
  wire [7:0] p7_array_index_1083530_comb;
  wire [7:0] p7_res7__393_comb;
  wire [127:0] p7_addedKey__38_comb;
  wire [7:0] p7_array_index_1083541_comb;
  wire [7:0] p7_res7__394_comb;
  wire [7:0] p7_array_index_1083777_comb;
  wire [7:0] p7_array_index_1083778_comb;
  wire [7:0] p7_array_index_1083779_comb;
  wire [7:0] p7_array_index_1083780_comb;
  wire [7:0] p7_array_index_1083781_comb;
  wire [7:0] p7_array_index_1083782_comb;
  wire [7:0] p7_array_index_1083784_comb;
  wire [7:0] p7_array_index_1083786_comb;
  wire [7:0] p7_array_index_1083787_comb;
  wire [7:0] p7_array_index_1083788_comb;
  wire [7:0] p7_array_index_1083789_comb;
  wire [7:0] p7_array_index_1083790_comb;
  wire [7:0] p7_array_index_1083791_comb;
  wire [7:0] p7_array_index_1083551_comb;
  wire [7:0] p7_array_index_1083793_comb;
  wire [7:0] p7_array_index_1083794_comb;
  wire [7:0] p7_array_index_1083795_comb;
  wire [7:0] p7_array_index_1083796_comb;
  wire [7:0] p7_array_index_1083797_comb;
  wire [7:0] p7_array_index_1083798_comb;
  wire [7:0] p7_array_index_1083799_comb;
  wire [7:0] p7_array_index_1083801_comb;
  wire [7:0] p7_res7__395_comb;
  wire [7:0] p7_res7__608_comb;
  wire [7:0] p7_array_index_1083810_comb;
  wire [7:0] p7_array_index_1083811_comb;
  wire [7:0] p7_array_index_1083812_comb;
  wire [7:0] p7_array_index_1083813_comb;
  wire [7:0] p7_array_index_1083814_comb;
  wire [7:0] p7_array_index_1083815_comb;
  wire [7:0] p7_res7__396_comb;
  wire [7:0] p7_res7__609_comb;
  wire [7:0] p7_array_index_1083825_comb;
  wire [7:0] p7_array_index_1083826_comb;
  wire [7:0] p7_array_index_1083827_comb;
  wire [7:0] p7_array_index_1083828_comb;
  wire [7:0] p7_array_index_1083829_comb;
  wire [7:0] p7_res7__397_comb;
  wire [7:0] p7_res7__610_comb;
  wire [7:0] p7_array_index_1083839_comb;
  wire [7:0] p7_array_index_1083840_comb;
  wire [7:0] p7_array_index_1083841_comb;
  wire [7:0] p7_array_index_1083842_comb;
  wire [7:0] p7_array_index_1083843_comb;
  wire [7:0] p7_res7__398_comb;
  wire [7:0] p7_res7__611_comb;
  wire [7:0] p7_array_index_1083854_comb;
  wire [7:0] p7_array_index_1083855_comb;
  wire [7:0] p7_array_index_1083856_comb;
  wire [7:0] p7_array_index_1083857_comb;
  wire [7:0] p7_res7__399_comb;
  wire [7:0] p7_res7__612_comb;
  wire [127:0] p7_res__24_comb;
  wire [7:0] p7_array_index_1083867_comb;
  wire [7:0] p7_array_index_1083868_comb;
  wire [7:0] p7_array_index_1083869_comb;
  wire [7:0] p7_array_index_1083870_comb;
  wire [127:0] p7_xor_1083591_comb;
  wire [7:0] p7_res7__613_comb;
  wire [127:0] p7_addedKey__66_comb;
  wire [7:0] p7_array_index_1083881_comb;
  wire [7:0] p7_array_index_1083882_comb;
  wire [7:0] p7_array_index_1083883_comb;
  wire [7:0] p7_res7__614_comb;
  wire [7:0] p7_array_index_1083607_comb;
  wire [7:0] p7_array_index_1083608_comb;
  wire [7:0] p7_array_index_1083609_comb;
  wire [7:0] p7_array_index_1083610_comb;
  wire [7:0] p7_array_index_1083611_comb;
  wire [7:0] p7_array_index_1083612_comb;
  wire [7:0] p7_array_index_1083614_comb;
  wire [7:0] p7_array_index_1083616_comb;
  wire [7:0] p7_array_index_1083617_comb;
  wire [7:0] p7_array_index_1083618_comb;
  wire [7:0] p7_array_index_1083619_comb;
  wire [7:0] p7_array_index_1083620_comb;
  wire [7:0] p7_array_index_1083621_comb;
  wire [7:0] p7_array_index_1083893_comb;
  wire [7:0] p7_array_index_1083894_comb;
  wire [7:0] p7_array_index_1083895_comb;
  wire [7:0] p7_array_index_1083623_comb;
  wire [7:0] p7_array_index_1083624_comb;
  wire [7:0] p7_array_index_1083625_comb;
  wire [7:0] p7_array_index_1083626_comb;
  wire [7:0] p7_array_index_1083627_comb;
  wire [7:0] p7_array_index_1083628_comb;
  wire [7:0] p7_array_index_1083629_comb;
  wire [7:0] p7_array_index_1083631_comb;
  wire [7:0] p7_res7__615_comb;
  wire [7:0] p7_res7__400_comb;
  wire [7:0] p7_array_index_1083906_comb;
  wire [7:0] p7_array_index_1083907_comb;
  wire [7:0] p7_array_index_1083640_comb;
  wire [7:0] p7_array_index_1083641_comb;
  wire [7:0] p7_array_index_1083642_comb;
  wire [7:0] p7_array_index_1083643_comb;
  wire [7:0] p7_array_index_1083644_comb;
  wire [7:0] p7_array_index_1083645_comb;
  wire [7:0] p7_res7__616_comb;
  wire [7:0] p7_res7__401_comb;
  wire [7:0] p7_array_index_1083917_comb;
  wire [7:0] p7_array_index_1083918_comb;
  wire [7:0] p7_array_index_1083655_comb;
  wire [7:0] p7_array_index_1083656_comb;
  wire [7:0] p7_array_index_1083657_comb;
  wire [7:0] p7_array_index_1083658_comb;
  wire [7:0] p7_array_index_1083659_comb;
  wire [7:0] p7_res7__617_comb;
  wire [7:0] p7_res7__402_comb;
  wire [7:0] p7_array_index_1083929_comb;
  wire [7:0] p7_array_index_1083669_comb;
  wire [7:0] p7_array_index_1083670_comb;
  wire [7:0] p7_array_index_1083671_comb;
  wire [7:0] p7_array_index_1083672_comb;
  wire [7:0] p7_array_index_1083673_comb;
  wire [7:0] p7_res7__618_comb;
  wire [7:0] p7_res7__403_comb;
  wire [7:0] p7_array_index_1083939_comb;
  wire [7:0] p7_array_index_1083684_comb;
  wire [7:0] p7_array_index_1083685_comb;
  wire [7:0] p7_array_index_1083686_comb;
  wire [7:0] p7_array_index_1083687_comb;
  wire [7:0] p7_res7__619_comb;
  wire [7:0] p7_res7__404_comb;
  wire [7:0] p7_array_index_1083697_comb;
  wire [7:0] p7_array_index_1083698_comb;
  wire [7:0] p7_array_index_1083699_comb;
  wire [7:0] p7_array_index_1083700_comb;
  wire [7:0] p7_res7__620_comb;
  wire [7:0] p7_res7__405_comb;
  wire [7:0] p7_array_index_1083711_comb;
  wire [7:0] p7_array_index_1083712_comb;
  wire [7:0] p7_array_index_1083713_comb;
  wire [7:0] p7_res7__621_comb;
  wire [7:0] p7_res7__406_comb;
  wire [7:0] p7_array_index_1083723_comb;
  wire [7:0] p7_array_index_1083724_comb;
  wire [7:0] p7_array_index_1083725_comb;
  wire [7:0] p7_res7__622_comb;
  wire [7:0] p7_res7__407_comb;
  wire [7:0] p7_array_index_1083736_comb;
  wire [7:0] p7_array_index_1083737_comb;
  wire [7:0] p7_res7__623_comb;
  wire [7:0] p7_res7__408_comb;
  wire [127:0] p7_res__38_comb;
  wire [7:0] p7_array_index_1083747_comb;
  wire [7:0] p7_array_index_1083748_comb;
  wire [127:0] p7_addedKey__39_comb;
  wire [7:0] p7_res7__409_comb;
  wire [7:0] p7_array_index_1083754_comb;
  wire [7:0] p7_array_index_1083755_comb;
  wire [7:0] p7_array_index_1083756_comb;
  wire [7:0] p7_array_index_1083757_comb;
  wire [7:0] p7_array_index_1083758_comb;
  wire [7:0] p7_array_index_1083759_comb;
  wire [7:0] p7_array_index_1083760_comb;
  wire [7:0] p7_array_index_1083761_comb;
  wire [7:0] p7_array_index_1083762_comb;
  wire [7:0] p7_array_index_1083993_comb;
  wire [7:0] p7_array_index_1083994_comb;
  wire [7:0] p7_array_index_1083995_comb;
  wire [7:0] p7_array_index_1083996_comb;
  wire [7:0] p7_array_index_1083997_comb;
  wire [7:0] p7_array_index_1083998_comb;
  wire [7:0] p7_array_index_1084000_comb;
  wire [7:0] p7_array_index_1084002_comb;
  wire [7:0] p7_array_index_1084003_comb;
  wire [7:0] p7_array_index_1084004_comb;
  wire [7:0] p7_array_index_1084005_comb;
  wire [7:0] p7_array_index_1084006_comb;
  wire [7:0] p7_array_index_1084007_comb;
  wire [7:0] p7_array_index_1084009_comb;
  wire [7:0] p7_array_index_1084010_comb;
  wire [7:0] p7_array_index_1084011_comb;
  assign p7_addedKey__63_comb = p6_xor_1082915 ^ 128'he65a_edb1_c831_097f_c9c0_34b3_188d_3e17;
  assign p7_array_index_1082953_comb = p6_arr[p7_addedKey__63_comb[127:120]];
  assign p7_array_index_1082954_comb = p6_arr[p7_addedKey__63_comb[119:112]];
  assign p7_array_index_1082955_comb = p6_arr[p7_addedKey__63_comb[111:104]];
  assign p7_array_index_1082956_comb = p6_arr[p7_addedKey__63_comb[103:96]];
  assign p7_array_index_1082957_comb = p6_arr[p7_addedKey__63_comb[95:88]];
  assign p7_array_index_1082958_comb = p6_arr[p7_addedKey__63_comb[87:80]];
  assign p7_array_index_1082960_comb = p6_arr[p7_addedKey__63_comb[71:64]];
  assign p7_array_index_1082962_comb = p6_arr[p7_addedKey__63_comb[55:48]];
  assign p7_array_index_1082963_comb = p6_arr[p7_addedKey__63_comb[47:40]];
  assign p7_array_index_1082964_comb = p6_arr[p7_addedKey__63_comb[39:32]];
  assign p7_array_index_1082965_comb = p6_arr[p7_addedKey__63_comb[31:24]];
  assign p7_array_index_1082966_comb = p6_arr[p7_addedKey__63_comb[23:16]];
  assign p7_array_index_1082967_comb = p6_arr[p7_addedKey__63_comb[15:8]];
  assign p7_array_index_1082969_comb = p6_literal_1076345[p7_array_index_1082953_comb];
  assign p7_array_index_1082970_comb = p6_literal_1076347[p7_array_index_1082954_comb];
  assign p7_array_index_1082971_comb = p6_literal_1076349[p7_array_index_1082955_comb];
  assign p7_array_index_1082972_comb = p6_literal_1076351[p7_array_index_1082956_comb];
  assign p7_array_index_1082973_comb = p6_literal_1076353[p7_array_index_1082957_comb];
  assign p7_array_index_1082974_comb = p6_literal_1076355[p7_array_index_1082958_comb];
  assign p7_array_index_1082975_comb = p6_arr[p7_addedKey__63_comb[79:72]];
  assign p7_array_index_1082977_comb = p6_arr[p7_addedKey__63_comb[63:56]];
  assign p7_res7__352_comb = p7_array_index_1082969_comb ^ p7_array_index_1082970_comb ^ p7_array_index_1082971_comb ^ p7_array_index_1082972_comb ^ p7_array_index_1082973_comb ^ p7_array_index_1082974_comb ^ p7_array_index_1082975_comb ^ p6_literal_1076358[p7_array_index_1082960_comb] ^ p7_array_index_1082977_comb ^ p6_literal_1076355[p7_array_index_1082962_comb] ^ p6_literal_1076353[p7_array_index_1082963_comb] ^ p6_literal_1076351[p7_array_index_1082964_comb] ^ p6_literal_1076349[p7_array_index_1082965_comb] ^ p6_literal_1076347[p7_array_index_1082966_comb] ^ p6_literal_1076345[p7_array_index_1082967_comb] ^ p6_arr[p7_addedKey__63_comb[7:0]];
  assign p7_array_index_1082986_comb = p6_literal_1076345[p7_res7__352_comb];
  assign p7_array_index_1082987_comb = p6_literal_1076347[p7_array_index_1082953_comb];
  assign p7_array_index_1082988_comb = p6_literal_1076349[p7_array_index_1082954_comb];
  assign p7_array_index_1082989_comb = p6_literal_1076351[p7_array_index_1082955_comb];
  assign p7_array_index_1082990_comb = p6_literal_1076353[p7_array_index_1082956_comb];
  assign p7_array_index_1082991_comb = p6_literal_1076355[p7_array_index_1082957_comb];
  assign p7_res7__353_comb = p7_array_index_1082986_comb ^ p7_array_index_1082987_comb ^ p7_array_index_1082988_comb ^ p7_array_index_1082989_comb ^ p7_array_index_1082990_comb ^ p7_array_index_1082991_comb ^ p7_array_index_1082958_comb ^ p6_literal_1076358[p7_array_index_1082975_comb] ^ p7_array_index_1082960_comb ^ p6_literal_1076355[p7_array_index_1082977_comb] ^ p6_literal_1076353[p7_array_index_1082962_comb] ^ p6_literal_1076351[p7_array_index_1082963_comb] ^ p6_literal_1076349[p7_array_index_1082964_comb] ^ p6_literal_1076347[p7_array_index_1082965_comb] ^ p6_literal_1076345[p7_array_index_1082966_comb] ^ p7_array_index_1082967_comb;
  assign p7_array_index_1083001_comb = p6_literal_1076347[p7_res7__352_comb];
  assign p7_array_index_1083002_comb = p6_literal_1076349[p7_array_index_1082953_comb];
  assign p7_array_index_1083003_comb = p6_literal_1076351[p7_array_index_1082954_comb];
  assign p7_array_index_1083004_comb = p6_literal_1076353[p7_array_index_1082955_comb];
  assign p7_array_index_1083005_comb = p6_literal_1076355[p7_array_index_1082956_comb];
  assign p7_res7__354_comb = p6_literal_1076345[p7_res7__353_comb] ^ p7_array_index_1083001_comb ^ p7_array_index_1083002_comb ^ p7_array_index_1083003_comb ^ p7_array_index_1083004_comb ^ p7_array_index_1083005_comb ^ p7_array_index_1082957_comb ^ p6_literal_1076358[p7_array_index_1082958_comb] ^ p7_array_index_1082975_comb ^ p6_literal_1076355[p7_array_index_1082960_comb] ^ p6_literal_1076353[p7_array_index_1082977_comb] ^ p6_literal_1076351[p7_array_index_1082962_comb] ^ p6_literal_1076349[p7_array_index_1082963_comb] ^ p6_literal_1076347[p7_array_index_1082964_comb] ^ p6_literal_1076345[p7_array_index_1082965_comb] ^ p7_array_index_1082966_comb;
  assign p7_array_index_1083015_comb = p6_literal_1076347[p7_res7__353_comb];
  assign p7_array_index_1083016_comb = p6_literal_1076349[p7_res7__352_comb];
  assign p7_array_index_1083017_comb = p6_literal_1076351[p7_array_index_1082953_comb];
  assign p7_array_index_1083018_comb = p6_literal_1076353[p7_array_index_1082954_comb];
  assign p7_array_index_1083019_comb = p6_literal_1076355[p7_array_index_1082955_comb];
  assign p7_res7__355_comb = p6_literal_1076345[p7_res7__354_comb] ^ p7_array_index_1083015_comb ^ p7_array_index_1083016_comb ^ p7_array_index_1083017_comb ^ p7_array_index_1083018_comb ^ p7_array_index_1083019_comb ^ p7_array_index_1082956_comb ^ p6_literal_1076358[p7_array_index_1082957_comb] ^ p7_array_index_1082958_comb ^ p6_literal_1076355[p7_array_index_1082975_comb] ^ p6_literal_1076353[p7_array_index_1082960_comb] ^ p6_literal_1076351[p7_array_index_1082977_comb] ^ p6_literal_1076349[p7_array_index_1082962_comb] ^ p6_literal_1076347[p7_array_index_1082963_comb] ^ p6_literal_1076345[p7_array_index_1082964_comb] ^ p7_array_index_1082965_comb;
  assign p7_array_index_1083030_comb = p6_literal_1076349[p7_res7__353_comb];
  assign p7_array_index_1083031_comb = p6_literal_1076351[p7_res7__352_comb];
  assign p7_array_index_1083032_comb = p6_literal_1076353[p7_array_index_1082953_comb];
  assign p7_array_index_1083033_comb = p6_literal_1076355[p7_array_index_1082954_comb];
  assign p7_res7__356_comb = p6_literal_1076345[p7_res7__355_comb] ^ p6_literal_1076347[p7_res7__354_comb] ^ p7_array_index_1083030_comb ^ p7_array_index_1083031_comb ^ p7_array_index_1083032_comb ^ p7_array_index_1083033_comb ^ p7_array_index_1082955_comb ^ p6_literal_1076358[p7_array_index_1082956_comb] ^ p7_array_index_1082957_comb ^ p7_array_index_1082974_comb ^ p6_literal_1076353[p7_array_index_1082975_comb] ^ p6_literal_1076351[p7_array_index_1082960_comb] ^ p6_literal_1076349[p7_array_index_1082977_comb] ^ p6_literal_1076347[p7_array_index_1082962_comb] ^ p6_literal_1076345[p7_array_index_1082963_comb] ^ p7_array_index_1082964_comb;
  assign p7_array_index_1083043_comb = p6_literal_1076349[p7_res7__354_comb];
  assign p7_array_index_1083044_comb = p6_literal_1076351[p7_res7__353_comb];
  assign p7_array_index_1083045_comb = p6_literal_1076353[p7_res7__352_comb];
  assign p7_array_index_1083046_comb = p6_literal_1076355[p7_array_index_1082953_comb];
  assign p7_res7__357_comb = p6_literal_1076345[p7_res7__356_comb] ^ p6_literal_1076347[p7_res7__355_comb] ^ p7_array_index_1083043_comb ^ p7_array_index_1083044_comb ^ p7_array_index_1083045_comb ^ p7_array_index_1083046_comb ^ p7_array_index_1082954_comb ^ p6_literal_1076358[p7_array_index_1082955_comb] ^ p7_array_index_1082956_comb ^ p7_array_index_1082991_comb ^ p6_literal_1076353[p7_array_index_1082958_comb] ^ p6_literal_1076351[p7_array_index_1082975_comb] ^ p6_literal_1076349[p7_array_index_1082960_comb] ^ p6_literal_1076347[p7_array_index_1082977_comb] ^ p6_literal_1076345[p7_array_index_1082962_comb] ^ p7_array_index_1082963_comb;
  assign p7_array_index_1083057_comb = p6_literal_1076351[p7_res7__354_comb];
  assign p7_array_index_1083058_comb = p6_literal_1076353[p7_res7__353_comb];
  assign p7_array_index_1083059_comb = p6_literal_1076355[p7_res7__352_comb];
  assign p7_res7__358_comb = p6_literal_1076345[p7_res7__357_comb] ^ p6_literal_1076347[p7_res7__356_comb] ^ p6_literal_1076349[p7_res7__355_comb] ^ p7_array_index_1083057_comb ^ p7_array_index_1083058_comb ^ p7_array_index_1083059_comb ^ p7_array_index_1082953_comb ^ p6_literal_1076358[p7_array_index_1082954_comb] ^ p7_array_index_1082955_comb ^ p7_array_index_1083005_comb ^ p7_array_index_1082973_comb ^ p6_literal_1076351[p7_array_index_1082958_comb] ^ p6_literal_1076349[p7_array_index_1082975_comb] ^ p6_literal_1076347[p7_array_index_1082960_comb] ^ p6_literal_1076345[p7_array_index_1082977_comb] ^ p7_array_index_1082962_comb;
  assign p7_array_index_1083069_comb = p6_literal_1076351[p7_res7__355_comb];
  assign p7_array_index_1083070_comb = p6_literal_1076353[p7_res7__354_comb];
  assign p7_array_index_1083071_comb = p6_literal_1076355[p7_res7__353_comb];
  assign p7_res7__359_comb = p6_literal_1076345[p7_res7__358_comb] ^ p6_literal_1076347[p7_res7__357_comb] ^ p6_literal_1076349[p7_res7__356_comb] ^ p7_array_index_1083069_comb ^ p7_array_index_1083070_comb ^ p7_array_index_1083071_comb ^ p7_res7__352_comb ^ p6_literal_1076358[p7_array_index_1082953_comb] ^ p7_array_index_1082954_comb ^ p7_array_index_1083019_comb ^ p7_array_index_1082990_comb ^ p6_literal_1076351[p7_array_index_1082957_comb] ^ p6_literal_1076349[p7_array_index_1082958_comb] ^ p6_literal_1076347[p7_array_index_1082975_comb] ^ p6_literal_1076345[p7_array_index_1082960_comb] ^ p7_array_index_1082977_comb;
  assign p7_array_index_1083082_comb = p6_literal_1076353[p7_res7__355_comb];
  assign p7_array_index_1083083_comb = p6_literal_1076355[p7_res7__354_comb];
  assign p7_res7__360_comb = p6_literal_1076345[p7_res7__359_comb] ^ p6_literal_1076347[p7_res7__358_comb] ^ p6_literal_1076349[p7_res7__357_comb] ^ p6_literal_1076351[p7_res7__356_comb] ^ p7_array_index_1083082_comb ^ p7_array_index_1083083_comb ^ p7_res7__353_comb ^ p6_literal_1076358[p7_res7__352_comb] ^ p7_array_index_1082953_comb ^ p7_array_index_1083033_comb ^ p7_array_index_1083004_comb ^ p7_array_index_1082972_comb ^ p6_literal_1076349[p7_array_index_1082957_comb] ^ p6_literal_1076347[p7_array_index_1082958_comb] ^ p6_literal_1076345[p7_array_index_1082975_comb] ^ p7_array_index_1082960_comb;
  assign p7_array_index_1083093_comb = p6_literal_1076353[p7_res7__356_comb];
  assign p7_array_index_1083094_comb = p6_literal_1076355[p7_res7__355_comb];
  assign p7_res7__361_comb = p6_literal_1076345[p7_res7__360_comb] ^ p6_literal_1076347[p7_res7__359_comb] ^ p6_literal_1076349[p7_res7__358_comb] ^ p6_literal_1076351[p7_res7__357_comb] ^ p7_array_index_1083093_comb ^ p7_array_index_1083094_comb ^ p7_res7__354_comb ^ p6_literal_1076358[p7_res7__353_comb] ^ p7_res7__352_comb ^ p7_array_index_1083046_comb ^ p7_array_index_1083018_comb ^ p7_array_index_1082989_comb ^ p6_literal_1076349[p7_array_index_1082956_comb] ^ p6_literal_1076347[p7_array_index_1082957_comb] ^ p6_literal_1076345[p7_array_index_1082958_comb] ^ p7_array_index_1082975_comb;
  assign p7_array_index_1083105_comb = p6_literal_1076355[p7_res7__356_comb];
  assign p7_res7__362_comb = p6_literal_1076345[p7_res7__361_comb] ^ p6_literal_1076347[p7_res7__360_comb] ^ p6_literal_1076349[p7_res7__359_comb] ^ p6_literal_1076351[p7_res7__358_comb] ^ p6_literal_1076353[p7_res7__357_comb] ^ p7_array_index_1083105_comb ^ p7_res7__355_comb ^ p6_literal_1076358[p7_res7__354_comb] ^ p7_res7__353_comb ^ p7_array_index_1083059_comb ^ p7_array_index_1083032_comb ^ p7_array_index_1083003_comb ^ p7_array_index_1082971_comb ^ p6_literal_1076347[p7_array_index_1082956_comb] ^ p6_literal_1076345[p7_array_index_1082957_comb] ^ p7_array_index_1082958_comb;
  assign p7_array_index_1083115_comb = p6_literal_1076355[p7_res7__357_comb];
  assign p7_res7__363_comb = p6_literal_1076345[p7_res7__362_comb] ^ p6_literal_1076347[p7_res7__361_comb] ^ p6_literal_1076349[p7_res7__360_comb] ^ p6_literal_1076351[p7_res7__359_comb] ^ p6_literal_1076353[p7_res7__358_comb] ^ p7_array_index_1083115_comb ^ p7_res7__356_comb ^ p6_literal_1076358[p7_res7__355_comb] ^ p7_res7__354_comb ^ p7_array_index_1083071_comb ^ p7_array_index_1083045_comb ^ p7_array_index_1083017_comb ^ p7_array_index_1082988_comb ^ p6_literal_1076347[p7_array_index_1082955_comb] ^ p6_literal_1076345[p7_array_index_1082956_comb] ^ p7_array_index_1082957_comb;
  assign p7_res7__364_comb = p6_literal_1076345[p7_res7__363_comb] ^ p6_literal_1076347[p7_res7__362_comb] ^ p6_literal_1076349[p7_res7__361_comb] ^ p6_literal_1076351[p7_res7__360_comb] ^ p6_literal_1076353[p7_res7__359_comb] ^ p6_literal_1076355[p7_res7__358_comb] ^ p7_res7__357_comb ^ p6_literal_1076358[p7_res7__356_comb] ^ p7_res7__355_comb ^ p7_array_index_1083083_comb ^ p7_array_index_1083058_comb ^ p7_array_index_1083031_comb ^ p7_array_index_1083002_comb ^ p7_array_index_1082970_comb ^ p6_literal_1076345[p7_array_index_1082955_comb] ^ p7_array_index_1082956_comb;
  assign p7_res7__365_comb = p6_literal_1076345[p7_res7__364_comb] ^ p6_literal_1076347[p7_res7__363_comb] ^ p6_literal_1076349[p7_res7__362_comb] ^ p6_literal_1076351[p7_res7__361_comb] ^ p6_literal_1076353[p7_res7__360_comb] ^ p6_literal_1076355[p7_res7__359_comb] ^ p7_res7__358_comb ^ p6_literal_1076358[p7_res7__357_comb] ^ p7_res7__356_comb ^ p7_array_index_1083094_comb ^ p7_array_index_1083070_comb ^ p7_array_index_1083044_comb ^ p7_array_index_1083016_comb ^ p7_array_index_1082987_comb ^ p6_literal_1076345[p7_array_index_1082954_comb] ^ p7_array_index_1082955_comb;
  assign p7_res7__366_comb = p6_literal_1076345[p7_res7__365_comb] ^ p6_literal_1076347[p7_res7__364_comb] ^ p6_literal_1076349[p7_res7__363_comb] ^ p6_literal_1076351[p7_res7__362_comb] ^ p6_literal_1076353[p7_res7__361_comb] ^ p6_literal_1076355[p7_res7__360_comb] ^ p7_res7__359_comb ^ p6_literal_1076358[p7_res7__358_comb] ^ p7_res7__357_comb ^ p7_array_index_1083105_comb ^ p7_array_index_1083082_comb ^ p7_array_index_1083057_comb ^ p7_array_index_1083030_comb ^ p7_array_index_1083001_comb ^ p7_array_index_1082969_comb ^ p7_array_index_1082954_comb;
  assign p7_res7__367_comb = p6_literal_1076345[p7_res7__366_comb] ^ p6_literal_1076347[p7_res7__365_comb] ^ p6_literal_1076349[p7_res7__364_comb] ^ p6_literal_1076351[p7_res7__363_comb] ^ p6_literal_1076353[p7_res7__362_comb] ^ p6_literal_1076355[p7_res7__361_comb] ^ p7_res7__360_comb ^ p6_literal_1076358[p7_res7__359_comb] ^ p7_res7__358_comb ^ p7_array_index_1083115_comb ^ p7_array_index_1083093_comb ^ p7_array_index_1083069_comb ^ p7_array_index_1083043_comb ^ p7_array_index_1083015_comb ^ p7_array_index_1082986_comb ^ p7_array_index_1082953_comb;
  assign p7_res__22_comb = {p7_res7__367_comb, p7_res7__366_comb, p7_res7__365_comb, p7_res7__364_comb, p7_res7__363_comb, p7_res7__362_comb, p7_res7__361_comb, p7_res7__360_comb, p7_res7__359_comb, p7_res7__358_comb, p7_res7__357_comb, p7_res7__356_comb, p7_res7__355_comb, p7_res7__354_comb, p7_res7__353_comb, p7_res7__352_comb};
  assign p7_k7_comb = p7_res__22_comb ^ p6_xor_1082697;
  assign p7_addedKey__64_comb = p7_k7_comb ^ 128'hd9eb_5a3a_e90f_fa58_34ce_2043_693d_7e18;
  assign p7_array_index_1083171_comb = p6_arr[p7_addedKey__64_comb[127:120]];
  assign p7_array_index_1083172_comb = p6_arr[p7_addedKey__64_comb[119:112]];
  assign p7_array_index_1083173_comb = p6_arr[p7_addedKey__64_comb[111:104]];
  assign p7_array_index_1083174_comb = p6_arr[p7_addedKey__64_comb[103:96]];
  assign p7_array_index_1083175_comb = p6_arr[p7_addedKey__64_comb[95:88]];
  assign p7_array_index_1083176_comb = p6_arr[p7_addedKey__64_comb[87:80]];
  assign p7_array_index_1083178_comb = p6_arr[p7_addedKey__64_comb[71:64]];
  assign p7_array_index_1083180_comb = p6_arr[p7_addedKey__64_comb[55:48]];
  assign p7_array_index_1083181_comb = p6_arr[p7_addedKey__64_comb[47:40]];
  assign p7_array_index_1083182_comb = p6_arr[p7_addedKey__64_comb[39:32]];
  assign p7_array_index_1083183_comb = p6_arr[p7_addedKey__64_comb[31:24]];
  assign p7_array_index_1083184_comb = p6_arr[p7_addedKey__64_comb[23:16]];
  assign p7_array_index_1083185_comb = p6_arr[p7_addedKey__64_comb[15:8]];
  assign p7_array_index_1083187_comb = p6_literal_1076345[p7_array_index_1083171_comb];
  assign p7_array_index_1083188_comb = p6_literal_1076347[p7_array_index_1083172_comb];
  assign p7_array_index_1083189_comb = p6_literal_1076349[p7_array_index_1083173_comb];
  assign p7_array_index_1083190_comb = p6_literal_1076351[p7_array_index_1083174_comb];
  assign p7_array_index_1083191_comb = p6_literal_1076353[p7_array_index_1083175_comb];
  assign p7_array_index_1083192_comb = p6_literal_1076355[p7_array_index_1083176_comb];
  assign p7_array_index_1083193_comb = p6_arr[p7_addedKey__64_comb[79:72]];
  assign p7_array_index_1083195_comb = p6_arr[p7_addedKey__64_comb[63:56]];
  assign p7_res7__368_comb = p7_array_index_1083187_comb ^ p7_array_index_1083188_comb ^ p7_array_index_1083189_comb ^ p7_array_index_1083190_comb ^ p7_array_index_1083191_comb ^ p7_array_index_1083192_comb ^ p7_array_index_1083193_comb ^ p6_literal_1076358[p7_array_index_1083178_comb] ^ p7_array_index_1083195_comb ^ p6_literal_1076355[p7_array_index_1083180_comb] ^ p6_literal_1076353[p7_array_index_1083181_comb] ^ p6_literal_1076351[p7_array_index_1083182_comb] ^ p6_literal_1076349[p7_array_index_1083183_comb] ^ p6_literal_1076347[p7_array_index_1083184_comb] ^ p6_literal_1076345[p7_array_index_1083185_comb] ^ p6_arr[p7_addedKey__64_comb[7:0]];
  assign p7_array_index_1083204_comb = p6_literal_1076345[p7_res7__368_comb];
  assign p7_array_index_1083205_comb = p6_literal_1076347[p7_array_index_1083171_comb];
  assign p7_array_index_1083206_comb = p6_literal_1076349[p7_array_index_1083172_comb];
  assign p7_array_index_1083207_comb = p6_literal_1076351[p7_array_index_1083173_comb];
  assign p7_array_index_1083208_comb = p6_literal_1076353[p7_array_index_1083174_comb];
  assign p7_array_index_1083209_comb = p6_literal_1076355[p7_array_index_1083175_comb];
  assign p7_res7__369_comb = p7_array_index_1083204_comb ^ p7_array_index_1083205_comb ^ p7_array_index_1083206_comb ^ p7_array_index_1083207_comb ^ p7_array_index_1083208_comb ^ p7_array_index_1083209_comb ^ p7_array_index_1083176_comb ^ p6_literal_1076358[p7_array_index_1083193_comb] ^ p7_array_index_1083178_comb ^ p6_literal_1076355[p7_array_index_1083195_comb] ^ p6_literal_1076353[p7_array_index_1083180_comb] ^ p6_literal_1076351[p7_array_index_1083181_comb] ^ p6_literal_1076349[p7_array_index_1083182_comb] ^ p6_literal_1076347[p7_array_index_1083183_comb] ^ p6_literal_1076345[p7_array_index_1083184_comb] ^ p7_array_index_1083185_comb;
  assign p7_array_index_1083219_comb = p6_literal_1076347[p7_res7__368_comb];
  assign p7_array_index_1083220_comb = p6_literal_1076349[p7_array_index_1083171_comb];
  assign p7_array_index_1083221_comb = p6_literal_1076351[p7_array_index_1083172_comb];
  assign p7_array_index_1083222_comb = p6_literal_1076353[p7_array_index_1083173_comb];
  assign p7_array_index_1083223_comb = p6_literal_1076355[p7_array_index_1083174_comb];
  assign p7_res7__370_comb = p6_literal_1076345[p7_res7__369_comb] ^ p7_array_index_1083219_comb ^ p7_array_index_1083220_comb ^ p7_array_index_1083221_comb ^ p7_array_index_1083222_comb ^ p7_array_index_1083223_comb ^ p7_array_index_1083175_comb ^ p6_literal_1076358[p7_array_index_1083176_comb] ^ p7_array_index_1083193_comb ^ p6_literal_1076355[p7_array_index_1083178_comb] ^ p6_literal_1076353[p7_array_index_1083195_comb] ^ p6_literal_1076351[p7_array_index_1083180_comb] ^ p6_literal_1076349[p7_array_index_1083181_comb] ^ p6_literal_1076347[p7_array_index_1083182_comb] ^ p6_literal_1076345[p7_array_index_1083183_comb] ^ p7_array_index_1083184_comb;
  assign p7_array_index_1083233_comb = p6_literal_1076347[p7_res7__369_comb];
  assign p7_array_index_1083234_comb = p6_literal_1076349[p7_res7__368_comb];
  assign p7_array_index_1083235_comb = p6_literal_1076351[p7_array_index_1083171_comb];
  assign p7_array_index_1083236_comb = p6_literal_1076353[p7_array_index_1083172_comb];
  assign p7_array_index_1083237_comb = p6_literal_1076355[p7_array_index_1083173_comb];
  assign p7_res7__371_comb = p6_literal_1076345[p7_res7__370_comb] ^ p7_array_index_1083233_comb ^ p7_array_index_1083234_comb ^ p7_array_index_1083235_comb ^ p7_array_index_1083236_comb ^ p7_array_index_1083237_comb ^ p7_array_index_1083174_comb ^ p6_literal_1076358[p7_array_index_1083175_comb] ^ p7_array_index_1083176_comb ^ p6_literal_1076355[p7_array_index_1083193_comb] ^ p6_literal_1076353[p7_array_index_1083178_comb] ^ p6_literal_1076351[p7_array_index_1083195_comb] ^ p6_literal_1076349[p7_array_index_1083180_comb] ^ p6_literal_1076347[p7_array_index_1083181_comb] ^ p6_literal_1076345[p7_array_index_1083182_comb] ^ p7_array_index_1083183_comb;
  assign p7_array_index_1083248_comb = p6_literal_1076349[p7_res7__369_comb];
  assign p7_array_index_1083249_comb = p6_literal_1076351[p7_res7__368_comb];
  assign p7_array_index_1083250_comb = p6_literal_1076353[p7_array_index_1083171_comb];
  assign p7_array_index_1083251_comb = p6_literal_1076355[p7_array_index_1083172_comb];
  assign p7_res7__372_comb = p6_literal_1076345[p7_res7__371_comb] ^ p6_literal_1076347[p7_res7__370_comb] ^ p7_array_index_1083248_comb ^ p7_array_index_1083249_comb ^ p7_array_index_1083250_comb ^ p7_array_index_1083251_comb ^ p7_array_index_1083173_comb ^ p6_literal_1076358[p7_array_index_1083174_comb] ^ p7_array_index_1083175_comb ^ p7_array_index_1083192_comb ^ p6_literal_1076353[p7_array_index_1083193_comb] ^ p6_literal_1076351[p7_array_index_1083178_comb] ^ p6_literal_1076349[p7_array_index_1083195_comb] ^ p6_literal_1076347[p7_array_index_1083180_comb] ^ p6_literal_1076345[p7_array_index_1083181_comb] ^ p7_array_index_1083182_comb;
  assign p7_array_index_1083261_comb = p6_literal_1076349[p7_res7__370_comb];
  assign p7_array_index_1083262_comb = p6_literal_1076351[p7_res7__369_comb];
  assign p7_array_index_1083263_comb = p6_literal_1076353[p7_res7__368_comb];
  assign p7_array_index_1083264_comb = p6_literal_1076355[p7_array_index_1083171_comb];
  assign p7_res7__373_comb = p6_literal_1076345[p7_res7__372_comb] ^ p6_literal_1076347[p7_res7__371_comb] ^ p7_array_index_1083261_comb ^ p7_array_index_1083262_comb ^ p7_array_index_1083263_comb ^ p7_array_index_1083264_comb ^ p7_array_index_1083172_comb ^ p6_literal_1076358[p7_array_index_1083173_comb] ^ p7_array_index_1083174_comb ^ p7_array_index_1083209_comb ^ p6_literal_1076353[p7_array_index_1083176_comb] ^ p6_literal_1076351[p7_array_index_1083193_comb] ^ p6_literal_1076349[p7_array_index_1083178_comb] ^ p6_literal_1076347[p7_array_index_1083195_comb] ^ p6_literal_1076345[p7_array_index_1083180_comb] ^ p7_array_index_1083181_comb;
  assign p7_array_index_1083275_comb = p6_literal_1076351[p7_res7__370_comb];
  assign p7_array_index_1083276_comb = p6_literal_1076353[p7_res7__369_comb];
  assign p7_array_index_1083277_comb = p6_literal_1076355[p7_res7__368_comb];
  assign p7_res7__374_comb = p6_literal_1076345[p7_res7__373_comb] ^ p6_literal_1076347[p7_res7__372_comb] ^ p6_literal_1076349[p7_res7__371_comb] ^ p7_array_index_1083275_comb ^ p7_array_index_1083276_comb ^ p7_array_index_1083277_comb ^ p7_array_index_1083171_comb ^ p6_literal_1076358[p7_array_index_1083172_comb] ^ p7_array_index_1083173_comb ^ p7_array_index_1083223_comb ^ p7_array_index_1083191_comb ^ p6_literal_1076351[p7_array_index_1083176_comb] ^ p6_literal_1076349[p7_array_index_1083193_comb] ^ p6_literal_1076347[p7_array_index_1083178_comb] ^ p6_literal_1076345[p7_array_index_1083195_comb] ^ p7_array_index_1083180_comb;
  assign p7_array_index_1083287_comb = p6_literal_1076351[p7_res7__371_comb];
  assign p7_array_index_1083288_comb = p6_literal_1076353[p7_res7__370_comb];
  assign p7_array_index_1083289_comb = p6_literal_1076355[p7_res7__369_comb];
  assign p7_res7__375_comb = p6_literal_1076345[p7_res7__374_comb] ^ p6_literal_1076347[p7_res7__373_comb] ^ p6_literal_1076349[p7_res7__372_comb] ^ p7_array_index_1083287_comb ^ p7_array_index_1083288_comb ^ p7_array_index_1083289_comb ^ p7_res7__368_comb ^ p6_literal_1076358[p7_array_index_1083171_comb] ^ p7_array_index_1083172_comb ^ p7_array_index_1083237_comb ^ p7_array_index_1083208_comb ^ p6_literal_1076351[p7_array_index_1083175_comb] ^ p6_literal_1076349[p7_array_index_1083176_comb] ^ p6_literal_1076347[p7_array_index_1083193_comb] ^ p6_literal_1076345[p7_array_index_1083178_comb] ^ p7_array_index_1083195_comb;
  assign p7_array_index_1083300_comb = p6_literal_1076353[p7_res7__371_comb];
  assign p7_array_index_1083301_comb = p6_literal_1076355[p7_res7__370_comb];
  assign p7_res7__376_comb = p6_literal_1076345[p7_res7__375_comb] ^ p6_literal_1076347[p7_res7__374_comb] ^ p6_literal_1076349[p7_res7__373_comb] ^ p6_literal_1076351[p7_res7__372_comb] ^ p7_array_index_1083300_comb ^ p7_array_index_1083301_comb ^ p7_res7__369_comb ^ p6_literal_1076358[p7_res7__368_comb] ^ p7_array_index_1083171_comb ^ p7_array_index_1083251_comb ^ p7_array_index_1083222_comb ^ p7_array_index_1083190_comb ^ p6_literal_1076349[p7_array_index_1083175_comb] ^ p6_literal_1076347[p7_array_index_1083176_comb] ^ p6_literal_1076345[p7_array_index_1083193_comb] ^ p7_array_index_1083178_comb;
  assign p7_array_index_1083311_comb = p6_literal_1076353[p7_res7__372_comb];
  assign p7_array_index_1083312_comb = p6_literal_1076355[p7_res7__371_comb];
  assign p7_res7__377_comb = p6_literal_1076345[p7_res7__376_comb] ^ p6_literal_1076347[p7_res7__375_comb] ^ p6_literal_1076349[p7_res7__374_comb] ^ p6_literal_1076351[p7_res7__373_comb] ^ p7_array_index_1083311_comb ^ p7_array_index_1083312_comb ^ p7_res7__370_comb ^ p6_literal_1076358[p7_res7__369_comb] ^ p7_res7__368_comb ^ p7_array_index_1083264_comb ^ p7_array_index_1083236_comb ^ p7_array_index_1083207_comb ^ p6_literal_1076349[p7_array_index_1083174_comb] ^ p6_literal_1076347[p7_array_index_1083175_comb] ^ p6_literal_1076345[p7_array_index_1083176_comb] ^ p7_array_index_1083193_comb;
  assign p7_array_index_1083323_comb = p6_literal_1076355[p7_res7__372_comb];
  assign p7_res7__378_comb = p6_literal_1076345[p7_res7__377_comb] ^ p6_literal_1076347[p7_res7__376_comb] ^ p6_literal_1076349[p7_res7__375_comb] ^ p6_literal_1076351[p7_res7__374_comb] ^ p6_literal_1076353[p7_res7__373_comb] ^ p7_array_index_1083323_comb ^ p7_res7__371_comb ^ p6_literal_1076358[p7_res7__370_comb] ^ p7_res7__369_comb ^ p7_array_index_1083277_comb ^ p7_array_index_1083250_comb ^ p7_array_index_1083221_comb ^ p7_array_index_1083189_comb ^ p6_literal_1076347[p7_array_index_1083174_comb] ^ p6_literal_1076345[p7_array_index_1083175_comb] ^ p7_array_index_1083176_comb;
  assign p7_array_index_1083333_comb = p6_literal_1076355[p7_res7__373_comb];
  assign p7_res7__379_comb = p6_literal_1076345[p7_res7__378_comb] ^ p6_literal_1076347[p7_res7__377_comb] ^ p6_literal_1076349[p7_res7__376_comb] ^ p6_literal_1076351[p7_res7__375_comb] ^ p6_literal_1076353[p7_res7__374_comb] ^ p7_array_index_1083333_comb ^ p7_res7__372_comb ^ p6_literal_1076358[p7_res7__371_comb] ^ p7_res7__370_comb ^ p7_array_index_1083289_comb ^ p7_array_index_1083263_comb ^ p7_array_index_1083235_comb ^ p7_array_index_1083206_comb ^ p6_literal_1076347[p7_array_index_1083173_comb] ^ p6_literal_1076345[p7_array_index_1083174_comb] ^ p7_array_index_1083175_comb;
  assign p7_res7__380_comb = p6_literal_1076345[p7_res7__379_comb] ^ p6_literal_1076347[p7_res7__378_comb] ^ p6_literal_1076349[p7_res7__377_comb] ^ p6_literal_1076351[p7_res7__376_comb] ^ p6_literal_1076353[p7_res7__375_comb] ^ p6_literal_1076355[p7_res7__374_comb] ^ p7_res7__373_comb ^ p6_literal_1076358[p7_res7__372_comb] ^ p7_res7__371_comb ^ p7_array_index_1083301_comb ^ p7_array_index_1083276_comb ^ p7_array_index_1083249_comb ^ p7_array_index_1083220_comb ^ p7_array_index_1083188_comb ^ p6_literal_1076345[p7_array_index_1083173_comb] ^ p7_array_index_1083174_comb;
  assign p7_res7__381_comb = p6_literal_1076345[p7_res7__380_comb] ^ p6_literal_1076347[p7_res7__379_comb] ^ p6_literal_1076349[p7_res7__378_comb] ^ p6_literal_1076351[p7_res7__377_comb] ^ p6_literal_1076353[p7_res7__376_comb] ^ p6_literal_1076355[p7_res7__375_comb] ^ p7_res7__374_comb ^ p6_literal_1076358[p7_res7__373_comb] ^ p7_res7__372_comb ^ p7_array_index_1083312_comb ^ p7_array_index_1083288_comb ^ p7_array_index_1083262_comb ^ p7_array_index_1083234_comb ^ p7_array_index_1083205_comb ^ p6_literal_1076345[p7_array_index_1083172_comb] ^ p7_array_index_1083173_comb;
  assign p7_res7__382_comb = p6_literal_1076345[p7_res7__381_comb] ^ p6_literal_1076347[p7_res7__380_comb] ^ p6_literal_1076349[p7_res7__379_comb] ^ p6_literal_1076351[p7_res7__378_comb] ^ p6_literal_1076353[p7_res7__377_comb] ^ p6_literal_1076355[p7_res7__376_comb] ^ p7_res7__375_comb ^ p6_literal_1076358[p7_res7__374_comb] ^ p7_res7__373_comb ^ p7_array_index_1083323_comb ^ p7_array_index_1083300_comb ^ p7_array_index_1083275_comb ^ p7_array_index_1083248_comb ^ p7_array_index_1083219_comb ^ p7_array_index_1083187_comb ^ p7_array_index_1083172_comb;
  assign p7_res7__383_comb = p6_literal_1076345[p7_res7__382_comb] ^ p6_literal_1076347[p7_res7__381_comb] ^ p6_literal_1076349[p7_res7__380_comb] ^ p6_literal_1076351[p7_res7__379_comb] ^ p6_literal_1076353[p7_res7__378_comb] ^ p6_literal_1076355[p7_res7__377_comb] ^ p7_res7__376_comb ^ p6_literal_1076358[p7_res7__375_comb] ^ p7_res7__374_comb ^ p7_array_index_1083333_comb ^ p7_array_index_1083311_comb ^ p7_array_index_1083287_comb ^ p7_array_index_1083261_comb ^ p7_array_index_1083233_comb ^ p7_array_index_1083204_comb ^ p7_array_index_1083171_comb;
  assign p7_res__23_comb = {p7_res7__383_comb, p7_res7__382_comb, p7_res7__381_comb, p7_res7__380_comb, p7_res7__379_comb, p7_res7__378_comb, p7_res7__377_comb, p7_res7__376_comb, p7_res7__375_comb, p7_res7__374_comb, p7_res7__373_comb, p7_res7__372_comb, p7_res7__371_comb, p7_res7__370_comb, p7_res7__369_comb, p7_res7__368_comb};
  assign p7_k6_comb = p7_res__23_comb ^ p6_xor_1082915;
  assign p7_addedKey__65_comb = p7_k6_comb ^ 128'hb749_2c48_8547_80e0_69e9_9d53_b4b9_ea19;
  assign p7_array_index_1083389_comb = p6_arr[p7_addedKey__65_comb[127:120]];
  assign p7_array_index_1083390_comb = p6_arr[p7_addedKey__65_comb[119:112]];
  assign p7_array_index_1083391_comb = p6_arr[p7_addedKey__65_comb[111:104]];
  assign p7_array_index_1083392_comb = p6_arr[p7_addedKey__65_comb[103:96]];
  assign p7_array_index_1083393_comb = p6_arr[p7_addedKey__65_comb[95:88]];
  assign p7_array_index_1083394_comb = p6_arr[p7_addedKey__65_comb[87:80]];
  assign p7_array_index_1083396_comb = p6_arr[p7_addedKey__65_comb[71:64]];
  assign p7_array_index_1083398_comb = p6_arr[p7_addedKey__65_comb[55:48]];
  assign p7_array_index_1083399_comb = p6_arr[p7_addedKey__65_comb[47:40]];
  assign p7_array_index_1083400_comb = p6_arr[p7_addedKey__65_comb[39:32]];
  assign p7_array_index_1083401_comb = p6_arr[p7_addedKey__65_comb[31:24]];
  assign p7_array_index_1083402_comb = p6_arr[p7_addedKey__65_comb[23:16]];
  assign p7_array_index_1083403_comb = p6_arr[p7_addedKey__65_comb[15:8]];
  assign p7_array_index_1083405_comb = p6_literal_1076345[p7_array_index_1083389_comb];
  assign p7_array_index_1083406_comb = p6_literal_1076347[p7_array_index_1083390_comb];
  assign p7_array_index_1083407_comb = p6_literal_1076349[p7_array_index_1083391_comb];
  assign p7_array_index_1083408_comb = p6_literal_1076351[p7_array_index_1083392_comb];
  assign p7_array_index_1083409_comb = p6_literal_1076353[p7_array_index_1083393_comb];
  assign p7_array_index_1083410_comb = p6_literal_1076355[p7_array_index_1083394_comb];
  assign p7_array_index_1083411_comb = p6_arr[p7_addedKey__65_comb[79:72]];
  assign p7_array_index_1083413_comb = p6_arr[p7_addedKey__65_comb[63:56]];
  assign p7_res7__384_comb = p7_array_index_1083405_comb ^ p7_array_index_1083406_comb ^ p7_array_index_1083407_comb ^ p7_array_index_1083408_comb ^ p7_array_index_1083409_comb ^ p7_array_index_1083410_comb ^ p7_array_index_1083411_comb ^ p6_literal_1076358[p7_array_index_1083396_comb] ^ p7_array_index_1083413_comb ^ p6_literal_1076355[p7_array_index_1083398_comb] ^ p6_literal_1076353[p7_array_index_1083399_comb] ^ p6_literal_1076351[p7_array_index_1083400_comb] ^ p6_literal_1076349[p7_array_index_1083401_comb] ^ p6_literal_1076347[p7_array_index_1083402_comb] ^ p6_literal_1076345[p7_array_index_1083403_comb] ^ p6_arr[p7_addedKey__65_comb[7:0]];
  assign p7_array_index_1083422_comb = p6_literal_1076345[p7_res7__384_comb];
  assign p7_array_index_1083423_comb = p6_literal_1076347[p7_array_index_1083389_comb];
  assign p7_array_index_1083424_comb = p6_literal_1076349[p7_array_index_1083390_comb];
  assign p7_array_index_1083425_comb = p6_literal_1076351[p7_array_index_1083391_comb];
  assign p7_array_index_1083426_comb = p6_literal_1076353[p7_array_index_1083392_comb];
  assign p7_array_index_1083427_comb = p6_literal_1076355[p7_array_index_1083393_comb];
  assign p7_res7__385_comb = p7_array_index_1083422_comb ^ p7_array_index_1083423_comb ^ p7_array_index_1083424_comb ^ p7_array_index_1083425_comb ^ p7_array_index_1083426_comb ^ p7_array_index_1083427_comb ^ p7_array_index_1083394_comb ^ p6_literal_1076358[p7_array_index_1083411_comb] ^ p7_array_index_1083396_comb ^ p6_literal_1076355[p7_array_index_1083413_comb] ^ p6_literal_1076353[p7_array_index_1083398_comb] ^ p6_literal_1076351[p7_array_index_1083399_comb] ^ p6_literal_1076349[p7_array_index_1083400_comb] ^ p6_literal_1076347[p7_array_index_1083401_comb] ^ p6_literal_1076345[p7_array_index_1083402_comb] ^ p7_array_index_1083403_comb;
  assign p7_array_index_1083437_comb = p6_literal_1076347[p7_res7__384_comb];
  assign p7_array_index_1083438_comb = p6_literal_1076349[p7_array_index_1083389_comb];
  assign p7_array_index_1083439_comb = p6_literal_1076351[p7_array_index_1083390_comb];
  assign p7_array_index_1083440_comb = p6_literal_1076353[p7_array_index_1083391_comb];
  assign p7_array_index_1083441_comb = p6_literal_1076355[p7_array_index_1083392_comb];
  assign p7_res7__386_comb = p6_literal_1076345[p7_res7__385_comb] ^ p7_array_index_1083437_comb ^ p7_array_index_1083438_comb ^ p7_array_index_1083439_comb ^ p7_array_index_1083440_comb ^ p7_array_index_1083441_comb ^ p7_array_index_1083393_comb ^ p6_literal_1076358[p7_array_index_1083394_comb] ^ p7_array_index_1083411_comb ^ p6_literal_1076355[p7_array_index_1083396_comb] ^ p6_literal_1076353[p7_array_index_1083413_comb] ^ p6_literal_1076351[p7_array_index_1083398_comb] ^ p6_literal_1076349[p7_array_index_1083399_comb] ^ p6_literal_1076347[p7_array_index_1083400_comb] ^ p6_literal_1076345[p7_array_index_1083401_comb] ^ p7_array_index_1083402_comb;
  assign p7_array_index_1083451_comb = p6_literal_1076347[p7_res7__385_comb];
  assign p7_array_index_1083452_comb = p6_literal_1076349[p7_res7__384_comb];
  assign p7_array_index_1083453_comb = p6_literal_1076351[p7_array_index_1083389_comb];
  assign p7_array_index_1083454_comb = p6_literal_1076353[p7_array_index_1083390_comb];
  assign p7_array_index_1083455_comb = p6_literal_1076355[p7_array_index_1083391_comb];
  assign p7_res7__387_comb = p6_literal_1076345[p7_res7__386_comb] ^ p7_array_index_1083451_comb ^ p7_array_index_1083452_comb ^ p7_array_index_1083453_comb ^ p7_array_index_1083454_comb ^ p7_array_index_1083455_comb ^ p7_array_index_1083392_comb ^ p6_literal_1076358[p7_array_index_1083393_comb] ^ p7_array_index_1083394_comb ^ p6_literal_1076355[p7_array_index_1083411_comb] ^ p6_literal_1076353[p7_array_index_1083396_comb] ^ p6_literal_1076351[p7_array_index_1083413_comb] ^ p6_literal_1076349[p7_array_index_1083398_comb] ^ p6_literal_1076347[p7_array_index_1083399_comb] ^ p6_literal_1076345[p7_array_index_1083400_comb] ^ p7_array_index_1083401_comb;
  assign p7_array_index_1083466_comb = p6_literal_1076349[p7_res7__385_comb];
  assign p7_array_index_1083467_comb = p6_literal_1076351[p7_res7__384_comb];
  assign p7_array_index_1083468_comb = p6_literal_1076353[p7_array_index_1083389_comb];
  assign p7_array_index_1083469_comb = p6_literal_1076355[p7_array_index_1083390_comb];
  assign p7_res7__388_comb = p6_literal_1076345[p7_res7__387_comb] ^ p6_literal_1076347[p7_res7__386_comb] ^ p7_array_index_1083466_comb ^ p7_array_index_1083467_comb ^ p7_array_index_1083468_comb ^ p7_array_index_1083469_comb ^ p7_array_index_1083391_comb ^ p6_literal_1076358[p7_array_index_1083392_comb] ^ p7_array_index_1083393_comb ^ p7_array_index_1083410_comb ^ p6_literal_1076353[p7_array_index_1083411_comb] ^ p6_literal_1076351[p7_array_index_1083396_comb] ^ p6_literal_1076349[p7_array_index_1083413_comb] ^ p6_literal_1076347[p7_array_index_1083398_comb] ^ p6_literal_1076345[p7_array_index_1083399_comb] ^ p7_array_index_1083400_comb;
  assign p7_array_index_1083479_comb = p6_literal_1076349[p7_res7__386_comb];
  assign p7_array_index_1083480_comb = p6_literal_1076351[p7_res7__385_comb];
  assign p7_array_index_1083481_comb = p6_literal_1076353[p7_res7__384_comb];
  assign p7_array_index_1083482_comb = p6_literal_1076355[p7_array_index_1083389_comb];
  assign p7_res7__389_comb = p6_literal_1076345[p7_res7__388_comb] ^ p6_literal_1076347[p7_res7__387_comb] ^ p7_array_index_1083479_comb ^ p7_array_index_1083480_comb ^ p7_array_index_1083481_comb ^ p7_array_index_1083482_comb ^ p7_array_index_1083390_comb ^ p6_literal_1076358[p7_array_index_1083391_comb] ^ p7_array_index_1083392_comb ^ p7_array_index_1083427_comb ^ p6_literal_1076353[p7_array_index_1083394_comb] ^ p6_literal_1076351[p7_array_index_1083411_comb] ^ p6_literal_1076349[p7_array_index_1083396_comb] ^ p6_literal_1076347[p7_array_index_1083413_comb] ^ p6_literal_1076345[p7_array_index_1083398_comb] ^ p7_array_index_1083399_comb;
  assign p7_array_index_1083493_comb = p6_literal_1076351[p7_res7__386_comb];
  assign p7_array_index_1083494_comb = p6_literal_1076353[p7_res7__385_comb];
  assign p7_array_index_1083495_comb = p6_literal_1076355[p7_res7__384_comb];
  assign p7_res7__390_comb = p6_literal_1076345[p7_res7__389_comb] ^ p6_literal_1076347[p7_res7__388_comb] ^ p6_literal_1076349[p7_res7__387_comb] ^ p7_array_index_1083493_comb ^ p7_array_index_1083494_comb ^ p7_array_index_1083495_comb ^ p7_array_index_1083389_comb ^ p6_literal_1076358[p7_array_index_1083390_comb] ^ p7_array_index_1083391_comb ^ p7_array_index_1083441_comb ^ p7_array_index_1083409_comb ^ p6_literal_1076351[p7_array_index_1083394_comb] ^ p6_literal_1076349[p7_array_index_1083411_comb] ^ p6_literal_1076347[p7_array_index_1083396_comb] ^ p6_literal_1076345[p7_array_index_1083413_comb] ^ p7_array_index_1083398_comb;
  assign p7_array_index_1083505_comb = p6_literal_1076351[p7_res7__387_comb];
  assign p7_array_index_1083506_comb = p6_literal_1076353[p7_res7__386_comb];
  assign p7_array_index_1083507_comb = p6_literal_1076355[p7_res7__385_comb];
  assign p7_res7__391_comb = p6_literal_1076345[p7_res7__390_comb] ^ p6_literal_1076347[p7_res7__389_comb] ^ p6_literal_1076349[p7_res7__388_comb] ^ p7_array_index_1083505_comb ^ p7_array_index_1083506_comb ^ p7_array_index_1083507_comb ^ p7_res7__384_comb ^ p6_literal_1076358[p7_array_index_1083389_comb] ^ p7_array_index_1083390_comb ^ p7_array_index_1083455_comb ^ p7_array_index_1083426_comb ^ p6_literal_1076351[p7_array_index_1083393_comb] ^ p6_literal_1076349[p7_array_index_1083394_comb] ^ p6_literal_1076347[p7_array_index_1083411_comb] ^ p6_literal_1076345[p7_array_index_1083396_comb] ^ p7_array_index_1083413_comb;
  assign p7_array_index_1083518_comb = p6_literal_1076353[p7_res7__387_comb];
  assign p7_array_index_1083519_comb = p6_literal_1076355[p7_res7__386_comb];
  assign p7_res7__392_comb = p6_literal_1076345[p7_res7__391_comb] ^ p6_literal_1076347[p7_res7__390_comb] ^ p6_literal_1076349[p7_res7__389_comb] ^ p6_literal_1076351[p7_res7__388_comb] ^ p7_array_index_1083518_comb ^ p7_array_index_1083519_comb ^ p7_res7__385_comb ^ p6_literal_1076358[p7_res7__384_comb] ^ p7_array_index_1083389_comb ^ p7_array_index_1083469_comb ^ p7_array_index_1083440_comb ^ p7_array_index_1083408_comb ^ p6_literal_1076349[p7_array_index_1083393_comb] ^ p6_literal_1076347[p7_array_index_1083394_comb] ^ p6_literal_1076345[p7_array_index_1083411_comb] ^ p7_array_index_1083396_comb;
  assign p7_array_index_1083529_comb = p6_literal_1076353[p7_res7__388_comb];
  assign p7_array_index_1083530_comb = p6_literal_1076355[p7_res7__387_comb];
  assign p7_res7__393_comb = p6_literal_1076345[p7_res7__392_comb] ^ p6_literal_1076347[p7_res7__391_comb] ^ p6_literal_1076349[p7_res7__390_comb] ^ p6_literal_1076351[p7_res7__389_comb] ^ p7_array_index_1083529_comb ^ p7_array_index_1083530_comb ^ p7_res7__386_comb ^ p6_literal_1076358[p7_res7__385_comb] ^ p7_res7__384_comb ^ p7_array_index_1083482_comb ^ p7_array_index_1083454_comb ^ p7_array_index_1083425_comb ^ p6_literal_1076349[p7_array_index_1083392_comb] ^ p6_literal_1076347[p7_array_index_1083393_comb] ^ p6_literal_1076345[p7_array_index_1083394_comb] ^ p7_array_index_1083411_comb;
  assign p7_addedKey__38_comb = p7_k6_comb ^ p6_res__37;
  assign p7_array_index_1083541_comb = p6_literal_1076355[p7_res7__388_comb];
  assign p7_res7__394_comb = p6_literal_1076345[p7_res7__393_comb] ^ p6_literal_1076347[p7_res7__392_comb] ^ p6_literal_1076349[p7_res7__391_comb] ^ p6_literal_1076351[p7_res7__390_comb] ^ p6_literal_1076353[p7_res7__389_comb] ^ p7_array_index_1083541_comb ^ p7_res7__387_comb ^ p6_literal_1076358[p7_res7__386_comb] ^ p7_res7__385_comb ^ p7_array_index_1083495_comb ^ p7_array_index_1083468_comb ^ p7_array_index_1083439_comb ^ p7_array_index_1083407_comb ^ p6_literal_1076347[p7_array_index_1083392_comb] ^ p6_literal_1076345[p7_array_index_1083393_comb] ^ p7_array_index_1083394_comb;
  assign p7_array_index_1083777_comb = p6_arr[p7_addedKey__38_comb[127:120]];
  assign p7_array_index_1083778_comb = p6_arr[p7_addedKey__38_comb[119:112]];
  assign p7_array_index_1083779_comb = p6_arr[p7_addedKey__38_comb[111:104]];
  assign p7_array_index_1083780_comb = p6_arr[p7_addedKey__38_comb[103:96]];
  assign p7_array_index_1083781_comb = p6_arr[p7_addedKey__38_comb[95:88]];
  assign p7_array_index_1083782_comb = p6_arr[p7_addedKey__38_comb[87:80]];
  assign p7_array_index_1083784_comb = p6_arr[p7_addedKey__38_comb[71:64]];
  assign p7_array_index_1083786_comb = p6_arr[p7_addedKey__38_comb[55:48]];
  assign p7_array_index_1083787_comb = p6_arr[p7_addedKey__38_comb[47:40]];
  assign p7_array_index_1083788_comb = p6_arr[p7_addedKey__38_comb[39:32]];
  assign p7_array_index_1083789_comb = p6_arr[p7_addedKey__38_comb[31:24]];
  assign p7_array_index_1083790_comb = p6_arr[p7_addedKey__38_comb[23:16]];
  assign p7_array_index_1083791_comb = p6_arr[p7_addedKey__38_comb[15:8]];
  assign p7_array_index_1083551_comb = p6_literal_1076355[p7_res7__389_comb];
  assign p7_array_index_1083793_comb = p6_literal_1076345[p7_array_index_1083777_comb];
  assign p7_array_index_1083794_comb = p6_literal_1076347[p7_array_index_1083778_comb];
  assign p7_array_index_1083795_comb = p6_literal_1076349[p7_array_index_1083779_comb];
  assign p7_array_index_1083796_comb = p6_literal_1076351[p7_array_index_1083780_comb];
  assign p7_array_index_1083797_comb = p6_literal_1076353[p7_array_index_1083781_comb];
  assign p7_array_index_1083798_comb = p6_literal_1076355[p7_array_index_1083782_comb];
  assign p7_array_index_1083799_comb = p6_arr[p7_addedKey__38_comb[79:72]];
  assign p7_array_index_1083801_comb = p6_arr[p7_addedKey__38_comb[63:56]];
  assign p7_res7__395_comb = p6_literal_1076345[p7_res7__394_comb] ^ p6_literal_1076347[p7_res7__393_comb] ^ p6_literal_1076349[p7_res7__392_comb] ^ p6_literal_1076351[p7_res7__391_comb] ^ p6_literal_1076353[p7_res7__390_comb] ^ p7_array_index_1083551_comb ^ p7_res7__388_comb ^ p6_literal_1076358[p7_res7__387_comb] ^ p7_res7__386_comb ^ p7_array_index_1083507_comb ^ p7_array_index_1083481_comb ^ p7_array_index_1083453_comb ^ p7_array_index_1083424_comb ^ p6_literal_1076347[p7_array_index_1083391_comb] ^ p6_literal_1076345[p7_array_index_1083392_comb] ^ p7_array_index_1083393_comb;
  assign p7_res7__608_comb = p7_array_index_1083793_comb ^ p7_array_index_1083794_comb ^ p7_array_index_1083795_comb ^ p7_array_index_1083796_comb ^ p7_array_index_1083797_comb ^ p7_array_index_1083798_comb ^ p7_array_index_1083799_comb ^ p6_literal_1076358[p7_array_index_1083784_comb] ^ p7_array_index_1083801_comb ^ p6_literal_1076355[p7_array_index_1083786_comb] ^ p6_literal_1076353[p7_array_index_1083787_comb] ^ p6_literal_1076351[p7_array_index_1083788_comb] ^ p6_literal_1076349[p7_array_index_1083789_comb] ^ p6_literal_1076347[p7_array_index_1083790_comb] ^ p6_literal_1076345[p7_array_index_1083791_comb] ^ p6_arr[p7_addedKey__38_comb[7:0]];
  assign p7_array_index_1083810_comb = p6_literal_1076345[p7_res7__608_comb];
  assign p7_array_index_1083811_comb = p6_literal_1076347[p7_array_index_1083777_comb];
  assign p7_array_index_1083812_comb = p6_literal_1076349[p7_array_index_1083778_comb];
  assign p7_array_index_1083813_comb = p6_literal_1076351[p7_array_index_1083779_comb];
  assign p7_array_index_1083814_comb = p6_literal_1076353[p7_array_index_1083780_comb];
  assign p7_array_index_1083815_comb = p6_literal_1076355[p7_array_index_1083781_comb];
  assign p7_res7__396_comb = p6_literal_1076345[p7_res7__395_comb] ^ p6_literal_1076347[p7_res7__394_comb] ^ p6_literal_1076349[p7_res7__393_comb] ^ p6_literal_1076351[p7_res7__392_comb] ^ p6_literal_1076353[p7_res7__391_comb] ^ p6_literal_1076355[p7_res7__390_comb] ^ p7_res7__389_comb ^ p6_literal_1076358[p7_res7__388_comb] ^ p7_res7__387_comb ^ p7_array_index_1083519_comb ^ p7_array_index_1083494_comb ^ p7_array_index_1083467_comb ^ p7_array_index_1083438_comb ^ p7_array_index_1083406_comb ^ p6_literal_1076345[p7_array_index_1083391_comb] ^ p7_array_index_1083392_comb;
  assign p7_res7__609_comb = p7_array_index_1083810_comb ^ p7_array_index_1083811_comb ^ p7_array_index_1083812_comb ^ p7_array_index_1083813_comb ^ p7_array_index_1083814_comb ^ p7_array_index_1083815_comb ^ p7_array_index_1083782_comb ^ p6_literal_1076358[p7_array_index_1083799_comb] ^ p7_array_index_1083784_comb ^ p6_literal_1076355[p7_array_index_1083801_comb] ^ p6_literal_1076353[p7_array_index_1083786_comb] ^ p6_literal_1076351[p7_array_index_1083787_comb] ^ p6_literal_1076349[p7_array_index_1083788_comb] ^ p6_literal_1076347[p7_array_index_1083789_comb] ^ p6_literal_1076345[p7_array_index_1083790_comb] ^ p7_array_index_1083791_comb;
  assign p7_array_index_1083825_comb = p6_literal_1076347[p7_res7__608_comb];
  assign p7_array_index_1083826_comb = p6_literal_1076349[p7_array_index_1083777_comb];
  assign p7_array_index_1083827_comb = p6_literal_1076351[p7_array_index_1083778_comb];
  assign p7_array_index_1083828_comb = p6_literal_1076353[p7_array_index_1083779_comb];
  assign p7_array_index_1083829_comb = p6_literal_1076355[p7_array_index_1083780_comb];
  assign p7_res7__397_comb = p6_literal_1076345[p7_res7__396_comb] ^ p6_literal_1076347[p7_res7__395_comb] ^ p6_literal_1076349[p7_res7__394_comb] ^ p6_literal_1076351[p7_res7__393_comb] ^ p6_literal_1076353[p7_res7__392_comb] ^ p6_literal_1076355[p7_res7__391_comb] ^ p7_res7__390_comb ^ p6_literal_1076358[p7_res7__389_comb] ^ p7_res7__388_comb ^ p7_array_index_1083530_comb ^ p7_array_index_1083506_comb ^ p7_array_index_1083480_comb ^ p7_array_index_1083452_comb ^ p7_array_index_1083423_comb ^ p6_literal_1076345[p7_array_index_1083390_comb] ^ p7_array_index_1083391_comb;
  assign p7_res7__610_comb = p6_literal_1076345[p7_res7__609_comb] ^ p7_array_index_1083825_comb ^ p7_array_index_1083826_comb ^ p7_array_index_1083827_comb ^ p7_array_index_1083828_comb ^ p7_array_index_1083829_comb ^ p7_array_index_1083781_comb ^ p6_literal_1076358[p7_array_index_1083782_comb] ^ p7_array_index_1083799_comb ^ p6_literal_1076355[p7_array_index_1083784_comb] ^ p6_literal_1076353[p7_array_index_1083801_comb] ^ p6_literal_1076351[p7_array_index_1083786_comb] ^ p6_literal_1076349[p7_array_index_1083787_comb] ^ p6_literal_1076347[p7_array_index_1083788_comb] ^ p6_literal_1076345[p7_array_index_1083789_comb] ^ p7_array_index_1083790_comb;
  assign p7_array_index_1083839_comb = p6_literal_1076347[p7_res7__609_comb];
  assign p7_array_index_1083840_comb = p6_literal_1076349[p7_res7__608_comb];
  assign p7_array_index_1083841_comb = p6_literal_1076351[p7_array_index_1083777_comb];
  assign p7_array_index_1083842_comb = p6_literal_1076353[p7_array_index_1083778_comb];
  assign p7_array_index_1083843_comb = p6_literal_1076355[p7_array_index_1083779_comb];
  assign p7_res7__398_comb = p6_literal_1076345[p7_res7__397_comb] ^ p6_literal_1076347[p7_res7__396_comb] ^ p6_literal_1076349[p7_res7__395_comb] ^ p6_literal_1076351[p7_res7__394_comb] ^ p6_literal_1076353[p7_res7__393_comb] ^ p6_literal_1076355[p7_res7__392_comb] ^ p7_res7__391_comb ^ p6_literal_1076358[p7_res7__390_comb] ^ p7_res7__389_comb ^ p7_array_index_1083541_comb ^ p7_array_index_1083518_comb ^ p7_array_index_1083493_comb ^ p7_array_index_1083466_comb ^ p7_array_index_1083437_comb ^ p7_array_index_1083405_comb ^ p7_array_index_1083390_comb;
  assign p7_res7__611_comb = p6_literal_1076345[p7_res7__610_comb] ^ p7_array_index_1083839_comb ^ p7_array_index_1083840_comb ^ p7_array_index_1083841_comb ^ p7_array_index_1083842_comb ^ p7_array_index_1083843_comb ^ p7_array_index_1083780_comb ^ p6_literal_1076358[p7_array_index_1083781_comb] ^ p7_array_index_1083782_comb ^ p6_literal_1076355[p7_array_index_1083799_comb] ^ p6_literal_1076353[p7_array_index_1083784_comb] ^ p6_literal_1076351[p7_array_index_1083801_comb] ^ p6_literal_1076349[p7_array_index_1083786_comb] ^ p6_literal_1076347[p7_array_index_1083787_comb] ^ p6_literal_1076345[p7_array_index_1083788_comb] ^ p7_array_index_1083789_comb;
  assign p7_array_index_1083854_comb = p6_literal_1076349[p7_res7__609_comb];
  assign p7_array_index_1083855_comb = p6_literal_1076351[p7_res7__608_comb];
  assign p7_array_index_1083856_comb = p6_literal_1076353[p7_array_index_1083777_comb];
  assign p7_array_index_1083857_comb = p6_literal_1076355[p7_array_index_1083778_comb];
  assign p7_res7__399_comb = p6_literal_1076345[p7_res7__398_comb] ^ p6_literal_1076347[p7_res7__397_comb] ^ p6_literal_1076349[p7_res7__396_comb] ^ p6_literal_1076351[p7_res7__395_comb] ^ p6_literal_1076353[p7_res7__394_comb] ^ p6_literal_1076355[p7_res7__393_comb] ^ p7_res7__392_comb ^ p6_literal_1076358[p7_res7__391_comb] ^ p7_res7__390_comb ^ p7_array_index_1083551_comb ^ p7_array_index_1083529_comb ^ p7_array_index_1083505_comb ^ p7_array_index_1083479_comb ^ p7_array_index_1083451_comb ^ p7_array_index_1083422_comb ^ p7_array_index_1083389_comb;
  assign p7_res7__612_comb = p6_literal_1076345[p7_res7__611_comb] ^ p6_literal_1076347[p7_res7__610_comb] ^ p7_array_index_1083854_comb ^ p7_array_index_1083855_comb ^ p7_array_index_1083856_comb ^ p7_array_index_1083857_comb ^ p7_array_index_1083779_comb ^ p6_literal_1076358[p7_array_index_1083780_comb] ^ p7_array_index_1083781_comb ^ p7_array_index_1083798_comb ^ p6_literal_1076353[p7_array_index_1083799_comb] ^ p6_literal_1076351[p7_array_index_1083784_comb] ^ p6_literal_1076349[p7_array_index_1083801_comb] ^ p6_literal_1076347[p7_array_index_1083786_comb] ^ p6_literal_1076345[p7_array_index_1083787_comb] ^ p7_array_index_1083788_comb;
  assign p7_res__24_comb = {p7_res7__399_comb, p7_res7__398_comb, p7_res7__397_comb, p7_res7__396_comb, p7_res7__395_comb, p7_res7__394_comb, p7_res7__393_comb, p7_res7__392_comb, p7_res7__391_comb, p7_res7__390_comb, p7_res7__389_comb, p7_res7__388_comb, p7_res7__387_comb, p7_res7__386_comb, p7_res7__385_comb, p7_res7__384_comb};
  assign p7_array_index_1083867_comb = p6_literal_1076349[p7_res7__610_comb];
  assign p7_array_index_1083868_comb = p6_literal_1076351[p7_res7__609_comb];
  assign p7_array_index_1083869_comb = p6_literal_1076353[p7_res7__608_comb];
  assign p7_array_index_1083870_comb = p6_literal_1076355[p7_array_index_1083777_comb];
  assign p7_xor_1083591_comb = p7_res__24_comb ^ p7_k7_comb;
  assign p7_res7__613_comb = p6_literal_1076345[p7_res7__612_comb] ^ p6_literal_1076347[p7_res7__611_comb] ^ p7_array_index_1083867_comb ^ p7_array_index_1083868_comb ^ p7_array_index_1083869_comb ^ p7_array_index_1083870_comb ^ p7_array_index_1083778_comb ^ p6_literal_1076358[p7_array_index_1083779_comb] ^ p7_array_index_1083780_comb ^ p7_array_index_1083815_comb ^ p6_literal_1076353[p7_array_index_1083782_comb] ^ p6_literal_1076351[p7_array_index_1083799_comb] ^ p6_literal_1076349[p7_array_index_1083784_comb] ^ p6_literal_1076347[p7_array_index_1083801_comb] ^ p6_literal_1076345[p7_array_index_1083786_comb] ^ p7_array_index_1083787_comb;
  assign p7_addedKey__66_comb = p7_xor_1083591_comb ^ 128'h056c_b6de_319f_0eeb_8e80_9963_10f6_951a;
  assign p7_array_index_1083881_comb = p6_literal_1076351[p7_res7__610_comb];
  assign p7_array_index_1083882_comb = p6_literal_1076353[p7_res7__609_comb];
  assign p7_array_index_1083883_comb = p6_literal_1076355[p7_res7__608_comb];
  assign p7_res7__614_comb = p6_literal_1076345[p7_res7__613_comb] ^ p6_literal_1076347[p7_res7__612_comb] ^ p6_literal_1076349[p7_res7__611_comb] ^ p7_array_index_1083881_comb ^ p7_array_index_1083882_comb ^ p7_array_index_1083883_comb ^ p7_array_index_1083777_comb ^ p6_literal_1076358[p7_array_index_1083778_comb] ^ p7_array_index_1083779_comb ^ p7_array_index_1083829_comb ^ p7_array_index_1083797_comb ^ p6_literal_1076351[p7_array_index_1083782_comb] ^ p6_literal_1076349[p7_array_index_1083799_comb] ^ p6_literal_1076347[p7_array_index_1083784_comb] ^ p6_literal_1076345[p7_array_index_1083801_comb] ^ p7_array_index_1083786_comb;
  assign p7_array_index_1083607_comb = p6_arr[p7_addedKey__66_comb[127:120]];
  assign p7_array_index_1083608_comb = p6_arr[p7_addedKey__66_comb[119:112]];
  assign p7_array_index_1083609_comb = p6_arr[p7_addedKey__66_comb[111:104]];
  assign p7_array_index_1083610_comb = p6_arr[p7_addedKey__66_comb[103:96]];
  assign p7_array_index_1083611_comb = p6_arr[p7_addedKey__66_comb[95:88]];
  assign p7_array_index_1083612_comb = p6_arr[p7_addedKey__66_comb[87:80]];
  assign p7_array_index_1083614_comb = p6_arr[p7_addedKey__66_comb[71:64]];
  assign p7_array_index_1083616_comb = p6_arr[p7_addedKey__66_comb[55:48]];
  assign p7_array_index_1083617_comb = p6_arr[p7_addedKey__66_comb[47:40]];
  assign p7_array_index_1083618_comb = p6_arr[p7_addedKey__66_comb[39:32]];
  assign p7_array_index_1083619_comb = p6_arr[p7_addedKey__66_comb[31:24]];
  assign p7_array_index_1083620_comb = p6_arr[p7_addedKey__66_comb[23:16]];
  assign p7_array_index_1083621_comb = p6_arr[p7_addedKey__66_comb[15:8]];
  assign p7_array_index_1083893_comb = p6_literal_1076351[p7_res7__611_comb];
  assign p7_array_index_1083894_comb = p6_literal_1076353[p7_res7__610_comb];
  assign p7_array_index_1083895_comb = p6_literal_1076355[p7_res7__609_comb];
  assign p7_array_index_1083623_comb = p6_literal_1076345[p7_array_index_1083607_comb];
  assign p7_array_index_1083624_comb = p6_literal_1076347[p7_array_index_1083608_comb];
  assign p7_array_index_1083625_comb = p6_literal_1076349[p7_array_index_1083609_comb];
  assign p7_array_index_1083626_comb = p6_literal_1076351[p7_array_index_1083610_comb];
  assign p7_array_index_1083627_comb = p6_literal_1076353[p7_array_index_1083611_comb];
  assign p7_array_index_1083628_comb = p6_literal_1076355[p7_array_index_1083612_comb];
  assign p7_array_index_1083629_comb = p6_arr[p7_addedKey__66_comb[79:72]];
  assign p7_array_index_1083631_comb = p6_arr[p7_addedKey__66_comb[63:56]];
  assign p7_res7__615_comb = p6_literal_1076345[p7_res7__614_comb] ^ p6_literal_1076347[p7_res7__613_comb] ^ p6_literal_1076349[p7_res7__612_comb] ^ p7_array_index_1083893_comb ^ p7_array_index_1083894_comb ^ p7_array_index_1083895_comb ^ p7_res7__608_comb ^ p6_literal_1076358[p7_array_index_1083777_comb] ^ p7_array_index_1083778_comb ^ p7_array_index_1083843_comb ^ p7_array_index_1083814_comb ^ p6_literal_1076351[p7_array_index_1083781_comb] ^ p6_literal_1076349[p7_array_index_1083782_comb] ^ p6_literal_1076347[p7_array_index_1083799_comb] ^ p6_literal_1076345[p7_array_index_1083784_comb] ^ p7_array_index_1083801_comb;
  assign p7_res7__400_comb = p7_array_index_1083623_comb ^ p7_array_index_1083624_comb ^ p7_array_index_1083625_comb ^ p7_array_index_1083626_comb ^ p7_array_index_1083627_comb ^ p7_array_index_1083628_comb ^ p7_array_index_1083629_comb ^ p6_literal_1076358[p7_array_index_1083614_comb] ^ p7_array_index_1083631_comb ^ p6_literal_1076355[p7_array_index_1083616_comb] ^ p6_literal_1076353[p7_array_index_1083617_comb] ^ p6_literal_1076351[p7_array_index_1083618_comb] ^ p6_literal_1076349[p7_array_index_1083619_comb] ^ p6_literal_1076347[p7_array_index_1083620_comb] ^ p6_literal_1076345[p7_array_index_1083621_comb] ^ p6_arr[p7_addedKey__66_comb[7:0]];
  assign p7_array_index_1083906_comb = p6_literal_1076353[p7_res7__611_comb];
  assign p7_array_index_1083907_comb = p6_literal_1076355[p7_res7__610_comb];
  assign p7_array_index_1083640_comb = p6_literal_1076345[p7_res7__400_comb];
  assign p7_array_index_1083641_comb = p6_literal_1076347[p7_array_index_1083607_comb];
  assign p7_array_index_1083642_comb = p6_literal_1076349[p7_array_index_1083608_comb];
  assign p7_array_index_1083643_comb = p6_literal_1076351[p7_array_index_1083609_comb];
  assign p7_array_index_1083644_comb = p6_literal_1076353[p7_array_index_1083610_comb];
  assign p7_array_index_1083645_comb = p6_literal_1076355[p7_array_index_1083611_comb];
  assign p7_res7__616_comb = p6_literal_1076345[p7_res7__615_comb] ^ p6_literal_1076347[p7_res7__614_comb] ^ p6_literal_1076349[p7_res7__613_comb] ^ p6_literal_1076351[p7_res7__612_comb] ^ p7_array_index_1083906_comb ^ p7_array_index_1083907_comb ^ p7_res7__609_comb ^ p6_literal_1076358[p7_res7__608_comb] ^ p7_array_index_1083777_comb ^ p7_array_index_1083857_comb ^ p7_array_index_1083828_comb ^ p7_array_index_1083796_comb ^ p6_literal_1076349[p7_array_index_1083781_comb] ^ p6_literal_1076347[p7_array_index_1083782_comb] ^ p6_literal_1076345[p7_array_index_1083799_comb] ^ p7_array_index_1083784_comb;
  assign p7_res7__401_comb = p7_array_index_1083640_comb ^ p7_array_index_1083641_comb ^ p7_array_index_1083642_comb ^ p7_array_index_1083643_comb ^ p7_array_index_1083644_comb ^ p7_array_index_1083645_comb ^ p7_array_index_1083612_comb ^ p6_literal_1076358[p7_array_index_1083629_comb] ^ p7_array_index_1083614_comb ^ p6_literal_1076355[p7_array_index_1083631_comb] ^ p6_literal_1076353[p7_array_index_1083616_comb] ^ p6_literal_1076351[p7_array_index_1083617_comb] ^ p6_literal_1076349[p7_array_index_1083618_comb] ^ p6_literal_1076347[p7_array_index_1083619_comb] ^ p6_literal_1076345[p7_array_index_1083620_comb] ^ p7_array_index_1083621_comb;
  assign p7_array_index_1083917_comb = p6_literal_1076353[p7_res7__612_comb];
  assign p7_array_index_1083918_comb = p6_literal_1076355[p7_res7__611_comb];
  assign p7_array_index_1083655_comb = p6_literal_1076347[p7_res7__400_comb];
  assign p7_array_index_1083656_comb = p6_literal_1076349[p7_array_index_1083607_comb];
  assign p7_array_index_1083657_comb = p6_literal_1076351[p7_array_index_1083608_comb];
  assign p7_array_index_1083658_comb = p6_literal_1076353[p7_array_index_1083609_comb];
  assign p7_array_index_1083659_comb = p6_literal_1076355[p7_array_index_1083610_comb];
  assign p7_res7__617_comb = p6_literal_1076345[p7_res7__616_comb] ^ p6_literal_1076347[p7_res7__615_comb] ^ p6_literal_1076349[p7_res7__614_comb] ^ p6_literal_1076351[p7_res7__613_comb] ^ p7_array_index_1083917_comb ^ p7_array_index_1083918_comb ^ p7_res7__610_comb ^ p6_literal_1076358[p7_res7__609_comb] ^ p7_res7__608_comb ^ p7_array_index_1083870_comb ^ p7_array_index_1083842_comb ^ p7_array_index_1083813_comb ^ p6_literal_1076349[p7_array_index_1083780_comb] ^ p6_literal_1076347[p7_array_index_1083781_comb] ^ p6_literal_1076345[p7_array_index_1083782_comb] ^ p7_array_index_1083799_comb;
  assign p7_res7__402_comb = p6_literal_1076345[p7_res7__401_comb] ^ p7_array_index_1083655_comb ^ p7_array_index_1083656_comb ^ p7_array_index_1083657_comb ^ p7_array_index_1083658_comb ^ p7_array_index_1083659_comb ^ p7_array_index_1083611_comb ^ p6_literal_1076358[p7_array_index_1083612_comb] ^ p7_array_index_1083629_comb ^ p6_literal_1076355[p7_array_index_1083614_comb] ^ p6_literal_1076353[p7_array_index_1083631_comb] ^ p6_literal_1076351[p7_array_index_1083616_comb] ^ p6_literal_1076349[p7_array_index_1083617_comb] ^ p6_literal_1076347[p7_array_index_1083618_comb] ^ p6_literal_1076345[p7_array_index_1083619_comb] ^ p7_array_index_1083620_comb;
  assign p7_array_index_1083929_comb = p6_literal_1076355[p7_res7__612_comb];
  assign p7_array_index_1083669_comb = p6_literal_1076347[p7_res7__401_comb];
  assign p7_array_index_1083670_comb = p6_literal_1076349[p7_res7__400_comb];
  assign p7_array_index_1083671_comb = p6_literal_1076351[p7_array_index_1083607_comb];
  assign p7_array_index_1083672_comb = p6_literal_1076353[p7_array_index_1083608_comb];
  assign p7_array_index_1083673_comb = p6_literal_1076355[p7_array_index_1083609_comb];
  assign p7_res7__618_comb = p6_literal_1076345[p7_res7__617_comb] ^ p6_literal_1076347[p7_res7__616_comb] ^ p6_literal_1076349[p7_res7__615_comb] ^ p6_literal_1076351[p7_res7__614_comb] ^ p6_literal_1076353[p7_res7__613_comb] ^ p7_array_index_1083929_comb ^ p7_res7__611_comb ^ p6_literal_1076358[p7_res7__610_comb] ^ p7_res7__609_comb ^ p7_array_index_1083883_comb ^ p7_array_index_1083856_comb ^ p7_array_index_1083827_comb ^ p7_array_index_1083795_comb ^ p6_literal_1076347[p7_array_index_1083780_comb] ^ p6_literal_1076345[p7_array_index_1083781_comb] ^ p7_array_index_1083782_comb;
  assign p7_res7__403_comb = p6_literal_1076345[p7_res7__402_comb] ^ p7_array_index_1083669_comb ^ p7_array_index_1083670_comb ^ p7_array_index_1083671_comb ^ p7_array_index_1083672_comb ^ p7_array_index_1083673_comb ^ p7_array_index_1083610_comb ^ p6_literal_1076358[p7_array_index_1083611_comb] ^ p7_array_index_1083612_comb ^ p6_literal_1076355[p7_array_index_1083629_comb] ^ p6_literal_1076353[p7_array_index_1083614_comb] ^ p6_literal_1076351[p7_array_index_1083631_comb] ^ p6_literal_1076349[p7_array_index_1083616_comb] ^ p6_literal_1076347[p7_array_index_1083617_comb] ^ p6_literal_1076345[p7_array_index_1083618_comb] ^ p7_array_index_1083619_comb;
  assign p7_array_index_1083939_comb = p6_literal_1076355[p7_res7__613_comb];
  assign p7_array_index_1083684_comb = p6_literal_1076349[p7_res7__401_comb];
  assign p7_array_index_1083685_comb = p6_literal_1076351[p7_res7__400_comb];
  assign p7_array_index_1083686_comb = p6_literal_1076353[p7_array_index_1083607_comb];
  assign p7_array_index_1083687_comb = p6_literal_1076355[p7_array_index_1083608_comb];
  assign p7_res7__619_comb = p6_literal_1076345[p7_res7__618_comb] ^ p6_literal_1076347[p7_res7__617_comb] ^ p6_literal_1076349[p7_res7__616_comb] ^ p6_literal_1076351[p7_res7__615_comb] ^ p6_literal_1076353[p7_res7__614_comb] ^ p7_array_index_1083939_comb ^ p7_res7__612_comb ^ p6_literal_1076358[p7_res7__611_comb] ^ p7_res7__610_comb ^ p7_array_index_1083895_comb ^ p7_array_index_1083869_comb ^ p7_array_index_1083841_comb ^ p7_array_index_1083812_comb ^ p6_literal_1076347[p7_array_index_1083779_comb] ^ p6_literal_1076345[p7_array_index_1083780_comb] ^ p7_array_index_1083781_comb;
  assign p7_res7__404_comb = p6_literal_1076345[p7_res7__403_comb] ^ p6_literal_1076347[p7_res7__402_comb] ^ p7_array_index_1083684_comb ^ p7_array_index_1083685_comb ^ p7_array_index_1083686_comb ^ p7_array_index_1083687_comb ^ p7_array_index_1083609_comb ^ p6_literal_1076358[p7_array_index_1083610_comb] ^ p7_array_index_1083611_comb ^ p7_array_index_1083628_comb ^ p6_literal_1076353[p7_array_index_1083629_comb] ^ p6_literal_1076351[p7_array_index_1083614_comb] ^ p6_literal_1076349[p7_array_index_1083631_comb] ^ p6_literal_1076347[p7_array_index_1083616_comb] ^ p6_literal_1076345[p7_array_index_1083617_comb] ^ p7_array_index_1083618_comb;
  assign p7_array_index_1083697_comb = p6_literal_1076349[p7_res7__402_comb];
  assign p7_array_index_1083698_comb = p6_literal_1076351[p7_res7__401_comb];
  assign p7_array_index_1083699_comb = p6_literal_1076353[p7_res7__400_comb];
  assign p7_array_index_1083700_comb = p6_literal_1076355[p7_array_index_1083607_comb];
  assign p7_res7__620_comb = p6_literal_1076345[p7_res7__619_comb] ^ p6_literal_1076347[p7_res7__618_comb] ^ p6_literal_1076349[p7_res7__617_comb] ^ p6_literal_1076351[p7_res7__616_comb] ^ p6_literal_1076353[p7_res7__615_comb] ^ p6_literal_1076355[p7_res7__614_comb] ^ p7_res7__613_comb ^ p6_literal_1076358[p7_res7__612_comb] ^ p7_res7__611_comb ^ p7_array_index_1083907_comb ^ p7_array_index_1083882_comb ^ p7_array_index_1083855_comb ^ p7_array_index_1083826_comb ^ p7_array_index_1083794_comb ^ p6_literal_1076345[p7_array_index_1083779_comb] ^ p7_array_index_1083780_comb;
  assign p7_res7__405_comb = p6_literal_1076345[p7_res7__404_comb] ^ p6_literal_1076347[p7_res7__403_comb] ^ p7_array_index_1083697_comb ^ p7_array_index_1083698_comb ^ p7_array_index_1083699_comb ^ p7_array_index_1083700_comb ^ p7_array_index_1083608_comb ^ p6_literal_1076358[p7_array_index_1083609_comb] ^ p7_array_index_1083610_comb ^ p7_array_index_1083645_comb ^ p6_literal_1076353[p7_array_index_1083612_comb] ^ p6_literal_1076351[p7_array_index_1083629_comb] ^ p6_literal_1076349[p7_array_index_1083614_comb] ^ p6_literal_1076347[p7_array_index_1083631_comb] ^ p6_literal_1076345[p7_array_index_1083616_comb] ^ p7_array_index_1083617_comb;
  assign p7_array_index_1083711_comb = p6_literal_1076351[p7_res7__402_comb];
  assign p7_array_index_1083712_comb = p6_literal_1076353[p7_res7__401_comb];
  assign p7_array_index_1083713_comb = p6_literal_1076355[p7_res7__400_comb];
  assign p7_res7__621_comb = p6_literal_1076345[p7_res7__620_comb] ^ p6_literal_1076347[p7_res7__619_comb] ^ p6_literal_1076349[p7_res7__618_comb] ^ p6_literal_1076351[p7_res7__617_comb] ^ p6_literal_1076353[p7_res7__616_comb] ^ p6_literal_1076355[p7_res7__615_comb] ^ p7_res7__614_comb ^ p6_literal_1076358[p7_res7__613_comb] ^ p7_res7__612_comb ^ p7_array_index_1083918_comb ^ p7_array_index_1083894_comb ^ p7_array_index_1083868_comb ^ p7_array_index_1083840_comb ^ p7_array_index_1083811_comb ^ p6_literal_1076345[p7_array_index_1083778_comb] ^ p7_array_index_1083779_comb;
  assign p7_res7__406_comb = p6_literal_1076345[p7_res7__405_comb] ^ p6_literal_1076347[p7_res7__404_comb] ^ p6_literal_1076349[p7_res7__403_comb] ^ p7_array_index_1083711_comb ^ p7_array_index_1083712_comb ^ p7_array_index_1083713_comb ^ p7_array_index_1083607_comb ^ p6_literal_1076358[p7_array_index_1083608_comb] ^ p7_array_index_1083609_comb ^ p7_array_index_1083659_comb ^ p7_array_index_1083627_comb ^ p6_literal_1076351[p7_array_index_1083612_comb] ^ p6_literal_1076349[p7_array_index_1083629_comb] ^ p6_literal_1076347[p7_array_index_1083614_comb] ^ p6_literal_1076345[p7_array_index_1083631_comb] ^ p7_array_index_1083616_comb;
  assign p7_array_index_1083723_comb = p6_literal_1076351[p7_res7__403_comb];
  assign p7_array_index_1083724_comb = p6_literal_1076353[p7_res7__402_comb];
  assign p7_array_index_1083725_comb = p6_literal_1076355[p7_res7__401_comb];
  assign p7_res7__622_comb = p6_literal_1076345[p7_res7__621_comb] ^ p6_literal_1076347[p7_res7__620_comb] ^ p6_literal_1076349[p7_res7__619_comb] ^ p6_literal_1076351[p7_res7__618_comb] ^ p6_literal_1076353[p7_res7__617_comb] ^ p6_literal_1076355[p7_res7__616_comb] ^ p7_res7__615_comb ^ p6_literal_1076358[p7_res7__614_comb] ^ p7_res7__613_comb ^ p7_array_index_1083929_comb ^ p7_array_index_1083906_comb ^ p7_array_index_1083881_comb ^ p7_array_index_1083854_comb ^ p7_array_index_1083825_comb ^ p7_array_index_1083793_comb ^ p7_array_index_1083778_comb;
  assign p7_res7__407_comb = p6_literal_1076345[p7_res7__406_comb] ^ p6_literal_1076347[p7_res7__405_comb] ^ p6_literal_1076349[p7_res7__404_comb] ^ p7_array_index_1083723_comb ^ p7_array_index_1083724_comb ^ p7_array_index_1083725_comb ^ p7_res7__400_comb ^ p6_literal_1076358[p7_array_index_1083607_comb] ^ p7_array_index_1083608_comb ^ p7_array_index_1083673_comb ^ p7_array_index_1083644_comb ^ p6_literal_1076351[p7_array_index_1083611_comb] ^ p6_literal_1076349[p7_array_index_1083612_comb] ^ p6_literal_1076347[p7_array_index_1083629_comb] ^ p6_literal_1076345[p7_array_index_1083614_comb] ^ p7_array_index_1083631_comb;
  assign p7_array_index_1083736_comb = p6_literal_1076353[p7_res7__403_comb];
  assign p7_array_index_1083737_comb = p6_literal_1076355[p7_res7__402_comb];
  assign p7_res7__623_comb = p6_literal_1076345[p7_res7__622_comb] ^ p6_literal_1076347[p7_res7__621_comb] ^ p6_literal_1076349[p7_res7__620_comb] ^ p6_literal_1076351[p7_res7__619_comb] ^ p6_literal_1076353[p7_res7__618_comb] ^ p6_literal_1076355[p7_res7__617_comb] ^ p7_res7__616_comb ^ p6_literal_1076358[p7_res7__615_comb] ^ p7_res7__614_comb ^ p7_array_index_1083939_comb ^ p7_array_index_1083917_comb ^ p7_array_index_1083893_comb ^ p7_array_index_1083867_comb ^ p7_array_index_1083839_comb ^ p7_array_index_1083810_comb ^ p7_array_index_1083777_comb;
  assign p7_res7__408_comb = p6_literal_1076345[p7_res7__407_comb] ^ p6_literal_1076347[p7_res7__406_comb] ^ p6_literal_1076349[p7_res7__405_comb] ^ p6_literal_1076351[p7_res7__404_comb] ^ p7_array_index_1083736_comb ^ p7_array_index_1083737_comb ^ p7_res7__401_comb ^ p6_literal_1076358[p7_res7__400_comb] ^ p7_array_index_1083607_comb ^ p7_array_index_1083687_comb ^ p7_array_index_1083658_comb ^ p7_array_index_1083626_comb ^ p6_literal_1076349[p7_array_index_1083611_comb] ^ p6_literal_1076347[p7_array_index_1083612_comb] ^ p6_literal_1076345[p7_array_index_1083629_comb] ^ p7_array_index_1083614_comb;
  assign p7_res__38_comb = {p7_res7__623_comb, p7_res7__622_comb, p7_res7__621_comb, p7_res7__620_comb, p7_res7__619_comb, p7_res7__618_comb, p7_res7__617_comb, p7_res7__616_comb, p7_res7__615_comb, p7_res7__614_comb, p7_res7__613_comb, p7_res7__612_comb, p7_res7__611_comb, p7_res7__610_comb, p7_res7__609_comb, p7_res7__608_comb};
  assign p7_array_index_1083747_comb = p6_literal_1076353[p7_res7__404_comb];
  assign p7_array_index_1083748_comb = p6_literal_1076355[p7_res7__403_comb];
  assign p7_addedKey__39_comb = p7_k7_comb ^ p7_res__38_comb;
  assign p7_res7__409_comb = p6_literal_1076345[p7_res7__408_comb] ^ p6_literal_1076347[p7_res7__407_comb] ^ p6_literal_1076349[p7_res7__406_comb] ^ p6_literal_1076351[p7_res7__405_comb] ^ p7_array_index_1083747_comb ^ p7_array_index_1083748_comb ^ p7_res7__402_comb ^ p6_literal_1076358[p7_res7__401_comb] ^ p7_res7__400_comb ^ p7_array_index_1083700_comb ^ p7_array_index_1083672_comb ^ p7_array_index_1083643_comb ^ p6_literal_1076349[p7_array_index_1083610_comb] ^ p6_literal_1076347[p7_array_index_1083611_comb] ^ p6_literal_1076345[p7_array_index_1083612_comb] ^ p7_array_index_1083629_comb;
  assign p7_array_index_1083754_comb = p6_literal_1076345[p7_res7__409_comb];
  assign p7_array_index_1083755_comb = p6_literal_1076347[p7_res7__408_comb];
  assign p7_array_index_1083756_comb = p6_literal_1076349[p7_res7__407_comb];
  assign p7_array_index_1083757_comb = p6_literal_1076351[p7_res7__406_comb];
  assign p7_array_index_1083758_comb = p6_literal_1076353[p7_res7__405_comb];
  assign p7_array_index_1083759_comb = p6_literal_1076355[p7_res7__404_comb];
  assign p7_array_index_1083760_comb = p6_literal_1076358[p7_res7__402_comb];
  assign p7_array_index_1083761_comb = p6_literal_1076347[p7_array_index_1083610_comb];
  assign p7_array_index_1083762_comb = p6_literal_1076345[p7_array_index_1083611_comb];
  assign p7_array_index_1083993_comb = p6_arr[p7_addedKey__39_comb[127:120]];
  assign p7_array_index_1083994_comb = p6_arr[p7_addedKey__39_comb[119:112]];
  assign p7_array_index_1083995_comb = p6_arr[p7_addedKey__39_comb[111:104]];
  assign p7_array_index_1083996_comb = p6_arr[p7_addedKey__39_comb[103:96]];
  assign p7_array_index_1083997_comb = p6_arr[p7_addedKey__39_comb[95:88]];
  assign p7_array_index_1083998_comb = p6_arr[p7_addedKey__39_comb[87:80]];
  assign p7_array_index_1084000_comb = p6_arr[p7_addedKey__39_comb[71:64]];
  assign p7_array_index_1084002_comb = p6_arr[p7_addedKey__39_comb[55:48]];
  assign p7_array_index_1084003_comb = p6_arr[p7_addedKey__39_comb[47:40]];
  assign p7_array_index_1084004_comb = p6_arr[p7_addedKey__39_comb[39:32]];
  assign p7_array_index_1084005_comb = p6_arr[p7_addedKey__39_comb[31:24]];
  assign p7_array_index_1084006_comb = p6_arr[p7_addedKey__39_comb[23:16]];
  assign p7_array_index_1084007_comb = p6_arr[p7_addedKey__39_comb[15:8]];
  assign p7_array_index_1084009_comb = p6_arr[p7_addedKey__39_comb[79:72]];
  assign p7_array_index_1084010_comb = p6_arr[p7_addedKey__39_comb[63:56]];
  assign p7_array_index_1084011_comb = p6_arr[p7_addedKey__39_comb[7:0]];

  // Registers for pipe stage 7:
  reg [127:0] p7_k6;
  reg [127:0] p7_xor_1083591;
  reg [7:0] p7_array_index_1083607;
  reg [7:0] p7_array_index_1083608;
  reg [7:0] p7_array_index_1083609;
  reg [7:0] p7_array_index_1083610;
  reg [7:0] p7_array_index_1083611;
  reg [7:0] p7_array_index_1083612;
  reg [7:0] p7_array_index_1083623;
  reg [7:0] p7_array_index_1083624;
  reg [7:0] p7_array_index_1083625;
  reg [7:0] p7_res7__400;
  reg [7:0] p7_array_index_1083640;
  reg [7:0] p7_array_index_1083641;
  reg [7:0] p7_array_index_1083642;
  reg [7:0] p7_res7__401;
  reg [7:0] p7_array_index_1083655;
  reg [7:0] p7_array_index_1083656;
  reg [7:0] p7_array_index_1083657;
  reg [7:0] p7_res7__402;
  reg [7:0] p7_array_index_1083669;
  reg [7:0] p7_array_index_1083670;
  reg [7:0] p7_array_index_1083671;
  reg [7:0] p7_res7__403;
  reg [7:0] p7_array_index_1083684;
  reg [7:0] p7_array_index_1083685;
  reg [7:0] p7_array_index_1083686;
  reg [7:0] p7_res7__404;
  reg [7:0] p7_array_index_1083697;
  reg [7:0] p7_array_index_1083698;
  reg [7:0] p7_array_index_1083699;
  reg [7:0] p7_res7__405;
  reg [7:0] p7_array_index_1083711;
  reg [7:0] p7_array_index_1083712;
  reg [7:0] p7_array_index_1083713;
  reg [7:0] p7_res7__406;
  reg [7:0] p7_array_index_1083723;
  reg [7:0] p7_array_index_1083724;
  reg [7:0] p7_array_index_1083725;
  reg [7:0] p7_res7__407;
  reg [7:0] p7_array_index_1083736;
  reg [7:0] p7_array_index_1083737;
  reg [7:0] p7_res7__408;
  reg [7:0] p7_array_index_1083747;
  reg [7:0] p7_array_index_1083748;
  reg [7:0] p7_res7__409;
  reg [7:0] p7_array_index_1083754;
  reg [7:0] p7_array_index_1083755;
  reg [7:0] p7_array_index_1083756;
  reg [7:0] p7_array_index_1083757;
  reg [7:0] p7_array_index_1083758;
  reg [7:0] p7_array_index_1083759;
  reg [7:0] p7_array_index_1083760;
  reg [7:0] p7_array_index_1083761;
  reg [7:0] p7_array_index_1083762;
  reg [7:0] p7_array_index_1083993;
  reg [7:0] p7_array_index_1083994;
  reg [7:0] p7_array_index_1083995;
  reg [7:0] p7_array_index_1083996;
  reg [7:0] p7_array_index_1083997;
  reg [7:0] p7_array_index_1083998;
  reg [7:0] p7_array_index_1084000;
  reg [7:0] p7_array_index_1084002;
  reg [7:0] p7_array_index_1084003;
  reg [7:0] p7_array_index_1084004;
  reg [7:0] p7_array_index_1084005;
  reg [7:0] p7_array_index_1084006;
  reg [7:0] p7_array_index_1084007;
  reg [7:0] p7_array_index_1084009;
  reg [7:0] p7_array_index_1084010;
  reg [7:0] p7_array_index_1084011;
  reg [7:0] p8_arr[256];
  reg [7:0] p8_literal_1076345[256];
  reg [7:0] p8_literal_1076347[256];
  reg [7:0] p8_literal_1076349[256];
  reg [7:0] p8_literal_1076351[256];
  reg [7:0] p8_literal_1076353[256];
  reg [7:0] p8_literal_1076355[256];
  reg [7:0] p8_literal_1076358[256];
  always_ff @ (posedge clk) begin
    p7_k6 <= p7_k6_comb;
    p7_xor_1083591 <= p7_xor_1083591_comb;
    p7_array_index_1083607 <= p7_array_index_1083607_comb;
    p7_array_index_1083608 <= p7_array_index_1083608_comb;
    p7_array_index_1083609 <= p7_array_index_1083609_comb;
    p7_array_index_1083610 <= p7_array_index_1083610_comb;
    p7_array_index_1083611 <= p7_array_index_1083611_comb;
    p7_array_index_1083612 <= p7_array_index_1083612_comb;
    p7_array_index_1083623 <= p7_array_index_1083623_comb;
    p7_array_index_1083624 <= p7_array_index_1083624_comb;
    p7_array_index_1083625 <= p7_array_index_1083625_comb;
    p7_res7__400 <= p7_res7__400_comb;
    p7_array_index_1083640 <= p7_array_index_1083640_comb;
    p7_array_index_1083641 <= p7_array_index_1083641_comb;
    p7_array_index_1083642 <= p7_array_index_1083642_comb;
    p7_res7__401 <= p7_res7__401_comb;
    p7_array_index_1083655 <= p7_array_index_1083655_comb;
    p7_array_index_1083656 <= p7_array_index_1083656_comb;
    p7_array_index_1083657 <= p7_array_index_1083657_comb;
    p7_res7__402 <= p7_res7__402_comb;
    p7_array_index_1083669 <= p7_array_index_1083669_comb;
    p7_array_index_1083670 <= p7_array_index_1083670_comb;
    p7_array_index_1083671 <= p7_array_index_1083671_comb;
    p7_res7__403 <= p7_res7__403_comb;
    p7_array_index_1083684 <= p7_array_index_1083684_comb;
    p7_array_index_1083685 <= p7_array_index_1083685_comb;
    p7_array_index_1083686 <= p7_array_index_1083686_comb;
    p7_res7__404 <= p7_res7__404_comb;
    p7_array_index_1083697 <= p7_array_index_1083697_comb;
    p7_array_index_1083698 <= p7_array_index_1083698_comb;
    p7_array_index_1083699 <= p7_array_index_1083699_comb;
    p7_res7__405 <= p7_res7__405_comb;
    p7_array_index_1083711 <= p7_array_index_1083711_comb;
    p7_array_index_1083712 <= p7_array_index_1083712_comb;
    p7_array_index_1083713 <= p7_array_index_1083713_comb;
    p7_res7__406 <= p7_res7__406_comb;
    p7_array_index_1083723 <= p7_array_index_1083723_comb;
    p7_array_index_1083724 <= p7_array_index_1083724_comb;
    p7_array_index_1083725 <= p7_array_index_1083725_comb;
    p7_res7__407 <= p7_res7__407_comb;
    p7_array_index_1083736 <= p7_array_index_1083736_comb;
    p7_array_index_1083737 <= p7_array_index_1083737_comb;
    p7_res7__408 <= p7_res7__408_comb;
    p7_array_index_1083747 <= p7_array_index_1083747_comb;
    p7_array_index_1083748 <= p7_array_index_1083748_comb;
    p7_res7__409 <= p7_res7__409_comb;
    p7_array_index_1083754 <= p7_array_index_1083754_comb;
    p7_array_index_1083755 <= p7_array_index_1083755_comb;
    p7_array_index_1083756 <= p7_array_index_1083756_comb;
    p7_array_index_1083757 <= p7_array_index_1083757_comb;
    p7_array_index_1083758 <= p7_array_index_1083758_comb;
    p7_array_index_1083759 <= p7_array_index_1083759_comb;
    p7_array_index_1083760 <= p7_array_index_1083760_comb;
    p7_array_index_1083761 <= p7_array_index_1083761_comb;
    p7_array_index_1083762 <= p7_array_index_1083762_comb;
    p7_array_index_1083993 <= p7_array_index_1083993_comb;
    p7_array_index_1083994 <= p7_array_index_1083994_comb;
    p7_array_index_1083995 <= p7_array_index_1083995_comb;
    p7_array_index_1083996 <= p7_array_index_1083996_comb;
    p7_array_index_1083997 <= p7_array_index_1083997_comb;
    p7_array_index_1083998 <= p7_array_index_1083998_comb;
    p7_array_index_1084000 <= p7_array_index_1084000_comb;
    p7_array_index_1084002 <= p7_array_index_1084002_comb;
    p7_array_index_1084003 <= p7_array_index_1084003_comb;
    p7_array_index_1084004 <= p7_array_index_1084004_comb;
    p7_array_index_1084005 <= p7_array_index_1084005_comb;
    p7_array_index_1084006 <= p7_array_index_1084006_comb;
    p7_array_index_1084007 <= p7_array_index_1084007_comb;
    p7_array_index_1084009 <= p7_array_index_1084009_comb;
    p7_array_index_1084010 <= p7_array_index_1084010_comb;
    p7_array_index_1084011 <= p7_array_index_1084011_comb;
    p8_arr <= p7_arr;
    p8_literal_1076345 <= p7_literal_1076345;
    p8_literal_1076347 <= p7_literal_1076347;
    p8_literal_1076349 <= p7_literal_1076349;
    p8_literal_1076351 <= p7_literal_1076351;
    p8_literal_1076353 <= p7_literal_1076353;
    p8_literal_1076355 <= p7_literal_1076355;
    p8_literal_1076358 <= p7_literal_1076358;
  end

  // ===== Pipe stage 8:
  wire [7:0] p8_res7__410_comb;
  wire [7:0] p8_array_index_1084176_comb;
  wire [7:0] p8_res7__411_comb;
  wire [7:0] p8_res7__412_comb;
  wire [7:0] p8_res7__413_comb;
  wire [7:0] p8_res7__414_comb;
  wire [7:0] p8_res7__415_comb;
  wire [127:0] p8_res__25_comb;
  wire [127:0] p8_xor_1084216_comb;
  wire [127:0] p8_addedKey__67_comb;
  wire [7:0] p8_array_index_1084232_comb;
  wire [7:0] p8_array_index_1084233_comb;
  wire [7:0] p8_array_index_1084234_comb;
  wire [7:0] p8_array_index_1084235_comb;
  wire [7:0] p8_array_index_1084236_comb;
  wire [7:0] p8_array_index_1084237_comb;
  wire [7:0] p8_array_index_1084239_comb;
  wire [7:0] p8_array_index_1084241_comb;
  wire [7:0] p8_array_index_1084242_comb;
  wire [7:0] p8_array_index_1084243_comb;
  wire [7:0] p8_array_index_1084244_comb;
  wire [7:0] p8_array_index_1084245_comb;
  wire [7:0] p8_array_index_1084246_comb;
  wire [7:0] p8_array_index_1084248_comb;
  wire [7:0] p8_array_index_1084249_comb;
  wire [7:0] p8_array_index_1084250_comb;
  wire [7:0] p8_array_index_1084251_comb;
  wire [7:0] p8_array_index_1084252_comb;
  wire [7:0] p8_array_index_1084253_comb;
  wire [7:0] p8_array_index_1084254_comb;
  wire [7:0] p8_array_index_1084256_comb;
  wire [7:0] p8_res7__416_comb;
  wire [7:0] p8_array_index_1084265_comb;
  wire [7:0] p8_array_index_1084266_comb;
  wire [7:0] p8_array_index_1084267_comb;
  wire [7:0] p8_array_index_1084268_comb;
  wire [7:0] p8_array_index_1084269_comb;
  wire [7:0] p8_array_index_1084270_comb;
  wire [7:0] p8_res7__417_comb;
  wire [7:0] p8_array_index_1084280_comb;
  wire [7:0] p8_array_index_1084281_comb;
  wire [7:0] p8_array_index_1084282_comb;
  wire [7:0] p8_array_index_1084283_comb;
  wire [7:0] p8_array_index_1084284_comb;
  wire [7:0] p8_res7__418_comb;
  wire [7:0] p8_array_index_1084294_comb;
  wire [7:0] p8_array_index_1084295_comb;
  wire [7:0] p8_array_index_1084296_comb;
  wire [7:0] p8_array_index_1084297_comb;
  wire [7:0] p8_array_index_1084298_comb;
  wire [7:0] p8_res7__419_comb;
  wire [7:0] p8_array_index_1084309_comb;
  wire [7:0] p8_array_index_1084310_comb;
  wire [7:0] p8_array_index_1084311_comb;
  wire [7:0] p8_array_index_1084312_comb;
  wire [7:0] p8_res7__420_comb;
  wire [7:0] p8_array_index_1084322_comb;
  wire [7:0] p8_array_index_1084323_comb;
  wire [7:0] p8_array_index_1084324_comb;
  wire [7:0] p8_array_index_1084325_comb;
  wire [7:0] p8_res7__421_comb;
  wire [7:0] p8_array_index_1084336_comb;
  wire [7:0] p8_array_index_1084337_comb;
  wire [7:0] p8_array_index_1084338_comb;
  wire [7:0] p8_res7__422_comb;
  wire [7:0] p8_array_index_1084348_comb;
  wire [7:0] p8_array_index_1084349_comb;
  wire [7:0] p8_array_index_1084350_comb;
  wire [7:0] p8_res7__423_comb;
  wire [7:0] p8_array_index_1084361_comb;
  wire [7:0] p8_array_index_1084362_comb;
  wire [7:0] p8_res7__424_comb;
  wire [7:0] p8_array_index_1084372_comb;
  wire [7:0] p8_array_index_1084373_comb;
  wire [7:0] p8_res7__425_comb;
  wire [7:0] p8_array_index_1084384_comb;
  wire [7:0] p8_res7__426_comb;
  wire [7:0] p8_array_index_1084394_comb;
  wire [7:0] p8_res7__427_comb;
  wire [7:0] p8_res7__428_comb;
  wire [7:0] p8_res7__429_comb;
  wire [7:0] p8_res7__430_comb;
  wire [7:0] p8_res7__431_comb;
  wire [127:0] p8_res__26_comb;
  wire [127:0] p8_xor_1084434_comb;
  wire [127:0] p8_addedKey__68_comb;
  wire [7:0] p8_array_index_1084450_comb;
  wire [7:0] p8_array_index_1084451_comb;
  wire [7:0] p8_array_index_1084452_comb;
  wire [7:0] p8_array_index_1084453_comb;
  wire [7:0] p8_array_index_1084454_comb;
  wire [7:0] p8_array_index_1084455_comb;
  wire [7:0] p8_array_index_1084457_comb;
  wire [7:0] p8_array_index_1084459_comb;
  wire [7:0] p8_array_index_1084460_comb;
  wire [7:0] p8_array_index_1084461_comb;
  wire [7:0] p8_array_index_1084462_comb;
  wire [7:0] p8_array_index_1084463_comb;
  wire [7:0] p8_array_index_1084464_comb;
  wire [7:0] p8_array_index_1084466_comb;
  wire [7:0] p8_array_index_1084467_comb;
  wire [7:0] p8_array_index_1084468_comb;
  wire [7:0] p8_array_index_1084469_comb;
  wire [7:0] p8_array_index_1084470_comb;
  wire [7:0] p8_array_index_1084471_comb;
  wire [7:0] p8_array_index_1084472_comb;
  wire [7:0] p8_array_index_1084474_comb;
  wire [7:0] p8_res7__432_comb;
  wire [7:0] p8_array_index_1084483_comb;
  wire [7:0] p8_array_index_1084484_comb;
  wire [7:0] p8_array_index_1084485_comb;
  wire [7:0] p8_array_index_1084486_comb;
  wire [7:0] p8_array_index_1084487_comb;
  wire [7:0] p8_array_index_1084488_comb;
  wire [7:0] p8_res7__433_comb;
  wire [7:0] p8_array_index_1084498_comb;
  wire [7:0] p8_array_index_1084499_comb;
  wire [7:0] p8_array_index_1084500_comb;
  wire [7:0] p8_array_index_1084501_comb;
  wire [7:0] p8_array_index_1084502_comb;
  wire [7:0] p8_res7__434_comb;
  wire [7:0] p8_array_index_1084512_comb;
  wire [7:0] p8_array_index_1084513_comb;
  wire [7:0] p8_array_index_1084514_comb;
  wire [7:0] p8_array_index_1084515_comb;
  wire [7:0] p8_array_index_1084516_comb;
  wire [7:0] p8_res7__435_comb;
  wire [7:0] p8_array_index_1084527_comb;
  wire [7:0] p8_array_index_1084528_comb;
  wire [7:0] p8_array_index_1084529_comb;
  wire [7:0] p8_array_index_1084530_comb;
  wire [7:0] p8_res7__436_comb;
  wire [7:0] p8_array_index_1084540_comb;
  wire [7:0] p8_array_index_1084541_comb;
  wire [7:0] p8_array_index_1084542_comb;
  wire [7:0] p8_array_index_1084543_comb;
  wire [7:0] p8_res7__437_comb;
  wire [7:0] p8_array_index_1084554_comb;
  wire [7:0] p8_array_index_1084555_comb;
  wire [7:0] p8_array_index_1084556_comb;
  wire [7:0] p8_res7__438_comb;
  wire [7:0] p8_array_index_1084566_comb;
  wire [7:0] p8_array_index_1084567_comb;
  wire [7:0] p8_array_index_1084568_comb;
  wire [7:0] p8_res7__439_comb;
  wire [7:0] p8_array_index_1084579_comb;
  wire [7:0] p8_array_index_1084580_comb;
  wire [7:0] p8_res7__440_comb;
  wire [7:0] p8_array_index_1084590_comb;
  wire [7:0] p8_array_index_1084591_comb;
  wire [7:0] p8_res7__441_comb;
  wire [7:0] p8_array_index_1084602_comb;
  wire [7:0] p8_res7__442_comb;
  wire [7:0] p8_array_index_1084612_comb;
  wire [7:0] p8_res7__443_comb;
  wire [7:0] p8_res7__444_comb;
  wire [7:0] p8_res7__445_comb;
  wire [7:0] p8_res7__446_comb;
  wire [7:0] p8_res7__447_comb;
  wire [127:0] p8_res__27_comb;
  wire [127:0] p8_xor_1084652_comb;
  wire [127:0] p8_addedKey__69_comb;
  wire [7:0] p8_array_index_1084668_comb;
  wire [7:0] p8_array_index_1084669_comb;
  wire [7:0] p8_array_index_1084670_comb;
  wire [7:0] p8_array_index_1084671_comb;
  wire [7:0] p8_array_index_1084672_comb;
  wire [7:0] p8_array_index_1084673_comb;
  wire [7:0] p8_array_index_1084675_comb;
  wire [7:0] p8_array_index_1084677_comb;
  wire [7:0] p8_array_index_1084678_comb;
  wire [7:0] p8_array_index_1084679_comb;
  wire [7:0] p8_array_index_1084680_comb;
  wire [7:0] p8_array_index_1084681_comb;
  wire [7:0] p8_array_index_1084682_comb;
  wire [7:0] p8_array_index_1084684_comb;
  wire [7:0] p8_array_index_1084685_comb;
  wire [7:0] p8_array_index_1084686_comb;
  wire [7:0] p8_array_index_1084687_comb;
  wire [7:0] p8_array_index_1084688_comb;
  wire [7:0] p8_array_index_1084689_comb;
  wire [7:0] p8_array_index_1084690_comb;
  wire [7:0] p8_array_index_1084692_comb;
  wire [7:0] p8_res7__448_comb;
  wire [7:0] p8_array_index_1084701_comb;
  wire [7:0] p8_array_index_1084702_comb;
  wire [7:0] p8_array_index_1084703_comb;
  wire [7:0] p8_array_index_1084704_comb;
  wire [7:0] p8_array_index_1084705_comb;
  wire [7:0] p8_array_index_1084706_comb;
  wire [7:0] p8_res7__449_comb;
  wire [7:0] p8_array_index_1084716_comb;
  wire [7:0] p8_array_index_1084717_comb;
  wire [7:0] p8_array_index_1084718_comb;
  wire [7:0] p8_array_index_1084719_comb;
  wire [7:0] p8_array_index_1084720_comb;
  wire [7:0] p8_res7__450_comb;
  wire [7:0] p8_array_index_1084730_comb;
  wire [7:0] p8_array_index_1084731_comb;
  wire [7:0] p8_array_index_1084732_comb;
  wire [7:0] p8_array_index_1084733_comb;
  wire [7:0] p8_array_index_1084734_comb;
  wire [7:0] p8_res7__451_comb;
  wire [7:0] p8_array_index_1084745_comb;
  wire [7:0] p8_array_index_1084746_comb;
  wire [7:0] p8_array_index_1084747_comb;
  wire [7:0] p8_array_index_1084748_comb;
  wire [7:0] p8_res7__452_comb;
  wire [7:0] p8_array_index_1084758_comb;
  wire [7:0] p8_array_index_1084759_comb;
  wire [7:0] p8_array_index_1084760_comb;
  wire [7:0] p8_array_index_1084761_comb;
  wire [7:0] p8_res7__453_comb;
  wire [7:0] p8_array_index_1084772_comb;
  wire [7:0] p8_array_index_1084773_comb;
  wire [7:0] p8_array_index_1084774_comb;
  wire [7:0] p8_res7__454_comb;
  wire [7:0] p8_array_index_1084784_comb;
  wire [7:0] p8_array_index_1084785_comb;
  wire [7:0] p8_array_index_1084786_comb;
  wire [7:0] p8_array_index_1084974_comb;
  wire [7:0] p8_array_index_1084975_comb;
  wire [7:0] p8_array_index_1084976_comb;
  wire [7:0] p8_array_index_1084977_comb;
  wire [7:0] p8_array_index_1084978_comb;
  wire [7:0] p8_array_index_1084979_comb;
  wire [7:0] p8_res7__455_comb;
  wire [7:0] p8_res7__624_comb;
  wire [7:0] p8_array_index_1084797_comb;
  wire [7:0] p8_array_index_1084798_comb;
  wire [7:0] p8_array_index_1084988_comb;
  wire [7:0] p8_array_index_1084989_comb;
  wire [7:0] p8_array_index_1084990_comb;
  wire [7:0] p8_array_index_1084991_comb;
  wire [7:0] p8_array_index_1084992_comb;
  wire [7:0] p8_array_index_1084993_comb;
  wire [7:0] p8_res7__456_comb;
  wire [7:0] p8_res7__625_comb;
  wire [7:0] p8_array_index_1084808_comb;
  wire [7:0] p8_array_index_1084809_comb;
  wire [7:0] p8_array_index_1085003_comb;
  wire [7:0] p8_array_index_1085004_comb;
  wire [7:0] p8_array_index_1085005_comb;
  wire [7:0] p8_array_index_1085006_comb;
  wire [7:0] p8_array_index_1085007_comb;
  wire [7:0] p8_res7__457_comb;
  wire [7:0] p8_res7__626_comb;
  wire [7:0] p8_array_index_1084820_comb;
  wire [7:0] p8_array_index_1085017_comb;
  wire [7:0] p8_array_index_1085018_comb;
  wire [7:0] p8_array_index_1085019_comb;
  wire [7:0] p8_array_index_1085020_comb;
  wire [7:0] p8_array_index_1085021_comb;
  wire [7:0] p8_res7__458_comb;
  wire [7:0] p8_res7__627_comb;
  wire [7:0] p8_array_index_1084830_comb;
  wire [7:0] p8_array_index_1085032_comb;
  wire [7:0] p8_array_index_1085033_comb;
  wire [7:0] p8_array_index_1085034_comb;
  wire [7:0] p8_array_index_1085035_comb;
  wire [7:0] p8_res7__459_comb;
  wire [7:0] p8_res7__628_comb;
  wire [7:0] p8_array_index_1085045_comb;
  wire [7:0] p8_array_index_1085046_comb;
  wire [7:0] p8_array_index_1085047_comb;
  wire [7:0] p8_array_index_1085048_comb;
  wire [7:0] p8_res7__460_comb;
  wire [7:0] p8_res7__629_comb;
  wire [7:0] p8_array_index_1085059_comb;
  wire [7:0] p8_array_index_1085060_comb;
  wire [7:0] p8_array_index_1085061_comb;
  wire [7:0] p8_res7__461_comb;
  wire [7:0] p8_res7__630_comb;
  wire [7:0] p8_array_index_1085071_comb;
  wire [7:0] p8_array_index_1085072_comb;
  wire [7:0] p8_array_index_1085073_comb;
  wire [7:0] p8_res7__462_comb;
  wire [7:0] p8_res7__631_comb;
  wire [7:0] p8_array_index_1085084_comb;
  wire [7:0] p8_array_index_1085085_comb;
  wire [7:0] p8_res7__463_comb;
  wire [7:0] p8_res7__632_comb;
  wire [127:0] p8_res__28_comb;
  wire [7:0] p8_array_index_1085095_comb;
  wire [7:0] p8_array_index_1085096_comb;
  wire [127:0] p8_xor_1084870_comb;
  wire [7:0] p8_res7__633_comb;
  wire [127:0] p8_addedKey__70_comb;
  wire [7:0] p8_array_index_1085107_comb;
  wire [7:0] p8_res7__634_comb;
  wire [7:0] p8_array_index_1084886_comb;
  wire [7:0] p8_array_index_1084887_comb;
  wire [7:0] p8_array_index_1084888_comb;
  wire [7:0] p8_array_index_1084889_comb;
  wire [7:0] p8_array_index_1084890_comb;
  wire [7:0] p8_array_index_1084891_comb;
  wire [7:0] p8_array_index_1084893_comb;
  wire [7:0] p8_array_index_1084895_comb;
  wire [7:0] p8_array_index_1084896_comb;
  wire [7:0] p8_array_index_1084897_comb;
  wire [7:0] p8_array_index_1084898_comb;
  wire [7:0] p8_array_index_1084899_comb;
  wire [7:0] p8_array_index_1084900_comb;
  wire [7:0] p8_array_index_1085117_comb;
  wire [7:0] p8_array_index_1084902_comb;
  wire [7:0] p8_array_index_1084903_comb;
  wire [7:0] p8_array_index_1084904_comb;
  wire [7:0] p8_array_index_1084905_comb;
  wire [7:0] p8_array_index_1084906_comb;
  wire [7:0] p8_array_index_1084907_comb;
  wire [7:0] p8_array_index_1084908_comb;
  wire [7:0] p8_array_index_1084910_comb;
  wire [7:0] p8_res7__635_comb;
  wire [7:0] p8_res7__464_comb;
  wire [7:0] p8_array_index_1084919_comb;
  wire [7:0] p8_array_index_1084920_comb;
  wire [7:0] p8_array_index_1084921_comb;
  wire [7:0] p8_array_index_1084922_comb;
  wire [7:0] p8_array_index_1084923_comb;
  wire [7:0] p8_array_index_1084924_comb;
  wire [7:0] p8_res7__636_comb;
  wire [7:0] p8_res7__465_comb;
  wire [7:0] p8_array_index_1084934_comb;
  wire [7:0] p8_array_index_1084935_comb;
  wire [7:0] p8_array_index_1084936_comb;
  wire [7:0] p8_array_index_1084937_comb;
  wire [7:0] p8_array_index_1084938_comb;
  wire [7:0] p8_res7__637_comb;
  wire [7:0] p8_res7__466_comb;
  wire [7:0] p8_array_index_1084948_comb;
  wire [7:0] p8_array_index_1084949_comb;
  wire [7:0] p8_array_index_1084950_comb;
  wire [7:0] p8_array_index_1084951_comb;
  wire [7:0] p8_array_index_1084952_comb;
  wire [7:0] p8_res7__638_comb;
  wire [7:0] p8_res7__467_comb;
  wire [7:0] p8_array_index_1084963_comb;
  wire [7:0] p8_array_index_1084964_comb;
  wire [7:0] p8_array_index_1084965_comb;
  wire [7:0] p8_array_index_1084966_comb;
  wire [7:0] p8_res7__639_comb;
  wire [7:0] p8_res7__468_comb;
  wire [127:0] p8_res__39_comb;
  assign p8_res7__410_comb = p7_array_index_1083754 ^ p7_array_index_1083755 ^ p7_array_index_1083756 ^ p7_array_index_1083757 ^ p7_array_index_1083758 ^ p7_array_index_1083759 ^ p7_res7__403 ^ p7_array_index_1083760 ^ p7_res7__401 ^ p7_array_index_1083713 ^ p7_array_index_1083686 ^ p7_array_index_1083657 ^ p7_array_index_1083625 ^ p7_array_index_1083761 ^ p7_array_index_1083762 ^ p7_array_index_1083612;
  assign p8_array_index_1084176_comb = p7_literal_1076355[p7_res7__405];
  assign p8_res7__411_comb = p7_literal_1076345[p8_res7__410_comb] ^ p7_literal_1076347[p7_res7__409] ^ p7_literal_1076349[p7_res7__408] ^ p7_literal_1076351[p7_res7__407] ^ p7_literal_1076353[p7_res7__406] ^ p8_array_index_1084176_comb ^ p7_res7__404 ^ p7_literal_1076358[p7_res7__403] ^ p7_res7__402 ^ p7_array_index_1083725 ^ p7_array_index_1083699 ^ p7_array_index_1083671 ^ p7_array_index_1083642 ^ p7_literal_1076347[p7_array_index_1083609] ^ p7_literal_1076345[p7_array_index_1083610] ^ p7_array_index_1083611;
  assign p8_res7__412_comb = p7_literal_1076345[p8_res7__411_comb] ^ p7_literal_1076347[p8_res7__410_comb] ^ p7_literal_1076349[p7_res7__409] ^ p7_literal_1076351[p7_res7__408] ^ p7_literal_1076353[p7_res7__407] ^ p7_literal_1076355[p7_res7__406] ^ p7_res7__405 ^ p7_literal_1076358[p7_res7__404] ^ p7_res7__403 ^ p7_array_index_1083737 ^ p7_array_index_1083712 ^ p7_array_index_1083685 ^ p7_array_index_1083656 ^ p7_array_index_1083624 ^ p7_literal_1076345[p7_array_index_1083609] ^ p7_array_index_1083610;
  assign p8_res7__413_comb = p7_literal_1076345[p8_res7__412_comb] ^ p7_literal_1076347[p8_res7__411_comb] ^ p7_literal_1076349[p8_res7__410_comb] ^ p7_literal_1076351[p7_res7__409] ^ p7_literal_1076353[p7_res7__408] ^ p7_literal_1076355[p7_res7__407] ^ p7_res7__406 ^ p7_literal_1076358[p7_res7__405] ^ p7_res7__404 ^ p7_array_index_1083748 ^ p7_array_index_1083724 ^ p7_array_index_1083698 ^ p7_array_index_1083670 ^ p7_array_index_1083641 ^ p7_literal_1076345[p7_array_index_1083608] ^ p7_array_index_1083609;
  assign p8_res7__414_comb = p7_literal_1076345[p8_res7__413_comb] ^ p7_literal_1076347[p8_res7__412_comb] ^ p7_literal_1076349[p8_res7__411_comb] ^ p7_literal_1076351[p8_res7__410_comb] ^ p7_literal_1076353[p7_res7__409] ^ p7_literal_1076355[p7_res7__408] ^ p7_res7__407 ^ p7_literal_1076358[p7_res7__406] ^ p7_res7__405 ^ p7_array_index_1083759 ^ p7_array_index_1083736 ^ p7_array_index_1083711 ^ p7_array_index_1083684 ^ p7_array_index_1083655 ^ p7_array_index_1083623 ^ p7_array_index_1083608;
  assign p8_res7__415_comb = p7_literal_1076345[p8_res7__414_comb] ^ p7_literal_1076347[p8_res7__413_comb] ^ p7_literal_1076349[p8_res7__412_comb] ^ p7_literal_1076351[p8_res7__411_comb] ^ p7_literal_1076353[p8_res7__410_comb] ^ p7_literal_1076355[p7_res7__409] ^ p7_res7__408 ^ p7_literal_1076358[p7_res7__407] ^ p7_res7__406 ^ p8_array_index_1084176_comb ^ p7_array_index_1083747 ^ p7_array_index_1083723 ^ p7_array_index_1083697 ^ p7_array_index_1083669 ^ p7_array_index_1083640 ^ p7_array_index_1083607;
  assign p8_res__25_comb = {p8_res7__415_comb, p8_res7__414_comb, p8_res7__413_comb, p8_res7__412_comb, p8_res7__411_comb, p8_res7__410_comb, p7_res7__409, p7_res7__408, p7_res7__407, p7_res7__406, p7_res7__405, p7_res7__404, p7_res7__403, p7_res7__402, p7_res7__401, p7_res7__400};
  assign p8_xor_1084216_comb = p8_res__25_comb ^ p7_k6;
  assign p8_addedKey__67_comb = p8_xor_1084216_comb ^ 128'h6bce_c0ac_5dd7_7453_d3a7_2473_cd72_011b;
  assign p8_array_index_1084232_comb = p7_arr[p8_addedKey__67_comb[127:120]];
  assign p8_array_index_1084233_comb = p7_arr[p8_addedKey__67_comb[119:112]];
  assign p8_array_index_1084234_comb = p7_arr[p8_addedKey__67_comb[111:104]];
  assign p8_array_index_1084235_comb = p7_arr[p8_addedKey__67_comb[103:96]];
  assign p8_array_index_1084236_comb = p7_arr[p8_addedKey__67_comb[95:88]];
  assign p8_array_index_1084237_comb = p7_arr[p8_addedKey__67_comb[87:80]];
  assign p8_array_index_1084239_comb = p7_arr[p8_addedKey__67_comb[71:64]];
  assign p8_array_index_1084241_comb = p7_arr[p8_addedKey__67_comb[55:48]];
  assign p8_array_index_1084242_comb = p7_arr[p8_addedKey__67_comb[47:40]];
  assign p8_array_index_1084243_comb = p7_arr[p8_addedKey__67_comb[39:32]];
  assign p8_array_index_1084244_comb = p7_arr[p8_addedKey__67_comb[31:24]];
  assign p8_array_index_1084245_comb = p7_arr[p8_addedKey__67_comb[23:16]];
  assign p8_array_index_1084246_comb = p7_arr[p8_addedKey__67_comb[15:8]];
  assign p8_array_index_1084248_comb = p7_literal_1076345[p8_array_index_1084232_comb];
  assign p8_array_index_1084249_comb = p7_literal_1076347[p8_array_index_1084233_comb];
  assign p8_array_index_1084250_comb = p7_literal_1076349[p8_array_index_1084234_comb];
  assign p8_array_index_1084251_comb = p7_literal_1076351[p8_array_index_1084235_comb];
  assign p8_array_index_1084252_comb = p7_literal_1076353[p8_array_index_1084236_comb];
  assign p8_array_index_1084253_comb = p7_literal_1076355[p8_array_index_1084237_comb];
  assign p8_array_index_1084254_comb = p7_arr[p8_addedKey__67_comb[79:72]];
  assign p8_array_index_1084256_comb = p7_arr[p8_addedKey__67_comb[63:56]];
  assign p8_res7__416_comb = p8_array_index_1084248_comb ^ p8_array_index_1084249_comb ^ p8_array_index_1084250_comb ^ p8_array_index_1084251_comb ^ p8_array_index_1084252_comb ^ p8_array_index_1084253_comb ^ p8_array_index_1084254_comb ^ p7_literal_1076358[p8_array_index_1084239_comb] ^ p8_array_index_1084256_comb ^ p7_literal_1076355[p8_array_index_1084241_comb] ^ p7_literal_1076353[p8_array_index_1084242_comb] ^ p7_literal_1076351[p8_array_index_1084243_comb] ^ p7_literal_1076349[p8_array_index_1084244_comb] ^ p7_literal_1076347[p8_array_index_1084245_comb] ^ p7_literal_1076345[p8_array_index_1084246_comb] ^ p7_arr[p8_addedKey__67_comb[7:0]];
  assign p8_array_index_1084265_comb = p7_literal_1076345[p8_res7__416_comb];
  assign p8_array_index_1084266_comb = p7_literal_1076347[p8_array_index_1084232_comb];
  assign p8_array_index_1084267_comb = p7_literal_1076349[p8_array_index_1084233_comb];
  assign p8_array_index_1084268_comb = p7_literal_1076351[p8_array_index_1084234_comb];
  assign p8_array_index_1084269_comb = p7_literal_1076353[p8_array_index_1084235_comb];
  assign p8_array_index_1084270_comb = p7_literal_1076355[p8_array_index_1084236_comb];
  assign p8_res7__417_comb = p8_array_index_1084265_comb ^ p8_array_index_1084266_comb ^ p8_array_index_1084267_comb ^ p8_array_index_1084268_comb ^ p8_array_index_1084269_comb ^ p8_array_index_1084270_comb ^ p8_array_index_1084237_comb ^ p7_literal_1076358[p8_array_index_1084254_comb] ^ p8_array_index_1084239_comb ^ p7_literal_1076355[p8_array_index_1084256_comb] ^ p7_literal_1076353[p8_array_index_1084241_comb] ^ p7_literal_1076351[p8_array_index_1084242_comb] ^ p7_literal_1076349[p8_array_index_1084243_comb] ^ p7_literal_1076347[p8_array_index_1084244_comb] ^ p7_literal_1076345[p8_array_index_1084245_comb] ^ p8_array_index_1084246_comb;
  assign p8_array_index_1084280_comb = p7_literal_1076347[p8_res7__416_comb];
  assign p8_array_index_1084281_comb = p7_literal_1076349[p8_array_index_1084232_comb];
  assign p8_array_index_1084282_comb = p7_literal_1076351[p8_array_index_1084233_comb];
  assign p8_array_index_1084283_comb = p7_literal_1076353[p8_array_index_1084234_comb];
  assign p8_array_index_1084284_comb = p7_literal_1076355[p8_array_index_1084235_comb];
  assign p8_res7__418_comb = p7_literal_1076345[p8_res7__417_comb] ^ p8_array_index_1084280_comb ^ p8_array_index_1084281_comb ^ p8_array_index_1084282_comb ^ p8_array_index_1084283_comb ^ p8_array_index_1084284_comb ^ p8_array_index_1084236_comb ^ p7_literal_1076358[p8_array_index_1084237_comb] ^ p8_array_index_1084254_comb ^ p7_literal_1076355[p8_array_index_1084239_comb] ^ p7_literal_1076353[p8_array_index_1084256_comb] ^ p7_literal_1076351[p8_array_index_1084241_comb] ^ p7_literal_1076349[p8_array_index_1084242_comb] ^ p7_literal_1076347[p8_array_index_1084243_comb] ^ p7_literal_1076345[p8_array_index_1084244_comb] ^ p8_array_index_1084245_comb;
  assign p8_array_index_1084294_comb = p7_literal_1076347[p8_res7__417_comb];
  assign p8_array_index_1084295_comb = p7_literal_1076349[p8_res7__416_comb];
  assign p8_array_index_1084296_comb = p7_literal_1076351[p8_array_index_1084232_comb];
  assign p8_array_index_1084297_comb = p7_literal_1076353[p8_array_index_1084233_comb];
  assign p8_array_index_1084298_comb = p7_literal_1076355[p8_array_index_1084234_comb];
  assign p8_res7__419_comb = p7_literal_1076345[p8_res7__418_comb] ^ p8_array_index_1084294_comb ^ p8_array_index_1084295_comb ^ p8_array_index_1084296_comb ^ p8_array_index_1084297_comb ^ p8_array_index_1084298_comb ^ p8_array_index_1084235_comb ^ p7_literal_1076358[p8_array_index_1084236_comb] ^ p8_array_index_1084237_comb ^ p7_literal_1076355[p8_array_index_1084254_comb] ^ p7_literal_1076353[p8_array_index_1084239_comb] ^ p7_literal_1076351[p8_array_index_1084256_comb] ^ p7_literal_1076349[p8_array_index_1084241_comb] ^ p7_literal_1076347[p8_array_index_1084242_comb] ^ p7_literal_1076345[p8_array_index_1084243_comb] ^ p8_array_index_1084244_comb;
  assign p8_array_index_1084309_comb = p7_literal_1076349[p8_res7__417_comb];
  assign p8_array_index_1084310_comb = p7_literal_1076351[p8_res7__416_comb];
  assign p8_array_index_1084311_comb = p7_literal_1076353[p8_array_index_1084232_comb];
  assign p8_array_index_1084312_comb = p7_literal_1076355[p8_array_index_1084233_comb];
  assign p8_res7__420_comb = p7_literal_1076345[p8_res7__419_comb] ^ p7_literal_1076347[p8_res7__418_comb] ^ p8_array_index_1084309_comb ^ p8_array_index_1084310_comb ^ p8_array_index_1084311_comb ^ p8_array_index_1084312_comb ^ p8_array_index_1084234_comb ^ p7_literal_1076358[p8_array_index_1084235_comb] ^ p8_array_index_1084236_comb ^ p8_array_index_1084253_comb ^ p7_literal_1076353[p8_array_index_1084254_comb] ^ p7_literal_1076351[p8_array_index_1084239_comb] ^ p7_literal_1076349[p8_array_index_1084256_comb] ^ p7_literal_1076347[p8_array_index_1084241_comb] ^ p7_literal_1076345[p8_array_index_1084242_comb] ^ p8_array_index_1084243_comb;
  assign p8_array_index_1084322_comb = p7_literal_1076349[p8_res7__418_comb];
  assign p8_array_index_1084323_comb = p7_literal_1076351[p8_res7__417_comb];
  assign p8_array_index_1084324_comb = p7_literal_1076353[p8_res7__416_comb];
  assign p8_array_index_1084325_comb = p7_literal_1076355[p8_array_index_1084232_comb];
  assign p8_res7__421_comb = p7_literal_1076345[p8_res7__420_comb] ^ p7_literal_1076347[p8_res7__419_comb] ^ p8_array_index_1084322_comb ^ p8_array_index_1084323_comb ^ p8_array_index_1084324_comb ^ p8_array_index_1084325_comb ^ p8_array_index_1084233_comb ^ p7_literal_1076358[p8_array_index_1084234_comb] ^ p8_array_index_1084235_comb ^ p8_array_index_1084270_comb ^ p7_literal_1076353[p8_array_index_1084237_comb] ^ p7_literal_1076351[p8_array_index_1084254_comb] ^ p7_literal_1076349[p8_array_index_1084239_comb] ^ p7_literal_1076347[p8_array_index_1084256_comb] ^ p7_literal_1076345[p8_array_index_1084241_comb] ^ p8_array_index_1084242_comb;
  assign p8_array_index_1084336_comb = p7_literal_1076351[p8_res7__418_comb];
  assign p8_array_index_1084337_comb = p7_literal_1076353[p8_res7__417_comb];
  assign p8_array_index_1084338_comb = p7_literal_1076355[p8_res7__416_comb];
  assign p8_res7__422_comb = p7_literal_1076345[p8_res7__421_comb] ^ p7_literal_1076347[p8_res7__420_comb] ^ p7_literal_1076349[p8_res7__419_comb] ^ p8_array_index_1084336_comb ^ p8_array_index_1084337_comb ^ p8_array_index_1084338_comb ^ p8_array_index_1084232_comb ^ p7_literal_1076358[p8_array_index_1084233_comb] ^ p8_array_index_1084234_comb ^ p8_array_index_1084284_comb ^ p8_array_index_1084252_comb ^ p7_literal_1076351[p8_array_index_1084237_comb] ^ p7_literal_1076349[p8_array_index_1084254_comb] ^ p7_literal_1076347[p8_array_index_1084239_comb] ^ p7_literal_1076345[p8_array_index_1084256_comb] ^ p8_array_index_1084241_comb;
  assign p8_array_index_1084348_comb = p7_literal_1076351[p8_res7__419_comb];
  assign p8_array_index_1084349_comb = p7_literal_1076353[p8_res7__418_comb];
  assign p8_array_index_1084350_comb = p7_literal_1076355[p8_res7__417_comb];
  assign p8_res7__423_comb = p7_literal_1076345[p8_res7__422_comb] ^ p7_literal_1076347[p8_res7__421_comb] ^ p7_literal_1076349[p8_res7__420_comb] ^ p8_array_index_1084348_comb ^ p8_array_index_1084349_comb ^ p8_array_index_1084350_comb ^ p8_res7__416_comb ^ p7_literal_1076358[p8_array_index_1084232_comb] ^ p8_array_index_1084233_comb ^ p8_array_index_1084298_comb ^ p8_array_index_1084269_comb ^ p7_literal_1076351[p8_array_index_1084236_comb] ^ p7_literal_1076349[p8_array_index_1084237_comb] ^ p7_literal_1076347[p8_array_index_1084254_comb] ^ p7_literal_1076345[p8_array_index_1084239_comb] ^ p8_array_index_1084256_comb;
  assign p8_array_index_1084361_comb = p7_literal_1076353[p8_res7__419_comb];
  assign p8_array_index_1084362_comb = p7_literal_1076355[p8_res7__418_comb];
  assign p8_res7__424_comb = p7_literal_1076345[p8_res7__423_comb] ^ p7_literal_1076347[p8_res7__422_comb] ^ p7_literal_1076349[p8_res7__421_comb] ^ p7_literal_1076351[p8_res7__420_comb] ^ p8_array_index_1084361_comb ^ p8_array_index_1084362_comb ^ p8_res7__417_comb ^ p7_literal_1076358[p8_res7__416_comb] ^ p8_array_index_1084232_comb ^ p8_array_index_1084312_comb ^ p8_array_index_1084283_comb ^ p8_array_index_1084251_comb ^ p7_literal_1076349[p8_array_index_1084236_comb] ^ p7_literal_1076347[p8_array_index_1084237_comb] ^ p7_literal_1076345[p8_array_index_1084254_comb] ^ p8_array_index_1084239_comb;
  assign p8_array_index_1084372_comb = p7_literal_1076353[p8_res7__420_comb];
  assign p8_array_index_1084373_comb = p7_literal_1076355[p8_res7__419_comb];
  assign p8_res7__425_comb = p7_literal_1076345[p8_res7__424_comb] ^ p7_literal_1076347[p8_res7__423_comb] ^ p7_literal_1076349[p8_res7__422_comb] ^ p7_literal_1076351[p8_res7__421_comb] ^ p8_array_index_1084372_comb ^ p8_array_index_1084373_comb ^ p8_res7__418_comb ^ p7_literal_1076358[p8_res7__417_comb] ^ p8_res7__416_comb ^ p8_array_index_1084325_comb ^ p8_array_index_1084297_comb ^ p8_array_index_1084268_comb ^ p7_literal_1076349[p8_array_index_1084235_comb] ^ p7_literal_1076347[p8_array_index_1084236_comb] ^ p7_literal_1076345[p8_array_index_1084237_comb] ^ p8_array_index_1084254_comb;
  assign p8_array_index_1084384_comb = p7_literal_1076355[p8_res7__420_comb];
  assign p8_res7__426_comb = p7_literal_1076345[p8_res7__425_comb] ^ p7_literal_1076347[p8_res7__424_comb] ^ p7_literal_1076349[p8_res7__423_comb] ^ p7_literal_1076351[p8_res7__422_comb] ^ p7_literal_1076353[p8_res7__421_comb] ^ p8_array_index_1084384_comb ^ p8_res7__419_comb ^ p7_literal_1076358[p8_res7__418_comb] ^ p8_res7__417_comb ^ p8_array_index_1084338_comb ^ p8_array_index_1084311_comb ^ p8_array_index_1084282_comb ^ p8_array_index_1084250_comb ^ p7_literal_1076347[p8_array_index_1084235_comb] ^ p7_literal_1076345[p8_array_index_1084236_comb] ^ p8_array_index_1084237_comb;
  assign p8_array_index_1084394_comb = p7_literal_1076355[p8_res7__421_comb];
  assign p8_res7__427_comb = p7_literal_1076345[p8_res7__426_comb] ^ p7_literal_1076347[p8_res7__425_comb] ^ p7_literal_1076349[p8_res7__424_comb] ^ p7_literal_1076351[p8_res7__423_comb] ^ p7_literal_1076353[p8_res7__422_comb] ^ p8_array_index_1084394_comb ^ p8_res7__420_comb ^ p7_literal_1076358[p8_res7__419_comb] ^ p8_res7__418_comb ^ p8_array_index_1084350_comb ^ p8_array_index_1084324_comb ^ p8_array_index_1084296_comb ^ p8_array_index_1084267_comb ^ p7_literal_1076347[p8_array_index_1084234_comb] ^ p7_literal_1076345[p8_array_index_1084235_comb] ^ p8_array_index_1084236_comb;
  assign p8_res7__428_comb = p7_literal_1076345[p8_res7__427_comb] ^ p7_literal_1076347[p8_res7__426_comb] ^ p7_literal_1076349[p8_res7__425_comb] ^ p7_literal_1076351[p8_res7__424_comb] ^ p7_literal_1076353[p8_res7__423_comb] ^ p7_literal_1076355[p8_res7__422_comb] ^ p8_res7__421_comb ^ p7_literal_1076358[p8_res7__420_comb] ^ p8_res7__419_comb ^ p8_array_index_1084362_comb ^ p8_array_index_1084337_comb ^ p8_array_index_1084310_comb ^ p8_array_index_1084281_comb ^ p8_array_index_1084249_comb ^ p7_literal_1076345[p8_array_index_1084234_comb] ^ p8_array_index_1084235_comb;
  assign p8_res7__429_comb = p7_literal_1076345[p8_res7__428_comb] ^ p7_literal_1076347[p8_res7__427_comb] ^ p7_literal_1076349[p8_res7__426_comb] ^ p7_literal_1076351[p8_res7__425_comb] ^ p7_literal_1076353[p8_res7__424_comb] ^ p7_literal_1076355[p8_res7__423_comb] ^ p8_res7__422_comb ^ p7_literal_1076358[p8_res7__421_comb] ^ p8_res7__420_comb ^ p8_array_index_1084373_comb ^ p8_array_index_1084349_comb ^ p8_array_index_1084323_comb ^ p8_array_index_1084295_comb ^ p8_array_index_1084266_comb ^ p7_literal_1076345[p8_array_index_1084233_comb] ^ p8_array_index_1084234_comb;
  assign p8_res7__430_comb = p7_literal_1076345[p8_res7__429_comb] ^ p7_literal_1076347[p8_res7__428_comb] ^ p7_literal_1076349[p8_res7__427_comb] ^ p7_literal_1076351[p8_res7__426_comb] ^ p7_literal_1076353[p8_res7__425_comb] ^ p7_literal_1076355[p8_res7__424_comb] ^ p8_res7__423_comb ^ p7_literal_1076358[p8_res7__422_comb] ^ p8_res7__421_comb ^ p8_array_index_1084384_comb ^ p8_array_index_1084361_comb ^ p8_array_index_1084336_comb ^ p8_array_index_1084309_comb ^ p8_array_index_1084280_comb ^ p8_array_index_1084248_comb ^ p8_array_index_1084233_comb;
  assign p8_res7__431_comb = p7_literal_1076345[p8_res7__430_comb] ^ p7_literal_1076347[p8_res7__429_comb] ^ p7_literal_1076349[p8_res7__428_comb] ^ p7_literal_1076351[p8_res7__427_comb] ^ p7_literal_1076353[p8_res7__426_comb] ^ p7_literal_1076355[p8_res7__425_comb] ^ p8_res7__424_comb ^ p7_literal_1076358[p8_res7__423_comb] ^ p8_res7__422_comb ^ p8_array_index_1084394_comb ^ p8_array_index_1084372_comb ^ p8_array_index_1084348_comb ^ p8_array_index_1084322_comb ^ p8_array_index_1084294_comb ^ p8_array_index_1084265_comb ^ p8_array_index_1084232_comb;
  assign p8_res__26_comb = {p8_res7__431_comb, p8_res7__430_comb, p8_res7__429_comb, p8_res7__428_comb, p8_res7__427_comb, p8_res7__426_comb, p8_res7__425_comb, p8_res7__424_comb, p8_res7__423_comb, p8_res7__422_comb, p8_res7__421_comb, p8_res7__420_comb, p8_res7__419_comb, p8_res7__418_comb, p8_res7__417_comb, p8_res7__416_comb};
  assign p8_xor_1084434_comb = p8_res__26_comb ^ p7_xor_1083591;
  assign p8_addedKey__68_comb = p8_xor_1084434_comb ^ 128'ha226_4131_9aec_d1fd_8352_9103_9b68_6b1c;
  assign p8_array_index_1084450_comb = p7_arr[p8_addedKey__68_comb[127:120]];
  assign p8_array_index_1084451_comb = p7_arr[p8_addedKey__68_comb[119:112]];
  assign p8_array_index_1084452_comb = p7_arr[p8_addedKey__68_comb[111:104]];
  assign p8_array_index_1084453_comb = p7_arr[p8_addedKey__68_comb[103:96]];
  assign p8_array_index_1084454_comb = p7_arr[p8_addedKey__68_comb[95:88]];
  assign p8_array_index_1084455_comb = p7_arr[p8_addedKey__68_comb[87:80]];
  assign p8_array_index_1084457_comb = p7_arr[p8_addedKey__68_comb[71:64]];
  assign p8_array_index_1084459_comb = p7_arr[p8_addedKey__68_comb[55:48]];
  assign p8_array_index_1084460_comb = p7_arr[p8_addedKey__68_comb[47:40]];
  assign p8_array_index_1084461_comb = p7_arr[p8_addedKey__68_comb[39:32]];
  assign p8_array_index_1084462_comb = p7_arr[p8_addedKey__68_comb[31:24]];
  assign p8_array_index_1084463_comb = p7_arr[p8_addedKey__68_comb[23:16]];
  assign p8_array_index_1084464_comb = p7_arr[p8_addedKey__68_comb[15:8]];
  assign p8_array_index_1084466_comb = p7_literal_1076345[p8_array_index_1084450_comb];
  assign p8_array_index_1084467_comb = p7_literal_1076347[p8_array_index_1084451_comb];
  assign p8_array_index_1084468_comb = p7_literal_1076349[p8_array_index_1084452_comb];
  assign p8_array_index_1084469_comb = p7_literal_1076351[p8_array_index_1084453_comb];
  assign p8_array_index_1084470_comb = p7_literal_1076353[p8_array_index_1084454_comb];
  assign p8_array_index_1084471_comb = p7_literal_1076355[p8_array_index_1084455_comb];
  assign p8_array_index_1084472_comb = p7_arr[p8_addedKey__68_comb[79:72]];
  assign p8_array_index_1084474_comb = p7_arr[p8_addedKey__68_comb[63:56]];
  assign p8_res7__432_comb = p8_array_index_1084466_comb ^ p8_array_index_1084467_comb ^ p8_array_index_1084468_comb ^ p8_array_index_1084469_comb ^ p8_array_index_1084470_comb ^ p8_array_index_1084471_comb ^ p8_array_index_1084472_comb ^ p7_literal_1076358[p8_array_index_1084457_comb] ^ p8_array_index_1084474_comb ^ p7_literal_1076355[p8_array_index_1084459_comb] ^ p7_literal_1076353[p8_array_index_1084460_comb] ^ p7_literal_1076351[p8_array_index_1084461_comb] ^ p7_literal_1076349[p8_array_index_1084462_comb] ^ p7_literal_1076347[p8_array_index_1084463_comb] ^ p7_literal_1076345[p8_array_index_1084464_comb] ^ p7_arr[p8_addedKey__68_comb[7:0]];
  assign p8_array_index_1084483_comb = p7_literal_1076345[p8_res7__432_comb];
  assign p8_array_index_1084484_comb = p7_literal_1076347[p8_array_index_1084450_comb];
  assign p8_array_index_1084485_comb = p7_literal_1076349[p8_array_index_1084451_comb];
  assign p8_array_index_1084486_comb = p7_literal_1076351[p8_array_index_1084452_comb];
  assign p8_array_index_1084487_comb = p7_literal_1076353[p8_array_index_1084453_comb];
  assign p8_array_index_1084488_comb = p7_literal_1076355[p8_array_index_1084454_comb];
  assign p8_res7__433_comb = p8_array_index_1084483_comb ^ p8_array_index_1084484_comb ^ p8_array_index_1084485_comb ^ p8_array_index_1084486_comb ^ p8_array_index_1084487_comb ^ p8_array_index_1084488_comb ^ p8_array_index_1084455_comb ^ p7_literal_1076358[p8_array_index_1084472_comb] ^ p8_array_index_1084457_comb ^ p7_literal_1076355[p8_array_index_1084474_comb] ^ p7_literal_1076353[p8_array_index_1084459_comb] ^ p7_literal_1076351[p8_array_index_1084460_comb] ^ p7_literal_1076349[p8_array_index_1084461_comb] ^ p7_literal_1076347[p8_array_index_1084462_comb] ^ p7_literal_1076345[p8_array_index_1084463_comb] ^ p8_array_index_1084464_comb;
  assign p8_array_index_1084498_comb = p7_literal_1076347[p8_res7__432_comb];
  assign p8_array_index_1084499_comb = p7_literal_1076349[p8_array_index_1084450_comb];
  assign p8_array_index_1084500_comb = p7_literal_1076351[p8_array_index_1084451_comb];
  assign p8_array_index_1084501_comb = p7_literal_1076353[p8_array_index_1084452_comb];
  assign p8_array_index_1084502_comb = p7_literal_1076355[p8_array_index_1084453_comb];
  assign p8_res7__434_comb = p7_literal_1076345[p8_res7__433_comb] ^ p8_array_index_1084498_comb ^ p8_array_index_1084499_comb ^ p8_array_index_1084500_comb ^ p8_array_index_1084501_comb ^ p8_array_index_1084502_comb ^ p8_array_index_1084454_comb ^ p7_literal_1076358[p8_array_index_1084455_comb] ^ p8_array_index_1084472_comb ^ p7_literal_1076355[p8_array_index_1084457_comb] ^ p7_literal_1076353[p8_array_index_1084474_comb] ^ p7_literal_1076351[p8_array_index_1084459_comb] ^ p7_literal_1076349[p8_array_index_1084460_comb] ^ p7_literal_1076347[p8_array_index_1084461_comb] ^ p7_literal_1076345[p8_array_index_1084462_comb] ^ p8_array_index_1084463_comb;
  assign p8_array_index_1084512_comb = p7_literal_1076347[p8_res7__433_comb];
  assign p8_array_index_1084513_comb = p7_literal_1076349[p8_res7__432_comb];
  assign p8_array_index_1084514_comb = p7_literal_1076351[p8_array_index_1084450_comb];
  assign p8_array_index_1084515_comb = p7_literal_1076353[p8_array_index_1084451_comb];
  assign p8_array_index_1084516_comb = p7_literal_1076355[p8_array_index_1084452_comb];
  assign p8_res7__435_comb = p7_literal_1076345[p8_res7__434_comb] ^ p8_array_index_1084512_comb ^ p8_array_index_1084513_comb ^ p8_array_index_1084514_comb ^ p8_array_index_1084515_comb ^ p8_array_index_1084516_comb ^ p8_array_index_1084453_comb ^ p7_literal_1076358[p8_array_index_1084454_comb] ^ p8_array_index_1084455_comb ^ p7_literal_1076355[p8_array_index_1084472_comb] ^ p7_literal_1076353[p8_array_index_1084457_comb] ^ p7_literal_1076351[p8_array_index_1084474_comb] ^ p7_literal_1076349[p8_array_index_1084459_comb] ^ p7_literal_1076347[p8_array_index_1084460_comb] ^ p7_literal_1076345[p8_array_index_1084461_comb] ^ p8_array_index_1084462_comb;
  assign p8_array_index_1084527_comb = p7_literal_1076349[p8_res7__433_comb];
  assign p8_array_index_1084528_comb = p7_literal_1076351[p8_res7__432_comb];
  assign p8_array_index_1084529_comb = p7_literal_1076353[p8_array_index_1084450_comb];
  assign p8_array_index_1084530_comb = p7_literal_1076355[p8_array_index_1084451_comb];
  assign p8_res7__436_comb = p7_literal_1076345[p8_res7__435_comb] ^ p7_literal_1076347[p8_res7__434_comb] ^ p8_array_index_1084527_comb ^ p8_array_index_1084528_comb ^ p8_array_index_1084529_comb ^ p8_array_index_1084530_comb ^ p8_array_index_1084452_comb ^ p7_literal_1076358[p8_array_index_1084453_comb] ^ p8_array_index_1084454_comb ^ p8_array_index_1084471_comb ^ p7_literal_1076353[p8_array_index_1084472_comb] ^ p7_literal_1076351[p8_array_index_1084457_comb] ^ p7_literal_1076349[p8_array_index_1084474_comb] ^ p7_literal_1076347[p8_array_index_1084459_comb] ^ p7_literal_1076345[p8_array_index_1084460_comb] ^ p8_array_index_1084461_comb;
  assign p8_array_index_1084540_comb = p7_literal_1076349[p8_res7__434_comb];
  assign p8_array_index_1084541_comb = p7_literal_1076351[p8_res7__433_comb];
  assign p8_array_index_1084542_comb = p7_literal_1076353[p8_res7__432_comb];
  assign p8_array_index_1084543_comb = p7_literal_1076355[p8_array_index_1084450_comb];
  assign p8_res7__437_comb = p7_literal_1076345[p8_res7__436_comb] ^ p7_literal_1076347[p8_res7__435_comb] ^ p8_array_index_1084540_comb ^ p8_array_index_1084541_comb ^ p8_array_index_1084542_comb ^ p8_array_index_1084543_comb ^ p8_array_index_1084451_comb ^ p7_literal_1076358[p8_array_index_1084452_comb] ^ p8_array_index_1084453_comb ^ p8_array_index_1084488_comb ^ p7_literal_1076353[p8_array_index_1084455_comb] ^ p7_literal_1076351[p8_array_index_1084472_comb] ^ p7_literal_1076349[p8_array_index_1084457_comb] ^ p7_literal_1076347[p8_array_index_1084474_comb] ^ p7_literal_1076345[p8_array_index_1084459_comb] ^ p8_array_index_1084460_comb;
  assign p8_array_index_1084554_comb = p7_literal_1076351[p8_res7__434_comb];
  assign p8_array_index_1084555_comb = p7_literal_1076353[p8_res7__433_comb];
  assign p8_array_index_1084556_comb = p7_literal_1076355[p8_res7__432_comb];
  assign p8_res7__438_comb = p7_literal_1076345[p8_res7__437_comb] ^ p7_literal_1076347[p8_res7__436_comb] ^ p7_literal_1076349[p8_res7__435_comb] ^ p8_array_index_1084554_comb ^ p8_array_index_1084555_comb ^ p8_array_index_1084556_comb ^ p8_array_index_1084450_comb ^ p7_literal_1076358[p8_array_index_1084451_comb] ^ p8_array_index_1084452_comb ^ p8_array_index_1084502_comb ^ p8_array_index_1084470_comb ^ p7_literal_1076351[p8_array_index_1084455_comb] ^ p7_literal_1076349[p8_array_index_1084472_comb] ^ p7_literal_1076347[p8_array_index_1084457_comb] ^ p7_literal_1076345[p8_array_index_1084474_comb] ^ p8_array_index_1084459_comb;
  assign p8_array_index_1084566_comb = p7_literal_1076351[p8_res7__435_comb];
  assign p8_array_index_1084567_comb = p7_literal_1076353[p8_res7__434_comb];
  assign p8_array_index_1084568_comb = p7_literal_1076355[p8_res7__433_comb];
  assign p8_res7__439_comb = p7_literal_1076345[p8_res7__438_comb] ^ p7_literal_1076347[p8_res7__437_comb] ^ p7_literal_1076349[p8_res7__436_comb] ^ p8_array_index_1084566_comb ^ p8_array_index_1084567_comb ^ p8_array_index_1084568_comb ^ p8_res7__432_comb ^ p7_literal_1076358[p8_array_index_1084450_comb] ^ p8_array_index_1084451_comb ^ p8_array_index_1084516_comb ^ p8_array_index_1084487_comb ^ p7_literal_1076351[p8_array_index_1084454_comb] ^ p7_literal_1076349[p8_array_index_1084455_comb] ^ p7_literal_1076347[p8_array_index_1084472_comb] ^ p7_literal_1076345[p8_array_index_1084457_comb] ^ p8_array_index_1084474_comb;
  assign p8_array_index_1084579_comb = p7_literal_1076353[p8_res7__435_comb];
  assign p8_array_index_1084580_comb = p7_literal_1076355[p8_res7__434_comb];
  assign p8_res7__440_comb = p7_literal_1076345[p8_res7__439_comb] ^ p7_literal_1076347[p8_res7__438_comb] ^ p7_literal_1076349[p8_res7__437_comb] ^ p7_literal_1076351[p8_res7__436_comb] ^ p8_array_index_1084579_comb ^ p8_array_index_1084580_comb ^ p8_res7__433_comb ^ p7_literal_1076358[p8_res7__432_comb] ^ p8_array_index_1084450_comb ^ p8_array_index_1084530_comb ^ p8_array_index_1084501_comb ^ p8_array_index_1084469_comb ^ p7_literal_1076349[p8_array_index_1084454_comb] ^ p7_literal_1076347[p8_array_index_1084455_comb] ^ p7_literal_1076345[p8_array_index_1084472_comb] ^ p8_array_index_1084457_comb;
  assign p8_array_index_1084590_comb = p7_literal_1076353[p8_res7__436_comb];
  assign p8_array_index_1084591_comb = p7_literal_1076355[p8_res7__435_comb];
  assign p8_res7__441_comb = p7_literal_1076345[p8_res7__440_comb] ^ p7_literal_1076347[p8_res7__439_comb] ^ p7_literal_1076349[p8_res7__438_comb] ^ p7_literal_1076351[p8_res7__437_comb] ^ p8_array_index_1084590_comb ^ p8_array_index_1084591_comb ^ p8_res7__434_comb ^ p7_literal_1076358[p8_res7__433_comb] ^ p8_res7__432_comb ^ p8_array_index_1084543_comb ^ p8_array_index_1084515_comb ^ p8_array_index_1084486_comb ^ p7_literal_1076349[p8_array_index_1084453_comb] ^ p7_literal_1076347[p8_array_index_1084454_comb] ^ p7_literal_1076345[p8_array_index_1084455_comb] ^ p8_array_index_1084472_comb;
  assign p8_array_index_1084602_comb = p7_literal_1076355[p8_res7__436_comb];
  assign p8_res7__442_comb = p7_literal_1076345[p8_res7__441_comb] ^ p7_literal_1076347[p8_res7__440_comb] ^ p7_literal_1076349[p8_res7__439_comb] ^ p7_literal_1076351[p8_res7__438_comb] ^ p7_literal_1076353[p8_res7__437_comb] ^ p8_array_index_1084602_comb ^ p8_res7__435_comb ^ p7_literal_1076358[p8_res7__434_comb] ^ p8_res7__433_comb ^ p8_array_index_1084556_comb ^ p8_array_index_1084529_comb ^ p8_array_index_1084500_comb ^ p8_array_index_1084468_comb ^ p7_literal_1076347[p8_array_index_1084453_comb] ^ p7_literal_1076345[p8_array_index_1084454_comb] ^ p8_array_index_1084455_comb;
  assign p8_array_index_1084612_comb = p7_literal_1076355[p8_res7__437_comb];
  assign p8_res7__443_comb = p7_literal_1076345[p8_res7__442_comb] ^ p7_literal_1076347[p8_res7__441_comb] ^ p7_literal_1076349[p8_res7__440_comb] ^ p7_literal_1076351[p8_res7__439_comb] ^ p7_literal_1076353[p8_res7__438_comb] ^ p8_array_index_1084612_comb ^ p8_res7__436_comb ^ p7_literal_1076358[p8_res7__435_comb] ^ p8_res7__434_comb ^ p8_array_index_1084568_comb ^ p8_array_index_1084542_comb ^ p8_array_index_1084514_comb ^ p8_array_index_1084485_comb ^ p7_literal_1076347[p8_array_index_1084452_comb] ^ p7_literal_1076345[p8_array_index_1084453_comb] ^ p8_array_index_1084454_comb;
  assign p8_res7__444_comb = p7_literal_1076345[p8_res7__443_comb] ^ p7_literal_1076347[p8_res7__442_comb] ^ p7_literal_1076349[p8_res7__441_comb] ^ p7_literal_1076351[p8_res7__440_comb] ^ p7_literal_1076353[p8_res7__439_comb] ^ p7_literal_1076355[p8_res7__438_comb] ^ p8_res7__437_comb ^ p7_literal_1076358[p8_res7__436_comb] ^ p8_res7__435_comb ^ p8_array_index_1084580_comb ^ p8_array_index_1084555_comb ^ p8_array_index_1084528_comb ^ p8_array_index_1084499_comb ^ p8_array_index_1084467_comb ^ p7_literal_1076345[p8_array_index_1084452_comb] ^ p8_array_index_1084453_comb;
  assign p8_res7__445_comb = p7_literal_1076345[p8_res7__444_comb] ^ p7_literal_1076347[p8_res7__443_comb] ^ p7_literal_1076349[p8_res7__442_comb] ^ p7_literal_1076351[p8_res7__441_comb] ^ p7_literal_1076353[p8_res7__440_comb] ^ p7_literal_1076355[p8_res7__439_comb] ^ p8_res7__438_comb ^ p7_literal_1076358[p8_res7__437_comb] ^ p8_res7__436_comb ^ p8_array_index_1084591_comb ^ p8_array_index_1084567_comb ^ p8_array_index_1084541_comb ^ p8_array_index_1084513_comb ^ p8_array_index_1084484_comb ^ p7_literal_1076345[p8_array_index_1084451_comb] ^ p8_array_index_1084452_comb;
  assign p8_res7__446_comb = p7_literal_1076345[p8_res7__445_comb] ^ p7_literal_1076347[p8_res7__444_comb] ^ p7_literal_1076349[p8_res7__443_comb] ^ p7_literal_1076351[p8_res7__442_comb] ^ p7_literal_1076353[p8_res7__441_comb] ^ p7_literal_1076355[p8_res7__440_comb] ^ p8_res7__439_comb ^ p7_literal_1076358[p8_res7__438_comb] ^ p8_res7__437_comb ^ p8_array_index_1084602_comb ^ p8_array_index_1084579_comb ^ p8_array_index_1084554_comb ^ p8_array_index_1084527_comb ^ p8_array_index_1084498_comb ^ p8_array_index_1084466_comb ^ p8_array_index_1084451_comb;
  assign p8_res7__447_comb = p7_literal_1076345[p8_res7__446_comb] ^ p7_literal_1076347[p8_res7__445_comb] ^ p7_literal_1076349[p8_res7__444_comb] ^ p7_literal_1076351[p8_res7__443_comb] ^ p7_literal_1076353[p8_res7__442_comb] ^ p7_literal_1076355[p8_res7__441_comb] ^ p8_res7__440_comb ^ p7_literal_1076358[p8_res7__439_comb] ^ p8_res7__438_comb ^ p8_array_index_1084612_comb ^ p8_array_index_1084590_comb ^ p8_array_index_1084566_comb ^ p8_array_index_1084540_comb ^ p8_array_index_1084512_comb ^ p8_array_index_1084483_comb ^ p8_array_index_1084450_comb;
  assign p8_res__27_comb = {p8_res7__447_comb, p8_res7__446_comb, p8_res7__445_comb, p8_res7__444_comb, p8_res7__443_comb, p8_res7__442_comb, p8_res7__441_comb, p8_res7__440_comb, p8_res7__439_comb, p8_res7__438_comb, p8_res7__437_comb, p8_res7__436_comb, p8_res7__435_comb, p8_res7__434_comb, p8_res7__433_comb, p8_res7__432_comb};
  assign p8_xor_1084652_comb = p8_res__27_comb ^ p8_xor_1084216_comb;
  assign p8_addedKey__69_comb = p8_xor_1084652_comb ^ 128'hcc84_3743_f6a4_ab45_de75_2c13_46ec_ff1d;
  assign p8_array_index_1084668_comb = p7_arr[p8_addedKey__69_comb[127:120]];
  assign p8_array_index_1084669_comb = p7_arr[p8_addedKey__69_comb[119:112]];
  assign p8_array_index_1084670_comb = p7_arr[p8_addedKey__69_comb[111:104]];
  assign p8_array_index_1084671_comb = p7_arr[p8_addedKey__69_comb[103:96]];
  assign p8_array_index_1084672_comb = p7_arr[p8_addedKey__69_comb[95:88]];
  assign p8_array_index_1084673_comb = p7_arr[p8_addedKey__69_comb[87:80]];
  assign p8_array_index_1084675_comb = p7_arr[p8_addedKey__69_comb[71:64]];
  assign p8_array_index_1084677_comb = p7_arr[p8_addedKey__69_comb[55:48]];
  assign p8_array_index_1084678_comb = p7_arr[p8_addedKey__69_comb[47:40]];
  assign p8_array_index_1084679_comb = p7_arr[p8_addedKey__69_comb[39:32]];
  assign p8_array_index_1084680_comb = p7_arr[p8_addedKey__69_comb[31:24]];
  assign p8_array_index_1084681_comb = p7_arr[p8_addedKey__69_comb[23:16]];
  assign p8_array_index_1084682_comb = p7_arr[p8_addedKey__69_comb[15:8]];
  assign p8_array_index_1084684_comb = p7_literal_1076345[p8_array_index_1084668_comb];
  assign p8_array_index_1084685_comb = p7_literal_1076347[p8_array_index_1084669_comb];
  assign p8_array_index_1084686_comb = p7_literal_1076349[p8_array_index_1084670_comb];
  assign p8_array_index_1084687_comb = p7_literal_1076351[p8_array_index_1084671_comb];
  assign p8_array_index_1084688_comb = p7_literal_1076353[p8_array_index_1084672_comb];
  assign p8_array_index_1084689_comb = p7_literal_1076355[p8_array_index_1084673_comb];
  assign p8_array_index_1084690_comb = p7_arr[p8_addedKey__69_comb[79:72]];
  assign p8_array_index_1084692_comb = p7_arr[p8_addedKey__69_comb[63:56]];
  assign p8_res7__448_comb = p8_array_index_1084684_comb ^ p8_array_index_1084685_comb ^ p8_array_index_1084686_comb ^ p8_array_index_1084687_comb ^ p8_array_index_1084688_comb ^ p8_array_index_1084689_comb ^ p8_array_index_1084690_comb ^ p7_literal_1076358[p8_array_index_1084675_comb] ^ p8_array_index_1084692_comb ^ p7_literal_1076355[p8_array_index_1084677_comb] ^ p7_literal_1076353[p8_array_index_1084678_comb] ^ p7_literal_1076351[p8_array_index_1084679_comb] ^ p7_literal_1076349[p8_array_index_1084680_comb] ^ p7_literal_1076347[p8_array_index_1084681_comb] ^ p7_literal_1076345[p8_array_index_1084682_comb] ^ p7_arr[p8_addedKey__69_comb[7:0]];
  assign p8_array_index_1084701_comb = p7_literal_1076345[p8_res7__448_comb];
  assign p8_array_index_1084702_comb = p7_literal_1076347[p8_array_index_1084668_comb];
  assign p8_array_index_1084703_comb = p7_literal_1076349[p8_array_index_1084669_comb];
  assign p8_array_index_1084704_comb = p7_literal_1076351[p8_array_index_1084670_comb];
  assign p8_array_index_1084705_comb = p7_literal_1076353[p8_array_index_1084671_comb];
  assign p8_array_index_1084706_comb = p7_literal_1076355[p8_array_index_1084672_comb];
  assign p8_res7__449_comb = p8_array_index_1084701_comb ^ p8_array_index_1084702_comb ^ p8_array_index_1084703_comb ^ p8_array_index_1084704_comb ^ p8_array_index_1084705_comb ^ p8_array_index_1084706_comb ^ p8_array_index_1084673_comb ^ p7_literal_1076358[p8_array_index_1084690_comb] ^ p8_array_index_1084675_comb ^ p7_literal_1076355[p8_array_index_1084692_comb] ^ p7_literal_1076353[p8_array_index_1084677_comb] ^ p7_literal_1076351[p8_array_index_1084678_comb] ^ p7_literal_1076349[p8_array_index_1084679_comb] ^ p7_literal_1076347[p8_array_index_1084680_comb] ^ p7_literal_1076345[p8_array_index_1084681_comb] ^ p8_array_index_1084682_comb;
  assign p8_array_index_1084716_comb = p7_literal_1076347[p8_res7__448_comb];
  assign p8_array_index_1084717_comb = p7_literal_1076349[p8_array_index_1084668_comb];
  assign p8_array_index_1084718_comb = p7_literal_1076351[p8_array_index_1084669_comb];
  assign p8_array_index_1084719_comb = p7_literal_1076353[p8_array_index_1084670_comb];
  assign p8_array_index_1084720_comb = p7_literal_1076355[p8_array_index_1084671_comb];
  assign p8_res7__450_comb = p7_literal_1076345[p8_res7__449_comb] ^ p8_array_index_1084716_comb ^ p8_array_index_1084717_comb ^ p8_array_index_1084718_comb ^ p8_array_index_1084719_comb ^ p8_array_index_1084720_comb ^ p8_array_index_1084672_comb ^ p7_literal_1076358[p8_array_index_1084673_comb] ^ p8_array_index_1084690_comb ^ p7_literal_1076355[p8_array_index_1084675_comb] ^ p7_literal_1076353[p8_array_index_1084692_comb] ^ p7_literal_1076351[p8_array_index_1084677_comb] ^ p7_literal_1076349[p8_array_index_1084678_comb] ^ p7_literal_1076347[p8_array_index_1084679_comb] ^ p7_literal_1076345[p8_array_index_1084680_comb] ^ p8_array_index_1084681_comb;
  assign p8_array_index_1084730_comb = p7_literal_1076347[p8_res7__449_comb];
  assign p8_array_index_1084731_comb = p7_literal_1076349[p8_res7__448_comb];
  assign p8_array_index_1084732_comb = p7_literal_1076351[p8_array_index_1084668_comb];
  assign p8_array_index_1084733_comb = p7_literal_1076353[p8_array_index_1084669_comb];
  assign p8_array_index_1084734_comb = p7_literal_1076355[p8_array_index_1084670_comb];
  assign p8_res7__451_comb = p7_literal_1076345[p8_res7__450_comb] ^ p8_array_index_1084730_comb ^ p8_array_index_1084731_comb ^ p8_array_index_1084732_comb ^ p8_array_index_1084733_comb ^ p8_array_index_1084734_comb ^ p8_array_index_1084671_comb ^ p7_literal_1076358[p8_array_index_1084672_comb] ^ p8_array_index_1084673_comb ^ p7_literal_1076355[p8_array_index_1084690_comb] ^ p7_literal_1076353[p8_array_index_1084675_comb] ^ p7_literal_1076351[p8_array_index_1084692_comb] ^ p7_literal_1076349[p8_array_index_1084677_comb] ^ p7_literal_1076347[p8_array_index_1084678_comb] ^ p7_literal_1076345[p8_array_index_1084679_comb] ^ p8_array_index_1084680_comb;
  assign p8_array_index_1084745_comb = p7_literal_1076349[p8_res7__449_comb];
  assign p8_array_index_1084746_comb = p7_literal_1076351[p8_res7__448_comb];
  assign p8_array_index_1084747_comb = p7_literal_1076353[p8_array_index_1084668_comb];
  assign p8_array_index_1084748_comb = p7_literal_1076355[p8_array_index_1084669_comb];
  assign p8_res7__452_comb = p7_literal_1076345[p8_res7__451_comb] ^ p7_literal_1076347[p8_res7__450_comb] ^ p8_array_index_1084745_comb ^ p8_array_index_1084746_comb ^ p8_array_index_1084747_comb ^ p8_array_index_1084748_comb ^ p8_array_index_1084670_comb ^ p7_literal_1076358[p8_array_index_1084671_comb] ^ p8_array_index_1084672_comb ^ p8_array_index_1084689_comb ^ p7_literal_1076353[p8_array_index_1084690_comb] ^ p7_literal_1076351[p8_array_index_1084675_comb] ^ p7_literal_1076349[p8_array_index_1084692_comb] ^ p7_literal_1076347[p8_array_index_1084677_comb] ^ p7_literal_1076345[p8_array_index_1084678_comb] ^ p8_array_index_1084679_comb;
  assign p8_array_index_1084758_comb = p7_literal_1076349[p8_res7__450_comb];
  assign p8_array_index_1084759_comb = p7_literal_1076351[p8_res7__449_comb];
  assign p8_array_index_1084760_comb = p7_literal_1076353[p8_res7__448_comb];
  assign p8_array_index_1084761_comb = p7_literal_1076355[p8_array_index_1084668_comb];
  assign p8_res7__453_comb = p7_literal_1076345[p8_res7__452_comb] ^ p7_literal_1076347[p8_res7__451_comb] ^ p8_array_index_1084758_comb ^ p8_array_index_1084759_comb ^ p8_array_index_1084760_comb ^ p8_array_index_1084761_comb ^ p8_array_index_1084669_comb ^ p7_literal_1076358[p8_array_index_1084670_comb] ^ p8_array_index_1084671_comb ^ p8_array_index_1084706_comb ^ p7_literal_1076353[p8_array_index_1084673_comb] ^ p7_literal_1076351[p8_array_index_1084690_comb] ^ p7_literal_1076349[p8_array_index_1084675_comb] ^ p7_literal_1076347[p8_array_index_1084692_comb] ^ p7_literal_1076345[p8_array_index_1084677_comb] ^ p8_array_index_1084678_comb;
  assign p8_array_index_1084772_comb = p7_literal_1076351[p8_res7__450_comb];
  assign p8_array_index_1084773_comb = p7_literal_1076353[p8_res7__449_comb];
  assign p8_array_index_1084774_comb = p7_literal_1076355[p8_res7__448_comb];
  assign p8_res7__454_comb = p7_literal_1076345[p8_res7__453_comb] ^ p7_literal_1076347[p8_res7__452_comb] ^ p7_literal_1076349[p8_res7__451_comb] ^ p8_array_index_1084772_comb ^ p8_array_index_1084773_comb ^ p8_array_index_1084774_comb ^ p8_array_index_1084668_comb ^ p7_literal_1076358[p8_array_index_1084669_comb] ^ p8_array_index_1084670_comb ^ p8_array_index_1084720_comb ^ p8_array_index_1084688_comb ^ p7_literal_1076351[p8_array_index_1084673_comb] ^ p7_literal_1076349[p8_array_index_1084690_comb] ^ p7_literal_1076347[p8_array_index_1084675_comb] ^ p7_literal_1076345[p8_array_index_1084692_comb] ^ p8_array_index_1084677_comb;
  assign p8_array_index_1084784_comb = p7_literal_1076351[p8_res7__451_comb];
  assign p8_array_index_1084785_comb = p7_literal_1076353[p8_res7__450_comb];
  assign p8_array_index_1084786_comb = p7_literal_1076355[p8_res7__449_comb];
  assign p8_array_index_1084974_comb = p7_literal_1076345[p7_array_index_1083993];
  assign p8_array_index_1084975_comb = p7_literal_1076347[p7_array_index_1083994];
  assign p8_array_index_1084976_comb = p7_literal_1076349[p7_array_index_1083995];
  assign p8_array_index_1084977_comb = p7_literal_1076351[p7_array_index_1083996];
  assign p8_array_index_1084978_comb = p7_literal_1076353[p7_array_index_1083997];
  assign p8_array_index_1084979_comb = p7_literal_1076355[p7_array_index_1083998];
  assign p8_res7__455_comb = p7_literal_1076345[p8_res7__454_comb] ^ p7_literal_1076347[p8_res7__453_comb] ^ p7_literal_1076349[p8_res7__452_comb] ^ p8_array_index_1084784_comb ^ p8_array_index_1084785_comb ^ p8_array_index_1084786_comb ^ p8_res7__448_comb ^ p7_literal_1076358[p8_array_index_1084668_comb] ^ p8_array_index_1084669_comb ^ p8_array_index_1084734_comb ^ p8_array_index_1084705_comb ^ p7_literal_1076351[p8_array_index_1084672_comb] ^ p7_literal_1076349[p8_array_index_1084673_comb] ^ p7_literal_1076347[p8_array_index_1084690_comb] ^ p7_literal_1076345[p8_array_index_1084675_comb] ^ p8_array_index_1084692_comb;
  assign p8_res7__624_comb = p8_array_index_1084974_comb ^ p8_array_index_1084975_comb ^ p8_array_index_1084976_comb ^ p8_array_index_1084977_comb ^ p8_array_index_1084978_comb ^ p8_array_index_1084979_comb ^ p7_array_index_1084009 ^ p7_literal_1076358[p7_array_index_1084000] ^ p7_array_index_1084010 ^ p7_literal_1076355[p7_array_index_1084002] ^ p7_literal_1076353[p7_array_index_1084003] ^ p7_literal_1076351[p7_array_index_1084004] ^ p7_literal_1076349[p7_array_index_1084005] ^ p7_literal_1076347[p7_array_index_1084006] ^ p7_literal_1076345[p7_array_index_1084007] ^ p7_array_index_1084011;
  assign p8_array_index_1084797_comb = p7_literal_1076353[p8_res7__451_comb];
  assign p8_array_index_1084798_comb = p7_literal_1076355[p8_res7__450_comb];
  assign p8_array_index_1084988_comb = p7_literal_1076345[p8_res7__624_comb];
  assign p8_array_index_1084989_comb = p7_literal_1076347[p7_array_index_1083993];
  assign p8_array_index_1084990_comb = p7_literal_1076349[p7_array_index_1083994];
  assign p8_array_index_1084991_comb = p7_literal_1076351[p7_array_index_1083995];
  assign p8_array_index_1084992_comb = p7_literal_1076353[p7_array_index_1083996];
  assign p8_array_index_1084993_comb = p7_literal_1076355[p7_array_index_1083997];
  assign p8_res7__456_comb = p7_literal_1076345[p8_res7__455_comb] ^ p7_literal_1076347[p8_res7__454_comb] ^ p7_literal_1076349[p8_res7__453_comb] ^ p7_literal_1076351[p8_res7__452_comb] ^ p8_array_index_1084797_comb ^ p8_array_index_1084798_comb ^ p8_res7__449_comb ^ p7_literal_1076358[p8_res7__448_comb] ^ p8_array_index_1084668_comb ^ p8_array_index_1084748_comb ^ p8_array_index_1084719_comb ^ p8_array_index_1084687_comb ^ p7_literal_1076349[p8_array_index_1084672_comb] ^ p7_literal_1076347[p8_array_index_1084673_comb] ^ p7_literal_1076345[p8_array_index_1084690_comb] ^ p8_array_index_1084675_comb;
  assign p8_res7__625_comb = p8_array_index_1084988_comb ^ p8_array_index_1084989_comb ^ p8_array_index_1084990_comb ^ p8_array_index_1084991_comb ^ p8_array_index_1084992_comb ^ p8_array_index_1084993_comb ^ p7_array_index_1083998 ^ p7_literal_1076358[p7_array_index_1084009] ^ p7_array_index_1084000 ^ p7_literal_1076355[p7_array_index_1084010] ^ p7_literal_1076353[p7_array_index_1084002] ^ p7_literal_1076351[p7_array_index_1084003] ^ p7_literal_1076349[p7_array_index_1084004] ^ p7_literal_1076347[p7_array_index_1084005] ^ p7_literal_1076345[p7_array_index_1084006] ^ p7_array_index_1084007;
  assign p8_array_index_1084808_comb = p7_literal_1076353[p8_res7__452_comb];
  assign p8_array_index_1084809_comb = p7_literal_1076355[p8_res7__451_comb];
  assign p8_array_index_1085003_comb = p7_literal_1076347[p8_res7__624_comb];
  assign p8_array_index_1085004_comb = p7_literal_1076349[p7_array_index_1083993];
  assign p8_array_index_1085005_comb = p7_literal_1076351[p7_array_index_1083994];
  assign p8_array_index_1085006_comb = p7_literal_1076353[p7_array_index_1083995];
  assign p8_array_index_1085007_comb = p7_literal_1076355[p7_array_index_1083996];
  assign p8_res7__457_comb = p7_literal_1076345[p8_res7__456_comb] ^ p7_literal_1076347[p8_res7__455_comb] ^ p7_literal_1076349[p8_res7__454_comb] ^ p7_literal_1076351[p8_res7__453_comb] ^ p8_array_index_1084808_comb ^ p8_array_index_1084809_comb ^ p8_res7__450_comb ^ p7_literal_1076358[p8_res7__449_comb] ^ p8_res7__448_comb ^ p8_array_index_1084761_comb ^ p8_array_index_1084733_comb ^ p8_array_index_1084704_comb ^ p7_literal_1076349[p8_array_index_1084671_comb] ^ p7_literal_1076347[p8_array_index_1084672_comb] ^ p7_literal_1076345[p8_array_index_1084673_comb] ^ p8_array_index_1084690_comb;
  assign p8_res7__626_comb = p7_literal_1076345[p8_res7__625_comb] ^ p8_array_index_1085003_comb ^ p8_array_index_1085004_comb ^ p8_array_index_1085005_comb ^ p8_array_index_1085006_comb ^ p8_array_index_1085007_comb ^ p7_array_index_1083997 ^ p7_literal_1076358[p7_array_index_1083998] ^ p7_array_index_1084009 ^ p7_literal_1076355[p7_array_index_1084000] ^ p7_literal_1076353[p7_array_index_1084010] ^ p7_literal_1076351[p7_array_index_1084002] ^ p7_literal_1076349[p7_array_index_1084003] ^ p7_literal_1076347[p7_array_index_1084004] ^ p7_literal_1076345[p7_array_index_1084005] ^ p7_array_index_1084006;
  assign p8_array_index_1084820_comb = p7_literal_1076355[p8_res7__452_comb];
  assign p8_array_index_1085017_comb = p7_literal_1076347[p8_res7__625_comb];
  assign p8_array_index_1085018_comb = p7_literal_1076349[p8_res7__624_comb];
  assign p8_array_index_1085019_comb = p7_literal_1076351[p7_array_index_1083993];
  assign p8_array_index_1085020_comb = p7_literal_1076353[p7_array_index_1083994];
  assign p8_array_index_1085021_comb = p7_literal_1076355[p7_array_index_1083995];
  assign p8_res7__458_comb = p7_literal_1076345[p8_res7__457_comb] ^ p7_literal_1076347[p8_res7__456_comb] ^ p7_literal_1076349[p8_res7__455_comb] ^ p7_literal_1076351[p8_res7__454_comb] ^ p7_literal_1076353[p8_res7__453_comb] ^ p8_array_index_1084820_comb ^ p8_res7__451_comb ^ p7_literal_1076358[p8_res7__450_comb] ^ p8_res7__449_comb ^ p8_array_index_1084774_comb ^ p8_array_index_1084747_comb ^ p8_array_index_1084718_comb ^ p8_array_index_1084686_comb ^ p7_literal_1076347[p8_array_index_1084671_comb] ^ p7_literal_1076345[p8_array_index_1084672_comb] ^ p8_array_index_1084673_comb;
  assign p8_res7__627_comb = p7_literal_1076345[p8_res7__626_comb] ^ p8_array_index_1085017_comb ^ p8_array_index_1085018_comb ^ p8_array_index_1085019_comb ^ p8_array_index_1085020_comb ^ p8_array_index_1085021_comb ^ p7_array_index_1083996 ^ p7_literal_1076358[p7_array_index_1083997] ^ p7_array_index_1083998 ^ p7_literal_1076355[p7_array_index_1084009] ^ p7_literal_1076353[p7_array_index_1084000] ^ p7_literal_1076351[p7_array_index_1084010] ^ p7_literal_1076349[p7_array_index_1084002] ^ p7_literal_1076347[p7_array_index_1084003] ^ p7_literal_1076345[p7_array_index_1084004] ^ p7_array_index_1084005;
  assign p8_array_index_1084830_comb = p7_literal_1076355[p8_res7__453_comb];
  assign p8_array_index_1085032_comb = p7_literal_1076349[p8_res7__625_comb];
  assign p8_array_index_1085033_comb = p7_literal_1076351[p8_res7__624_comb];
  assign p8_array_index_1085034_comb = p7_literal_1076353[p7_array_index_1083993];
  assign p8_array_index_1085035_comb = p7_literal_1076355[p7_array_index_1083994];
  assign p8_res7__459_comb = p7_literal_1076345[p8_res7__458_comb] ^ p7_literal_1076347[p8_res7__457_comb] ^ p7_literal_1076349[p8_res7__456_comb] ^ p7_literal_1076351[p8_res7__455_comb] ^ p7_literal_1076353[p8_res7__454_comb] ^ p8_array_index_1084830_comb ^ p8_res7__452_comb ^ p7_literal_1076358[p8_res7__451_comb] ^ p8_res7__450_comb ^ p8_array_index_1084786_comb ^ p8_array_index_1084760_comb ^ p8_array_index_1084732_comb ^ p8_array_index_1084703_comb ^ p7_literal_1076347[p8_array_index_1084670_comb] ^ p7_literal_1076345[p8_array_index_1084671_comb] ^ p8_array_index_1084672_comb;
  assign p8_res7__628_comb = p7_literal_1076345[p8_res7__627_comb] ^ p7_literal_1076347[p8_res7__626_comb] ^ p8_array_index_1085032_comb ^ p8_array_index_1085033_comb ^ p8_array_index_1085034_comb ^ p8_array_index_1085035_comb ^ p7_array_index_1083995 ^ p7_literal_1076358[p7_array_index_1083996] ^ p7_array_index_1083997 ^ p8_array_index_1084979_comb ^ p7_literal_1076353[p7_array_index_1084009] ^ p7_literal_1076351[p7_array_index_1084000] ^ p7_literal_1076349[p7_array_index_1084010] ^ p7_literal_1076347[p7_array_index_1084002] ^ p7_literal_1076345[p7_array_index_1084003] ^ p7_array_index_1084004;
  assign p8_array_index_1085045_comb = p7_literal_1076349[p8_res7__626_comb];
  assign p8_array_index_1085046_comb = p7_literal_1076351[p8_res7__625_comb];
  assign p8_array_index_1085047_comb = p7_literal_1076353[p8_res7__624_comb];
  assign p8_array_index_1085048_comb = p7_literal_1076355[p7_array_index_1083993];
  assign p8_res7__460_comb = p7_literal_1076345[p8_res7__459_comb] ^ p7_literal_1076347[p8_res7__458_comb] ^ p7_literal_1076349[p8_res7__457_comb] ^ p7_literal_1076351[p8_res7__456_comb] ^ p7_literal_1076353[p8_res7__455_comb] ^ p7_literal_1076355[p8_res7__454_comb] ^ p8_res7__453_comb ^ p7_literal_1076358[p8_res7__452_comb] ^ p8_res7__451_comb ^ p8_array_index_1084798_comb ^ p8_array_index_1084773_comb ^ p8_array_index_1084746_comb ^ p8_array_index_1084717_comb ^ p8_array_index_1084685_comb ^ p7_literal_1076345[p8_array_index_1084670_comb] ^ p8_array_index_1084671_comb;
  assign p8_res7__629_comb = p7_literal_1076345[p8_res7__628_comb] ^ p7_literal_1076347[p8_res7__627_comb] ^ p8_array_index_1085045_comb ^ p8_array_index_1085046_comb ^ p8_array_index_1085047_comb ^ p8_array_index_1085048_comb ^ p7_array_index_1083994 ^ p7_literal_1076358[p7_array_index_1083995] ^ p7_array_index_1083996 ^ p8_array_index_1084993_comb ^ p7_literal_1076353[p7_array_index_1083998] ^ p7_literal_1076351[p7_array_index_1084009] ^ p7_literal_1076349[p7_array_index_1084000] ^ p7_literal_1076347[p7_array_index_1084010] ^ p7_literal_1076345[p7_array_index_1084002] ^ p7_array_index_1084003;
  assign p8_array_index_1085059_comb = p7_literal_1076351[p8_res7__626_comb];
  assign p8_array_index_1085060_comb = p7_literal_1076353[p8_res7__625_comb];
  assign p8_array_index_1085061_comb = p7_literal_1076355[p8_res7__624_comb];
  assign p8_res7__461_comb = p7_literal_1076345[p8_res7__460_comb] ^ p7_literal_1076347[p8_res7__459_comb] ^ p7_literal_1076349[p8_res7__458_comb] ^ p7_literal_1076351[p8_res7__457_comb] ^ p7_literal_1076353[p8_res7__456_comb] ^ p7_literal_1076355[p8_res7__455_comb] ^ p8_res7__454_comb ^ p7_literal_1076358[p8_res7__453_comb] ^ p8_res7__452_comb ^ p8_array_index_1084809_comb ^ p8_array_index_1084785_comb ^ p8_array_index_1084759_comb ^ p8_array_index_1084731_comb ^ p8_array_index_1084702_comb ^ p7_literal_1076345[p8_array_index_1084669_comb] ^ p8_array_index_1084670_comb;
  assign p8_res7__630_comb = p7_literal_1076345[p8_res7__629_comb] ^ p7_literal_1076347[p8_res7__628_comb] ^ p7_literal_1076349[p8_res7__627_comb] ^ p8_array_index_1085059_comb ^ p8_array_index_1085060_comb ^ p8_array_index_1085061_comb ^ p7_array_index_1083993 ^ p7_literal_1076358[p7_array_index_1083994] ^ p7_array_index_1083995 ^ p8_array_index_1085007_comb ^ p8_array_index_1084978_comb ^ p7_literal_1076351[p7_array_index_1083998] ^ p7_literal_1076349[p7_array_index_1084009] ^ p7_literal_1076347[p7_array_index_1084000] ^ p7_literal_1076345[p7_array_index_1084010] ^ p7_array_index_1084002;
  assign p8_array_index_1085071_comb = p7_literal_1076351[p8_res7__627_comb];
  assign p8_array_index_1085072_comb = p7_literal_1076353[p8_res7__626_comb];
  assign p8_array_index_1085073_comb = p7_literal_1076355[p8_res7__625_comb];
  assign p8_res7__462_comb = p7_literal_1076345[p8_res7__461_comb] ^ p7_literal_1076347[p8_res7__460_comb] ^ p7_literal_1076349[p8_res7__459_comb] ^ p7_literal_1076351[p8_res7__458_comb] ^ p7_literal_1076353[p8_res7__457_comb] ^ p7_literal_1076355[p8_res7__456_comb] ^ p8_res7__455_comb ^ p7_literal_1076358[p8_res7__454_comb] ^ p8_res7__453_comb ^ p8_array_index_1084820_comb ^ p8_array_index_1084797_comb ^ p8_array_index_1084772_comb ^ p8_array_index_1084745_comb ^ p8_array_index_1084716_comb ^ p8_array_index_1084684_comb ^ p8_array_index_1084669_comb;
  assign p8_res7__631_comb = p7_literal_1076345[p8_res7__630_comb] ^ p7_literal_1076347[p8_res7__629_comb] ^ p7_literal_1076349[p8_res7__628_comb] ^ p8_array_index_1085071_comb ^ p8_array_index_1085072_comb ^ p8_array_index_1085073_comb ^ p8_res7__624_comb ^ p7_literal_1076358[p7_array_index_1083993] ^ p7_array_index_1083994 ^ p8_array_index_1085021_comb ^ p8_array_index_1084992_comb ^ p7_literal_1076351[p7_array_index_1083997] ^ p7_literal_1076349[p7_array_index_1083998] ^ p7_literal_1076347[p7_array_index_1084009] ^ p7_literal_1076345[p7_array_index_1084000] ^ p7_array_index_1084010;
  assign p8_array_index_1085084_comb = p7_literal_1076353[p8_res7__627_comb];
  assign p8_array_index_1085085_comb = p7_literal_1076355[p8_res7__626_comb];
  assign p8_res7__463_comb = p7_literal_1076345[p8_res7__462_comb] ^ p7_literal_1076347[p8_res7__461_comb] ^ p7_literal_1076349[p8_res7__460_comb] ^ p7_literal_1076351[p8_res7__459_comb] ^ p7_literal_1076353[p8_res7__458_comb] ^ p7_literal_1076355[p8_res7__457_comb] ^ p8_res7__456_comb ^ p7_literal_1076358[p8_res7__455_comb] ^ p8_res7__454_comb ^ p8_array_index_1084830_comb ^ p8_array_index_1084808_comb ^ p8_array_index_1084784_comb ^ p8_array_index_1084758_comb ^ p8_array_index_1084730_comb ^ p8_array_index_1084701_comb ^ p8_array_index_1084668_comb;
  assign p8_res7__632_comb = p7_literal_1076345[p8_res7__631_comb] ^ p7_literal_1076347[p8_res7__630_comb] ^ p7_literal_1076349[p8_res7__629_comb] ^ p7_literal_1076351[p8_res7__628_comb] ^ p8_array_index_1085084_comb ^ p8_array_index_1085085_comb ^ p8_res7__625_comb ^ p7_literal_1076358[p8_res7__624_comb] ^ p7_array_index_1083993 ^ p8_array_index_1085035_comb ^ p8_array_index_1085006_comb ^ p8_array_index_1084977_comb ^ p7_literal_1076349[p7_array_index_1083997] ^ p7_literal_1076347[p7_array_index_1083998] ^ p7_literal_1076345[p7_array_index_1084009] ^ p7_array_index_1084000;
  assign p8_res__28_comb = {p8_res7__463_comb, p8_res7__462_comb, p8_res7__461_comb, p8_res7__460_comb, p8_res7__459_comb, p8_res7__458_comb, p8_res7__457_comb, p8_res7__456_comb, p8_res7__455_comb, p8_res7__454_comb, p8_res7__453_comb, p8_res7__452_comb, p8_res7__451_comb, p8_res7__450_comb, p8_res7__449_comb, p8_res7__448_comb};
  assign p8_array_index_1085095_comb = p7_literal_1076353[p8_res7__628_comb];
  assign p8_array_index_1085096_comb = p7_literal_1076355[p8_res7__627_comb];
  assign p8_xor_1084870_comb = p8_res__28_comb ^ p8_xor_1084434_comb;
  assign p8_res7__633_comb = p7_literal_1076345[p8_res7__632_comb] ^ p7_literal_1076347[p8_res7__631_comb] ^ p7_literal_1076349[p8_res7__630_comb] ^ p7_literal_1076351[p8_res7__629_comb] ^ p8_array_index_1085095_comb ^ p8_array_index_1085096_comb ^ p8_res7__626_comb ^ p7_literal_1076358[p8_res7__625_comb] ^ p8_res7__624_comb ^ p8_array_index_1085048_comb ^ p8_array_index_1085020_comb ^ p8_array_index_1084991_comb ^ p7_literal_1076349[p7_array_index_1083996] ^ p7_literal_1076347[p7_array_index_1083997] ^ p7_literal_1076345[p7_array_index_1083998] ^ p7_array_index_1084009;
  assign p8_addedKey__70_comb = p8_xor_1084870_comb ^ 128'h7ea1_add5_427c_254e_391c_2823_e2a3_801e;
  assign p8_array_index_1085107_comb = p7_literal_1076355[p8_res7__628_comb];
  assign p8_res7__634_comb = p7_literal_1076345[p8_res7__633_comb] ^ p7_literal_1076347[p8_res7__632_comb] ^ p7_literal_1076349[p8_res7__631_comb] ^ p7_literal_1076351[p8_res7__630_comb] ^ p7_literal_1076353[p8_res7__629_comb] ^ p8_array_index_1085107_comb ^ p8_res7__627_comb ^ p7_literal_1076358[p8_res7__626_comb] ^ p8_res7__625_comb ^ p8_array_index_1085061_comb ^ p8_array_index_1085034_comb ^ p8_array_index_1085005_comb ^ p8_array_index_1084976_comb ^ p7_literal_1076347[p7_array_index_1083996] ^ p7_literal_1076345[p7_array_index_1083997] ^ p7_array_index_1083998;
  assign p8_array_index_1084886_comb = p7_arr[p8_addedKey__70_comb[127:120]];
  assign p8_array_index_1084887_comb = p7_arr[p8_addedKey__70_comb[119:112]];
  assign p8_array_index_1084888_comb = p7_arr[p8_addedKey__70_comb[111:104]];
  assign p8_array_index_1084889_comb = p7_arr[p8_addedKey__70_comb[103:96]];
  assign p8_array_index_1084890_comb = p7_arr[p8_addedKey__70_comb[95:88]];
  assign p8_array_index_1084891_comb = p7_arr[p8_addedKey__70_comb[87:80]];
  assign p8_array_index_1084893_comb = p7_arr[p8_addedKey__70_comb[71:64]];
  assign p8_array_index_1084895_comb = p7_arr[p8_addedKey__70_comb[55:48]];
  assign p8_array_index_1084896_comb = p7_arr[p8_addedKey__70_comb[47:40]];
  assign p8_array_index_1084897_comb = p7_arr[p8_addedKey__70_comb[39:32]];
  assign p8_array_index_1084898_comb = p7_arr[p8_addedKey__70_comb[31:24]];
  assign p8_array_index_1084899_comb = p7_arr[p8_addedKey__70_comb[23:16]];
  assign p8_array_index_1084900_comb = p7_arr[p8_addedKey__70_comb[15:8]];
  assign p8_array_index_1085117_comb = p7_literal_1076355[p8_res7__629_comb];
  assign p8_array_index_1084902_comb = p7_literal_1076345[p8_array_index_1084886_comb];
  assign p8_array_index_1084903_comb = p7_literal_1076347[p8_array_index_1084887_comb];
  assign p8_array_index_1084904_comb = p7_literal_1076349[p8_array_index_1084888_comb];
  assign p8_array_index_1084905_comb = p7_literal_1076351[p8_array_index_1084889_comb];
  assign p8_array_index_1084906_comb = p7_literal_1076353[p8_array_index_1084890_comb];
  assign p8_array_index_1084907_comb = p7_literal_1076355[p8_array_index_1084891_comb];
  assign p8_array_index_1084908_comb = p7_arr[p8_addedKey__70_comb[79:72]];
  assign p8_array_index_1084910_comb = p7_arr[p8_addedKey__70_comb[63:56]];
  assign p8_res7__635_comb = p7_literal_1076345[p8_res7__634_comb] ^ p7_literal_1076347[p8_res7__633_comb] ^ p7_literal_1076349[p8_res7__632_comb] ^ p7_literal_1076351[p8_res7__631_comb] ^ p7_literal_1076353[p8_res7__630_comb] ^ p8_array_index_1085117_comb ^ p8_res7__628_comb ^ p7_literal_1076358[p8_res7__627_comb] ^ p8_res7__626_comb ^ p8_array_index_1085073_comb ^ p8_array_index_1085047_comb ^ p8_array_index_1085019_comb ^ p8_array_index_1084990_comb ^ p7_literal_1076347[p7_array_index_1083995] ^ p7_literal_1076345[p7_array_index_1083996] ^ p7_array_index_1083997;
  assign p8_res7__464_comb = p8_array_index_1084902_comb ^ p8_array_index_1084903_comb ^ p8_array_index_1084904_comb ^ p8_array_index_1084905_comb ^ p8_array_index_1084906_comb ^ p8_array_index_1084907_comb ^ p8_array_index_1084908_comb ^ p7_literal_1076358[p8_array_index_1084893_comb] ^ p8_array_index_1084910_comb ^ p7_literal_1076355[p8_array_index_1084895_comb] ^ p7_literal_1076353[p8_array_index_1084896_comb] ^ p7_literal_1076351[p8_array_index_1084897_comb] ^ p7_literal_1076349[p8_array_index_1084898_comb] ^ p7_literal_1076347[p8_array_index_1084899_comb] ^ p7_literal_1076345[p8_array_index_1084900_comb] ^ p7_arr[p8_addedKey__70_comb[7:0]];
  assign p8_array_index_1084919_comb = p7_literal_1076345[p8_res7__464_comb];
  assign p8_array_index_1084920_comb = p7_literal_1076347[p8_array_index_1084886_comb];
  assign p8_array_index_1084921_comb = p7_literal_1076349[p8_array_index_1084887_comb];
  assign p8_array_index_1084922_comb = p7_literal_1076351[p8_array_index_1084888_comb];
  assign p8_array_index_1084923_comb = p7_literal_1076353[p8_array_index_1084889_comb];
  assign p8_array_index_1084924_comb = p7_literal_1076355[p8_array_index_1084890_comb];
  assign p8_res7__636_comb = p7_literal_1076345[p8_res7__635_comb] ^ p7_literal_1076347[p8_res7__634_comb] ^ p7_literal_1076349[p8_res7__633_comb] ^ p7_literal_1076351[p8_res7__632_comb] ^ p7_literal_1076353[p8_res7__631_comb] ^ p7_literal_1076355[p8_res7__630_comb] ^ p8_res7__629_comb ^ p7_literal_1076358[p8_res7__628_comb] ^ p8_res7__627_comb ^ p8_array_index_1085085_comb ^ p8_array_index_1085060_comb ^ p8_array_index_1085033_comb ^ p8_array_index_1085004_comb ^ p8_array_index_1084975_comb ^ p7_literal_1076345[p7_array_index_1083995] ^ p7_array_index_1083996;
  assign p8_res7__465_comb = p8_array_index_1084919_comb ^ p8_array_index_1084920_comb ^ p8_array_index_1084921_comb ^ p8_array_index_1084922_comb ^ p8_array_index_1084923_comb ^ p8_array_index_1084924_comb ^ p8_array_index_1084891_comb ^ p7_literal_1076358[p8_array_index_1084908_comb] ^ p8_array_index_1084893_comb ^ p7_literal_1076355[p8_array_index_1084910_comb] ^ p7_literal_1076353[p8_array_index_1084895_comb] ^ p7_literal_1076351[p8_array_index_1084896_comb] ^ p7_literal_1076349[p8_array_index_1084897_comb] ^ p7_literal_1076347[p8_array_index_1084898_comb] ^ p7_literal_1076345[p8_array_index_1084899_comb] ^ p8_array_index_1084900_comb;
  assign p8_array_index_1084934_comb = p7_literal_1076347[p8_res7__464_comb];
  assign p8_array_index_1084935_comb = p7_literal_1076349[p8_array_index_1084886_comb];
  assign p8_array_index_1084936_comb = p7_literal_1076351[p8_array_index_1084887_comb];
  assign p8_array_index_1084937_comb = p7_literal_1076353[p8_array_index_1084888_comb];
  assign p8_array_index_1084938_comb = p7_literal_1076355[p8_array_index_1084889_comb];
  assign p8_res7__637_comb = p7_literal_1076345[p8_res7__636_comb] ^ p7_literal_1076347[p8_res7__635_comb] ^ p7_literal_1076349[p8_res7__634_comb] ^ p7_literal_1076351[p8_res7__633_comb] ^ p7_literal_1076353[p8_res7__632_comb] ^ p7_literal_1076355[p8_res7__631_comb] ^ p8_res7__630_comb ^ p7_literal_1076358[p8_res7__629_comb] ^ p8_res7__628_comb ^ p8_array_index_1085096_comb ^ p8_array_index_1085072_comb ^ p8_array_index_1085046_comb ^ p8_array_index_1085018_comb ^ p8_array_index_1084989_comb ^ p7_literal_1076345[p7_array_index_1083994] ^ p7_array_index_1083995;
  assign p8_res7__466_comb = p7_literal_1076345[p8_res7__465_comb] ^ p8_array_index_1084934_comb ^ p8_array_index_1084935_comb ^ p8_array_index_1084936_comb ^ p8_array_index_1084937_comb ^ p8_array_index_1084938_comb ^ p8_array_index_1084890_comb ^ p7_literal_1076358[p8_array_index_1084891_comb] ^ p8_array_index_1084908_comb ^ p7_literal_1076355[p8_array_index_1084893_comb] ^ p7_literal_1076353[p8_array_index_1084910_comb] ^ p7_literal_1076351[p8_array_index_1084895_comb] ^ p7_literal_1076349[p8_array_index_1084896_comb] ^ p7_literal_1076347[p8_array_index_1084897_comb] ^ p7_literal_1076345[p8_array_index_1084898_comb] ^ p8_array_index_1084899_comb;
  assign p8_array_index_1084948_comb = p7_literal_1076347[p8_res7__465_comb];
  assign p8_array_index_1084949_comb = p7_literal_1076349[p8_res7__464_comb];
  assign p8_array_index_1084950_comb = p7_literal_1076351[p8_array_index_1084886_comb];
  assign p8_array_index_1084951_comb = p7_literal_1076353[p8_array_index_1084887_comb];
  assign p8_array_index_1084952_comb = p7_literal_1076355[p8_array_index_1084888_comb];
  assign p8_res7__638_comb = p7_literal_1076345[p8_res7__637_comb] ^ p7_literal_1076347[p8_res7__636_comb] ^ p7_literal_1076349[p8_res7__635_comb] ^ p7_literal_1076351[p8_res7__634_comb] ^ p7_literal_1076353[p8_res7__633_comb] ^ p7_literal_1076355[p8_res7__632_comb] ^ p8_res7__631_comb ^ p7_literal_1076358[p8_res7__630_comb] ^ p8_res7__629_comb ^ p8_array_index_1085107_comb ^ p8_array_index_1085084_comb ^ p8_array_index_1085059_comb ^ p8_array_index_1085032_comb ^ p8_array_index_1085003_comb ^ p8_array_index_1084974_comb ^ p7_array_index_1083994;
  assign p8_res7__467_comb = p7_literal_1076345[p8_res7__466_comb] ^ p8_array_index_1084948_comb ^ p8_array_index_1084949_comb ^ p8_array_index_1084950_comb ^ p8_array_index_1084951_comb ^ p8_array_index_1084952_comb ^ p8_array_index_1084889_comb ^ p7_literal_1076358[p8_array_index_1084890_comb] ^ p8_array_index_1084891_comb ^ p7_literal_1076355[p8_array_index_1084908_comb] ^ p7_literal_1076353[p8_array_index_1084893_comb] ^ p7_literal_1076351[p8_array_index_1084910_comb] ^ p7_literal_1076349[p8_array_index_1084895_comb] ^ p7_literal_1076347[p8_array_index_1084896_comb] ^ p7_literal_1076345[p8_array_index_1084897_comb] ^ p8_array_index_1084898_comb;
  assign p8_array_index_1084963_comb = p7_literal_1076349[p8_res7__465_comb];
  assign p8_array_index_1084964_comb = p7_literal_1076351[p8_res7__464_comb];
  assign p8_array_index_1084965_comb = p7_literal_1076353[p8_array_index_1084886_comb];
  assign p8_array_index_1084966_comb = p7_literal_1076355[p8_array_index_1084887_comb];
  assign p8_res7__639_comb = p7_literal_1076345[p8_res7__638_comb] ^ p7_literal_1076347[p8_res7__637_comb] ^ p7_literal_1076349[p8_res7__636_comb] ^ p7_literal_1076351[p8_res7__635_comb] ^ p7_literal_1076353[p8_res7__634_comb] ^ p7_literal_1076355[p8_res7__633_comb] ^ p8_res7__632_comb ^ p7_literal_1076358[p8_res7__631_comb] ^ p8_res7__630_comb ^ p8_array_index_1085117_comb ^ p8_array_index_1085095_comb ^ p8_array_index_1085071_comb ^ p8_array_index_1085045_comb ^ p8_array_index_1085017_comb ^ p8_array_index_1084988_comb ^ p7_array_index_1083993;
  assign p8_res7__468_comb = p7_literal_1076345[p8_res7__467_comb] ^ p7_literal_1076347[p8_res7__466_comb] ^ p8_array_index_1084963_comb ^ p8_array_index_1084964_comb ^ p8_array_index_1084965_comb ^ p8_array_index_1084966_comb ^ p8_array_index_1084888_comb ^ p7_literal_1076358[p8_array_index_1084889_comb] ^ p8_array_index_1084890_comb ^ p8_array_index_1084907_comb ^ p7_literal_1076353[p8_array_index_1084908_comb] ^ p7_literal_1076351[p8_array_index_1084893_comb] ^ p7_literal_1076349[p8_array_index_1084910_comb] ^ p7_literal_1076347[p8_array_index_1084895_comb] ^ p7_literal_1076345[p8_array_index_1084896_comb] ^ p8_array_index_1084897_comb;
  assign p8_res__39_comb = {p8_res7__639_comb, p8_res7__638_comb, p8_res7__637_comb, p8_res7__636_comb, p8_res7__635_comb, p8_res7__634_comb, p8_res7__633_comb, p8_res7__632_comb, p8_res7__631_comb, p8_res7__630_comb, p8_res7__629_comb, p8_res7__628_comb, p8_res7__627_comb, p8_res7__626_comb, p8_res7__625_comb, p8_res7__624_comb};

  // Registers for pipe stage 8:
  reg [127:0] p8_xor_1084652;
  reg [127:0] p8_xor_1084870;
  reg [7:0] p8_array_index_1084886;
  reg [7:0] p8_array_index_1084887;
  reg [7:0] p8_array_index_1084888;
  reg [7:0] p8_array_index_1084889;
  reg [7:0] p8_array_index_1084890;
  reg [7:0] p8_array_index_1084891;
  reg [7:0] p8_array_index_1084893;
  reg [7:0] p8_array_index_1084895;
  reg [7:0] p8_array_index_1084896;
  reg [7:0] p8_array_index_1084902;
  reg [7:0] p8_array_index_1084903;
  reg [7:0] p8_array_index_1084904;
  reg [7:0] p8_array_index_1084905;
  reg [7:0] p8_array_index_1084906;
  reg [7:0] p8_array_index_1084908;
  reg [7:0] p8_array_index_1084910;
  reg [7:0] p8_res7__464;
  reg [7:0] p8_array_index_1084919;
  reg [7:0] p8_array_index_1084920;
  reg [7:0] p8_array_index_1084921;
  reg [7:0] p8_array_index_1084922;
  reg [7:0] p8_array_index_1084923;
  reg [7:0] p8_array_index_1084924;
  reg [7:0] p8_res7__465;
  reg [7:0] p8_array_index_1084934;
  reg [7:0] p8_array_index_1084935;
  reg [7:0] p8_array_index_1084936;
  reg [7:0] p8_array_index_1084937;
  reg [7:0] p8_array_index_1084938;
  reg [7:0] p8_res7__466;
  reg [7:0] p8_array_index_1084948;
  reg [7:0] p8_array_index_1084949;
  reg [7:0] p8_array_index_1084950;
  reg [7:0] p8_array_index_1084951;
  reg [7:0] p8_array_index_1084952;
  reg [7:0] p8_res7__467;
  reg [7:0] p8_array_index_1084963;
  reg [7:0] p8_array_index_1084964;
  reg [7:0] p8_array_index_1084965;
  reg [7:0] p8_array_index_1084966;
  reg [7:0] p8_res7__468;
  reg [127:0] p8_res__39;
  always_ff @ (posedge clk) begin
    p8_xor_1084652 <= p8_xor_1084652_comb;
    p8_xor_1084870 <= p8_xor_1084870_comb;
    p8_array_index_1084886 <= p8_array_index_1084886_comb;
    p8_array_index_1084887 <= p8_array_index_1084887_comb;
    p8_array_index_1084888 <= p8_array_index_1084888_comb;
    p8_array_index_1084889 <= p8_array_index_1084889_comb;
    p8_array_index_1084890 <= p8_array_index_1084890_comb;
    p8_array_index_1084891 <= p8_array_index_1084891_comb;
    p8_array_index_1084893 <= p8_array_index_1084893_comb;
    p8_array_index_1084895 <= p8_array_index_1084895_comb;
    p8_array_index_1084896 <= p8_array_index_1084896_comb;
    p8_array_index_1084902 <= p8_array_index_1084902_comb;
    p8_array_index_1084903 <= p8_array_index_1084903_comb;
    p8_array_index_1084904 <= p8_array_index_1084904_comb;
    p8_array_index_1084905 <= p8_array_index_1084905_comb;
    p8_array_index_1084906 <= p8_array_index_1084906_comb;
    p8_array_index_1084908 <= p8_array_index_1084908_comb;
    p8_array_index_1084910 <= p8_array_index_1084910_comb;
    p8_res7__464 <= p8_res7__464_comb;
    p8_array_index_1084919 <= p8_array_index_1084919_comb;
    p8_array_index_1084920 <= p8_array_index_1084920_comb;
    p8_array_index_1084921 <= p8_array_index_1084921_comb;
    p8_array_index_1084922 <= p8_array_index_1084922_comb;
    p8_array_index_1084923 <= p8_array_index_1084923_comb;
    p8_array_index_1084924 <= p8_array_index_1084924_comb;
    p8_res7__465 <= p8_res7__465_comb;
    p8_array_index_1084934 <= p8_array_index_1084934_comb;
    p8_array_index_1084935 <= p8_array_index_1084935_comb;
    p8_array_index_1084936 <= p8_array_index_1084936_comb;
    p8_array_index_1084937 <= p8_array_index_1084937_comb;
    p8_array_index_1084938 <= p8_array_index_1084938_comb;
    p8_res7__466 <= p8_res7__466_comb;
    p8_array_index_1084948 <= p8_array_index_1084948_comb;
    p8_array_index_1084949 <= p8_array_index_1084949_comb;
    p8_array_index_1084950 <= p8_array_index_1084950_comb;
    p8_array_index_1084951 <= p8_array_index_1084951_comb;
    p8_array_index_1084952 <= p8_array_index_1084952_comb;
    p8_res7__467 <= p8_res7__467_comb;
    p8_array_index_1084963 <= p8_array_index_1084963_comb;
    p8_array_index_1084964 <= p8_array_index_1084964_comb;
    p8_array_index_1084965 <= p8_array_index_1084965_comb;
    p8_array_index_1084966 <= p8_array_index_1084966_comb;
    p8_res7__468 <= p8_res7__468_comb;
    p8_res__39 <= p8_res__39_comb;
  end

  // ===== Pipe stage 9:
  wire [7:0] p9_array_index_1085263_comb;
  wire [7:0] p9_array_index_1085264_comb;
  wire [7:0] p9_array_index_1085265_comb;
  wire [7:0] p9_array_index_1085266_comb;
  wire [7:0] p9_res7__469_comb;
  wire [7:0] p9_array_index_1085277_comb;
  wire [7:0] p9_array_index_1085278_comb;
  wire [7:0] p9_array_index_1085279_comb;
  wire [7:0] p9_res7__470_comb;
  wire [7:0] p9_array_index_1085289_comb;
  wire [7:0] p9_array_index_1085290_comb;
  wire [7:0] p9_array_index_1085291_comb;
  wire [7:0] p9_res7__471_comb;
  wire [7:0] p9_array_index_1085302_comb;
  wire [7:0] p9_array_index_1085303_comb;
  wire [7:0] p9_res7__472_comb;
  wire [7:0] p9_array_index_1085313_comb;
  wire [7:0] p9_array_index_1085314_comb;
  wire [7:0] p9_res7__473_comb;
  wire [7:0] p9_array_index_1085325_comb;
  wire [7:0] p9_res7__474_comb;
  wire [7:0] p9_array_index_1085335_comb;
  wire [7:0] p9_res7__475_comb;
  wire [7:0] p9_res7__476_comb;
  wire [7:0] p9_res7__477_comb;
  wire [7:0] p9_res7__478_comb;
  wire [7:0] p9_res7__479_comb;
  wire [127:0] p9_res__29_comb;
  wire [127:0] p9_xor_1085375_comb;
  wire [127:0] p9_addedKey__71_comb;
  wire [7:0] p9_array_index_1085391_comb;
  wire [7:0] p9_array_index_1085392_comb;
  wire [7:0] p9_array_index_1085393_comb;
  wire [7:0] p9_array_index_1085394_comb;
  wire [7:0] p9_array_index_1085395_comb;
  wire [7:0] p9_array_index_1085396_comb;
  wire [7:0] p9_array_index_1085398_comb;
  wire [7:0] p9_array_index_1085400_comb;
  wire [7:0] p9_array_index_1085401_comb;
  wire [7:0] p9_array_index_1085402_comb;
  wire [7:0] p9_array_index_1085403_comb;
  wire [7:0] p9_array_index_1085404_comb;
  wire [7:0] p9_array_index_1085405_comb;
  wire [7:0] p9_array_index_1085407_comb;
  wire [7:0] p9_array_index_1085408_comb;
  wire [7:0] p9_array_index_1085409_comb;
  wire [7:0] p9_array_index_1085410_comb;
  wire [7:0] p9_array_index_1085411_comb;
  wire [7:0] p9_array_index_1085412_comb;
  wire [7:0] p9_array_index_1085413_comb;
  wire [7:0] p9_array_index_1085415_comb;
  wire [7:0] p9_res7__480_comb;
  wire [7:0] p9_array_index_1085424_comb;
  wire [7:0] p9_array_index_1085425_comb;
  wire [7:0] p9_array_index_1085426_comb;
  wire [7:0] p9_array_index_1085427_comb;
  wire [7:0] p9_array_index_1085428_comb;
  wire [7:0] p9_array_index_1085429_comb;
  wire [7:0] p9_res7__481_comb;
  wire [7:0] p9_array_index_1085439_comb;
  wire [7:0] p9_array_index_1085440_comb;
  wire [7:0] p9_array_index_1085441_comb;
  wire [7:0] p9_array_index_1085442_comb;
  wire [7:0] p9_array_index_1085443_comb;
  wire [7:0] p9_res7__482_comb;
  wire [7:0] p9_array_index_1085453_comb;
  wire [7:0] p9_array_index_1085454_comb;
  wire [7:0] p9_array_index_1085455_comb;
  wire [7:0] p9_array_index_1085456_comb;
  wire [7:0] p9_array_index_1085457_comb;
  wire [7:0] p9_res7__483_comb;
  wire [7:0] p9_array_index_1085468_comb;
  wire [7:0] p9_array_index_1085469_comb;
  wire [7:0] p9_array_index_1085470_comb;
  wire [7:0] p9_array_index_1085471_comb;
  wire [7:0] p9_res7__484_comb;
  wire [7:0] p9_array_index_1085481_comb;
  wire [7:0] p9_array_index_1085482_comb;
  wire [7:0] p9_array_index_1085483_comb;
  wire [7:0] p9_array_index_1085484_comb;
  wire [7:0] p9_res7__485_comb;
  wire [7:0] p9_array_index_1085495_comb;
  wire [7:0] p9_array_index_1085496_comb;
  wire [7:0] p9_array_index_1085497_comb;
  wire [7:0] p9_res7__486_comb;
  wire [7:0] p9_array_index_1085507_comb;
  wire [7:0] p9_array_index_1085508_comb;
  wire [7:0] p9_array_index_1085509_comb;
  wire [7:0] p9_res7__487_comb;
  wire [7:0] p9_array_index_1085520_comb;
  wire [7:0] p9_array_index_1085521_comb;
  wire [7:0] p9_res7__488_comb;
  wire [7:0] p9_array_index_1085531_comb;
  wire [7:0] p9_array_index_1085532_comb;
  wire [7:0] p9_res7__489_comb;
  wire [7:0] p9_array_index_1085543_comb;
  wire [7:0] p9_res7__490_comb;
  wire [7:0] p9_array_index_1085553_comb;
  wire [7:0] p9_res7__491_comb;
  wire [7:0] p9_res7__492_comb;
  wire [7:0] p9_res7__493_comb;
  wire [7:0] p9_res7__494_comb;
  wire [7:0] p9_res7__495_comb;
  wire [127:0] p9_res__30_comb;
  wire [127:0] p9_k9_comb;
  wire [127:0] p9_addedKey__72_comb;
  wire [7:0] p9_array_index_1085609_comb;
  wire [7:0] p9_array_index_1085610_comb;
  wire [7:0] p9_array_index_1085611_comb;
  wire [7:0] p9_array_index_1085612_comb;
  wire [7:0] p9_array_index_1085613_comb;
  wire [7:0] p9_array_index_1085614_comb;
  wire [7:0] p9_array_index_1085616_comb;
  wire [7:0] p9_array_index_1085618_comb;
  wire [7:0] p9_array_index_1085619_comb;
  wire [7:0] p9_array_index_1085620_comb;
  wire [7:0] p9_array_index_1085621_comb;
  wire [7:0] p9_array_index_1085622_comb;
  wire [7:0] p9_array_index_1085623_comb;
  wire [7:0] p9_array_index_1085625_comb;
  wire [7:0] p9_array_index_1085626_comb;
  wire [7:0] p9_array_index_1085627_comb;
  wire [7:0] p9_array_index_1085628_comb;
  wire [7:0] p9_array_index_1085629_comb;
  wire [7:0] p9_array_index_1085630_comb;
  wire [7:0] p9_array_index_1085631_comb;
  wire [7:0] p9_array_index_1085633_comb;
  wire [7:0] p9_res7__496_comb;
  wire [7:0] p9_array_index_1085642_comb;
  wire [7:0] p9_array_index_1085643_comb;
  wire [7:0] p9_array_index_1085644_comb;
  wire [7:0] p9_array_index_1085645_comb;
  wire [7:0] p9_array_index_1085646_comb;
  wire [7:0] p9_array_index_1085647_comb;
  wire [7:0] p9_res7__497_comb;
  wire [7:0] p9_array_index_1085657_comb;
  wire [7:0] p9_array_index_1085658_comb;
  wire [7:0] p9_array_index_1085659_comb;
  wire [7:0] p9_array_index_1085660_comb;
  wire [7:0] p9_array_index_1085661_comb;
  wire [7:0] p9_res7__498_comb;
  wire [7:0] p9_array_index_1085671_comb;
  wire [7:0] p9_array_index_1085672_comb;
  wire [7:0] p9_array_index_1085673_comb;
  wire [7:0] p9_array_index_1085674_comb;
  wire [7:0] p9_array_index_1085675_comb;
  wire [7:0] p9_res7__499_comb;
  wire [7:0] p9_array_index_1085686_comb;
  wire [7:0] p9_array_index_1085687_comb;
  wire [7:0] p9_array_index_1085688_comb;
  wire [7:0] p9_array_index_1085689_comb;
  wire [7:0] p9_res7__500_comb;
  wire [7:0] p9_array_index_1085699_comb;
  wire [7:0] p9_array_index_1085700_comb;
  wire [7:0] p9_array_index_1085701_comb;
  wire [7:0] p9_array_index_1085702_comb;
  wire [7:0] p9_res7__501_comb;
  wire [7:0] p9_array_index_1085713_comb;
  wire [7:0] p9_array_index_1085714_comb;
  wire [7:0] p9_array_index_1085715_comb;
  wire [7:0] p9_res7__502_comb;
  wire [7:0] p9_array_index_1085725_comb;
  wire [7:0] p9_array_index_1085726_comb;
  wire [7:0] p9_array_index_1085727_comb;
  wire [7:0] p9_res7__503_comb;
  wire [7:0] p9_array_index_1085738_comb;
  wire [7:0] p9_array_index_1085739_comb;
  wire [7:0] p9_res7__504_comb;
  wire [7:0] p9_array_index_1085749_comb;
  wire [7:0] p9_array_index_1085750_comb;
  wire [7:0] p9_res7__505_comb;
  wire [7:0] p9_array_index_1085761_comb;
  wire [7:0] p9_res7__506_comb;
  wire [7:0] p9_array_index_1085771_comb;
  wire [7:0] p9_res7__507_comb;
  wire [7:0] p9_res7__508_comb;
  wire [7:0] p9_res7__509_comb;
  wire [7:0] p9_res7__510_comb;
  wire [7:0] p9_res7__511_comb;
  wire [127:0] p9_res__31_comb;
  wire [127:0] p9_addedKey__40_comb;
  wire [7:0] p9_array_index_1085825_comb;
  wire [7:0] p9_array_index_1085826_comb;
  wire [7:0] p9_array_index_1085827_comb;
  wire [7:0] p9_array_index_1085828_comb;
  wire [7:0] p9_array_index_1085829_comb;
  wire [7:0] p9_array_index_1085830_comb;
  wire [7:0] p9_array_index_1085832_comb;
  wire [7:0] p9_array_index_1085834_comb;
  wire [7:0] p9_array_index_1085835_comb;
  wire [7:0] p9_array_index_1085836_comb;
  wire [7:0] p9_array_index_1085837_comb;
  wire [7:0] p9_array_index_1085838_comb;
  wire [7:0] p9_array_index_1085839_comb;
  wire [7:0] p9_array_index_1085841_comb;
  wire [7:0] p9_array_index_1085842_comb;
  wire [7:0] p9_array_index_1085843_comb;
  wire [7:0] p9_array_index_1085844_comb;
  wire [7:0] p9_array_index_1085845_comb;
  wire [7:0] p9_array_index_1085846_comb;
  wire [7:0] p9_array_index_1085847_comb;
  wire [7:0] p9_array_index_1085849_comb;
  wire [7:0] p9_res7__640_comb;
  wire [7:0] p9_array_index_1085858_comb;
  wire [7:0] p9_array_index_1085859_comb;
  wire [7:0] p9_array_index_1085860_comb;
  wire [7:0] p9_array_index_1085861_comb;
  wire [7:0] p9_array_index_1085862_comb;
  wire [7:0] p9_array_index_1085863_comb;
  wire [7:0] p9_res7__641_comb;
  wire [7:0] p9_array_index_1085873_comb;
  wire [7:0] p9_array_index_1085874_comb;
  wire [7:0] p9_array_index_1085875_comb;
  wire [7:0] p9_array_index_1085876_comb;
  wire [7:0] p9_array_index_1085877_comb;
  wire [7:0] p9_res7__642_comb;
  wire [7:0] p9_array_index_1085887_comb;
  wire [7:0] p9_array_index_1085888_comb;
  wire [7:0] p9_array_index_1085889_comb;
  wire [7:0] p9_array_index_1085890_comb;
  wire [7:0] p9_array_index_1085891_comb;
  wire [7:0] p9_res7__643_comb;
  wire [7:0] p9_array_index_1085902_comb;
  wire [7:0] p9_array_index_1085903_comb;
  wire [7:0] p9_array_index_1085904_comb;
  wire [7:0] p9_array_index_1085905_comb;
  wire [7:0] p9_res7__644_comb;
  wire [7:0] p9_array_index_1085915_comb;
  wire [7:0] p9_array_index_1085916_comb;
  wire [7:0] p9_array_index_1085917_comb;
  wire [7:0] p9_array_index_1085918_comb;
  wire [7:0] p9_res7__645_comb;
  wire [7:0] p9_array_index_1085929_comb;
  wire [7:0] p9_array_index_1085930_comb;
  wire [7:0] p9_array_index_1085931_comb;
  wire [7:0] p9_res7__646_comb;
  wire [7:0] p9_array_index_1085941_comb;
  wire [7:0] p9_array_index_1085942_comb;
  wire [7:0] p9_array_index_1085943_comb;
  wire [7:0] p9_res7__647_comb;
  wire [7:0] p9_array_index_1085954_comb;
  wire [7:0] p9_array_index_1085955_comb;
  wire [7:0] p9_res7__648_comb;
  wire [7:0] p9_array_index_1085965_comb;
  wire [7:0] p9_array_index_1085966_comb;
  wire [7:0] p9_res7__649_comb;
  wire [7:0] p9_array_index_1085977_comb;
  wire [7:0] p9_res7__650_comb;
  wire [7:0] p9_array_index_1085987_comb;
  wire [7:0] p9_res7__651_comb;
  wire [7:0] p9_res7__652_comb;
  wire [7:0] p9_res7__653_comb;
  wire [7:0] p9_res7__654_comb;
  wire [7:0] p9_res7__655_comb;
  wire [127:0] p9_newValue_comb;
  wire [127:0] p9_xor_1086027_comb;
  assign p9_array_index_1085263_comb = p8_literal_1076349[p8_res7__466];
  assign p9_array_index_1085264_comb = p8_literal_1076351[p8_res7__465];
  assign p9_array_index_1085265_comb = p8_literal_1076353[p8_res7__464];
  assign p9_array_index_1085266_comb = p8_literal_1076355[p8_array_index_1084886];
  assign p9_res7__469_comb = p8_literal_1076345[p8_res7__468] ^ p8_literal_1076347[p8_res7__467] ^ p9_array_index_1085263_comb ^ p9_array_index_1085264_comb ^ p9_array_index_1085265_comb ^ p9_array_index_1085266_comb ^ p8_array_index_1084887 ^ p8_literal_1076358[p8_array_index_1084888] ^ p8_array_index_1084889 ^ p8_array_index_1084924 ^ p8_literal_1076353[p8_array_index_1084891] ^ p8_literal_1076351[p8_array_index_1084908] ^ p8_literal_1076349[p8_array_index_1084893] ^ p8_literal_1076347[p8_array_index_1084910] ^ p8_literal_1076345[p8_array_index_1084895] ^ p8_array_index_1084896;
  assign p9_array_index_1085277_comb = p8_literal_1076351[p8_res7__466];
  assign p9_array_index_1085278_comb = p8_literal_1076353[p8_res7__465];
  assign p9_array_index_1085279_comb = p8_literal_1076355[p8_res7__464];
  assign p9_res7__470_comb = p8_literal_1076345[p9_res7__469_comb] ^ p8_literal_1076347[p8_res7__468] ^ p8_literal_1076349[p8_res7__467] ^ p9_array_index_1085277_comb ^ p9_array_index_1085278_comb ^ p9_array_index_1085279_comb ^ p8_array_index_1084886 ^ p8_literal_1076358[p8_array_index_1084887] ^ p8_array_index_1084888 ^ p8_array_index_1084938 ^ p8_array_index_1084906 ^ p8_literal_1076351[p8_array_index_1084891] ^ p8_literal_1076349[p8_array_index_1084908] ^ p8_literal_1076347[p8_array_index_1084893] ^ p8_literal_1076345[p8_array_index_1084910] ^ p8_array_index_1084895;
  assign p9_array_index_1085289_comb = p8_literal_1076351[p8_res7__467];
  assign p9_array_index_1085290_comb = p8_literal_1076353[p8_res7__466];
  assign p9_array_index_1085291_comb = p8_literal_1076355[p8_res7__465];
  assign p9_res7__471_comb = p8_literal_1076345[p9_res7__470_comb] ^ p8_literal_1076347[p9_res7__469_comb] ^ p8_literal_1076349[p8_res7__468] ^ p9_array_index_1085289_comb ^ p9_array_index_1085290_comb ^ p9_array_index_1085291_comb ^ p8_res7__464 ^ p8_literal_1076358[p8_array_index_1084886] ^ p8_array_index_1084887 ^ p8_array_index_1084952 ^ p8_array_index_1084923 ^ p8_literal_1076351[p8_array_index_1084890] ^ p8_literal_1076349[p8_array_index_1084891] ^ p8_literal_1076347[p8_array_index_1084908] ^ p8_literal_1076345[p8_array_index_1084893] ^ p8_array_index_1084910;
  assign p9_array_index_1085302_comb = p8_literal_1076353[p8_res7__467];
  assign p9_array_index_1085303_comb = p8_literal_1076355[p8_res7__466];
  assign p9_res7__472_comb = p8_literal_1076345[p9_res7__471_comb] ^ p8_literal_1076347[p9_res7__470_comb] ^ p8_literal_1076349[p9_res7__469_comb] ^ p8_literal_1076351[p8_res7__468] ^ p9_array_index_1085302_comb ^ p9_array_index_1085303_comb ^ p8_res7__465 ^ p8_literal_1076358[p8_res7__464] ^ p8_array_index_1084886 ^ p8_array_index_1084966 ^ p8_array_index_1084937 ^ p8_array_index_1084905 ^ p8_literal_1076349[p8_array_index_1084890] ^ p8_literal_1076347[p8_array_index_1084891] ^ p8_literal_1076345[p8_array_index_1084908] ^ p8_array_index_1084893;
  assign p9_array_index_1085313_comb = p8_literal_1076353[p8_res7__468];
  assign p9_array_index_1085314_comb = p8_literal_1076355[p8_res7__467];
  assign p9_res7__473_comb = p8_literal_1076345[p9_res7__472_comb] ^ p8_literal_1076347[p9_res7__471_comb] ^ p8_literal_1076349[p9_res7__470_comb] ^ p8_literal_1076351[p9_res7__469_comb] ^ p9_array_index_1085313_comb ^ p9_array_index_1085314_comb ^ p8_res7__466 ^ p8_literal_1076358[p8_res7__465] ^ p8_res7__464 ^ p9_array_index_1085266_comb ^ p8_array_index_1084951 ^ p8_array_index_1084922 ^ p8_literal_1076349[p8_array_index_1084889] ^ p8_literal_1076347[p8_array_index_1084890] ^ p8_literal_1076345[p8_array_index_1084891] ^ p8_array_index_1084908;
  assign p9_array_index_1085325_comb = p8_literal_1076355[p8_res7__468];
  assign p9_res7__474_comb = p8_literal_1076345[p9_res7__473_comb] ^ p8_literal_1076347[p9_res7__472_comb] ^ p8_literal_1076349[p9_res7__471_comb] ^ p8_literal_1076351[p9_res7__470_comb] ^ p8_literal_1076353[p9_res7__469_comb] ^ p9_array_index_1085325_comb ^ p8_res7__467 ^ p8_literal_1076358[p8_res7__466] ^ p8_res7__465 ^ p9_array_index_1085279_comb ^ p8_array_index_1084965 ^ p8_array_index_1084936 ^ p8_array_index_1084904 ^ p8_literal_1076347[p8_array_index_1084889] ^ p8_literal_1076345[p8_array_index_1084890] ^ p8_array_index_1084891;
  assign p9_array_index_1085335_comb = p8_literal_1076355[p9_res7__469_comb];
  assign p9_res7__475_comb = p8_literal_1076345[p9_res7__474_comb] ^ p8_literal_1076347[p9_res7__473_comb] ^ p8_literal_1076349[p9_res7__472_comb] ^ p8_literal_1076351[p9_res7__471_comb] ^ p8_literal_1076353[p9_res7__470_comb] ^ p9_array_index_1085335_comb ^ p8_res7__468 ^ p8_literal_1076358[p8_res7__467] ^ p8_res7__466 ^ p9_array_index_1085291_comb ^ p9_array_index_1085265_comb ^ p8_array_index_1084950 ^ p8_array_index_1084921 ^ p8_literal_1076347[p8_array_index_1084888] ^ p8_literal_1076345[p8_array_index_1084889] ^ p8_array_index_1084890;
  assign p9_res7__476_comb = p8_literal_1076345[p9_res7__475_comb] ^ p8_literal_1076347[p9_res7__474_comb] ^ p8_literal_1076349[p9_res7__473_comb] ^ p8_literal_1076351[p9_res7__472_comb] ^ p8_literal_1076353[p9_res7__471_comb] ^ p8_literal_1076355[p9_res7__470_comb] ^ p9_res7__469_comb ^ p8_literal_1076358[p8_res7__468] ^ p8_res7__467 ^ p9_array_index_1085303_comb ^ p9_array_index_1085278_comb ^ p8_array_index_1084964 ^ p8_array_index_1084935 ^ p8_array_index_1084903 ^ p8_literal_1076345[p8_array_index_1084888] ^ p8_array_index_1084889;
  assign p9_res7__477_comb = p8_literal_1076345[p9_res7__476_comb] ^ p8_literal_1076347[p9_res7__475_comb] ^ p8_literal_1076349[p9_res7__474_comb] ^ p8_literal_1076351[p9_res7__473_comb] ^ p8_literal_1076353[p9_res7__472_comb] ^ p8_literal_1076355[p9_res7__471_comb] ^ p9_res7__470_comb ^ p8_literal_1076358[p9_res7__469_comb] ^ p8_res7__468 ^ p9_array_index_1085314_comb ^ p9_array_index_1085290_comb ^ p9_array_index_1085264_comb ^ p8_array_index_1084949 ^ p8_array_index_1084920 ^ p8_literal_1076345[p8_array_index_1084887] ^ p8_array_index_1084888;
  assign p9_res7__478_comb = p8_literal_1076345[p9_res7__477_comb] ^ p8_literal_1076347[p9_res7__476_comb] ^ p8_literal_1076349[p9_res7__475_comb] ^ p8_literal_1076351[p9_res7__474_comb] ^ p8_literal_1076353[p9_res7__473_comb] ^ p8_literal_1076355[p9_res7__472_comb] ^ p9_res7__471_comb ^ p8_literal_1076358[p9_res7__470_comb] ^ p9_res7__469_comb ^ p9_array_index_1085325_comb ^ p9_array_index_1085302_comb ^ p9_array_index_1085277_comb ^ p8_array_index_1084963 ^ p8_array_index_1084934 ^ p8_array_index_1084902 ^ p8_array_index_1084887;
  assign p9_res7__479_comb = p8_literal_1076345[p9_res7__478_comb] ^ p8_literal_1076347[p9_res7__477_comb] ^ p8_literal_1076349[p9_res7__476_comb] ^ p8_literal_1076351[p9_res7__475_comb] ^ p8_literal_1076353[p9_res7__474_comb] ^ p8_literal_1076355[p9_res7__473_comb] ^ p9_res7__472_comb ^ p8_literal_1076358[p9_res7__471_comb] ^ p9_res7__470_comb ^ p9_array_index_1085335_comb ^ p9_array_index_1085313_comb ^ p9_array_index_1085289_comb ^ p9_array_index_1085263_comb ^ p8_array_index_1084948 ^ p8_array_index_1084919 ^ p8_array_index_1084886;
  assign p9_res__29_comb = {p9_res7__479_comb, p9_res7__478_comb, p9_res7__477_comb, p9_res7__476_comb, p9_res7__475_comb, p9_res7__474_comb, p9_res7__473_comb, p9_res7__472_comb, p9_res7__471_comb, p9_res7__470_comb, p9_res7__469_comb, p8_res7__468, p8_res7__467, p8_res7__466, p8_res7__465, p8_res7__464};
  assign p9_xor_1085375_comb = p9_res__29_comb ^ p8_xor_1084652;
  assign p9_addedKey__71_comb = p9_xor_1085375_comb ^ 128'h1003_dba7_2e34_5ff6_643b_9533_3f27_141f;
  assign p9_array_index_1085391_comb = p8_arr[p9_addedKey__71_comb[127:120]];
  assign p9_array_index_1085392_comb = p8_arr[p9_addedKey__71_comb[119:112]];
  assign p9_array_index_1085393_comb = p8_arr[p9_addedKey__71_comb[111:104]];
  assign p9_array_index_1085394_comb = p8_arr[p9_addedKey__71_comb[103:96]];
  assign p9_array_index_1085395_comb = p8_arr[p9_addedKey__71_comb[95:88]];
  assign p9_array_index_1085396_comb = p8_arr[p9_addedKey__71_comb[87:80]];
  assign p9_array_index_1085398_comb = p8_arr[p9_addedKey__71_comb[71:64]];
  assign p9_array_index_1085400_comb = p8_arr[p9_addedKey__71_comb[55:48]];
  assign p9_array_index_1085401_comb = p8_arr[p9_addedKey__71_comb[47:40]];
  assign p9_array_index_1085402_comb = p8_arr[p9_addedKey__71_comb[39:32]];
  assign p9_array_index_1085403_comb = p8_arr[p9_addedKey__71_comb[31:24]];
  assign p9_array_index_1085404_comb = p8_arr[p9_addedKey__71_comb[23:16]];
  assign p9_array_index_1085405_comb = p8_arr[p9_addedKey__71_comb[15:8]];
  assign p9_array_index_1085407_comb = p8_literal_1076345[p9_array_index_1085391_comb];
  assign p9_array_index_1085408_comb = p8_literal_1076347[p9_array_index_1085392_comb];
  assign p9_array_index_1085409_comb = p8_literal_1076349[p9_array_index_1085393_comb];
  assign p9_array_index_1085410_comb = p8_literal_1076351[p9_array_index_1085394_comb];
  assign p9_array_index_1085411_comb = p8_literal_1076353[p9_array_index_1085395_comb];
  assign p9_array_index_1085412_comb = p8_literal_1076355[p9_array_index_1085396_comb];
  assign p9_array_index_1085413_comb = p8_arr[p9_addedKey__71_comb[79:72]];
  assign p9_array_index_1085415_comb = p8_arr[p9_addedKey__71_comb[63:56]];
  assign p9_res7__480_comb = p9_array_index_1085407_comb ^ p9_array_index_1085408_comb ^ p9_array_index_1085409_comb ^ p9_array_index_1085410_comb ^ p9_array_index_1085411_comb ^ p9_array_index_1085412_comb ^ p9_array_index_1085413_comb ^ p8_literal_1076358[p9_array_index_1085398_comb] ^ p9_array_index_1085415_comb ^ p8_literal_1076355[p9_array_index_1085400_comb] ^ p8_literal_1076353[p9_array_index_1085401_comb] ^ p8_literal_1076351[p9_array_index_1085402_comb] ^ p8_literal_1076349[p9_array_index_1085403_comb] ^ p8_literal_1076347[p9_array_index_1085404_comb] ^ p8_literal_1076345[p9_array_index_1085405_comb] ^ p8_arr[p9_addedKey__71_comb[7:0]];
  assign p9_array_index_1085424_comb = p8_literal_1076345[p9_res7__480_comb];
  assign p9_array_index_1085425_comb = p8_literal_1076347[p9_array_index_1085391_comb];
  assign p9_array_index_1085426_comb = p8_literal_1076349[p9_array_index_1085392_comb];
  assign p9_array_index_1085427_comb = p8_literal_1076351[p9_array_index_1085393_comb];
  assign p9_array_index_1085428_comb = p8_literal_1076353[p9_array_index_1085394_comb];
  assign p9_array_index_1085429_comb = p8_literal_1076355[p9_array_index_1085395_comb];
  assign p9_res7__481_comb = p9_array_index_1085424_comb ^ p9_array_index_1085425_comb ^ p9_array_index_1085426_comb ^ p9_array_index_1085427_comb ^ p9_array_index_1085428_comb ^ p9_array_index_1085429_comb ^ p9_array_index_1085396_comb ^ p8_literal_1076358[p9_array_index_1085413_comb] ^ p9_array_index_1085398_comb ^ p8_literal_1076355[p9_array_index_1085415_comb] ^ p8_literal_1076353[p9_array_index_1085400_comb] ^ p8_literal_1076351[p9_array_index_1085401_comb] ^ p8_literal_1076349[p9_array_index_1085402_comb] ^ p8_literal_1076347[p9_array_index_1085403_comb] ^ p8_literal_1076345[p9_array_index_1085404_comb] ^ p9_array_index_1085405_comb;
  assign p9_array_index_1085439_comb = p8_literal_1076347[p9_res7__480_comb];
  assign p9_array_index_1085440_comb = p8_literal_1076349[p9_array_index_1085391_comb];
  assign p9_array_index_1085441_comb = p8_literal_1076351[p9_array_index_1085392_comb];
  assign p9_array_index_1085442_comb = p8_literal_1076353[p9_array_index_1085393_comb];
  assign p9_array_index_1085443_comb = p8_literal_1076355[p9_array_index_1085394_comb];
  assign p9_res7__482_comb = p8_literal_1076345[p9_res7__481_comb] ^ p9_array_index_1085439_comb ^ p9_array_index_1085440_comb ^ p9_array_index_1085441_comb ^ p9_array_index_1085442_comb ^ p9_array_index_1085443_comb ^ p9_array_index_1085395_comb ^ p8_literal_1076358[p9_array_index_1085396_comb] ^ p9_array_index_1085413_comb ^ p8_literal_1076355[p9_array_index_1085398_comb] ^ p8_literal_1076353[p9_array_index_1085415_comb] ^ p8_literal_1076351[p9_array_index_1085400_comb] ^ p8_literal_1076349[p9_array_index_1085401_comb] ^ p8_literal_1076347[p9_array_index_1085402_comb] ^ p8_literal_1076345[p9_array_index_1085403_comb] ^ p9_array_index_1085404_comb;
  assign p9_array_index_1085453_comb = p8_literal_1076347[p9_res7__481_comb];
  assign p9_array_index_1085454_comb = p8_literal_1076349[p9_res7__480_comb];
  assign p9_array_index_1085455_comb = p8_literal_1076351[p9_array_index_1085391_comb];
  assign p9_array_index_1085456_comb = p8_literal_1076353[p9_array_index_1085392_comb];
  assign p9_array_index_1085457_comb = p8_literal_1076355[p9_array_index_1085393_comb];
  assign p9_res7__483_comb = p8_literal_1076345[p9_res7__482_comb] ^ p9_array_index_1085453_comb ^ p9_array_index_1085454_comb ^ p9_array_index_1085455_comb ^ p9_array_index_1085456_comb ^ p9_array_index_1085457_comb ^ p9_array_index_1085394_comb ^ p8_literal_1076358[p9_array_index_1085395_comb] ^ p9_array_index_1085396_comb ^ p8_literal_1076355[p9_array_index_1085413_comb] ^ p8_literal_1076353[p9_array_index_1085398_comb] ^ p8_literal_1076351[p9_array_index_1085415_comb] ^ p8_literal_1076349[p9_array_index_1085400_comb] ^ p8_literal_1076347[p9_array_index_1085401_comb] ^ p8_literal_1076345[p9_array_index_1085402_comb] ^ p9_array_index_1085403_comb;
  assign p9_array_index_1085468_comb = p8_literal_1076349[p9_res7__481_comb];
  assign p9_array_index_1085469_comb = p8_literal_1076351[p9_res7__480_comb];
  assign p9_array_index_1085470_comb = p8_literal_1076353[p9_array_index_1085391_comb];
  assign p9_array_index_1085471_comb = p8_literal_1076355[p9_array_index_1085392_comb];
  assign p9_res7__484_comb = p8_literal_1076345[p9_res7__483_comb] ^ p8_literal_1076347[p9_res7__482_comb] ^ p9_array_index_1085468_comb ^ p9_array_index_1085469_comb ^ p9_array_index_1085470_comb ^ p9_array_index_1085471_comb ^ p9_array_index_1085393_comb ^ p8_literal_1076358[p9_array_index_1085394_comb] ^ p9_array_index_1085395_comb ^ p9_array_index_1085412_comb ^ p8_literal_1076353[p9_array_index_1085413_comb] ^ p8_literal_1076351[p9_array_index_1085398_comb] ^ p8_literal_1076349[p9_array_index_1085415_comb] ^ p8_literal_1076347[p9_array_index_1085400_comb] ^ p8_literal_1076345[p9_array_index_1085401_comb] ^ p9_array_index_1085402_comb;
  assign p9_array_index_1085481_comb = p8_literal_1076349[p9_res7__482_comb];
  assign p9_array_index_1085482_comb = p8_literal_1076351[p9_res7__481_comb];
  assign p9_array_index_1085483_comb = p8_literal_1076353[p9_res7__480_comb];
  assign p9_array_index_1085484_comb = p8_literal_1076355[p9_array_index_1085391_comb];
  assign p9_res7__485_comb = p8_literal_1076345[p9_res7__484_comb] ^ p8_literal_1076347[p9_res7__483_comb] ^ p9_array_index_1085481_comb ^ p9_array_index_1085482_comb ^ p9_array_index_1085483_comb ^ p9_array_index_1085484_comb ^ p9_array_index_1085392_comb ^ p8_literal_1076358[p9_array_index_1085393_comb] ^ p9_array_index_1085394_comb ^ p9_array_index_1085429_comb ^ p8_literal_1076353[p9_array_index_1085396_comb] ^ p8_literal_1076351[p9_array_index_1085413_comb] ^ p8_literal_1076349[p9_array_index_1085398_comb] ^ p8_literal_1076347[p9_array_index_1085415_comb] ^ p8_literal_1076345[p9_array_index_1085400_comb] ^ p9_array_index_1085401_comb;
  assign p9_array_index_1085495_comb = p8_literal_1076351[p9_res7__482_comb];
  assign p9_array_index_1085496_comb = p8_literal_1076353[p9_res7__481_comb];
  assign p9_array_index_1085497_comb = p8_literal_1076355[p9_res7__480_comb];
  assign p9_res7__486_comb = p8_literal_1076345[p9_res7__485_comb] ^ p8_literal_1076347[p9_res7__484_comb] ^ p8_literal_1076349[p9_res7__483_comb] ^ p9_array_index_1085495_comb ^ p9_array_index_1085496_comb ^ p9_array_index_1085497_comb ^ p9_array_index_1085391_comb ^ p8_literal_1076358[p9_array_index_1085392_comb] ^ p9_array_index_1085393_comb ^ p9_array_index_1085443_comb ^ p9_array_index_1085411_comb ^ p8_literal_1076351[p9_array_index_1085396_comb] ^ p8_literal_1076349[p9_array_index_1085413_comb] ^ p8_literal_1076347[p9_array_index_1085398_comb] ^ p8_literal_1076345[p9_array_index_1085415_comb] ^ p9_array_index_1085400_comb;
  assign p9_array_index_1085507_comb = p8_literal_1076351[p9_res7__483_comb];
  assign p9_array_index_1085508_comb = p8_literal_1076353[p9_res7__482_comb];
  assign p9_array_index_1085509_comb = p8_literal_1076355[p9_res7__481_comb];
  assign p9_res7__487_comb = p8_literal_1076345[p9_res7__486_comb] ^ p8_literal_1076347[p9_res7__485_comb] ^ p8_literal_1076349[p9_res7__484_comb] ^ p9_array_index_1085507_comb ^ p9_array_index_1085508_comb ^ p9_array_index_1085509_comb ^ p9_res7__480_comb ^ p8_literal_1076358[p9_array_index_1085391_comb] ^ p9_array_index_1085392_comb ^ p9_array_index_1085457_comb ^ p9_array_index_1085428_comb ^ p8_literal_1076351[p9_array_index_1085395_comb] ^ p8_literal_1076349[p9_array_index_1085396_comb] ^ p8_literal_1076347[p9_array_index_1085413_comb] ^ p8_literal_1076345[p9_array_index_1085398_comb] ^ p9_array_index_1085415_comb;
  assign p9_array_index_1085520_comb = p8_literal_1076353[p9_res7__483_comb];
  assign p9_array_index_1085521_comb = p8_literal_1076355[p9_res7__482_comb];
  assign p9_res7__488_comb = p8_literal_1076345[p9_res7__487_comb] ^ p8_literal_1076347[p9_res7__486_comb] ^ p8_literal_1076349[p9_res7__485_comb] ^ p8_literal_1076351[p9_res7__484_comb] ^ p9_array_index_1085520_comb ^ p9_array_index_1085521_comb ^ p9_res7__481_comb ^ p8_literal_1076358[p9_res7__480_comb] ^ p9_array_index_1085391_comb ^ p9_array_index_1085471_comb ^ p9_array_index_1085442_comb ^ p9_array_index_1085410_comb ^ p8_literal_1076349[p9_array_index_1085395_comb] ^ p8_literal_1076347[p9_array_index_1085396_comb] ^ p8_literal_1076345[p9_array_index_1085413_comb] ^ p9_array_index_1085398_comb;
  assign p9_array_index_1085531_comb = p8_literal_1076353[p9_res7__484_comb];
  assign p9_array_index_1085532_comb = p8_literal_1076355[p9_res7__483_comb];
  assign p9_res7__489_comb = p8_literal_1076345[p9_res7__488_comb] ^ p8_literal_1076347[p9_res7__487_comb] ^ p8_literal_1076349[p9_res7__486_comb] ^ p8_literal_1076351[p9_res7__485_comb] ^ p9_array_index_1085531_comb ^ p9_array_index_1085532_comb ^ p9_res7__482_comb ^ p8_literal_1076358[p9_res7__481_comb] ^ p9_res7__480_comb ^ p9_array_index_1085484_comb ^ p9_array_index_1085456_comb ^ p9_array_index_1085427_comb ^ p8_literal_1076349[p9_array_index_1085394_comb] ^ p8_literal_1076347[p9_array_index_1085395_comb] ^ p8_literal_1076345[p9_array_index_1085396_comb] ^ p9_array_index_1085413_comb;
  assign p9_array_index_1085543_comb = p8_literal_1076355[p9_res7__484_comb];
  assign p9_res7__490_comb = p8_literal_1076345[p9_res7__489_comb] ^ p8_literal_1076347[p9_res7__488_comb] ^ p8_literal_1076349[p9_res7__487_comb] ^ p8_literal_1076351[p9_res7__486_comb] ^ p8_literal_1076353[p9_res7__485_comb] ^ p9_array_index_1085543_comb ^ p9_res7__483_comb ^ p8_literal_1076358[p9_res7__482_comb] ^ p9_res7__481_comb ^ p9_array_index_1085497_comb ^ p9_array_index_1085470_comb ^ p9_array_index_1085441_comb ^ p9_array_index_1085409_comb ^ p8_literal_1076347[p9_array_index_1085394_comb] ^ p8_literal_1076345[p9_array_index_1085395_comb] ^ p9_array_index_1085396_comb;
  assign p9_array_index_1085553_comb = p8_literal_1076355[p9_res7__485_comb];
  assign p9_res7__491_comb = p8_literal_1076345[p9_res7__490_comb] ^ p8_literal_1076347[p9_res7__489_comb] ^ p8_literal_1076349[p9_res7__488_comb] ^ p8_literal_1076351[p9_res7__487_comb] ^ p8_literal_1076353[p9_res7__486_comb] ^ p9_array_index_1085553_comb ^ p9_res7__484_comb ^ p8_literal_1076358[p9_res7__483_comb] ^ p9_res7__482_comb ^ p9_array_index_1085509_comb ^ p9_array_index_1085483_comb ^ p9_array_index_1085455_comb ^ p9_array_index_1085426_comb ^ p8_literal_1076347[p9_array_index_1085393_comb] ^ p8_literal_1076345[p9_array_index_1085394_comb] ^ p9_array_index_1085395_comb;
  assign p9_res7__492_comb = p8_literal_1076345[p9_res7__491_comb] ^ p8_literal_1076347[p9_res7__490_comb] ^ p8_literal_1076349[p9_res7__489_comb] ^ p8_literal_1076351[p9_res7__488_comb] ^ p8_literal_1076353[p9_res7__487_comb] ^ p8_literal_1076355[p9_res7__486_comb] ^ p9_res7__485_comb ^ p8_literal_1076358[p9_res7__484_comb] ^ p9_res7__483_comb ^ p9_array_index_1085521_comb ^ p9_array_index_1085496_comb ^ p9_array_index_1085469_comb ^ p9_array_index_1085440_comb ^ p9_array_index_1085408_comb ^ p8_literal_1076345[p9_array_index_1085393_comb] ^ p9_array_index_1085394_comb;
  assign p9_res7__493_comb = p8_literal_1076345[p9_res7__492_comb] ^ p8_literal_1076347[p9_res7__491_comb] ^ p8_literal_1076349[p9_res7__490_comb] ^ p8_literal_1076351[p9_res7__489_comb] ^ p8_literal_1076353[p9_res7__488_comb] ^ p8_literal_1076355[p9_res7__487_comb] ^ p9_res7__486_comb ^ p8_literal_1076358[p9_res7__485_comb] ^ p9_res7__484_comb ^ p9_array_index_1085532_comb ^ p9_array_index_1085508_comb ^ p9_array_index_1085482_comb ^ p9_array_index_1085454_comb ^ p9_array_index_1085425_comb ^ p8_literal_1076345[p9_array_index_1085392_comb] ^ p9_array_index_1085393_comb;
  assign p9_res7__494_comb = p8_literal_1076345[p9_res7__493_comb] ^ p8_literal_1076347[p9_res7__492_comb] ^ p8_literal_1076349[p9_res7__491_comb] ^ p8_literal_1076351[p9_res7__490_comb] ^ p8_literal_1076353[p9_res7__489_comb] ^ p8_literal_1076355[p9_res7__488_comb] ^ p9_res7__487_comb ^ p8_literal_1076358[p9_res7__486_comb] ^ p9_res7__485_comb ^ p9_array_index_1085543_comb ^ p9_array_index_1085520_comb ^ p9_array_index_1085495_comb ^ p9_array_index_1085468_comb ^ p9_array_index_1085439_comb ^ p9_array_index_1085407_comb ^ p9_array_index_1085392_comb;
  assign p9_res7__495_comb = p8_literal_1076345[p9_res7__494_comb] ^ p8_literal_1076347[p9_res7__493_comb] ^ p8_literal_1076349[p9_res7__492_comb] ^ p8_literal_1076351[p9_res7__491_comb] ^ p8_literal_1076353[p9_res7__490_comb] ^ p8_literal_1076355[p9_res7__489_comb] ^ p9_res7__488_comb ^ p8_literal_1076358[p9_res7__487_comb] ^ p9_res7__486_comb ^ p9_array_index_1085553_comb ^ p9_array_index_1085531_comb ^ p9_array_index_1085507_comb ^ p9_array_index_1085481_comb ^ p9_array_index_1085453_comb ^ p9_array_index_1085424_comb ^ p9_array_index_1085391_comb;
  assign p9_res__30_comb = {p9_res7__495_comb, p9_res7__494_comb, p9_res7__493_comb, p9_res7__492_comb, p9_res7__491_comb, p9_res7__490_comb, p9_res7__489_comb, p9_res7__488_comb, p9_res7__487_comb, p9_res7__486_comb, p9_res7__485_comb, p9_res7__484_comb, p9_res7__483_comb, p9_res7__482_comb, p9_res7__481_comb, p9_res7__480_comb};
  assign p9_k9_comb = p9_res__30_comb ^ p8_xor_1084870;
  assign p9_addedKey__72_comb = p9_k9_comb ^ 128'h5ea7_d858_1e14_9b61_f16a_c145_9ced_a820;
  assign p9_array_index_1085609_comb = p8_arr[p9_addedKey__72_comb[127:120]];
  assign p9_array_index_1085610_comb = p8_arr[p9_addedKey__72_comb[119:112]];
  assign p9_array_index_1085611_comb = p8_arr[p9_addedKey__72_comb[111:104]];
  assign p9_array_index_1085612_comb = p8_arr[p9_addedKey__72_comb[103:96]];
  assign p9_array_index_1085613_comb = p8_arr[p9_addedKey__72_comb[95:88]];
  assign p9_array_index_1085614_comb = p8_arr[p9_addedKey__72_comb[87:80]];
  assign p9_array_index_1085616_comb = p8_arr[p9_addedKey__72_comb[71:64]];
  assign p9_array_index_1085618_comb = p8_arr[p9_addedKey__72_comb[55:48]];
  assign p9_array_index_1085619_comb = p8_arr[p9_addedKey__72_comb[47:40]];
  assign p9_array_index_1085620_comb = p8_arr[p9_addedKey__72_comb[39:32]];
  assign p9_array_index_1085621_comb = p8_arr[p9_addedKey__72_comb[31:24]];
  assign p9_array_index_1085622_comb = p8_arr[p9_addedKey__72_comb[23:16]];
  assign p9_array_index_1085623_comb = p8_arr[p9_addedKey__72_comb[15:8]];
  assign p9_array_index_1085625_comb = p8_literal_1076345[p9_array_index_1085609_comb];
  assign p9_array_index_1085626_comb = p8_literal_1076347[p9_array_index_1085610_comb];
  assign p9_array_index_1085627_comb = p8_literal_1076349[p9_array_index_1085611_comb];
  assign p9_array_index_1085628_comb = p8_literal_1076351[p9_array_index_1085612_comb];
  assign p9_array_index_1085629_comb = p8_literal_1076353[p9_array_index_1085613_comb];
  assign p9_array_index_1085630_comb = p8_literal_1076355[p9_array_index_1085614_comb];
  assign p9_array_index_1085631_comb = p8_arr[p9_addedKey__72_comb[79:72]];
  assign p9_array_index_1085633_comb = p8_arr[p9_addedKey__72_comb[63:56]];
  assign p9_res7__496_comb = p9_array_index_1085625_comb ^ p9_array_index_1085626_comb ^ p9_array_index_1085627_comb ^ p9_array_index_1085628_comb ^ p9_array_index_1085629_comb ^ p9_array_index_1085630_comb ^ p9_array_index_1085631_comb ^ p8_literal_1076358[p9_array_index_1085616_comb] ^ p9_array_index_1085633_comb ^ p8_literal_1076355[p9_array_index_1085618_comb] ^ p8_literal_1076353[p9_array_index_1085619_comb] ^ p8_literal_1076351[p9_array_index_1085620_comb] ^ p8_literal_1076349[p9_array_index_1085621_comb] ^ p8_literal_1076347[p9_array_index_1085622_comb] ^ p8_literal_1076345[p9_array_index_1085623_comb] ^ p8_arr[p9_addedKey__72_comb[7:0]];
  assign p9_array_index_1085642_comb = p8_literal_1076345[p9_res7__496_comb];
  assign p9_array_index_1085643_comb = p8_literal_1076347[p9_array_index_1085609_comb];
  assign p9_array_index_1085644_comb = p8_literal_1076349[p9_array_index_1085610_comb];
  assign p9_array_index_1085645_comb = p8_literal_1076351[p9_array_index_1085611_comb];
  assign p9_array_index_1085646_comb = p8_literal_1076353[p9_array_index_1085612_comb];
  assign p9_array_index_1085647_comb = p8_literal_1076355[p9_array_index_1085613_comb];
  assign p9_res7__497_comb = p9_array_index_1085642_comb ^ p9_array_index_1085643_comb ^ p9_array_index_1085644_comb ^ p9_array_index_1085645_comb ^ p9_array_index_1085646_comb ^ p9_array_index_1085647_comb ^ p9_array_index_1085614_comb ^ p8_literal_1076358[p9_array_index_1085631_comb] ^ p9_array_index_1085616_comb ^ p8_literal_1076355[p9_array_index_1085633_comb] ^ p8_literal_1076353[p9_array_index_1085618_comb] ^ p8_literal_1076351[p9_array_index_1085619_comb] ^ p8_literal_1076349[p9_array_index_1085620_comb] ^ p8_literal_1076347[p9_array_index_1085621_comb] ^ p8_literal_1076345[p9_array_index_1085622_comb] ^ p9_array_index_1085623_comb;
  assign p9_array_index_1085657_comb = p8_literal_1076347[p9_res7__496_comb];
  assign p9_array_index_1085658_comb = p8_literal_1076349[p9_array_index_1085609_comb];
  assign p9_array_index_1085659_comb = p8_literal_1076351[p9_array_index_1085610_comb];
  assign p9_array_index_1085660_comb = p8_literal_1076353[p9_array_index_1085611_comb];
  assign p9_array_index_1085661_comb = p8_literal_1076355[p9_array_index_1085612_comb];
  assign p9_res7__498_comb = p8_literal_1076345[p9_res7__497_comb] ^ p9_array_index_1085657_comb ^ p9_array_index_1085658_comb ^ p9_array_index_1085659_comb ^ p9_array_index_1085660_comb ^ p9_array_index_1085661_comb ^ p9_array_index_1085613_comb ^ p8_literal_1076358[p9_array_index_1085614_comb] ^ p9_array_index_1085631_comb ^ p8_literal_1076355[p9_array_index_1085616_comb] ^ p8_literal_1076353[p9_array_index_1085633_comb] ^ p8_literal_1076351[p9_array_index_1085618_comb] ^ p8_literal_1076349[p9_array_index_1085619_comb] ^ p8_literal_1076347[p9_array_index_1085620_comb] ^ p8_literal_1076345[p9_array_index_1085621_comb] ^ p9_array_index_1085622_comb;
  assign p9_array_index_1085671_comb = p8_literal_1076347[p9_res7__497_comb];
  assign p9_array_index_1085672_comb = p8_literal_1076349[p9_res7__496_comb];
  assign p9_array_index_1085673_comb = p8_literal_1076351[p9_array_index_1085609_comb];
  assign p9_array_index_1085674_comb = p8_literal_1076353[p9_array_index_1085610_comb];
  assign p9_array_index_1085675_comb = p8_literal_1076355[p9_array_index_1085611_comb];
  assign p9_res7__499_comb = p8_literal_1076345[p9_res7__498_comb] ^ p9_array_index_1085671_comb ^ p9_array_index_1085672_comb ^ p9_array_index_1085673_comb ^ p9_array_index_1085674_comb ^ p9_array_index_1085675_comb ^ p9_array_index_1085612_comb ^ p8_literal_1076358[p9_array_index_1085613_comb] ^ p9_array_index_1085614_comb ^ p8_literal_1076355[p9_array_index_1085631_comb] ^ p8_literal_1076353[p9_array_index_1085616_comb] ^ p8_literal_1076351[p9_array_index_1085633_comb] ^ p8_literal_1076349[p9_array_index_1085618_comb] ^ p8_literal_1076347[p9_array_index_1085619_comb] ^ p8_literal_1076345[p9_array_index_1085620_comb] ^ p9_array_index_1085621_comb;
  assign p9_array_index_1085686_comb = p8_literal_1076349[p9_res7__497_comb];
  assign p9_array_index_1085687_comb = p8_literal_1076351[p9_res7__496_comb];
  assign p9_array_index_1085688_comb = p8_literal_1076353[p9_array_index_1085609_comb];
  assign p9_array_index_1085689_comb = p8_literal_1076355[p9_array_index_1085610_comb];
  assign p9_res7__500_comb = p8_literal_1076345[p9_res7__499_comb] ^ p8_literal_1076347[p9_res7__498_comb] ^ p9_array_index_1085686_comb ^ p9_array_index_1085687_comb ^ p9_array_index_1085688_comb ^ p9_array_index_1085689_comb ^ p9_array_index_1085611_comb ^ p8_literal_1076358[p9_array_index_1085612_comb] ^ p9_array_index_1085613_comb ^ p9_array_index_1085630_comb ^ p8_literal_1076353[p9_array_index_1085631_comb] ^ p8_literal_1076351[p9_array_index_1085616_comb] ^ p8_literal_1076349[p9_array_index_1085633_comb] ^ p8_literal_1076347[p9_array_index_1085618_comb] ^ p8_literal_1076345[p9_array_index_1085619_comb] ^ p9_array_index_1085620_comb;
  assign p9_array_index_1085699_comb = p8_literal_1076349[p9_res7__498_comb];
  assign p9_array_index_1085700_comb = p8_literal_1076351[p9_res7__497_comb];
  assign p9_array_index_1085701_comb = p8_literal_1076353[p9_res7__496_comb];
  assign p9_array_index_1085702_comb = p8_literal_1076355[p9_array_index_1085609_comb];
  assign p9_res7__501_comb = p8_literal_1076345[p9_res7__500_comb] ^ p8_literal_1076347[p9_res7__499_comb] ^ p9_array_index_1085699_comb ^ p9_array_index_1085700_comb ^ p9_array_index_1085701_comb ^ p9_array_index_1085702_comb ^ p9_array_index_1085610_comb ^ p8_literal_1076358[p9_array_index_1085611_comb] ^ p9_array_index_1085612_comb ^ p9_array_index_1085647_comb ^ p8_literal_1076353[p9_array_index_1085614_comb] ^ p8_literal_1076351[p9_array_index_1085631_comb] ^ p8_literal_1076349[p9_array_index_1085616_comb] ^ p8_literal_1076347[p9_array_index_1085633_comb] ^ p8_literal_1076345[p9_array_index_1085618_comb] ^ p9_array_index_1085619_comb;
  assign p9_array_index_1085713_comb = p8_literal_1076351[p9_res7__498_comb];
  assign p9_array_index_1085714_comb = p8_literal_1076353[p9_res7__497_comb];
  assign p9_array_index_1085715_comb = p8_literal_1076355[p9_res7__496_comb];
  assign p9_res7__502_comb = p8_literal_1076345[p9_res7__501_comb] ^ p8_literal_1076347[p9_res7__500_comb] ^ p8_literal_1076349[p9_res7__499_comb] ^ p9_array_index_1085713_comb ^ p9_array_index_1085714_comb ^ p9_array_index_1085715_comb ^ p9_array_index_1085609_comb ^ p8_literal_1076358[p9_array_index_1085610_comb] ^ p9_array_index_1085611_comb ^ p9_array_index_1085661_comb ^ p9_array_index_1085629_comb ^ p8_literal_1076351[p9_array_index_1085614_comb] ^ p8_literal_1076349[p9_array_index_1085631_comb] ^ p8_literal_1076347[p9_array_index_1085616_comb] ^ p8_literal_1076345[p9_array_index_1085633_comb] ^ p9_array_index_1085618_comb;
  assign p9_array_index_1085725_comb = p8_literal_1076351[p9_res7__499_comb];
  assign p9_array_index_1085726_comb = p8_literal_1076353[p9_res7__498_comb];
  assign p9_array_index_1085727_comb = p8_literal_1076355[p9_res7__497_comb];
  assign p9_res7__503_comb = p8_literal_1076345[p9_res7__502_comb] ^ p8_literal_1076347[p9_res7__501_comb] ^ p8_literal_1076349[p9_res7__500_comb] ^ p9_array_index_1085725_comb ^ p9_array_index_1085726_comb ^ p9_array_index_1085727_comb ^ p9_res7__496_comb ^ p8_literal_1076358[p9_array_index_1085609_comb] ^ p9_array_index_1085610_comb ^ p9_array_index_1085675_comb ^ p9_array_index_1085646_comb ^ p8_literal_1076351[p9_array_index_1085613_comb] ^ p8_literal_1076349[p9_array_index_1085614_comb] ^ p8_literal_1076347[p9_array_index_1085631_comb] ^ p8_literal_1076345[p9_array_index_1085616_comb] ^ p9_array_index_1085633_comb;
  assign p9_array_index_1085738_comb = p8_literal_1076353[p9_res7__499_comb];
  assign p9_array_index_1085739_comb = p8_literal_1076355[p9_res7__498_comb];
  assign p9_res7__504_comb = p8_literal_1076345[p9_res7__503_comb] ^ p8_literal_1076347[p9_res7__502_comb] ^ p8_literal_1076349[p9_res7__501_comb] ^ p8_literal_1076351[p9_res7__500_comb] ^ p9_array_index_1085738_comb ^ p9_array_index_1085739_comb ^ p9_res7__497_comb ^ p8_literal_1076358[p9_res7__496_comb] ^ p9_array_index_1085609_comb ^ p9_array_index_1085689_comb ^ p9_array_index_1085660_comb ^ p9_array_index_1085628_comb ^ p8_literal_1076349[p9_array_index_1085613_comb] ^ p8_literal_1076347[p9_array_index_1085614_comb] ^ p8_literal_1076345[p9_array_index_1085631_comb] ^ p9_array_index_1085616_comb;
  assign p9_array_index_1085749_comb = p8_literal_1076353[p9_res7__500_comb];
  assign p9_array_index_1085750_comb = p8_literal_1076355[p9_res7__499_comb];
  assign p9_res7__505_comb = p8_literal_1076345[p9_res7__504_comb] ^ p8_literal_1076347[p9_res7__503_comb] ^ p8_literal_1076349[p9_res7__502_comb] ^ p8_literal_1076351[p9_res7__501_comb] ^ p9_array_index_1085749_comb ^ p9_array_index_1085750_comb ^ p9_res7__498_comb ^ p8_literal_1076358[p9_res7__497_comb] ^ p9_res7__496_comb ^ p9_array_index_1085702_comb ^ p9_array_index_1085674_comb ^ p9_array_index_1085645_comb ^ p8_literal_1076349[p9_array_index_1085612_comb] ^ p8_literal_1076347[p9_array_index_1085613_comb] ^ p8_literal_1076345[p9_array_index_1085614_comb] ^ p9_array_index_1085631_comb;
  assign p9_array_index_1085761_comb = p8_literal_1076355[p9_res7__500_comb];
  assign p9_res7__506_comb = p8_literal_1076345[p9_res7__505_comb] ^ p8_literal_1076347[p9_res7__504_comb] ^ p8_literal_1076349[p9_res7__503_comb] ^ p8_literal_1076351[p9_res7__502_comb] ^ p8_literal_1076353[p9_res7__501_comb] ^ p9_array_index_1085761_comb ^ p9_res7__499_comb ^ p8_literal_1076358[p9_res7__498_comb] ^ p9_res7__497_comb ^ p9_array_index_1085715_comb ^ p9_array_index_1085688_comb ^ p9_array_index_1085659_comb ^ p9_array_index_1085627_comb ^ p8_literal_1076347[p9_array_index_1085612_comb] ^ p8_literal_1076345[p9_array_index_1085613_comb] ^ p9_array_index_1085614_comb;
  assign p9_array_index_1085771_comb = p8_literal_1076355[p9_res7__501_comb];
  assign p9_res7__507_comb = p8_literal_1076345[p9_res7__506_comb] ^ p8_literal_1076347[p9_res7__505_comb] ^ p8_literal_1076349[p9_res7__504_comb] ^ p8_literal_1076351[p9_res7__503_comb] ^ p8_literal_1076353[p9_res7__502_comb] ^ p9_array_index_1085771_comb ^ p9_res7__500_comb ^ p8_literal_1076358[p9_res7__499_comb] ^ p9_res7__498_comb ^ p9_array_index_1085727_comb ^ p9_array_index_1085701_comb ^ p9_array_index_1085673_comb ^ p9_array_index_1085644_comb ^ p8_literal_1076347[p9_array_index_1085611_comb] ^ p8_literal_1076345[p9_array_index_1085612_comb] ^ p9_array_index_1085613_comb;
  assign p9_res7__508_comb = p8_literal_1076345[p9_res7__507_comb] ^ p8_literal_1076347[p9_res7__506_comb] ^ p8_literal_1076349[p9_res7__505_comb] ^ p8_literal_1076351[p9_res7__504_comb] ^ p8_literal_1076353[p9_res7__503_comb] ^ p8_literal_1076355[p9_res7__502_comb] ^ p9_res7__501_comb ^ p8_literal_1076358[p9_res7__500_comb] ^ p9_res7__499_comb ^ p9_array_index_1085739_comb ^ p9_array_index_1085714_comb ^ p9_array_index_1085687_comb ^ p9_array_index_1085658_comb ^ p9_array_index_1085626_comb ^ p8_literal_1076345[p9_array_index_1085611_comb] ^ p9_array_index_1085612_comb;
  assign p9_res7__509_comb = p8_literal_1076345[p9_res7__508_comb] ^ p8_literal_1076347[p9_res7__507_comb] ^ p8_literal_1076349[p9_res7__506_comb] ^ p8_literal_1076351[p9_res7__505_comb] ^ p8_literal_1076353[p9_res7__504_comb] ^ p8_literal_1076355[p9_res7__503_comb] ^ p9_res7__502_comb ^ p8_literal_1076358[p9_res7__501_comb] ^ p9_res7__500_comb ^ p9_array_index_1085750_comb ^ p9_array_index_1085726_comb ^ p9_array_index_1085700_comb ^ p9_array_index_1085672_comb ^ p9_array_index_1085643_comb ^ p8_literal_1076345[p9_array_index_1085610_comb] ^ p9_array_index_1085611_comb;
  assign p9_res7__510_comb = p8_literal_1076345[p9_res7__509_comb] ^ p8_literal_1076347[p9_res7__508_comb] ^ p8_literal_1076349[p9_res7__507_comb] ^ p8_literal_1076351[p9_res7__506_comb] ^ p8_literal_1076353[p9_res7__505_comb] ^ p8_literal_1076355[p9_res7__504_comb] ^ p9_res7__503_comb ^ p8_literal_1076358[p9_res7__502_comb] ^ p9_res7__501_comb ^ p9_array_index_1085761_comb ^ p9_array_index_1085738_comb ^ p9_array_index_1085713_comb ^ p9_array_index_1085686_comb ^ p9_array_index_1085657_comb ^ p9_array_index_1085625_comb ^ p9_array_index_1085610_comb;
  assign p9_res7__511_comb = p8_literal_1076345[p9_res7__510_comb] ^ p8_literal_1076347[p9_res7__509_comb] ^ p8_literal_1076349[p9_res7__508_comb] ^ p8_literal_1076351[p9_res7__507_comb] ^ p8_literal_1076353[p9_res7__506_comb] ^ p8_literal_1076355[p9_res7__505_comb] ^ p9_res7__504_comb ^ p8_literal_1076358[p9_res7__503_comb] ^ p9_res7__502_comb ^ p9_array_index_1085771_comb ^ p9_array_index_1085749_comb ^ p9_array_index_1085725_comb ^ p9_array_index_1085699_comb ^ p9_array_index_1085671_comb ^ p9_array_index_1085642_comb ^ p9_array_index_1085609_comb;
  assign p9_res__31_comb = {p9_res7__511_comb, p9_res7__510_comb, p9_res7__509_comb, p9_res7__508_comb, p9_res7__507_comb, p9_res7__506_comb, p9_res7__505_comb, p9_res7__504_comb, p9_res7__503_comb, p9_res7__502_comb, p9_res7__501_comb, p9_res7__500_comb, p9_res7__499_comb, p9_res7__498_comb, p9_res7__497_comb, p9_res7__496_comb};
  assign p9_addedKey__40_comb = p9_res__31_comb ^ p9_xor_1085375_comb ^ p8_res__39;
  assign p9_array_index_1085825_comb = p8_arr[p9_addedKey__40_comb[127:120]];
  assign p9_array_index_1085826_comb = p8_arr[p9_addedKey__40_comb[119:112]];
  assign p9_array_index_1085827_comb = p8_arr[p9_addedKey__40_comb[111:104]];
  assign p9_array_index_1085828_comb = p8_arr[p9_addedKey__40_comb[103:96]];
  assign p9_array_index_1085829_comb = p8_arr[p9_addedKey__40_comb[95:88]];
  assign p9_array_index_1085830_comb = p8_arr[p9_addedKey__40_comb[87:80]];
  assign p9_array_index_1085832_comb = p8_arr[p9_addedKey__40_comb[71:64]];
  assign p9_array_index_1085834_comb = p8_arr[p9_addedKey__40_comb[55:48]];
  assign p9_array_index_1085835_comb = p8_arr[p9_addedKey__40_comb[47:40]];
  assign p9_array_index_1085836_comb = p8_arr[p9_addedKey__40_comb[39:32]];
  assign p9_array_index_1085837_comb = p8_arr[p9_addedKey__40_comb[31:24]];
  assign p9_array_index_1085838_comb = p8_arr[p9_addedKey__40_comb[23:16]];
  assign p9_array_index_1085839_comb = p8_arr[p9_addedKey__40_comb[15:8]];
  assign p9_array_index_1085841_comb = p8_literal_1076345[p9_array_index_1085825_comb];
  assign p9_array_index_1085842_comb = p8_literal_1076347[p9_array_index_1085826_comb];
  assign p9_array_index_1085843_comb = p8_literal_1076349[p9_array_index_1085827_comb];
  assign p9_array_index_1085844_comb = p8_literal_1076351[p9_array_index_1085828_comb];
  assign p9_array_index_1085845_comb = p8_literal_1076353[p9_array_index_1085829_comb];
  assign p9_array_index_1085846_comb = p8_literal_1076355[p9_array_index_1085830_comb];
  assign p9_array_index_1085847_comb = p8_arr[p9_addedKey__40_comb[79:72]];
  assign p9_array_index_1085849_comb = p8_arr[p9_addedKey__40_comb[63:56]];
  assign p9_res7__640_comb = p9_array_index_1085841_comb ^ p9_array_index_1085842_comb ^ p9_array_index_1085843_comb ^ p9_array_index_1085844_comb ^ p9_array_index_1085845_comb ^ p9_array_index_1085846_comb ^ p9_array_index_1085847_comb ^ p8_literal_1076358[p9_array_index_1085832_comb] ^ p9_array_index_1085849_comb ^ p8_literal_1076355[p9_array_index_1085834_comb] ^ p8_literal_1076353[p9_array_index_1085835_comb] ^ p8_literal_1076351[p9_array_index_1085836_comb] ^ p8_literal_1076349[p9_array_index_1085837_comb] ^ p8_literal_1076347[p9_array_index_1085838_comb] ^ p8_literal_1076345[p9_array_index_1085839_comb] ^ p8_arr[p9_addedKey__40_comb[7:0]];
  assign p9_array_index_1085858_comb = p8_literal_1076345[p9_res7__640_comb];
  assign p9_array_index_1085859_comb = p8_literal_1076347[p9_array_index_1085825_comb];
  assign p9_array_index_1085860_comb = p8_literal_1076349[p9_array_index_1085826_comb];
  assign p9_array_index_1085861_comb = p8_literal_1076351[p9_array_index_1085827_comb];
  assign p9_array_index_1085862_comb = p8_literal_1076353[p9_array_index_1085828_comb];
  assign p9_array_index_1085863_comb = p8_literal_1076355[p9_array_index_1085829_comb];
  assign p9_res7__641_comb = p9_array_index_1085858_comb ^ p9_array_index_1085859_comb ^ p9_array_index_1085860_comb ^ p9_array_index_1085861_comb ^ p9_array_index_1085862_comb ^ p9_array_index_1085863_comb ^ p9_array_index_1085830_comb ^ p8_literal_1076358[p9_array_index_1085847_comb] ^ p9_array_index_1085832_comb ^ p8_literal_1076355[p9_array_index_1085849_comb] ^ p8_literal_1076353[p9_array_index_1085834_comb] ^ p8_literal_1076351[p9_array_index_1085835_comb] ^ p8_literal_1076349[p9_array_index_1085836_comb] ^ p8_literal_1076347[p9_array_index_1085837_comb] ^ p8_literal_1076345[p9_array_index_1085838_comb] ^ p9_array_index_1085839_comb;
  assign p9_array_index_1085873_comb = p8_literal_1076347[p9_res7__640_comb];
  assign p9_array_index_1085874_comb = p8_literal_1076349[p9_array_index_1085825_comb];
  assign p9_array_index_1085875_comb = p8_literal_1076351[p9_array_index_1085826_comb];
  assign p9_array_index_1085876_comb = p8_literal_1076353[p9_array_index_1085827_comb];
  assign p9_array_index_1085877_comb = p8_literal_1076355[p9_array_index_1085828_comb];
  assign p9_res7__642_comb = p8_literal_1076345[p9_res7__641_comb] ^ p9_array_index_1085873_comb ^ p9_array_index_1085874_comb ^ p9_array_index_1085875_comb ^ p9_array_index_1085876_comb ^ p9_array_index_1085877_comb ^ p9_array_index_1085829_comb ^ p8_literal_1076358[p9_array_index_1085830_comb] ^ p9_array_index_1085847_comb ^ p8_literal_1076355[p9_array_index_1085832_comb] ^ p8_literal_1076353[p9_array_index_1085849_comb] ^ p8_literal_1076351[p9_array_index_1085834_comb] ^ p8_literal_1076349[p9_array_index_1085835_comb] ^ p8_literal_1076347[p9_array_index_1085836_comb] ^ p8_literal_1076345[p9_array_index_1085837_comb] ^ p9_array_index_1085838_comb;
  assign p9_array_index_1085887_comb = p8_literal_1076347[p9_res7__641_comb];
  assign p9_array_index_1085888_comb = p8_literal_1076349[p9_res7__640_comb];
  assign p9_array_index_1085889_comb = p8_literal_1076351[p9_array_index_1085825_comb];
  assign p9_array_index_1085890_comb = p8_literal_1076353[p9_array_index_1085826_comb];
  assign p9_array_index_1085891_comb = p8_literal_1076355[p9_array_index_1085827_comb];
  assign p9_res7__643_comb = p8_literal_1076345[p9_res7__642_comb] ^ p9_array_index_1085887_comb ^ p9_array_index_1085888_comb ^ p9_array_index_1085889_comb ^ p9_array_index_1085890_comb ^ p9_array_index_1085891_comb ^ p9_array_index_1085828_comb ^ p8_literal_1076358[p9_array_index_1085829_comb] ^ p9_array_index_1085830_comb ^ p8_literal_1076355[p9_array_index_1085847_comb] ^ p8_literal_1076353[p9_array_index_1085832_comb] ^ p8_literal_1076351[p9_array_index_1085849_comb] ^ p8_literal_1076349[p9_array_index_1085834_comb] ^ p8_literal_1076347[p9_array_index_1085835_comb] ^ p8_literal_1076345[p9_array_index_1085836_comb] ^ p9_array_index_1085837_comb;
  assign p9_array_index_1085902_comb = p8_literal_1076349[p9_res7__641_comb];
  assign p9_array_index_1085903_comb = p8_literal_1076351[p9_res7__640_comb];
  assign p9_array_index_1085904_comb = p8_literal_1076353[p9_array_index_1085825_comb];
  assign p9_array_index_1085905_comb = p8_literal_1076355[p9_array_index_1085826_comb];
  assign p9_res7__644_comb = p8_literal_1076345[p9_res7__643_comb] ^ p8_literal_1076347[p9_res7__642_comb] ^ p9_array_index_1085902_comb ^ p9_array_index_1085903_comb ^ p9_array_index_1085904_comb ^ p9_array_index_1085905_comb ^ p9_array_index_1085827_comb ^ p8_literal_1076358[p9_array_index_1085828_comb] ^ p9_array_index_1085829_comb ^ p9_array_index_1085846_comb ^ p8_literal_1076353[p9_array_index_1085847_comb] ^ p8_literal_1076351[p9_array_index_1085832_comb] ^ p8_literal_1076349[p9_array_index_1085849_comb] ^ p8_literal_1076347[p9_array_index_1085834_comb] ^ p8_literal_1076345[p9_array_index_1085835_comb] ^ p9_array_index_1085836_comb;
  assign p9_array_index_1085915_comb = p8_literal_1076349[p9_res7__642_comb];
  assign p9_array_index_1085916_comb = p8_literal_1076351[p9_res7__641_comb];
  assign p9_array_index_1085917_comb = p8_literal_1076353[p9_res7__640_comb];
  assign p9_array_index_1085918_comb = p8_literal_1076355[p9_array_index_1085825_comb];
  assign p9_res7__645_comb = p8_literal_1076345[p9_res7__644_comb] ^ p8_literal_1076347[p9_res7__643_comb] ^ p9_array_index_1085915_comb ^ p9_array_index_1085916_comb ^ p9_array_index_1085917_comb ^ p9_array_index_1085918_comb ^ p9_array_index_1085826_comb ^ p8_literal_1076358[p9_array_index_1085827_comb] ^ p9_array_index_1085828_comb ^ p9_array_index_1085863_comb ^ p8_literal_1076353[p9_array_index_1085830_comb] ^ p8_literal_1076351[p9_array_index_1085847_comb] ^ p8_literal_1076349[p9_array_index_1085832_comb] ^ p8_literal_1076347[p9_array_index_1085849_comb] ^ p8_literal_1076345[p9_array_index_1085834_comb] ^ p9_array_index_1085835_comb;
  assign p9_array_index_1085929_comb = p8_literal_1076351[p9_res7__642_comb];
  assign p9_array_index_1085930_comb = p8_literal_1076353[p9_res7__641_comb];
  assign p9_array_index_1085931_comb = p8_literal_1076355[p9_res7__640_comb];
  assign p9_res7__646_comb = p8_literal_1076345[p9_res7__645_comb] ^ p8_literal_1076347[p9_res7__644_comb] ^ p8_literal_1076349[p9_res7__643_comb] ^ p9_array_index_1085929_comb ^ p9_array_index_1085930_comb ^ p9_array_index_1085931_comb ^ p9_array_index_1085825_comb ^ p8_literal_1076358[p9_array_index_1085826_comb] ^ p9_array_index_1085827_comb ^ p9_array_index_1085877_comb ^ p9_array_index_1085845_comb ^ p8_literal_1076351[p9_array_index_1085830_comb] ^ p8_literal_1076349[p9_array_index_1085847_comb] ^ p8_literal_1076347[p9_array_index_1085832_comb] ^ p8_literal_1076345[p9_array_index_1085849_comb] ^ p9_array_index_1085834_comb;
  assign p9_array_index_1085941_comb = p8_literal_1076351[p9_res7__643_comb];
  assign p9_array_index_1085942_comb = p8_literal_1076353[p9_res7__642_comb];
  assign p9_array_index_1085943_comb = p8_literal_1076355[p9_res7__641_comb];
  assign p9_res7__647_comb = p8_literal_1076345[p9_res7__646_comb] ^ p8_literal_1076347[p9_res7__645_comb] ^ p8_literal_1076349[p9_res7__644_comb] ^ p9_array_index_1085941_comb ^ p9_array_index_1085942_comb ^ p9_array_index_1085943_comb ^ p9_res7__640_comb ^ p8_literal_1076358[p9_array_index_1085825_comb] ^ p9_array_index_1085826_comb ^ p9_array_index_1085891_comb ^ p9_array_index_1085862_comb ^ p8_literal_1076351[p9_array_index_1085829_comb] ^ p8_literal_1076349[p9_array_index_1085830_comb] ^ p8_literal_1076347[p9_array_index_1085847_comb] ^ p8_literal_1076345[p9_array_index_1085832_comb] ^ p9_array_index_1085849_comb;
  assign p9_array_index_1085954_comb = p8_literal_1076353[p9_res7__643_comb];
  assign p9_array_index_1085955_comb = p8_literal_1076355[p9_res7__642_comb];
  assign p9_res7__648_comb = p8_literal_1076345[p9_res7__647_comb] ^ p8_literal_1076347[p9_res7__646_comb] ^ p8_literal_1076349[p9_res7__645_comb] ^ p8_literal_1076351[p9_res7__644_comb] ^ p9_array_index_1085954_comb ^ p9_array_index_1085955_comb ^ p9_res7__641_comb ^ p8_literal_1076358[p9_res7__640_comb] ^ p9_array_index_1085825_comb ^ p9_array_index_1085905_comb ^ p9_array_index_1085876_comb ^ p9_array_index_1085844_comb ^ p8_literal_1076349[p9_array_index_1085829_comb] ^ p8_literal_1076347[p9_array_index_1085830_comb] ^ p8_literal_1076345[p9_array_index_1085847_comb] ^ p9_array_index_1085832_comb;
  assign p9_array_index_1085965_comb = p8_literal_1076353[p9_res7__644_comb];
  assign p9_array_index_1085966_comb = p8_literal_1076355[p9_res7__643_comb];
  assign p9_res7__649_comb = p8_literal_1076345[p9_res7__648_comb] ^ p8_literal_1076347[p9_res7__647_comb] ^ p8_literal_1076349[p9_res7__646_comb] ^ p8_literal_1076351[p9_res7__645_comb] ^ p9_array_index_1085965_comb ^ p9_array_index_1085966_comb ^ p9_res7__642_comb ^ p8_literal_1076358[p9_res7__641_comb] ^ p9_res7__640_comb ^ p9_array_index_1085918_comb ^ p9_array_index_1085890_comb ^ p9_array_index_1085861_comb ^ p8_literal_1076349[p9_array_index_1085828_comb] ^ p8_literal_1076347[p9_array_index_1085829_comb] ^ p8_literal_1076345[p9_array_index_1085830_comb] ^ p9_array_index_1085847_comb;
  assign p9_array_index_1085977_comb = p8_literal_1076355[p9_res7__644_comb];
  assign p9_res7__650_comb = p8_literal_1076345[p9_res7__649_comb] ^ p8_literal_1076347[p9_res7__648_comb] ^ p8_literal_1076349[p9_res7__647_comb] ^ p8_literal_1076351[p9_res7__646_comb] ^ p8_literal_1076353[p9_res7__645_comb] ^ p9_array_index_1085977_comb ^ p9_res7__643_comb ^ p8_literal_1076358[p9_res7__642_comb] ^ p9_res7__641_comb ^ p9_array_index_1085931_comb ^ p9_array_index_1085904_comb ^ p9_array_index_1085875_comb ^ p9_array_index_1085843_comb ^ p8_literal_1076347[p9_array_index_1085828_comb] ^ p8_literal_1076345[p9_array_index_1085829_comb] ^ p9_array_index_1085830_comb;
  assign p9_array_index_1085987_comb = p8_literal_1076355[p9_res7__645_comb];
  assign p9_res7__651_comb = p8_literal_1076345[p9_res7__650_comb] ^ p8_literal_1076347[p9_res7__649_comb] ^ p8_literal_1076349[p9_res7__648_comb] ^ p8_literal_1076351[p9_res7__647_comb] ^ p8_literal_1076353[p9_res7__646_comb] ^ p9_array_index_1085987_comb ^ p9_res7__644_comb ^ p8_literal_1076358[p9_res7__643_comb] ^ p9_res7__642_comb ^ p9_array_index_1085943_comb ^ p9_array_index_1085917_comb ^ p9_array_index_1085889_comb ^ p9_array_index_1085860_comb ^ p8_literal_1076347[p9_array_index_1085827_comb] ^ p8_literal_1076345[p9_array_index_1085828_comb] ^ p9_array_index_1085829_comb;
  assign p9_res7__652_comb = p8_literal_1076345[p9_res7__651_comb] ^ p8_literal_1076347[p9_res7__650_comb] ^ p8_literal_1076349[p9_res7__649_comb] ^ p8_literal_1076351[p9_res7__648_comb] ^ p8_literal_1076353[p9_res7__647_comb] ^ p8_literal_1076355[p9_res7__646_comb] ^ p9_res7__645_comb ^ p8_literal_1076358[p9_res7__644_comb] ^ p9_res7__643_comb ^ p9_array_index_1085955_comb ^ p9_array_index_1085930_comb ^ p9_array_index_1085903_comb ^ p9_array_index_1085874_comb ^ p9_array_index_1085842_comb ^ p8_literal_1076345[p9_array_index_1085827_comb] ^ p9_array_index_1085828_comb;
  assign p9_res7__653_comb = p8_literal_1076345[p9_res7__652_comb] ^ p8_literal_1076347[p9_res7__651_comb] ^ p8_literal_1076349[p9_res7__650_comb] ^ p8_literal_1076351[p9_res7__649_comb] ^ p8_literal_1076353[p9_res7__648_comb] ^ p8_literal_1076355[p9_res7__647_comb] ^ p9_res7__646_comb ^ p8_literal_1076358[p9_res7__645_comb] ^ p9_res7__644_comb ^ p9_array_index_1085966_comb ^ p9_array_index_1085942_comb ^ p9_array_index_1085916_comb ^ p9_array_index_1085888_comb ^ p9_array_index_1085859_comb ^ p8_literal_1076345[p9_array_index_1085826_comb] ^ p9_array_index_1085827_comb;
  assign p9_res7__654_comb = p8_literal_1076345[p9_res7__653_comb] ^ p8_literal_1076347[p9_res7__652_comb] ^ p8_literal_1076349[p9_res7__651_comb] ^ p8_literal_1076351[p9_res7__650_comb] ^ p8_literal_1076353[p9_res7__649_comb] ^ p8_literal_1076355[p9_res7__648_comb] ^ p9_res7__647_comb ^ p8_literal_1076358[p9_res7__646_comb] ^ p9_res7__645_comb ^ p9_array_index_1085977_comb ^ p9_array_index_1085954_comb ^ p9_array_index_1085929_comb ^ p9_array_index_1085902_comb ^ p9_array_index_1085873_comb ^ p9_array_index_1085841_comb ^ p9_array_index_1085826_comb;
  assign p9_res7__655_comb = p8_literal_1076345[p9_res7__654_comb] ^ p8_literal_1076347[p9_res7__653_comb] ^ p8_literal_1076349[p9_res7__652_comb] ^ p8_literal_1076351[p9_res7__651_comb] ^ p8_literal_1076353[p9_res7__650_comb] ^ p8_literal_1076355[p9_res7__649_comb] ^ p9_res7__648_comb ^ p8_literal_1076358[p9_res7__647_comb] ^ p9_res7__646_comb ^ p9_array_index_1085987_comb ^ p9_array_index_1085965_comb ^ p9_array_index_1085941_comb ^ p9_array_index_1085915_comb ^ p9_array_index_1085887_comb ^ p9_array_index_1085858_comb ^ p9_array_index_1085825_comb;
  assign p9_newValue_comb = {p9_res7__655_comb, p9_res7__654_comb, p9_res7__653_comb, p9_res7__652_comb, p9_res7__651_comb, p9_res7__650_comb, p9_res7__649_comb, p9_res7__648_comb, p9_res7__647_comb, p9_res7__646_comb, p9_res7__645_comb, p9_res7__644_comb, p9_res7__643_comb, p9_res7__642_comb, p9_res7__641_comb, p9_res7__640_comb};
  assign p9_xor_1086027_comb = p9_newValue_comb ^ p9_k9_comb;

  // Registers for pipe stage 9:
  reg [127:0] p9_xor_1086027;
  always_ff @ (posedge clk) begin
    p9_xor_1086027 <= p9_xor_1086027_comb;
  end
  assign out = p9_xor_1086027;
endmodule
