module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , 
 n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , 
 n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , 
 n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , 
 n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , 
 n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , 
 n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , 
 n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , 
 n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , 
 n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , 
 n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , 
 n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , 
 n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , 
 n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , 
 n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , 
 n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , 
 n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
 n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
 n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , 
 n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , 
 n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , 
 n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , 
 n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , 
 n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , 
 n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , 
 n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , 
 n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , 
 n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , 
 n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , 
 n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , 
 n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , 
 n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , 
 n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , 
 n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , 
 n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , 
 n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , 
 n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , 
 n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , 
 n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , 
 n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , 
 n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , 
 n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , 
 n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , 
 n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
 n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
 n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
 n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , 
 n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , 
 n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , 
 n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , 
 n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , 
 n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , 
 n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , 
 n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , 
 n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , 
 n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , 
 n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , 
 n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , 
 n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , 
 n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , 
 n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , 
 n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , 
 n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , 
 n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , 
 n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , 
 n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , 
 n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , 
 n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , 
 n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , 
 n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , 
 n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , 
 n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
 n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
 n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
 n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
 n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
 n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
 n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
 n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
 n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
 n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
 n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
 n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
 n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
 n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , 
 n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , 
 n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , 
 n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , 
 n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , 
 n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , 
 n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , 
 n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , 
 n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , 
 n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , 
 n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , 
 n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
 n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
 n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , 
 n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , 
 n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , 
 n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , 
 n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
 n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , 
 n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , 
 n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , 
 n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , 
 n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , 
 n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , 
 n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , 
 n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , 
 n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , 
 n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , 
 n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , 
 n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , 
 n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , 
 n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , 
 n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , 
 n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , 
 n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , 
 n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , 
 n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , 
 n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , 
 n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , 
 n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , 
 n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , 
 n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , 
 n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , 
 n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , 
 n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , 
 n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , 
 n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , 
 n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , 
 n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , 
 n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , 
 n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , 
 n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , 
 n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , 
 n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , 
 n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , 
 n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , 
 n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , 
 n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
 n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
 n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , 
 n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , 
 n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , 
 n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , 
 n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , 
 n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , 
 n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , 
 n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , 
 n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , 
 n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , 
 n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , 
 n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , 
 n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , 
 n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , 
 n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , 
 n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
 n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , 
 n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , 
 n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , 
 n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , 
 n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , 
 n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , 
 n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , 
 n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , 
 n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , 
 n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , 
 n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , 
 n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , 
 n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , 
 n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , 
 n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , 
 n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , 
 n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , 
 n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , 
 n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , 
 n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , 
 n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , 
 n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , 
 n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , 
 n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , 
 n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , 
 n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , 
 n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , 
 n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , 
 n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , 
 n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , 
 n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , 
 n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , 
 n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , 
 n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , 
 n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , 
 n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , 
 n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , 
 n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , 
 n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , 
 n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , 
 n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , 
 n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , 
 n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , 
 n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , 
 n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , 
 n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , 
 n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , 
 n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , 
 n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , 
 n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , 
 n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , 
 n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , 
 n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , 
 n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , 
 n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , 
 n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , 
 n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , 
 n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , 
 n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , 
 n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , 
 n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , 
 n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , 
 n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , 
 n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , 
 n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , 
 n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , 
 n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , 
 n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , 
 n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , 
 n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , 
 n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , 
 n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , 
 n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , 
 n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , 
 n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , 
 n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , 
 n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , 
 n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , 
 n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , 
 n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , 
 n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , 
 n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , 
 n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , 
 n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , 
 n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , 
 n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , 
 n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , 
 n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , 
 n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , 
 n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , 
 n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , 
 n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , 
 n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , 
 n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , 
 n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , 
 n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , 
 n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , 
 n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , 
 n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , 
 n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , 
 n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , 
 n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , 
 n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , 
 n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , 
 n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , 
 n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , 
 n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , 
 n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , 
 n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , 
 n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
 n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , 
 n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , 
 n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , 
 n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , 
 n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , 
 n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , 
 n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , 
 n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , 
 n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , 
 n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , 
 n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , 
 n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , 
 n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , 
 n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , 
 n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , 
 n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , 
 n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , 
 n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , 
 n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , 
 n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , 
 n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , 
 n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , 
 n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , 
 n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , 
 n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , 
 n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , 
 n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , 
 n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , 
 n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , 
 n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , 
 n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , 
 n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
 n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , 
 n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , 
 n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , 
 n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , 
 n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , 
 n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , 
 n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , 
 n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , 
 n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , 
 n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , 
 n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , 
 n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
 n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , 
 n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , 
 n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , 
 n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , 
 n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , 
 n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , 
 n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , 
 n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , 
 n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , 
 n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , 
 n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , 
 n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , 
 n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , 
 n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
 n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
 n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
 n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , 
 n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , 
 n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , 
 n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , 
 n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , 
 n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , 
 n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , 
 n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , 
 n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , 
 n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , 
 n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , 
 n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , 
 n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , 
 n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , 
 n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , 
 n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , 
 n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , 
 n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , 
 n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , 
 n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , 
 n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , 
 n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , 
 n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , 
 n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , 
 n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , 
 n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , 
 n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , 
 n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , 
 n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , 
 n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , 
 n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , 
 n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , 
 n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , 
 n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , 
 n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , 
 n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , 
 n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , 
 n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , 
 n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , 
 n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , 
 n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , 
 n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , 
 n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , 
 n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , 
 n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , 
 n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , 
 n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , 
 n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , 
 n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , 
 n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , 
 n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , 
 n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , 
 n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , 
 n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , 
 n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , 
 n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , 
 n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , 
 n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , 
 n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , 
 n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , 
 n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , 
 n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , 
 n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , 
 n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , 
 n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , 
 n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , 
 n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , 
 n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , 
 n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , 
 n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , 
 n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , 
 n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , 
 n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , 
 n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , 
 n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , 
 n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , 
 n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , 
 n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , 
 n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , 
 n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , 
 n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , 
 n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , 
 n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , 
 n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , 
 n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , 
 n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , 
 n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , 
 n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , 
 n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
 n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
 n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , 
 n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , 
 n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , 
 n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , 
 n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , 
 n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , 
 n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , 
 n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , 
 n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , 
 n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , 
 n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , 
 n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , 
 n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
 n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , 
 n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , 
 n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , 
 n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , 
 n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , 
 n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , 
 n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , 
 n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , 
 n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , 
 n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , 
 n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , 
 n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , 
 n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , 
 n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , 
 n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , 
 n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , 
 n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
 n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , 
 n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , 
 n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , 
 n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , 
 n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
 n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
 n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
 n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
 n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
 n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
 n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
 n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
 n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
 n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
 n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
 n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
 n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
 n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
 n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
 n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
 n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
 n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
 n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
 n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
 n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
 n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
 n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
 n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
 n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
 n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
 n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
 n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , 
 n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
 n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
 n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
 n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
 n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
 n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
 n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , 
 n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , 
 n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , 
 n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , 
 n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , 
 n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , 
 n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , 
 n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , 
 n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , 
 n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , 
 n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , 
 n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , 
 n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , 
 n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , 
 n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , 
 n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , 
 n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , 
 n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , 
 n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , 
 n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , 
 n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
 n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
 n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , 
 n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , 
 n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , 
 n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , 
 n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , 
 n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , 
 n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , 
 n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , 
 n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , 
 n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , 
 n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , 
 n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , 
 n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
 n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , 
 n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , 
 n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , 
 n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , 
 n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , 
 n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , 
 n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , 
 n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , 
 n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , 
 n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , 
 n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , 
 n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , 
 n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , 
 n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , 
 n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , 
 n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , 
 n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , 
 n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , 
 n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , 
 n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , 
 n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , 
 n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , 
 n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , 
 n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , 
 n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , 
 n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , 
 n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , 
 n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , 
 n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , 
 n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , 
 n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , 
 n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , 
 n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , 
 n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , 
 n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , 
 n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
 n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , 
 n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
 n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
 n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
 n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
 n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
 n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
 n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
 n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
 n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
 n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , 
 n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , 
 n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
 n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
 n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
 n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
 n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , 
 n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , 
 n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , 
 n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , 
 n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , 
 n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , 
 n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , 
 n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , 
 n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , 
 n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , 
 n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , 
 n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , 
 n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , 
 n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , 
 n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , 
 n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , 
 n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , 
 n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , 
 n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , 
 n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , 
 n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , 
 n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , 
 n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , 
 n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , 
 n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , 
 n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , 
 n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , 
 n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , 
 n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , 
 n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , 
 n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , 
 n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , 
 n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , 
 n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , 
 n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , 
 n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , 
 n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , 
 n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , 
 n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , 
 n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , 
 n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , 
 n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , 
 n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , 
 n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , 
 n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , 
 n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , 
 n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , 
 n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , 
 n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , 
 n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
 n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
 n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
 n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
 n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
 n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , 
 n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , 
 n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , 
 n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , 
 n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , 
 n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , 
 n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , 
 n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , 
 n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , 
 n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , 
 n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , 
 n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , 
 n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , 
 n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , 
 n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , 
 n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , 
 n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , 
 n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , 
 n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , 
 n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , 
 n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , 
 n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , 
 n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , 
 n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , 
 n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , 
 n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , 
 n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , 
 n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , 
 n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , 
 n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , 
 n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , 
 n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , 
 n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , 
 n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , 
 n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , 
 n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , 
 n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , 
 n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , 
 n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , 
 n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , 
 n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , 
 n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , 
 n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , 
 n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , 
 n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , 
 n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , 
 n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , 
 n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
 n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , 
 n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , 
 n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , 
 n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , 
 n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , 
 n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , 
 n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , 
 n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , 
 n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , 
 n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , 
 n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , 
 n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , 
 n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , 
 n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , 
 n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
 n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , 
 n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , 
 n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , 
 n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , 
 n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , 
 n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , 
 n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , 
 n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , 
 n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , 
 n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , 
 n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , 
 n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , 
 n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , 
 n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , 
 n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , 
 n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , 
 n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , 
 n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , 
 n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , 
 n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , 
 n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , 
 n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , 
 n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , 
 n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , 
 n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , 
 n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , 
 n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , 
 n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , 
 n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , 
 n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , 
 n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , 
 n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , 
 n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , 
 n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , 
 n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , 
 n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , 
 n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , 
 n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , 
 n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , 
 n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , 
 n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , 
 n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , 
 n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , 
 n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , 
 n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , 
 n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , 
 n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , 
 n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , 
 n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , 
 n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , 
 n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , 
 n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , 
 n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , 
 n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , 
 n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , 
 n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , 
 n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , 
 n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , 
 n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , 
 n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , 
 n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , 
 n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , 
 n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , 
 n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
 n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , 
 n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , 
 n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , 
 n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , 
 n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , 
 n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , 
 n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , 
 n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , 
 n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , 
 n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , 
 n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , 
 n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , 
 n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , 
 n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , 
 n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , 
 n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , 
 n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , 
 n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , 
 n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , 
 n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , 
 n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , 
 n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , 
 n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , 
 n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , 
 n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , 
 n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , 
 n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , 
 n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , 
 n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , 
 n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , 
 n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , 
 n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , 
 n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , 
 n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , 
 n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , 
 n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , 
 n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , 
 n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , 
 n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , 
 n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , 
 n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , 
 n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , 
 n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , 
 n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , 
 n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , 
 n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , 
 n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , 
 n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , 
 n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , 
 n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , 
 n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , 
 n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , 
 n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , 
 n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , 
 n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , 
 n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , 
 n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , 
 n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , 
 n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , 
 n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , 
 n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , 
 n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , 
 n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , 
 n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , 
 n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , 
 n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , 
 n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , 
 n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , 
 n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , 
 n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , 
 n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , 
 n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , 
 n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , 
 n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , 
 n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , 
 n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , 
 n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , 
 n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , 
 n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , 
 n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , 
 n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , 
 n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , 
 n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , 
 n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , 
 n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , 
 n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , 
 n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , 
 n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , 
 n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , 
 n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , 
 n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , 
 n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , 
 n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , 
 n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , 
 n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , 
 n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , 
 n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , 
 n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , 
 n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , 
 n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , 
 n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , 
 n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , 
 n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , 
 n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , 
 n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , 
 n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , 
 n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , 
 n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , 
 n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
 n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
 n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , 
 n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , 
 n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , 
 n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , 
 n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , 
 n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , 
 n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , 
 n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , 
 n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , 
 n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , 
 n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , 
 n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , 
 n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , 
 n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , 
 n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , 
 n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , 
 n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , 
 n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , 
 n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , 
 n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , 
 n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , 
 n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , 
 n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , 
 n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , 
 n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , 
 n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , 
 n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , 
 n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , 
 n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
 n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
 n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , 
 n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , 
 n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , 
 n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , 
 n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , 
 n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , 
 n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , 
 n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , 
 n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , 
 n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , 
 n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , 
 n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , 
 n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , 
 n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , 
 n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , 
 n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , 
 n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , 
 n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
 n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , 
 n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , 
 n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , 
 n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , 
 n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , 
 n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , 
 n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , 
 n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , 
 n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , 
 n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , 
 n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , 
 n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , 
 n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , 
 n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , 
 n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , 
 n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , 
 n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , 
 n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , 
 n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , 
 n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , 
 n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , 
 n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , 
 n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , 
 n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , 
 n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , 
 n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , 
 n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , 
 n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , 
 n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , 
 n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , 
 n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , 
 n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , 
 n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , 
 n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , 
 n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , 
 n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , 
 n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , 
 n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , 
 n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , 
 n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , 
 n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , 
 n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , 
 n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , 
 n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , 
 n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , 
 n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , 
 n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , 
 n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , 
 n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , 
 n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , 
 n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , 
 n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , 
 n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , 
 n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , 
 n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , 
 n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , 
 n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , 
 n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , 
 n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , 
 n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , 
 n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , 
 n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , 
 n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , 
 n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , 
 n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , 
 n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , 
 n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , 
 n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , 
 n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , 
 n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , 
 n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , 
 n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , 
 n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , 
 n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , 
 n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , 
 n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , 
 n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , 
 n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , 
 n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , 
 n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , 
 n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , 
 n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , 
 n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
 n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , 
 n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , 
 n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , 
 n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , 
 n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , 
 n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , 
 n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , 
 n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , 
 n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , 
 n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , 
 n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , 
 n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , 
 n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , 
 n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , 
 n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , 
 n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , 
 n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , 
 n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , 
 n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , 
 n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , 
 n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , 
 n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , 
 n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , 
 n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , 
 n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , 
 n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , 
 n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , 
 n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , 
 n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , 
 n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , 
 n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , 
 n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , 
 n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , 
 n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , 
 n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , 
 n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , 
 n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , 
 n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , 
 n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , 
 n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , 
 n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , 
 n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , 
 n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , 
 n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , 
 n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , 
 n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , 
 n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , 
 n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , 
 n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , 
 n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , 
 n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , 
 n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , 
 n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , 
 n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , 
 n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , 
 n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , 
 n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , 
 n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , 
 n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , 
 n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , 
 n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , 
 n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , 
 n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , 
 n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , 
 n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , 
 n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , 
 n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , 
 n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , 
 n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , 
 n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , 
 n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , 
 n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , 
 n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , 
 n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , 
 n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , 
 n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , 
 n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , 
 n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , 
 n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , 
 n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , 
 n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , 
 n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , 
 n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , 
 n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , 
 n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , 
 n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , 
 n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , 
 n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , 
 n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
 n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
 n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , 
 n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , 
 n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , 
 n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , 
 n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , 
 n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , 
 n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , 
 n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , 
 n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , 
 n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , 
 n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , 
 n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , 
 n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , 
 n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , 
 n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , 
 n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , 
 n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , 
 n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , 
 n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , 
 n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , 
 n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
 n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , 
 n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , 
 n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , 
 n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , 
 n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , 
 n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , 
 n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , 
 n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , 
 n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
 n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
 n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , 
 n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , 
 n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , 
 n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , 
 n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , 
 n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , 
 n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , 
 n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , 
 n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , 
 n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , 
 n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , 
 n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , 
 n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , 
 n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , 
 n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , 
 n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
 n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , 
 n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , 
 n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , 
 n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , 
 n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , 
 n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , 
 n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , 
 n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , 
 n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , 
 n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , 
 n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , 
 n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , 
 n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , 
 n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , 
 n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , 
 n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , 
 n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , 
 n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , 
 n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , 
 n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , 
 n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , 
 n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , 
 n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , 
 n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , 
 n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , 
 n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , 
 n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , 
 n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , 
 n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
 n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
 n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
 n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
 n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
 n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
 n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
 n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
 n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , 
 n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , 
 n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , 
 n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , 
 n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , 
 n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , 
 n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , 
 n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , 
 n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
 n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , 
 n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , 
 n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
 n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , 
 n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , 
 n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , 
 n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , 
 n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , 
 n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , 
 n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , 
 n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , 
 n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , 
 n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , 
 n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , 
 n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , 
 n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , 
 n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , 
 n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , 
 n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , 
 n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , 
 n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , 
 n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , 
 n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , 
 n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , 
 n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , 
 n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , 
 n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , 
 n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , 
 n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , 
 n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , 
 n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , 
 n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , 
 n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , 
 n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , 
 n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , 
 n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
 n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , 
 n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , 
 n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , 
 n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , 
 n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , 
 n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , 
 n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , 
 n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , 
 n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , 
 n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , 
 n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , 
 n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , 
 n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , 
 n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , 
 n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , 
 n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
 n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , 
 n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , 
 n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , 
 n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , 
 n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , 
 n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , 
 n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , 
 n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , 
 n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , 
 n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , 
 n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , 
 n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , 
 n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , 
 n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , 
 n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
 n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , 
 n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , 
 n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , 
 n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , 
 n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , 
 n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , 
 n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , 
 n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , 
 n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , 
 n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , 
 n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , 
 n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , 
 n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , 
 n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , 
 n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , 
 n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , 
 n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , 
 n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , 
 n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , 
 n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , 
 n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , 
 n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , 
 n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , 
 n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , 
 n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , 
 n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , 
 n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , 
 n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , 
 n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
 n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
 n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , 
 n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , 
 n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , 
 n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , 
 n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , 
 n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , 
 n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , 
 n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , 
 n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , 
 n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , 
 n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , 
 n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , 
 n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , 
 n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , 
 n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , 
 n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , 
 n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , 
 n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , 
 n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , 
 n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , 
 n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , 
 n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , 
 n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , 
 n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , 
 n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , 
 n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , 
 n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , 
 n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , 
 n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , 
 n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , 
 n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , 
 n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , 
 n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , 
 n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , 
 n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , 
 n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , 
 n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , 
 n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , 
 n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , 
 n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , 
 n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , 
 n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , 
 n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , 
 n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , 
 n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , 
 n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , 
 n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , 
 n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , 
 n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , 
 n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , 
 n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , 
 n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , 
 n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , 
 n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , 
 n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , 
 n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , 
 n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , 
 n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , 
 n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , 
 n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , 
 n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , 
 n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , 
 n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , 
 n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , 
 n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , 
 n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
 n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
 n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
 n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , 
 n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
 n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
 n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , 
 n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , 
 n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , 
 n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , 
 n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , 
 n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , 
 n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , 
 n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , 
 n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , 
 n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , 
 n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , 
 n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , 
 n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , 
 n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , 
 n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , 
 n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , 
 n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , 
 n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , 
 n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , 
 n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , 
 n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , 
 n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , 
 n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , 
 n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , 
 n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , 
 n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , 
 n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , 
 n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , 
 n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , 
 n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , C0n , C0 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , n17538 );
buf ( n570 , n17437 );
buf ( n571 , n17320 );
buf ( n572 , n17209 );
buf ( n573 , n17060 );
buf ( n574 , n16904 );
buf ( n575 , n16722 );
buf ( n576 , n16527 );
buf ( n577 , n16318 );
buf ( n578 , n16099 );
buf ( n579 , n15870 );
buf ( n580 , n15630 );
buf ( n581 , n15367 );
buf ( n582 , n15080 );
buf ( n583 , n14772 );
buf ( n584 , n14459 );
buf ( n585 , n14133 );
buf ( n586 , n13787 );
buf ( n587 , n13422 );
buf ( n588 , n13056 );
buf ( n589 , n12664 );
buf ( n590 , n12273 );
buf ( n591 , n11860 );
buf ( n592 , n11450 );
buf ( n593 , n11023 );
buf ( n594 , n10595 );
buf ( n595 , n10154 );
buf ( n596 , n9716 );
buf ( n597 , n9247 );
buf ( n598 , n8803 );
buf ( n599 , n8338 );
buf ( n600 , n7905 );
buf ( n601 , n7472 );
buf ( n602 , n7046 );
buf ( n603 , n6659 );
buf ( n604 , n6287 );
buf ( n605 , n5949 );
buf ( n606 , n5634 );
buf ( n607 , n5354 );
buf ( n608 , n5082 );
buf ( n609 , n4861 );
buf ( n610 , n4661 );
buf ( n611 , n4501 );
buf ( n612 , n17821 );
buf ( n613 , n17813 );
buf ( n614 , n17805 );
buf ( n615 , n17797 );
buf ( n616 , n17789 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , n17781 );
buf ( n634 , n17762 );
buf ( n635 , n17727 );
buf ( n636 , n17682 );
buf ( n637 , n17627 );
buf ( n638 , n17560 );
buf ( n639 , n17461 );
buf ( n640 , n17351 );
buf ( n641 , n17233 );
buf ( n642 , n17089 );
buf ( n643 , n16929 );
buf ( n644 , n16751 );
buf ( n645 , n16558 );
buf ( n646 , n16351 );
buf ( n647 , n16130 );
buf ( n648 , n15899 );
buf ( n649 , n15654 );
buf ( n650 , n15397 );
buf ( n651 , n15107 );
buf ( n652 , n14805 );
buf ( n653 , n14490 );
buf ( n654 , n14162 );
buf ( n655 , n13811 );
buf ( n656 , n13451 );
buf ( n657 , n13080 );
buf ( n658 , n12693 );
buf ( n659 , n12298 );
buf ( n660 , n11889 );
buf ( n661 , n11475 );
buf ( n662 , n11052 );
buf ( n663 , n10619 );
buf ( n664 , n10183 );
buf ( n665 , n9740 );
buf ( n666 , n9276 );
buf ( n667 , n8827 );
buf ( n668 , n8367 );
buf ( n669 , n7934 );
buf ( n670 , n7501 );
buf ( n671 , n7075 );
buf ( n672 , n6688 );
buf ( n673 , n6316 );
buf ( n674 , n5978 );
buf ( n675 , n5655 );
buf ( n676 , n5370 );
buf ( n677 , n5104 );
buf ( n678 , n4877 );
buf ( n679 , n4670 );
buf ( n680 , n4513 );
buf ( n681 , n520 );
buf ( n682 , n681 );
buf ( n683 , n501 );
buf ( n684 , n683 );
buf ( n685 , n502 );
buf ( n686 , n685 );
xor ( n687 , n684 , n686 );
buf ( n688 , n503 );
buf ( n689 , n688 );
xor ( n690 , n686 , n689 );
not ( n691 , n690 );
and ( n692 , n687 , n691 );
and ( n693 , n682 , n692 );
buf ( n694 , n519 );
buf ( n695 , n694 );
and ( n696 , n695 , n690 );
nor ( n697 , n693 , n696 );
and ( n698 , n686 , n689 );
not ( n699 , n698 );
and ( n700 , n684 , n699 );
xnor ( n701 , n697 , n700 );
buf ( n702 , n518 );
buf ( n703 , n702 );
buf ( n704 , n504 );
buf ( n705 , n704 );
xor ( n706 , n689 , n705 );
not ( n707 , n705 );
and ( n708 , n706 , n707 );
and ( n709 , n703 , n708 );
buf ( n710 , n517 );
buf ( n711 , n710 );
and ( n712 , n711 , n705 );
nor ( n713 , n709 , n712 );
xnor ( n714 , n713 , n689 );
and ( n715 , n682 , n690 );
not ( n716 , n715 );
and ( n717 , n716 , n700 );
xnor ( n718 , n714 , n717 );
xnor ( n719 , n701 , n718 );
and ( n720 , n695 , n708 );
and ( n721 , n703 , n705 );
nor ( n722 , n720 , n721 );
xnor ( n723 , n722 , n689 );
and ( n724 , n723 , n715 );
xor ( n725 , n723 , n715 );
and ( n726 , n682 , n708 );
and ( n727 , n695 , n705 );
nor ( n728 , n726 , n727 );
xnor ( n729 , n728 , n689 );
and ( n730 , n682 , n705 );
not ( n731 , n730 );
and ( n732 , n731 , n689 );
and ( n733 , n729 , n732 );
and ( n734 , n725 , n733 );
or ( n735 , n724 , n734 );
xor ( n736 , n719 , n735 );
buf ( n737 , n736 );
not ( n738 , n456 );
and ( n739 , n738 , n488 );
and ( n740 , n472 , n456 );
or ( n741 , n739 , n740 );
buf ( n742 , n741 );
buf ( n743 , n742 );
buf ( n744 , n501 );
buf ( n745 , n744 );
buf ( n746 , n502 );
buf ( n747 , n746 );
xor ( n748 , n745 , n747 );
buf ( n749 , n503 );
buf ( n750 , n749 );
xor ( n751 , n747 , n750 );
not ( n752 , n751 );
and ( n753 , n748 , n752 );
and ( n754 , n743 , n753 );
not ( n755 , n456 );
and ( n756 , n755 , n487 );
and ( n757 , n471 , n456 );
or ( n758 , n756 , n757 );
buf ( n759 , n758 );
buf ( n760 , n759 );
and ( n761 , n760 , n751 );
nor ( n762 , n754 , n761 );
and ( n763 , n747 , n750 );
not ( n764 , n763 );
and ( n765 , n745 , n764 );
xnor ( n766 , n762 , n765 );
not ( n767 , n456 );
and ( n768 , n767 , n486 );
and ( n769 , n470 , n456 );
or ( n770 , n768 , n769 );
buf ( n771 , n770 );
buf ( n772 , n771 );
buf ( n773 , n504 );
buf ( n774 , n773 );
xor ( n775 , n750 , n774 );
not ( n776 , n774 );
and ( n777 , n775 , n776 );
and ( n778 , n772 , n777 );
not ( n779 , n456 );
and ( n780 , n779 , n485 );
and ( n781 , n469 , n456 );
or ( n782 , n780 , n781 );
buf ( n783 , n782 );
buf ( n784 , n783 );
and ( n785 , n784 , n774 );
nor ( n786 , n778 , n785 );
xnor ( n787 , n786 , n750 );
and ( n788 , n743 , n751 );
not ( n789 , n788 );
and ( n790 , n789 , n765 );
xor ( n791 , n787 , n790 );
xor ( n792 , n766 , n791 );
and ( n793 , n760 , n777 );
and ( n794 , n772 , n774 );
nor ( n795 , n793 , n794 );
xnor ( n796 , n795 , n750 );
and ( n797 , n796 , n788 );
xor ( n798 , n796 , n788 );
and ( n799 , n743 , n777 );
and ( n800 , n760 , n774 );
nor ( n801 , n799 , n800 );
xnor ( n802 , n801 , n750 );
and ( n803 , n743 , n774 );
not ( n804 , n803 );
and ( n805 , n804 , n750 );
and ( n806 , n802 , n805 );
and ( n807 , n798 , n806 );
or ( n808 , n797 , n807 );
xor ( n809 , n792 , n808 );
buf ( n810 , n809 );
not ( n811 , n455 );
and ( n812 , n811 , n737 );
and ( n813 , n810 , n455 );
or ( n814 , n812 , n813 );
and ( n815 , n711 , n708 );
buf ( n816 , n516 );
buf ( n817 , n816 );
and ( n818 , n817 , n705 );
nor ( n819 , n815 , n818 );
xnor ( n820 , n819 , n689 );
and ( n821 , n695 , n692 );
and ( n822 , n703 , n690 );
nor ( n823 , n821 , n822 );
xnor ( n824 , n823 , n700 );
xor ( n825 , n820 , n824 );
buf ( n826 , n500 );
buf ( n827 , n826 );
xor ( n828 , n827 , n684 );
and ( n829 , n682 , n828 );
xor ( n830 , n825 , n829 );
or ( n831 , n714 , n717 );
xor ( n832 , n830 , n831 );
or ( n833 , n701 , n718 );
xor ( n834 , n832 , n833 );
not ( n835 , n834 );
and ( n836 , n719 , n735 );
xor ( n837 , n835 , n836 );
buf ( n838 , n837 );
and ( n839 , n784 , n777 );
not ( n840 , n456 );
and ( n841 , n840 , n484 );
and ( n842 , n468 , n456 );
or ( n843 , n841 , n842 );
buf ( n844 , n843 );
buf ( n845 , n844 );
and ( n846 , n845 , n774 );
nor ( n847 , n839 , n846 );
xnor ( n848 , n847 , n750 );
and ( n849 , n760 , n753 );
and ( n850 , n772 , n751 );
nor ( n851 , n849 , n850 );
xnor ( n852 , n851 , n765 );
xor ( n853 , n848 , n852 );
buf ( n854 , n500 );
buf ( n855 , n854 );
xor ( n856 , n855 , n745 );
and ( n857 , n743 , n856 );
xor ( n858 , n853 , n857 );
and ( n859 , n787 , n790 );
xor ( n860 , n858 , n859 );
and ( n861 , n766 , n791 );
and ( n862 , n792 , n808 );
or ( n863 , n861 , n862 );
xor ( n864 , n860 , n863 );
buf ( n865 , n864 );
not ( n866 , n455 );
and ( n867 , n866 , n838 );
and ( n868 , n865 , n455 );
or ( n869 , n867 , n868 );
and ( n870 , n820 , n824 );
and ( n871 , n824 , n829 );
and ( n872 , n820 , n829 );
or ( n873 , n870 , n871 , n872 );
and ( n874 , n817 , n708 );
buf ( n875 , n515 );
buf ( n876 , n875 );
and ( n877 , n876 , n705 );
nor ( n878 , n874 , n877 );
xnor ( n879 , n878 , n689 );
not ( n880 , n829 );
buf ( n881 , n499 );
buf ( n882 , n881 );
and ( n883 , n827 , n684 );
not ( n884 , n883 );
and ( n885 , n882 , n884 );
and ( n886 , n880 , n885 );
xor ( n887 , n879 , n886 );
and ( n888 , n703 , n692 );
and ( n889 , n711 , n690 );
nor ( n890 , n888 , n889 );
xnor ( n891 , n890 , n700 );
xor ( n892 , n887 , n891 );
xor ( n893 , n882 , n827 );
not ( n894 , n828 );
and ( n895 , n893 , n894 );
and ( n896 , n682 , n895 );
and ( n897 , n695 , n828 );
nor ( n898 , n896 , n897 );
xnor ( n899 , n898 , n885 );
xor ( n900 , n892 , n899 );
xor ( n901 , n873 , n900 );
and ( n902 , n830 , n831 );
and ( n903 , n831 , n833 );
and ( n904 , n830 , n833 );
or ( n905 , n902 , n903 , n904 );
xor ( n906 , n901 , n905 );
not ( n907 , n906 );
and ( n908 , n835 , n836 );
or ( n909 , n834 , n908 );
xor ( n910 , n907 , n909 );
buf ( n911 , n910 );
and ( n912 , n848 , n852 );
and ( n913 , n852 , n857 );
and ( n914 , n848 , n857 );
or ( n915 , n912 , n913 , n914 );
and ( n916 , n772 , n753 );
and ( n917 , n784 , n751 );
nor ( n918 , n916 , n917 );
xnor ( n919 , n918 , n765 );
buf ( n920 , n499 );
buf ( n921 , n920 );
xor ( n922 , n921 , n855 );
not ( n923 , n856 );
and ( n924 , n922 , n923 );
and ( n925 , n743 , n924 );
and ( n926 , n760 , n856 );
nor ( n927 , n925 , n926 );
and ( n928 , n855 , n745 );
not ( n929 , n928 );
and ( n930 , n921 , n929 );
xnor ( n931 , n927 , n930 );
xor ( n932 , n919 , n931 );
and ( n933 , n845 , n777 );
not ( n934 , n456 );
and ( n935 , n934 , n483 );
and ( n936 , n467 , n456 );
or ( n937 , n935 , n936 );
buf ( n938 , n937 );
buf ( n939 , n938 );
and ( n940 , n939 , n774 );
nor ( n941 , n933 , n940 );
xnor ( n942 , n941 , n750 );
not ( n943 , n857 );
and ( n944 , n943 , n930 );
xor ( n945 , n942 , n944 );
xor ( n946 , n932 , n945 );
xor ( n947 , n915 , n946 );
and ( n948 , n858 , n859 );
and ( n949 , n860 , n863 );
or ( n950 , n948 , n949 );
xor ( n951 , n947 , n950 );
buf ( n952 , n951 );
not ( n953 , n455 );
and ( n954 , n953 , n911 );
and ( n955 , n952 , n455 );
or ( n956 , n954 , n955 );
and ( n957 , n879 , n886 );
and ( n958 , n695 , n895 );
and ( n959 , n703 , n828 );
nor ( n960 , n958 , n959 );
xnor ( n961 , n960 , n885 );
xor ( n962 , n957 , n961 );
and ( n963 , n876 , n708 );
buf ( n964 , n514 );
buf ( n965 , n964 );
and ( n966 , n965 , n705 );
nor ( n967 , n963 , n966 );
xnor ( n968 , n967 , n689 );
and ( n969 , n711 , n692 );
and ( n970 , n817 , n690 );
nor ( n971 , n969 , n970 );
xnor ( n972 , n971 , n700 );
xor ( n973 , n968 , n972 );
buf ( n974 , n498 );
buf ( n975 , n974 );
xor ( n976 , n975 , n882 );
and ( n977 , n682 , n976 );
xor ( n978 , n973 , n977 );
xor ( n979 , n962 , n978 );
and ( n980 , n887 , n891 );
and ( n981 , n891 , n899 );
and ( n982 , n887 , n899 );
or ( n983 , n980 , n981 , n982 );
xor ( n984 , n979 , n983 );
and ( n985 , n873 , n900 );
and ( n986 , n900 , n905 );
and ( n987 , n873 , n905 );
or ( n988 , n985 , n986 , n987 );
xor ( n989 , n984 , n988 );
not ( n990 , n989 );
and ( n991 , n907 , n909 );
or ( n992 , n906 , n991 );
xor ( n993 , n990 , n992 );
buf ( n994 , n993 );
and ( n995 , n919 , n931 );
and ( n996 , n931 , n945 );
and ( n997 , n919 , n945 );
or ( n998 , n995 , n996 , n997 );
and ( n999 , n784 , n753 );
and ( n1000 , n845 , n751 );
nor ( n1001 , n999 , n1000 );
xnor ( n1002 , n1001 , n765 );
and ( n1003 , n939 , n777 );
not ( n1004 , n456 );
and ( n1005 , n1004 , n482 );
and ( n1006 , n466 , n456 );
or ( n1007 , n1005 , n1006 );
buf ( n1008 , n1007 );
buf ( n1009 , n1008 );
and ( n1010 , n1009 , n774 );
nor ( n1011 , n1003 , n1010 );
xnor ( n1012 , n1011 , n750 );
buf ( n1013 , n498 );
buf ( n1014 , n1013 );
xor ( n1015 , n1014 , n921 );
and ( n1016 , n743 , n1015 );
xor ( n1017 , n1012 , n1016 );
xor ( n1018 , n1002 , n1017 );
and ( n1019 , n942 , n944 );
and ( n1020 , n760 , n924 );
and ( n1021 , n772 , n856 );
nor ( n1022 , n1020 , n1021 );
xnor ( n1023 , n1022 , n930 );
xor ( n1024 , n1019 , n1023 );
xor ( n1025 , n1018 , n1024 );
xor ( n1026 , n998 , n1025 );
and ( n1027 , n915 , n946 );
and ( n1028 , n947 , n950 );
or ( n1029 , n1027 , n1028 );
xor ( n1030 , n1026 , n1029 );
buf ( n1031 , n1030 );
not ( n1032 , n455 );
and ( n1033 , n1032 , n994 );
and ( n1034 , n1031 , n455 );
or ( n1035 , n1033 , n1034 );
and ( n1036 , n965 , n708 );
buf ( n1037 , n513 );
buf ( n1038 , n1037 );
and ( n1039 , n1038 , n705 );
nor ( n1040 , n1036 , n1039 );
xnor ( n1041 , n1040 , n689 );
not ( n1042 , n977 );
buf ( n1043 , n497 );
buf ( n1044 , n1043 );
and ( n1045 , n975 , n882 );
not ( n1046 , n1045 );
and ( n1047 , n1044 , n1046 );
and ( n1048 , n1042 , n1047 );
xor ( n1049 , n1041 , n1048 );
and ( n1050 , n968 , n972 );
and ( n1051 , n972 , n977 );
and ( n1052 , n968 , n977 );
or ( n1053 , n1050 , n1051 , n1052 );
xor ( n1054 , n1049 , n1053 );
and ( n1055 , n817 , n692 );
and ( n1056 , n876 , n690 );
nor ( n1057 , n1055 , n1056 );
xnor ( n1058 , n1057 , n700 );
and ( n1059 , n703 , n895 );
and ( n1060 , n711 , n828 );
nor ( n1061 , n1059 , n1060 );
xnor ( n1062 , n1061 , n885 );
xor ( n1063 , n1058 , n1062 );
xor ( n1064 , n1044 , n975 );
not ( n1065 , n976 );
and ( n1066 , n1064 , n1065 );
and ( n1067 , n682 , n1066 );
and ( n1068 , n695 , n976 );
nor ( n1069 , n1067 , n1068 );
xnor ( n1070 , n1069 , n1047 );
xor ( n1071 , n1063 , n1070 );
xor ( n1072 , n1054 , n1071 );
and ( n1073 , n957 , n961 );
and ( n1074 , n961 , n978 );
and ( n1075 , n957 , n978 );
or ( n1076 , n1073 , n1074 , n1075 );
xor ( n1077 , n1072 , n1076 );
and ( n1078 , n979 , n983 );
and ( n1079 , n983 , n988 );
and ( n1080 , n979 , n988 );
or ( n1081 , n1078 , n1079 , n1080 );
xor ( n1082 , n1077 , n1081 );
not ( n1083 , n1082 );
and ( n1084 , n990 , n992 );
or ( n1085 , n989 , n1084 );
xor ( n1086 , n1083 , n1085 );
buf ( n1087 , n1086 );
and ( n1088 , n1002 , n1017 );
and ( n1089 , n1017 , n1024 );
and ( n1090 , n1002 , n1024 );
or ( n1091 , n1088 , n1089 , n1090 );
and ( n1092 , n1012 , n1016 );
and ( n1093 , n1019 , n1023 );
xor ( n1094 , n1092 , n1093 );
and ( n1095 , n772 , n924 );
and ( n1096 , n784 , n856 );
nor ( n1097 , n1095 , n1096 );
xnor ( n1098 , n1097 , n930 );
and ( n1099 , n845 , n753 );
and ( n1100 , n939 , n751 );
nor ( n1101 , n1099 , n1100 );
xnor ( n1102 , n1101 , n765 );
buf ( n1103 , n497 );
buf ( n1104 , n1103 );
xor ( n1105 , n1104 , n1014 );
not ( n1106 , n1015 );
and ( n1107 , n1105 , n1106 );
and ( n1108 , n743 , n1107 );
and ( n1109 , n760 , n1015 );
nor ( n1110 , n1108 , n1109 );
and ( n1111 , n1014 , n921 );
not ( n1112 , n1111 );
and ( n1113 , n1104 , n1112 );
xnor ( n1114 , n1110 , n1113 );
xor ( n1115 , n1102 , n1114 );
xor ( n1116 , n1098 , n1115 );
and ( n1117 , n1009 , n777 );
not ( n1118 , n456 );
and ( n1119 , n1118 , n481 );
and ( n1120 , n465 , n456 );
or ( n1121 , n1119 , n1120 );
buf ( n1122 , n1121 );
buf ( n1123 , n1122 );
and ( n1124 , n1123 , n774 );
nor ( n1125 , n1117 , n1124 );
xnor ( n1126 , n1125 , n750 );
not ( n1127 , n1016 );
and ( n1128 , n1127 , n1113 );
xor ( n1129 , n1126 , n1128 );
xor ( n1130 , n1116 , n1129 );
xor ( n1131 , n1094 , n1130 );
xor ( n1132 , n1091 , n1131 );
and ( n1133 , n998 , n1025 );
and ( n1134 , n1026 , n1029 );
or ( n1135 , n1133 , n1134 );
xor ( n1136 , n1132 , n1135 );
buf ( n1137 , n1136 );
not ( n1138 , n455 );
and ( n1139 , n1138 , n1087 );
and ( n1140 , n1137 , n455 );
or ( n1141 , n1139 , n1140 );
and ( n1142 , n1049 , n1053 );
and ( n1143 , n1053 , n1071 );
and ( n1144 , n1049 , n1071 );
or ( n1145 , n1142 , n1143 , n1144 );
and ( n1146 , n1041 , n1048 );
and ( n1147 , n876 , n692 );
and ( n1148 , n965 , n690 );
nor ( n1149 , n1147 , n1148 );
xnor ( n1150 , n1149 , n700 );
xor ( n1151 , n1146 , n1150 );
and ( n1152 , n711 , n895 );
and ( n1153 , n817 , n828 );
nor ( n1154 , n1152 , n1153 );
xnor ( n1155 , n1154 , n885 );
xor ( n1156 , n1151 , n1155 );
not ( n1157 , n1156 );
and ( n1158 , n1058 , n1062 );
and ( n1159 , n1062 , n1070 );
and ( n1160 , n1058 , n1070 );
or ( n1161 , n1158 , n1159 , n1160 );
and ( n1162 , n1038 , n708 );
buf ( n1163 , n512 );
buf ( n1164 , n1163 );
and ( n1165 , n1164 , n705 );
nor ( n1166 , n1162 , n1165 );
xnor ( n1167 , n1166 , n689 );
and ( n1168 , n695 , n1066 );
and ( n1169 , n703 , n976 );
nor ( n1170 , n1168 , n1169 );
xnor ( n1171 , n1170 , n1047 );
xor ( n1172 , n1167 , n1171 );
buf ( n1173 , n496 );
buf ( n1174 , n1173 );
xor ( n1175 , n1174 , n1044 );
and ( n1176 , n682 , n1175 );
xor ( n1177 , n1172 , n1176 );
xor ( n1178 , n1161 , n1177 );
xor ( n1179 , n1157 , n1178 );
xor ( n1180 , n1145 , n1179 );
and ( n1181 , n1072 , n1076 );
and ( n1182 , n1076 , n1081 );
and ( n1183 , n1072 , n1081 );
or ( n1184 , n1181 , n1182 , n1183 );
xor ( n1185 , n1180 , n1184 );
and ( n1186 , n1083 , n1085 );
or ( n1187 , n1082 , n1186 );
xor ( n1188 , n1185 , n1187 );
buf ( n1189 , n1188 );
and ( n1190 , n760 , n1107 );
and ( n1191 , n772 , n1015 );
nor ( n1192 , n1190 , n1191 );
xnor ( n1193 , n1192 , n1113 );
buf ( n1194 , n496 );
buf ( n1195 , n1194 );
xor ( n1196 , n1195 , n1104 );
and ( n1197 , n743 , n1196 );
xor ( n1198 , n1193 , n1197 );
and ( n1199 , n1102 , n1114 );
xor ( n1200 , n1198 , n1199 );
and ( n1201 , n1092 , n1093 );
and ( n1202 , n1093 , n1130 );
and ( n1203 , n1092 , n1130 );
or ( n1204 , n1201 , n1202 , n1203 );
xor ( n1205 , n1200 , n1204 );
and ( n1206 , n1126 , n1128 );
and ( n1207 , n1123 , n777 );
not ( n1208 , n456 );
and ( n1209 , n1208 , n480 );
and ( n1210 , n464 , n456 );
or ( n1211 , n1209 , n1210 );
buf ( n1212 , n1211 );
buf ( n1213 , n1212 );
and ( n1214 , n1213 , n774 );
nor ( n1215 , n1207 , n1214 );
xnor ( n1216 , n1215 , n750 );
and ( n1217 , n939 , n753 );
and ( n1218 , n1009 , n751 );
nor ( n1219 , n1217 , n1218 );
xnor ( n1220 , n1219 , n765 );
xor ( n1221 , n1216 , n1220 );
and ( n1222 , n784 , n924 );
and ( n1223 , n845 , n856 );
nor ( n1224 , n1222 , n1223 );
xnor ( n1225 , n1224 , n930 );
xor ( n1226 , n1221 , n1225 );
xor ( n1227 , n1206 , n1226 );
and ( n1228 , n1098 , n1115 );
and ( n1229 , n1115 , n1129 );
and ( n1230 , n1098 , n1129 );
or ( n1231 , n1228 , n1229 , n1230 );
xor ( n1232 , n1227 , n1231 );
xor ( n1233 , n1205 , n1232 );
and ( n1234 , n1091 , n1131 );
and ( n1235 , n1132 , n1135 );
or ( n1236 , n1234 , n1235 );
xor ( n1237 , n1233 , n1236 );
buf ( n1238 , n1237 );
not ( n1239 , n455 );
and ( n1240 , n1239 , n1189 );
and ( n1241 , n1238 , n455 );
or ( n1242 , n1240 , n1241 );
buf ( n1243 , n1156 );
and ( n1244 , n1161 , n1177 );
and ( n1245 , n1146 , n1150 );
and ( n1246 , n1150 , n1155 );
and ( n1247 , n1146 , n1155 );
or ( n1248 , n1245 , n1246 , n1247 );
and ( n1249 , n1164 , n708 );
buf ( n1250 , n511 );
buf ( n1251 , n1250 );
and ( n1252 , n1251 , n705 );
nor ( n1253 , n1249 , n1252 );
xnor ( n1254 , n1253 , n689 );
and ( n1255 , n703 , n1066 );
and ( n1256 , n711 , n976 );
nor ( n1257 , n1255 , n1256 );
xnor ( n1258 , n1257 , n1047 );
xor ( n1259 , n1254 , n1258 );
buf ( n1260 , n495 );
buf ( n1261 , n1260 );
xor ( n1262 , n1261 , n1174 );
not ( n1263 , n1175 );
and ( n1264 , n1262 , n1263 );
and ( n1265 , n682 , n1264 );
and ( n1266 , n695 , n1175 );
nor ( n1267 , n1265 , n1266 );
and ( n1268 , n1174 , n1044 );
not ( n1269 , n1268 );
and ( n1270 , n1261 , n1269 );
xnor ( n1271 , n1267 , n1270 );
xor ( n1272 , n1259 , n1271 );
xor ( n1273 , n1248 , n1272 );
and ( n1274 , n965 , n692 );
and ( n1275 , n1038 , n690 );
nor ( n1276 , n1274 , n1275 );
xnor ( n1277 , n1276 , n700 );
not ( n1278 , n1176 );
and ( n1279 , n1278 , n1270 );
xor ( n1280 , n1277 , n1279 );
and ( n1281 , n1167 , n1171 );
and ( n1282 , n1171 , n1176 );
and ( n1283 , n1167 , n1176 );
or ( n1284 , n1281 , n1282 , n1283 );
xor ( n1285 , n1280 , n1284 );
and ( n1286 , n817 , n895 );
and ( n1287 , n876 , n828 );
nor ( n1288 , n1286 , n1287 );
xnor ( n1289 , n1288 , n885 );
xor ( n1290 , n1285 , n1289 );
xor ( n1291 , n1273 , n1290 );
xor ( n1292 , n1244 , n1291 );
and ( n1293 , n1157 , n1178 );
xor ( n1294 , n1292 , n1293 );
xor ( n1295 , n1243 , n1294 );
and ( n1296 , n1145 , n1179 );
and ( n1297 , n1179 , n1184 );
and ( n1298 , n1145 , n1184 );
or ( n1299 , n1296 , n1297 , n1298 );
xor ( n1300 , n1295 , n1299 );
not ( n1301 , n1300 );
and ( n1302 , n1185 , n1187 );
xor ( n1303 , n1301 , n1302 );
buf ( n1304 , n1303 );
and ( n1305 , n1200 , n1204 );
and ( n1306 , n1204 , n1232 );
and ( n1307 , n1200 , n1232 );
or ( n1308 , n1305 , n1306 , n1307 );
and ( n1309 , n1193 , n1197 );
and ( n1310 , n1197 , n1199 );
and ( n1311 , n1193 , n1199 );
or ( n1312 , n1309 , n1310 , n1311 );
and ( n1313 , n1216 , n1220 );
and ( n1314 , n1220 , n1225 );
and ( n1315 , n1216 , n1225 );
or ( n1316 , n1313 , n1314 , n1315 );
and ( n1317 , n1213 , n777 );
not ( n1318 , n456 );
and ( n1319 , n1318 , n479 );
and ( n1320 , n463 , n456 );
or ( n1321 , n1319 , n1320 );
buf ( n1322 , n1321 );
buf ( n1323 , n1322 );
and ( n1324 , n1323 , n774 );
nor ( n1325 , n1317 , n1324 );
xnor ( n1326 , n1325 , n750 );
and ( n1327 , n1009 , n753 );
and ( n1328 , n1123 , n751 );
nor ( n1329 , n1327 , n1328 );
xnor ( n1330 , n1329 , n765 );
xor ( n1331 , n1326 , n1330 );
and ( n1332 , n845 , n924 );
and ( n1333 , n939 , n856 );
nor ( n1334 , n1332 , n1333 );
xnor ( n1335 , n1334 , n930 );
xor ( n1336 , n1331 , n1335 );
xor ( n1337 , n1316 , n1336 );
and ( n1338 , n772 , n1107 );
and ( n1339 , n784 , n1015 );
nor ( n1340 , n1338 , n1339 );
xnor ( n1341 , n1340 , n1113 );
buf ( n1342 , n495 );
buf ( n1343 , n1342 );
xor ( n1344 , n1343 , n1195 );
not ( n1345 , n1196 );
and ( n1346 , n1344 , n1345 );
and ( n1347 , n743 , n1346 );
and ( n1348 , n760 , n1196 );
nor ( n1349 , n1347 , n1348 );
and ( n1350 , n1195 , n1104 );
not ( n1351 , n1350 );
and ( n1352 , n1343 , n1351 );
xnor ( n1353 , n1349 , n1352 );
xor ( n1354 , n1341 , n1353 );
not ( n1355 , n1197 );
and ( n1356 , n1355 , n1352 );
xor ( n1357 , n1354 , n1356 );
xor ( n1358 , n1337 , n1357 );
xor ( n1359 , n1312 , n1358 );
and ( n1360 , n1206 , n1226 );
and ( n1361 , n1226 , n1231 );
and ( n1362 , n1206 , n1231 );
or ( n1363 , n1360 , n1361 , n1362 );
xor ( n1364 , n1359 , n1363 );
xor ( n1365 , n1308 , n1364 );
and ( n1366 , n1233 , n1236 );
xor ( n1367 , n1365 , n1366 );
buf ( n1368 , n1367 );
not ( n1369 , n455 );
and ( n1370 , n1369 , n1304 );
and ( n1371 , n1368 , n455 );
or ( n1372 , n1370 , n1371 );
and ( n1373 , n1280 , n1284 );
and ( n1374 , n1284 , n1289 );
and ( n1375 , n1280 , n1289 );
or ( n1376 , n1373 , n1374 , n1375 );
and ( n1377 , n1251 , n708 );
buf ( n1378 , n510 );
buf ( n1379 , n1378 );
and ( n1380 , n1379 , n705 );
nor ( n1381 , n1377 , n1380 );
xnor ( n1382 , n1381 , n689 );
and ( n1383 , n876 , n895 );
and ( n1384 , n965 , n828 );
nor ( n1385 , n1383 , n1384 );
xnor ( n1386 , n1385 , n885 );
xor ( n1387 , n1382 , n1386 );
and ( n1388 , n695 , n1264 );
and ( n1389 , n703 , n1175 );
nor ( n1390 , n1388 , n1389 );
xnor ( n1391 , n1390 , n1270 );
xor ( n1392 , n1387 , n1391 );
xor ( n1393 , n1376 , n1392 );
and ( n1394 , n1254 , n1258 );
and ( n1395 , n1258 , n1271 );
and ( n1396 , n1254 , n1271 );
or ( n1397 , n1394 , n1395 , n1396 );
and ( n1398 , n1277 , n1279 );
xor ( n1399 , n1397 , n1398 );
and ( n1400 , n1038 , n692 );
and ( n1401 , n1164 , n690 );
nor ( n1402 , n1400 , n1401 );
xnor ( n1403 , n1402 , n700 );
and ( n1404 , n711 , n1066 );
and ( n1405 , n817 , n976 );
nor ( n1406 , n1404 , n1405 );
xnor ( n1407 , n1406 , n1047 );
xor ( n1408 , n1403 , n1407 );
buf ( n1409 , n494 );
buf ( n1410 , n1409 );
xor ( n1411 , n1410 , n1261 );
and ( n1412 , n682 , n1411 );
xor ( n1413 , n1408 , n1412 );
xor ( n1414 , n1399 , n1413 );
xor ( n1415 , n1393 , n1414 );
and ( n1416 , n1248 , n1272 );
and ( n1417 , n1272 , n1290 );
and ( n1418 , n1248 , n1290 );
or ( n1419 , n1416 , n1417 , n1418 );
xor ( n1420 , n1415 , n1419 );
and ( n1421 , n1244 , n1291 );
and ( n1422 , n1291 , n1293 );
and ( n1423 , n1244 , n1293 );
or ( n1424 , n1421 , n1422 , n1423 );
xor ( n1425 , n1420 , n1424 );
and ( n1426 , n1243 , n1294 );
and ( n1427 , n1294 , n1299 );
and ( n1428 , n1243 , n1299 );
or ( n1429 , n1426 , n1427 , n1428 );
xnor ( n1430 , n1425 , n1429 );
and ( n1431 , n1301 , n1302 );
or ( n1432 , n1300 , n1431 );
xor ( n1433 , n1430 , n1432 );
buf ( n1434 , n1433 );
and ( n1435 , n784 , n1107 );
and ( n1436 , n845 , n1015 );
nor ( n1437 , n1435 , n1436 );
xnor ( n1438 , n1437 , n1113 );
and ( n1439 , n760 , n1346 );
and ( n1440 , n772 , n1196 );
nor ( n1441 , n1439 , n1440 );
xnor ( n1442 , n1441 , n1352 );
xor ( n1443 , n1438 , n1442 );
buf ( n1444 , n494 );
buf ( n1445 , n1444 );
xor ( n1446 , n1445 , n1343 );
and ( n1447 , n743 , n1446 );
xor ( n1448 , n1443 , n1447 );
and ( n1449 , n1316 , n1336 );
and ( n1450 , n1336 , n1357 );
and ( n1451 , n1316 , n1357 );
or ( n1452 , n1449 , n1450 , n1451 );
xor ( n1453 , n1448 , n1452 );
and ( n1454 , n1326 , n1330 );
and ( n1455 , n1330 , n1335 );
and ( n1456 , n1326 , n1335 );
or ( n1457 , n1454 , n1455 , n1456 );
and ( n1458 , n1341 , n1353 );
and ( n1459 , n1353 , n1356 );
and ( n1460 , n1341 , n1356 );
or ( n1461 , n1458 , n1459 , n1460 );
xor ( n1462 , n1457 , n1461 );
and ( n1463 , n1323 , n777 );
not ( n1464 , n456 );
and ( n1465 , n1464 , n478 );
and ( n1466 , n462 , n456 );
or ( n1467 , n1465 , n1466 );
buf ( n1468 , n1467 );
buf ( n1469 , n1468 );
and ( n1470 , n1469 , n774 );
nor ( n1471 , n1463 , n1470 );
xnor ( n1472 , n1471 , n750 );
and ( n1473 , n1123 , n753 );
and ( n1474 , n1213 , n751 );
nor ( n1475 , n1473 , n1474 );
xnor ( n1476 , n1475 , n765 );
xor ( n1477 , n1472 , n1476 );
and ( n1478 , n939 , n924 );
and ( n1479 , n1009 , n856 );
nor ( n1480 , n1478 , n1479 );
xnor ( n1481 , n1480 , n930 );
xor ( n1482 , n1477 , n1481 );
xor ( n1483 , n1462 , n1482 );
xor ( n1484 , n1453 , n1483 );
and ( n1485 , n1312 , n1358 );
and ( n1486 , n1358 , n1363 );
and ( n1487 , n1312 , n1363 );
or ( n1488 , n1485 , n1486 , n1487 );
xor ( n1489 , n1484 , n1488 );
and ( n1490 , n1308 , n1364 );
and ( n1491 , n1365 , n1366 );
or ( n1492 , n1490 , n1491 );
xor ( n1493 , n1489 , n1492 );
buf ( n1494 , n1493 );
not ( n1495 , n455 );
and ( n1496 , n1495 , n1434 );
and ( n1497 , n1494 , n455 );
or ( n1498 , n1496 , n1497 );
and ( n1499 , n1397 , n1398 );
and ( n1500 , n1398 , n1413 );
and ( n1501 , n1397 , n1413 );
or ( n1502 , n1499 , n1500 , n1501 );
and ( n1503 , n1164 , n692 );
and ( n1504 , n1251 , n690 );
nor ( n1505 , n1503 , n1504 );
xnor ( n1506 , n1505 , n700 );
not ( n1507 , n1412 );
buf ( n1508 , n493 );
buf ( n1509 , n1508 );
and ( n1510 , n1410 , n1261 );
not ( n1511 , n1510 );
and ( n1512 , n1509 , n1511 );
and ( n1513 , n1507 , n1512 );
xor ( n1514 , n1506 , n1513 );
and ( n1515 , n965 , n895 );
and ( n1516 , n1038 , n828 );
nor ( n1517 , n1515 , n1516 );
xnor ( n1518 , n1517 , n885 );
xor ( n1519 , n1514 , n1518 );
xor ( n1520 , n1509 , n1410 );
not ( n1521 , n1411 );
and ( n1522 , n1520 , n1521 );
and ( n1523 , n682 , n1522 );
and ( n1524 , n695 , n1411 );
nor ( n1525 , n1523 , n1524 );
xnor ( n1526 , n1525 , n1512 );
xor ( n1527 , n1519 , n1526 );
xor ( n1528 , n1502 , n1527 );
and ( n1529 , n1403 , n1407 );
and ( n1530 , n1407 , n1412 );
and ( n1531 , n1403 , n1412 );
or ( n1532 , n1529 , n1530 , n1531 );
and ( n1533 , n1382 , n1386 );
and ( n1534 , n1386 , n1391 );
and ( n1535 , n1382 , n1391 );
or ( n1536 , n1533 , n1534 , n1535 );
xor ( n1537 , n1532 , n1536 );
and ( n1538 , n1379 , n708 );
buf ( n1539 , n509 );
buf ( n1540 , n1539 );
and ( n1541 , n1540 , n705 );
nor ( n1542 , n1538 , n1541 );
xnor ( n1543 , n1542 , n689 );
and ( n1544 , n817 , n1066 );
and ( n1545 , n876 , n976 );
nor ( n1546 , n1544 , n1545 );
xnor ( n1547 , n1546 , n1047 );
xor ( n1548 , n1543 , n1547 );
and ( n1549 , n703 , n1264 );
and ( n1550 , n711 , n1175 );
nor ( n1551 , n1549 , n1550 );
xnor ( n1552 , n1551 , n1270 );
xor ( n1553 , n1548 , n1552 );
xor ( n1554 , n1537 , n1553 );
xor ( n1555 , n1528 , n1554 );
and ( n1556 , n1376 , n1392 );
and ( n1557 , n1392 , n1414 );
and ( n1558 , n1376 , n1414 );
or ( n1559 , n1556 , n1557 , n1558 );
xor ( n1560 , n1555 , n1559 );
and ( n1561 , n1415 , n1419 );
and ( n1562 , n1419 , n1424 );
and ( n1563 , n1415 , n1424 );
or ( n1564 , n1561 , n1562 , n1563 );
xor ( n1565 , n1560 , n1564 );
or ( n1566 , n1425 , n1429 );
xnor ( n1567 , n1565 , n1566 );
and ( n1568 , n1430 , n1432 );
xor ( n1569 , n1567 , n1568 );
buf ( n1570 , n1569 );
and ( n1571 , n845 , n1107 );
and ( n1572 , n939 , n1015 );
nor ( n1573 , n1571 , n1572 );
xnor ( n1574 , n1573 , n1113 );
and ( n1575 , n772 , n1346 );
and ( n1576 , n784 , n1196 );
nor ( n1577 , n1575 , n1576 );
xnor ( n1578 , n1577 , n1352 );
xor ( n1579 , n1574 , n1578 );
and ( n1580 , n1009 , n924 );
and ( n1581 , n1123 , n856 );
nor ( n1582 , n1580 , n1581 );
xnor ( n1583 , n1582 , n930 );
buf ( n1584 , n493 );
buf ( n1585 , n1584 );
xor ( n1586 , n1585 , n1445 );
not ( n1587 , n1446 );
and ( n1588 , n1586 , n1587 );
and ( n1589 , n743 , n1588 );
and ( n1590 , n760 , n1446 );
nor ( n1591 , n1589 , n1590 );
and ( n1592 , n1445 , n1343 );
not ( n1593 , n1592 );
and ( n1594 , n1585 , n1593 );
xnor ( n1595 , n1591 , n1594 );
xor ( n1596 , n1583 , n1595 );
xor ( n1597 , n1579 , n1596 );
and ( n1598 , n1472 , n1476 );
and ( n1599 , n1476 , n1481 );
and ( n1600 , n1472 , n1481 );
or ( n1601 , n1598 , n1599 , n1600 );
xor ( n1602 , n1597 , n1601 );
and ( n1603 , n1448 , n1452 );
and ( n1604 , n1452 , n1483 );
and ( n1605 , n1448 , n1483 );
or ( n1606 , n1603 , n1604 , n1605 );
xor ( n1607 , n1602 , n1606 );
and ( n1608 , n1438 , n1442 );
and ( n1609 , n1442 , n1447 );
and ( n1610 , n1438 , n1447 );
or ( n1611 , n1608 , n1609 , n1610 );
and ( n1612 , n1469 , n777 );
not ( n1613 , n456 );
and ( n1614 , n1613 , n477 );
and ( n1615 , n461 , n456 );
or ( n1616 , n1614 , n1615 );
buf ( n1617 , n1616 );
buf ( n1618 , n1617 );
and ( n1619 , n1618 , n774 );
nor ( n1620 , n1612 , n1619 );
xnor ( n1621 , n1620 , n750 );
and ( n1622 , n1213 , n753 );
and ( n1623 , n1323 , n751 );
nor ( n1624 , n1622 , n1623 );
xnor ( n1625 , n1624 , n765 );
xor ( n1626 , n1621 , n1625 );
not ( n1627 , n1447 );
and ( n1628 , n1627 , n1594 );
xor ( n1629 , n1626 , n1628 );
xor ( n1630 , n1611 , n1629 );
and ( n1631 , n1457 , n1461 );
and ( n1632 , n1461 , n1482 );
and ( n1633 , n1457 , n1482 );
or ( n1634 , n1631 , n1632 , n1633 );
xor ( n1635 , n1630 , n1634 );
xor ( n1636 , n1607 , n1635 );
and ( n1637 , n1484 , n1488 );
and ( n1638 , n1489 , n1492 );
or ( n1639 , n1637 , n1638 );
xor ( n1640 , n1636 , n1639 );
buf ( n1641 , n1640 );
not ( n1642 , n455 );
and ( n1643 , n1642 , n1570 );
and ( n1644 , n1641 , n455 );
or ( n1645 , n1643 , n1644 );
and ( n1646 , n1502 , n1527 );
and ( n1647 , n1527 , n1554 );
and ( n1648 , n1502 , n1554 );
or ( n1649 , n1646 , n1647 , n1648 );
and ( n1650 , n1532 , n1536 );
and ( n1651 , n1536 , n1553 );
and ( n1652 , n1532 , n1553 );
or ( n1653 , n1650 , n1651 , n1652 );
and ( n1654 , n1543 , n1547 );
and ( n1655 , n1547 , n1552 );
and ( n1656 , n1543 , n1552 );
or ( n1657 , n1654 , n1655 , n1656 );
and ( n1658 , n1506 , n1513 );
xor ( n1659 , n1657 , n1658 );
and ( n1660 , n1038 , n895 );
and ( n1661 , n1164 , n828 );
nor ( n1662 , n1660 , n1661 );
xnor ( n1663 , n1662 , n885 );
xor ( n1664 , n1659 , n1663 );
xor ( n1665 , n1653 , n1664 );
and ( n1666 , n1514 , n1518 );
and ( n1667 , n1518 , n1526 );
and ( n1668 , n1514 , n1526 );
or ( n1669 , n1666 , n1667 , n1668 );
and ( n1670 , n1540 , n708 );
buf ( n1671 , n508 );
buf ( n1672 , n1671 );
and ( n1673 , n1672 , n705 );
nor ( n1674 , n1670 , n1673 );
xnor ( n1675 , n1674 , n689 );
and ( n1676 , n711 , n1264 );
and ( n1677 , n817 , n1175 );
nor ( n1678 , n1676 , n1677 );
xnor ( n1679 , n1678 , n1270 );
xor ( n1680 , n1675 , n1679 );
and ( n1681 , n695 , n1522 );
and ( n1682 , n703 , n1411 );
nor ( n1683 , n1681 , n1682 );
xnor ( n1684 , n1683 , n1512 );
xor ( n1685 , n1680 , n1684 );
xor ( n1686 , n1669 , n1685 );
and ( n1687 , n1251 , n692 );
and ( n1688 , n1379 , n690 );
nor ( n1689 , n1687 , n1688 );
xnor ( n1690 , n1689 , n700 );
and ( n1691 , n876 , n1066 );
and ( n1692 , n965 , n976 );
nor ( n1693 , n1691 , n1692 );
xnor ( n1694 , n1693 , n1047 );
xor ( n1695 , n1690 , n1694 );
buf ( n1696 , n492 );
buf ( n1697 , n1696 );
xor ( n1698 , n1697 , n1509 );
and ( n1699 , n682 , n1698 );
xor ( n1700 , n1695 , n1699 );
xor ( n1701 , n1686 , n1700 );
xor ( n1702 , n1665 , n1701 );
xor ( n1703 , n1649 , n1702 );
and ( n1704 , n1555 , n1559 );
and ( n1705 , n1559 , n1564 );
and ( n1706 , n1555 , n1564 );
or ( n1707 , n1704 , n1705 , n1706 );
xor ( n1708 , n1703 , n1707 );
or ( n1709 , n1565 , n1566 );
xnor ( n1710 , n1708 , n1709 );
and ( n1711 , n1567 , n1568 );
xor ( n1712 , n1710 , n1711 );
buf ( n1713 , n1712 );
and ( n1714 , n1611 , n1629 );
and ( n1715 , n1629 , n1634 );
and ( n1716 , n1611 , n1634 );
or ( n1717 , n1714 , n1715 , n1716 );
and ( n1718 , n1579 , n1596 );
and ( n1719 , n1596 , n1601 );
and ( n1720 , n1579 , n1601 );
or ( n1721 , n1718 , n1719 , n1720 );
buf ( n1722 , n492 );
buf ( n1723 , n1722 );
xor ( n1724 , n1723 , n1585 );
and ( n1725 , n743 , n1724 );
and ( n1726 , n1618 , n777 );
not ( n1727 , n456 );
and ( n1728 , n1727 , n476 );
and ( n1729 , n460 , n456 );
or ( n1730 , n1728 , n1729 );
buf ( n1731 , n1730 );
buf ( n1732 , n1731 );
and ( n1733 , n1732 , n774 );
nor ( n1734 , n1726 , n1733 );
xnor ( n1735 , n1734 , n750 );
and ( n1736 , n784 , n1346 );
and ( n1737 , n845 , n1196 );
nor ( n1738 , n1736 , n1737 );
xnor ( n1739 , n1738 , n1352 );
xor ( n1740 , n1735 , n1739 );
and ( n1741 , n760 , n1588 );
and ( n1742 , n772 , n1446 );
nor ( n1743 , n1741 , n1742 );
xnor ( n1744 , n1743 , n1594 );
xor ( n1745 , n1740 , n1744 );
xor ( n1746 , n1725 , n1745 );
and ( n1747 , n1574 , n1578 );
xor ( n1748 , n1746 , n1747 );
xor ( n1749 , n1721 , n1748 );
and ( n1750 , n1583 , n1595 );
and ( n1751 , n1621 , n1625 );
and ( n1752 , n1625 , n1628 );
and ( n1753 , n1621 , n1628 );
or ( n1754 , n1751 , n1752 , n1753 );
xor ( n1755 , n1750 , n1754 );
and ( n1756 , n1323 , n753 );
and ( n1757 , n1469 , n751 );
nor ( n1758 , n1756 , n1757 );
xnor ( n1759 , n1758 , n765 );
and ( n1760 , n1123 , n924 );
and ( n1761 , n1213 , n856 );
nor ( n1762 , n1760 , n1761 );
xnor ( n1763 , n1762 , n930 );
xor ( n1764 , n1759 , n1763 );
and ( n1765 , n939 , n1107 );
and ( n1766 , n1009 , n1015 );
nor ( n1767 , n1765 , n1766 );
xnor ( n1768 , n1767 , n1113 );
xor ( n1769 , n1764 , n1768 );
xor ( n1770 , n1755 , n1769 );
xor ( n1771 , n1749 , n1770 );
xor ( n1772 , n1717 , n1771 );
and ( n1773 , n1602 , n1606 );
and ( n1774 , n1606 , n1635 );
and ( n1775 , n1602 , n1635 );
or ( n1776 , n1773 , n1774 , n1775 );
xor ( n1777 , n1772 , n1776 );
and ( n1778 , n1636 , n1639 );
xor ( n1779 , n1777 , n1778 );
buf ( n1780 , n1779 );
not ( n1781 , n455 );
and ( n1782 , n1781 , n1713 );
and ( n1783 , n1780 , n455 );
or ( n1784 , n1782 , n1783 );
and ( n1785 , n1669 , n1685 );
and ( n1786 , n1685 , n1700 );
and ( n1787 , n1669 , n1700 );
or ( n1788 , n1785 , n1786 , n1787 );
and ( n1789 , n1672 , n708 );
buf ( n1790 , n507 );
buf ( n1791 , n1790 );
and ( n1792 , n1791 , n705 );
nor ( n1793 , n1789 , n1792 );
xnor ( n1794 , n1793 , n689 );
not ( n1795 , n1699 );
buf ( n1796 , n491 );
buf ( n1797 , n1796 );
and ( n1798 , n1697 , n1509 );
not ( n1799 , n1798 );
and ( n1800 , n1797 , n1799 );
and ( n1801 , n1795 , n1800 );
xor ( n1802 , n1794 , n1801 );
and ( n1803 , n1675 , n1679 );
and ( n1804 , n1679 , n1684 );
and ( n1805 , n1675 , n1684 );
or ( n1806 , n1803 , n1804 , n1805 );
xor ( n1807 , n1802 , n1806 );
and ( n1808 , n1690 , n1694 );
and ( n1809 , n1694 , n1699 );
and ( n1810 , n1690 , n1699 );
or ( n1811 , n1808 , n1809 , n1810 );
xor ( n1812 , n1807 , n1811 );
xor ( n1813 , n1788 , n1812 );
and ( n1814 , n1657 , n1658 );
and ( n1815 , n1658 , n1663 );
and ( n1816 , n1657 , n1663 );
or ( n1817 , n1814 , n1815 , n1816 );
and ( n1818 , n1164 , n895 );
and ( n1819 , n1251 , n828 );
nor ( n1820 , n1818 , n1819 );
xnor ( n1821 , n1820 , n885 );
and ( n1822 , n703 , n1522 );
and ( n1823 , n711 , n1411 );
nor ( n1824 , n1822 , n1823 );
xnor ( n1825 , n1824 , n1512 );
xor ( n1826 , n1821 , n1825 );
xor ( n1827 , n1797 , n1697 );
not ( n1828 , n1698 );
and ( n1829 , n1827 , n1828 );
and ( n1830 , n682 , n1829 );
and ( n1831 , n695 , n1698 );
nor ( n1832 , n1830 , n1831 );
xnor ( n1833 , n1832 , n1800 );
xor ( n1834 , n1826 , n1833 );
xor ( n1835 , n1817 , n1834 );
and ( n1836 , n1379 , n692 );
and ( n1837 , n1540 , n690 );
nor ( n1838 , n1836 , n1837 );
xnor ( n1839 , n1838 , n700 );
and ( n1840 , n965 , n1066 );
and ( n1841 , n1038 , n976 );
nor ( n1842 , n1840 , n1841 );
xnor ( n1843 , n1842 , n1047 );
xor ( n1844 , n1839 , n1843 );
and ( n1845 , n817 , n1264 );
and ( n1846 , n876 , n1175 );
nor ( n1847 , n1845 , n1846 );
xnor ( n1848 , n1847 , n1270 );
xor ( n1849 , n1844 , n1848 );
xor ( n1850 , n1835 , n1849 );
xor ( n1851 , n1813 , n1850 );
and ( n1852 , n1653 , n1664 );
and ( n1853 , n1664 , n1701 );
and ( n1854 , n1653 , n1701 );
or ( n1855 , n1852 , n1853 , n1854 );
xor ( n1856 , n1851 , n1855 );
and ( n1857 , n1649 , n1702 );
and ( n1858 , n1702 , n1707 );
and ( n1859 , n1649 , n1707 );
or ( n1860 , n1857 , n1858 , n1859 );
xor ( n1861 , n1856 , n1860 );
or ( n1862 , n1708 , n1709 );
xnor ( n1863 , n1861 , n1862 );
and ( n1864 , n1710 , n1711 );
xor ( n1865 , n1863 , n1864 );
buf ( n1866 , n1865 );
and ( n1867 , n1469 , n753 );
and ( n1868 , n1618 , n751 );
nor ( n1869 , n1867 , n1868 );
xnor ( n1870 , n1869 , n765 );
and ( n1871 , n1213 , n924 );
and ( n1872 , n1323 , n856 );
nor ( n1873 , n1871 , n1872 );
xnor ( n1874 , n1873 , n930 );
xor ( n1875 , n1870 , n1874 );
and ( n1876 , n1009 , n1107 );
and ( n1877 , n1123 , n1015 );
nor ( n1878 , n1876 , n1877 );
xnor ( n1879 , n1878 , n1113 );
xor ( n1880 , n1875 , n1879 );
and ( n1881 , n845 , n1346 );
and ( n1882 , n939 , n1196 );
nor ( n1883 , n1881 , n1882 );
xnor ( n1884 , n1883 , n1352 );
and ( n1885 , n772 , n1588 );
and ( n1886 , n784 , n1446 );
nor ( n1887 , n1885 , n1886 );
xnor ( n1888 , n1887 , n1594 );
xor ( n1889 , n1884 , n1888 );
buf ( n1890 , n491 );
buf ( n1891 , n1890 );
xor ( n1892 , n1891 , n1723 );
not ( n1893 , n1724 );
and ( n1894 , n1892 , n1893 );
and ( n1895 , n743 , n1894 );
and ( n1896 , n760 , n1724 );
nor ( n1897 , n1895 , n1896 );
and ( n1898 , n1723 , n1585 );
not ( n1899 , n1898 );
and ( n1900 , n1891 , n1899 );
xnor ( n1901 , n1897 , n1900 );
xor ( n1902 , n1889 , n1901 );
xor ( n1903 , n1880 , n1902 );
and ( n1904 , n1725 , n1745 );
and ( n1905 , n1745 , n1747 );
and ( n1906 , n1725 , n1747 );
or ( n1907 , n1904 , n1905 , n1906 );
xor ( n1908 , n1903 , n1907 );
and ( n1909 , n1750 , n1754 );
and ( n1910 , n1754 , n1769 );
and ( n1911 , n1750 , n1769 );
or ( n1912 , n1909 , n1910 , n1911 );
and ( n1913 , n1732 , n777 );
not ( n1914 , n456 );
and ( n1915 , n1914 , n475 );
and ( n1916 , n459 , n456 );
or ( n1917 , n1915 , n1916 );
buf ( n1918 , n1917 );
buf ( n1919 , n1918 );
and ( n1920 , n1919 , n774 );
nor ( n1921 , n1913 , n1920 );
xnor ( n1922 , n1921 , n750 );
not ( n1923 , n1725 );
and ( n1924 , n1923 , n1900 );
xor ( n1925 , n1922 , n1924 );
and ( n1926 , n1735 , n1739 );
and ( n1927 , n1739 , n1744 );
and ( n1928 , n1735 , n1744 );
or ( n1929 , n1926 , n1927 , n1928 );
xor ( n1930 , n1925 , n1929 );
and ( n1931 , n1759 , n1763 );
and ( n1932 , n1763 , n1768 );
and ( n1933 , n1759 , n1768 );
or ( n1934 , n1931 , n1932 , n1933 );
xor ( n1935 , n1930 , n1934 );
xor ( n1936 , n1912 , n1935 );
and ( n1937 , n1721 , n1748 );
and ( n1938 , n1748 , n1770 );
and ( n1939 , n1721 , n1770 );
or ( n1940 , n1937 , n1938 , n1939 );
xor ( n1941 , n1936 , n1940 );
xor ( n1942 , n1908 , n1941 );
and ( n1943 , n1717 , n1771 );
and ( n1944 , n1771 , n1776 );
and ( n1945 , n1717 , n1776 );
or ( n1946 , n1943 , n1944 , n1945 );
xor ( n1947 , n1942 , n1946 );
and ( n1948 , n1777 , n1778 );
xor ( n1949 , n1947 , n1948 );
buf ( n1950 , n1949 );
not ( n1951 , n455 );
and ( n1952 , n1951 , n1866 );
and ( n1953 , n1950 , n455 );
or ( n1954 , n1952 , n1953 );
and ( n1955 , n1817 , n1834 );
and ( n1956 , n1834 , n1849 );
and ( n1957 , n1817 , n1849 );
or ( n1958 , n1955 , n1956 , n1957 );
and ( n1959 , n1821 , n1825 );
and ( n1960 , n1825 , n1833 );
and ( n1961 , n1821 , n1833 );
or ( n1962 , n1959 , n1960 , n1961 );
and ( n1963 , n1839 , n1843 );
and ( n1964 , n1843 , n1848 );
and ( n1965 , n1839 , n1848 );
or ( n1966 , n1963 , n1964 , n1965 );
xor ( n1967 , n1962 , n1966 );
and ( n1968 , n1791 , n708 );
buf ( n1969 , n506 );
buf ( n1970 , n1969 );
and ( n1971 , n1970 , n705 );
nor ( n1972 , n1968 , n1971 );
xnor ( n1973 , n1972 , n689 );
and ( n1974 , n1540 , n692 );
and ( n1975 , n1672 , n690 );
nor ( n1976 , n1974 , n1975 );
xnor ( n1977 , n1976 , n700 );
xor ( n1978 , n1973 , n1977 );
buf ( n1979 , n490 );
buf ( n1980 , n1979 );
xor ( n1981 , n1980 , n1797 );
and ( n1982 , n682 , n1981 );
xor ( n1983 , n1978 , n1982 );
xor ( n1984 , n1967 , n1983 );
xor ( n1985 , n1958 , n1984 );
and ( n1986 , n1802 , n1806 );
and ( n1987 , n1806 , n1811 );
and ( n1988 , n1802 , n1811 );
or ( n1989 , n1986 , n1987 , n1988 );
and ( n1990 , n1251 , n895 );
and ( n1991 , n1379 , n828 );
nor ( n1992 , n1990 , n1991 );
xnor ( n1993 , n1992 , n885 );
and ( n1994 , n1038 , n1066 );
and ( n1995 , n1164 , n976 );
nor ( n1996 , n1994 , n1995 );
xnor ( n1997 , n1996 , n1047 );
xor ( n1998 , n1993 , n1997 );
and ( n1999 , n876 , n1264 );
and ( n2000 , n965 , n1175 );
nor ( n2001 , n1999 , n2000 );
xnor ( n2002 , n2001 , n1270 );
xor ( n2003 , n1998 , n2002 );
xor ( n2004 , n1989 , n2003 );
and ( n2005 , n1794 , n1801 );
and ( n2006 , n711 , n1522 );
and ( n2007 , n817 , n1411 );
nor ( n2008 , n2006 , n2007 );
xnor ( n2009 , n2008 , n1512 );
xor ( n2010 , n2005 , n2009 );
and ( n2011 , n695 , n1829 );
and ( n2012 , n703 , n1698 );
nor ( n2013 , n2011 , n2012 );
xnor ( n2014 , n2013 , n1800 );
xor ( n2015 , n2010 , n2014 );
xor ( n2016 , n2004 , n2015 );
xor ( n2017 , n1985 , n2016 );
and ( n2018 , n1788 , n1812 );
and ( n2019 , n1812 , n1850 );
and ( n2020 , n1788 , n1850 );
or ( n2021 , n2018 , n2019 , n2020 );
xor ( n2022 , n2017 , n2021 );
and ( n2023 , n1851 , n1855 );
and ( n2024 , n1855 , n1860 );
and ( n2025 , n1851 , n1860 );
or ( n2026 , n2023 , n2024 , n2025 );
xor ( n2027 , n2022 , n2026 );
or ( n2028 , n1861 , n1862 );
xnor ( n2029 , n2027 , n2028 );
and ( n2030 , n1863 , n1864 );
xor ( n2031 , n2029 , n2030 );
buf ( n2032 , n2031 );
and ( n2033 , n1884 , n1888 );
and ( n2034 , n1888 , n1901 );
and ( n2035 , n1884 , n1901 );
or ( n2036 , n2033 , n2034 , n2035 );
and ( n2037 , n1618 , n753 );
and ( n2038 , n1732 , n751 );
nor ( n2039 , n2037 , n2038 );
xnor ( n2040 , n2039 , n765 );
and ( n2041 , n1323 , n924 );
and ( n2042 , n1469 , n856 );
nor ( n2043 , n2041 , n2042 );
xnor ( n2044 , n2043 , n930 );
xor ( n2045 , n2040 , n2044 );
and ( n2046 , n1123 , n1107 );
and ( n2047 , n1213 , n1015 );
nor ( n2048 , n2046 , n2047 );
xnor ( n2049 , n2048 , n1113 );
xor ( n2050 , n2045 , n2049 );
xor ( n2051 , n2036 , n2050 );
and ( n2052 , n1922 , n1924 );
and ( n2053 , n784 , n1588 );
and ( n2054 , n845 , n1446 );
nor ( n2055 , n2053 , n2054 );
xnor ( n2056 , n2055 , n1594 );
xor ( n2057 , n2052 , n2056 );
and ( n2058 , n760 , n1894 );
and ( n2059 , n772 , n1724 );
nor ( n2060 , n2058 , n2059 );
xnor ( n2061 , n2060 , n1900 );
xor ( n2062 , n2057 , n2061 );
xor ( n2063 , n2051 , n2062 );
and ( n2064 , n1912 , n1935 );
and ( n2065 , n1935 , n1940 );
and ( n2066 , n1912 , n1940 );
or ( n2067 , n2064 , n2065 , n2066 );
xor ( n2068 , n2063 , n2067 );
and ( n2069 , n1925 , n1929 );
and ( n2070 , n1929 , n1934 );
and ( n2071 , n1925 , n1934 );
or ( n2072 , n2069 , n2070 , n2071 );
and ( n2073 , n939 , n1346 );
and ( n2074 , n1009 , n1196 );
nor ( n2075 , n2073 , n2074 );
xnor ( n2076 , n2075 , n1352 );
and ( n2077 , n1919 , n777 );
not ( n2078 , n456 );
and ( n2079 , n2078 , n474 );
and ( n2080 , n458 , n456 );
or ( n2081 , n2079 , n2080 );
buf ( n2082 , n2081 );
buf ( n2083 , n2082 );
and ( n2084 , n2083 , n774 );
nor ( n2085 , n2077 , n2084 );
xnor ( n2086 , n2085 , n750 );
buf ( n2087 , n490 );
buf ( n2088 , n2087 );
xor ( n2089 , n2088 , n1891 );
and ( n2090 , n743 , n2089 );
xor ( n2091 , n2086 , n2090 );
xor ( n2092 , n2076 , n2091 );
and ( n2093 , n1870 , n1874 );
and ( n2094 , n1874 , n1879 );
and ( n2095 , n1870 , n1879 );
or ( n2096 , n2093 , n2094 , n2095 );
xor ( n2097 , n2092 , n2096 );
xor ( n2098 , n2072 , n2097 );
and ( n2099 , n1880 , n1902 );
and ( n2100 , n1902 , n1907 );
and ( n2101 , n1880 , n1907 );
or ( n2102 , n2099 , n2100 , n2101 );
xor ( n2103 , n2098 , n2102 );
xor ( n2104 , n2068 , n2103 );
and ( n2105 , n1908 , n1941 );
and ( n2106 , n1941 , n1946 );
and ( n2107 , n1908 , n1946 );
or ( n2108 , n2105 , n2106 , n2107 );
xor ( n2109 , n2104 , n2108 );
and ( n2110 , n1947 , n1948 );
xor ( n2111 , n2109 , n2110 );
buf ( n2112 , n2111 );
not ( n2113 , n455 );
and ( n2114 , n2113 , n2032 );
and ( n2115 , n2112 , n455 );
or ( n2116 , n2114 , n2115 );
and ( n2117 , n1989 , n2003 );
and ( n2118 , n2003 , n2015 );
and ( n2119 , n1989 , n2015 );
or ( n2120 , n2117 , n2118 , n2119 );
and ( n2121 , n1993 , n1997 );
and ( n2122 , n1997 , n2002 );
and ( n2123 , n1993 , n2002 );
or ( n2124 , n2121 , n2122 , n2123 );
and ( n2125 , n1672 , n692 );
and ( n2126 , n1791 , n690 );
nor ( n2127 , n2125 , n2126 );
xnor ( n2128 , n2127 , n700 );
and ( n2129 , n1164 , n1066 );
and ( n2130 , n1251 , n976 );
nor ( n2131 , n2129 , n2130 );
xnor ( n2132 , n2131 , n1047 );
xor ( n2133 , n2128 , n2132 );
buf ( n2134 , n489 );
buf ( n2135 , n2134 );
xor ( n2136 , n2135 , n1980 );
not ( n2137 , n1981 );
and ( n2138 , n2136 , n2137 );
and ( n2139 , n682 , n2138 );
and ( n2140 , n695 , n1981 );
nor ( n2141 , n2139 , n2140 );
and ( n2142 , n1980 , n1797 );
not ( n2143 , n2142 );
and ( n2144 , n2135 , n2143 );
xnor ( n2145 , n2141 , n2144 );
xor ( n2146 , n2133 , n2145 );
xor ( n2147 , n2124 , n2146 );
and ( n2148 , n1379 , n895 );
and ( n2149 , n1540 , n828 );
nor ( n2150 , n2148 , n2149 );
xnor ( n2151 , n2150 , n885 );
and ( n2152 , n965 , n1264 );
and ( n2153 , n1038 , n1175 );
nor ( n2154 , n2152 , n2153 );
xnor ( n2155 , n2154 , n1270 );
xor ( n2156 , n2151 , n2155 );
and ( n2157 , n817 , n1522 );
and ( n2158 , n876 , n1411 );
nor ( n2159 , n2157 , n2158 );
xnor ( n2160 , n2159 , n1512 );
xor ( n2161 , n2156 , n2160 );
xor ( n2162 , n2147 , n2161 );
xor ( n2163 , n2120 , n2162 );
and ( n2164 , n2005 , n2009 );
and ( n2165 , n2009 , n2014 );
and ( n2166 , n2005 , n2014 );
or ( n2167 , n2164 , n2165 , n2166 );
and ( n2168 , n1962 , n1966 );
and ( n2169 , n1966 , n1983 );
and ( n2170 , n1962 , n1983 );
or ( n2171 , n2168 , n2169 , n2170 );
xor ( n2172 , n2167 , n2171 );
and ( n2173 , n1970 , n708 );
buf ( n2174 , n505 );
buf ( n2175 , n2174 );
and ( n2176 , n2175 , n705 );
nor ( n2177 , n2173 , n2176 );
xnor ( n2178 , n2177 , n689 );
not ( n2179 , n1982 );
and ( n2180 , n2179 , n2144 );
xor ( n2181 , n2178 , n2180 );
and ( n2182 , n1973 , n1977 );
and ( n2183 , n1977 , n1982 );
and ( n2184 , n1973 , n1982 );
or ( n2185 , n2182 , n2183 , n2184 );
xor ( n2186 , n2181 , n2185 );
and ( n2187 , n703 , n1829 );
and ( n2188 , n711 , n1698 );
nor ( n2189 , n2187 , n2188 );
xnor ( n2190 , n2189 , n1800 );
xor ( n2191 , n2186 , n2190 );
xor ( n2192 , n2172 , n2191 );
xor ( n2193 , n2163 , n2192 );
and ( n2194 , n1958 , n1984 );
and ( n2195 , n1984 , n2016 );
and ( n2196 , n1958 , n2016 );
or ( n2197 , n2194 , n2195 , n2196 );
xor ( n2198 , n2193 , n2197 );
and ( n2199 , n2017 , n2021 );
and ( n2200 , n2021 , n2026 );
and ( n2201 , n2017 , n2026 );
or ( n2202 , n2199 , n2200 , n2201 );
xor ( n2203 , n2198 , n2202 );
or ( n2204 , n2027 , n2028 );
xnor ( n2205 , n2203 , n2204 );
and ( n2206 , n2029 , n2030 );
xor ( n2207 , n2205 , n2206 );
buf ( n2208 , n2207 );
and ( n2209 , n2063 , n2067 );
and ( n2210 , n2067 , n2103 );
and ( n2211 , n2063 , n2103 );
or ( n2212 , n2209 , n2210 , n2211 );
and ( n2213 , n2083 , n777 );
not ( n2214 , n456 );
and ( n2215 , n2214 , n473 );
and ( n2216 , n457 , n456 );
or ( n2217 , n2215 , n2216 );
buf ( n2218 , n2217 );
buf ( n2219 , n2218 );
and ( n2220 , n2219 , n774 );
nor ( n2221 , n2213 , n2220 );
xnor ( n2222 , n2221 , n750 );
and ( n2223 , n1469 , n924 );
and ( n2224 , n1618 , n856 );
nor ( n2225 , n2223 , n2224 );
xnor ( n2226 , n2225 , n930 );
xor ( n2227 , n2222 , n2226 );
and ( n2228 , n1009 , n1346 );
and ( n2229 , n1123 , n1196 );
nor ( n2230 , n2228 , n2229 );
xnor ( n2231 , n2230 , n1352 );
xor ( n2232 , n2227 , n2231 );
and ( n2233 , n845 , n1588 );
and ( n2234 , n939 , n1446 );
nor ( n2235 , n2233 , n2234 );
xnor ( n2236 , n2235 , n1594 );
and ( n2237 , n772 , n1894 );
and ( n2238 , n784 , n1724 );
nor ( n2239 , n2237 , n2238 );
xnor ( n2240 , n2239 , n1900 );
xor ( n2241 , n2236 , n2240 );
not ( n2242 , n2090 );
buf ( n2243 , n489 );
buf ( n2244 , n2243 );
and ( n2245 , n2088 , n1891 );
not ( n2246 , n2245 );
and ( n2247 , n2244 , n2246 );
and ( n2248 , n2242 , n2247 );
xor ( n2249 , n2241 , n2248 );
xor ( n2250 , n2232 , n2249 );
and ( n2251 , n2052 , n2056 );
and ( n2252 , n2056 , n2061 );
and ( n2253 , n2052 , n2061 );
or ( n2254 , n2251 , n2252 , n2253 );
xor ( n2255 , n2250 , n2254 );
and ( n2256 , n2072 , n2097 );
and ( n2257 , n2097 , n2102 );
and ( n2258 , n2072 , n2102 );
or ( n2259 , n2256 , n2257 , n2258 );
xor ( n2260 , n2255 , n2259 );
and ( n2261 , n2076 , n2091 );
and ( n2262 , n2091 , n2096 );
and ( n2263 , n2076 , n2096 );
or ( n2264 , n2261 , n2262 , n2263 );
and ( n2265 , n1732 , n753 );
and ( n2266 , n1919 , n751 );
nor ( n2267 , n2265 , n2266 );
xnor ( n2268 , n2267 , n765 );
and ( n2269 , n1213 , n1107 );
and ( n2270 , n1323 , n1015 );
nor ( n2271 , n2269 , n2270 );
xnor ( n2272 , n2271 , n1113 );
xor ( n2273 , n2268 , n2272 );
xor ( n2274 , n2244 , n2088 );
not ( n2275 , n2089 );
and ( n2276 , n2274 , n2275 );
and ( n2277 , n743 , n2276 );
and ( n2278 , n760 , n2089 );
nor ( n2279 , n2277 , n2278 );
xnor ( n2280 , n2279 , n2247 );
xor ( n2281 , n2273 , n2280 );
and ( n2282 , n2086 , n2090 );
xor ( n2283 , n2281 , n2282 );
and ( n2284 , n2040 , n2044 );
and ( n2285 , n2044 , n2049 );
and ( n2286 , n2040 , n2049 );
or ( n2287 , n2284 , n2285 , n2286 );
xor ( n2288 , n2283 , n2287 );
xor ( n2289 , n2264 , n2288 );
and ( n2290 , n2036 , n2050 );
and ( n2291 , n2050 , n2062 );
and ( n2292 , n2036 , n2062 );
or ( n2293 , n2290 , n2291 , n2292 );
xor ( n2294 , n2289 , n2293 );
xor ( n2295 , n2260 , n2294 );
xor ( n2296 , n2212 , n2295 );
and ( n2297 , n2104 , n2108 );
and ( n2298 , n2109 , n2110 );
or ( n2299 , n2297 , n2298 );
xor ( n2300 , n2296 , n2299 );
buf ( n2301 , n2300 );
not ( n2302 , n455 );
and ( n2303 , n2302 , n2208 );
and ( n2304 , n2301 , n455 );
or ( n2305 , n2303 , n2304 );
and ( n2306 , n2167 , n2171 );
and ( n2307 , n2171 , n2191 );
and ( n2308 , n2167 , n2191 );
or ( n2309 , n2306 , n2307 , n2308 );
and ( n2310 , n1540 , n895 );
and ( n2311 , n1672 , n828 );
nor ( n2312 , n2310 , n2311 );
xnor ( n2313 , n2312 , n885 );
and ( n2314 , n876 , n1522 );
and ( n2315 , n965 , n1411 );
nor ( n2316 , n2314 , n2315 );
xnor ( n2317 , n2316 , n1512 );
xor ( n2318 , n2313 , n2317 );
and ( n2319 , n711 , n1829 );
and ( n2320 , n817 , n1698 );
nor ( n2321 , n2319 , n2320 );
xnor ( n2322 , n2321 , n1800 );
xor ( n2323 , n2318 , n2322 );
and ( n2324 , n2175 , n708 );
not ( n2325 , n2324 );
xnor ( n2326 , n2325 , n689 );
and ( n2327 , n1791 , n692 );
and ( n2328 , n1970 , n690 );
nor ( n2329 , n2327 , n2328 );
xnor ( n2330 , n2329 , n700 );
xor ( n2331 , n2326 , n2330 );
and ( n2332 , n682 , n2135 );
xor ( n2333 , n2331 , n2332 );
xor ( n2334 , n2323 , n2333 );
and ( n2335 , n1251 , n1066 );
and ( n2336 , n1379 , n976 );
nor ( n2337 , n2335 , n2336 );
xnor ( n2338 , n2337 , n1047 );
and ( n2339 , n1038 , n1264 );
and ( n2340 , n1164 , n1175 );
nor ( n2341 , n2339 , n2340 );
xnor ( n2342 , n2341 , n1270 );
xor ( n2343 , n2338 , n2342 );
and ( n2344 , n695 , n2138 );
and ( n2345 , n703 , n1981 );
nor ( n2346 , n2344 , n2345 );
xnor ( n2347 , n2346 , n2144 );
xor ( n2348 , n2343 , n2347 );
xor ( n2349 , n2334 , n2348 );
xor ( n2350 , n2309 , n2349 );
and ( n2351 , n2181 , n2185 );
and ( n2352 , n2185 , n2190 );
and ( n2353 , n2181 , n2190 );
or ( n2354 , n2351 , n2352 , n2353 );
and ( n2355 , n2124 , n2146 );
and ( n2356 , n2146 , n2161 );
and ( n2357 , n2124 , n2161 );
or ( n2358 , n2355 , n2356 , n2357 );
xor ( n2359 , n2354 , n2358 );
and ( n2360 , n2128 , n2132 );
and ( n2361 , n2132 , n2145 );
and ( n2362 , n2128 , n2145 );
or ( n2363 , n2360 , n2361 , n2362 );
and ( n2364 , n2151 , n2155 );
and ( n2365 , n2155 , n2160 );
and ( n2366 , n2151 , n2160 );
or ( n2367 , n2364 , n2365 , n2366 );
xor ( n2368 , n2363 , n2367 );
and ( n2369 , n2178 , n2180 );
xor ( n2370 , n2368 , n2369 );
xor ( n2371 , n2359 , n2370 );
xor ( n2372 , n2350 , n2371 );
and ( n2373 , n2120 , n2162 );
and ( n2374 , n2162 , n2192 );
and ( n2375 , n2120 , n2192 );
or ( n2376 , n2373 , n2374 , n2375 );
xor ( n2377 , n2372 , n2376 );
and ( n2378 , n2193 , n2197 );
and ( n2379 , n2197 , n2202 );
and ( n2380 , n2193 , n2202 );
or ( n2381 , n2378 , n2379 , n2380 );
xor ( n2382 , n2377 , n2381 );
or ( n2383 , n2203 , n2204 );
xnor ( n2384 , n2382 , n2383 );
and ( n2385 , n2205 , n2206 );
xor ( n2386 , n2384 , n2385 );
buf ( n2387 , n2386 );
and ( n2388 , n2255 , n2259 );
and ( n2389 , n2259 , n2294 );
and ( n2390 , n2255 , n2294 );
or ( n2391 , n2388 , n2389 , n2390 );
and ( n2392 , n2232 , n2249 );
and ( n2393 , n2249 , n2254 );
and ( n2394 , n2232 , n2254 );
or ( n2395 , n2392 , n2393 , n2394 );
and ( n2396 , n2281 , n2282 );
and ( n2397 , n2282 , n2287 );
and ( n2398 , n2281 , n2287 );
or ( n2399 , n2396 , n2397 , n2398 );
and ( n2400 , n2268 , n2272 );
and ( n2401 , n2272 , n2280 );
and ( n2402 , n2268 , n2280 );
or ( n2403 , n2400 , n2401 , n2402 );
and ( n2404 , n2222 , n2226 );
and ( n2405 , n2226 , n2231 );
and ( n2406 , n2222 , n2231 );
or ( n2407 , n2404 , n2405 , n2406 );
xor ( n2408 , n2403 , n2407 );
and ( n2409 , n2236 , n2240 );
and ( n2410 , n2240 , n2248 );
and ( n2411 , n2236 , n2248 );
or ( n2412 , n2409 , n2410 , n2411 );
xor ( n2413 , n2408 , n2412 );
xor ( n2414 , n2399 , n2413 );
and ( n2415 , n2219 , n777 );
not ( n2416 , n2415 );
xnor ( n2417 , n2416 , n750 );
and ( n2418 , n1919 , n753 );
and ( n2419 , n2083 , n751 );
nor ( n2420 , n2418 , n2419 );
xnor ( n2421 , n2420 , n765 );
xor ( n2422 , n2417 , n2421 );
and ( n2423 , n1618 , n924 );
and ( n2424 , n1732 , n856 );
nor ( n2425 , n2423 , n2424 );
xnor ( n2426 , n2425 , n930 );
xor ( n2427 , n2422 , n2426 );
and ( n2428 , n1323 , n1107 );
and ( n2429 , n1469 , n1015 );
nor ( n2430 , n2428 , n2429 );
xnor ( n2431 , n2430 , n1113 );
and ( n2432 , n1123 , n1346 );
and ( n2433 , n1213 , n1196 );
nor ( n2434 , n2432 , n2433 );
xnor ( n2435 , n2434 , n1352 );
xor ( n2436 , n2431 , n2435 );
and ( n2437 , n939 , n1588 );
and ( n2438 , n1009 , n1446 );
nor ( n2439 , n2437 , n2438 );
xnor ( n2440 , n2439 , n1594 );
xor ( n2441 , n2436 , n2440 );
xor ( n2442 , n2427 , n2441 );
and ( n2443 , n784 , n1894 );
and ( n2444 , n845 , n1724 );
nor ( n2445 , n2443 , n2444 );
xnor ( n2446 , n2445 , n1900 );
and ( n2447 , n760 , n2276 );
and ( n2448 , n772 , n2089 );
nor ( n2449 , n2447 , n2448 );
xnor ( n2450 , n2449 , n2247 );
xor ( n2451 , n2446 , n2450 );
and ( n2452 , n743 , n2244 );
xor ( n2453 , n2451 , n2452 );
xor ( n2454 , n2442 , n2453 );
xor ( n2455 , n2414 , n2454 );
xor ( n2456 , n2395 , n2455 );
and ( n2457 , n2264 , n2288 );
and ( n2458 , n2288 , n2293 );
and ( n2459 , n2264 , n2293 );
or ( n2460 , n2457 , n2458 , n2459 );
xor ( n2461 , n2456 , n2460 );
xor ( n2462 , n2391 , n2461 );
and ( n2463 , n2212 , n2295 );
and ( n2464 , n2296 , n2299 );
or ( n2465 , n2463 , n2464 );
xor ( n2466 , n2462 , n2465 );
buf ( n2467 , n2466 );
not ( n2468 , n455 );
and ( n2469 , n2468 , n2387 );
and ( n2470 , n2467 , n455 );
or ( n2471 , n2469 , n2470 );
and ( n2472 , n2354 , n2358 );
and ( n2473 , n2358 , n2370 );
and ( n2474 , n2354 , n2370 );
or ( n2475 , n2472 , n2473 , n2474 );
and ( n2476 , n2363 , n2367 );
and ( n2477 , n2367 , n2369 );
and ( n2478 , n2363 , n2369 );
or ( n2479 , n2476 , n2477 , n2478 );
not ( n2480 , n689 );
and ( n2481 , n703 , n2138 );
and ( n2482 , n711 , n1981 );
nor ( n2483 , n2481 , n2482 );
xnor ( n2484 , n2483 , n2144 );
xor ( n2485 , n2480 , n2484 );
and ( n2486 , n695 , n2135 );
xor ( n2487 , n2485 , n2486 );
xor ( n2488 , n2479 , n2487 );
and ( n2489 , n1970 , n692 );
and ( n2490 , n2175 , n690 );
nor ( n2491 , n2489 , n2490 );
xnor ( n2492 , n2491 , n700 );
and ( n2493 , n1672 , n895 );
and ( n2494 , n1791 , n828 );
nor ( n2495 , n2493 , n2494 );
xnor ( n2496 , n2495 , n885 );
xor ( n2497 , n2492 , n2496 );
and ( n2498 , n1164 , n1264 );
and ( n2499 , n1251 , n1175 );
nor ( n2500 , n2498 , n2499 );
xnor ( n2501 , n2500 , n1270 );
xor ( n2502 , n2497 , n2501 );
xor ( n2503 , n2488 , n2502 );
xor ( n2504 , n2475 , n2503 );
and ( n2505 , n2323 , n2333 );
and ( n2506 , n2333 , n2348 );
and ( n2507 , n2323 , n2348 );
or ( n2508 , n2505 , n2506 , n2507 );
and ( n2509 , n2313 , n2317 );
and ( n2510 , n2317 , n2322 );
and ( n2511 , n2313 , n2322 );
or ( n2512 , n2509 , n2510 , n2511 );
and ( n2513 , n2326 , n2330 );
and ( n2514 , n2330 , n2332 );
and ( n2515 , n2326 , n2332 );
or ( n2516 , n2513 , n2514 , n2515 );
xor ( n2517 , n2512 , n2516 );
and ( n2518 , n2338 , n2342 );
and ( n2519 , n2342 , n2347 );
and ( n2520 , n2338 , n2347 );
or ( n2521 , n2518 , n2519 , n2520 );
xor ( n2522 , n2517 , n2521 );
xor ( n2523 , n2508 , n2522 );
and ( n2524 , n1379 , n1066 );
and ( n2525 , n1540 , n976 );
nor ( n2526 , n2524 , n2525 );
xnor ( n2527 , n2526 , n1047 );
not ( n2528 , n2527 );
and ( n2529 , n965 , n1522 );
and ( n2530 , n1038 , n1411 );
nor ( n2531 , n2529 , n2530 );
xnor ( n2532 , n2531 , n1512 );
xor ( n2533 , n2528 , n2532 );
and ( n2534 , n817 , n1829 );
and ( n2535 , n876 , n1698 );
nor ( n2536 , n2534 , n2535 );
xnor ( n2537 , n2536 , n1800 );
xor ( n2538 , n2533 , n2537 );
xor ( n2539 , n2523 , n2538 );
xor ( n2540 , n2504 , n2539 );
and ( n2541 , n2309 , n2349 );
and ( n2542 , n2349 , n2371 );
and ( n2543 , n2309 , n2371 );
or ( n2544 , n2541 , n2542 , n2543 );
xor ( n2545 , n2540 , n2544 );
and ( n2546 , n2372 , n2376 );
and ( n2547 , n2376 , n2381 );
and ( n2548 , n2372 , n2381 );
or ( n2549 , n2546 , n2547 , n2548 );
xor ( n2550 , n2545 , n2549 );
or ( n2551 , n2382 , n2383 );
xnor ( n2552 , n2550 , n2551 );
and ( n2553 , n2384 , n2385 );
xor ( n2554 , n2552 , n2553 );
buf ( n2555 , n2554 );
and ( n2556 , n2399 , n2413 );
and ( n2557 , n2413 , n2454 );
and ( n2558 , n2399 , n2454 );
or ( n2559 , n2556 , n2557 , n2558 );
and ( n2560 , n2083 , n753 );
and ( n2561 , n2219 , n751 );
nor ( n2562 , n2560 , n2561 );
xnor ( n2563 , n2562 , n765 );
and ( n2564 , n1732 , n924 );
and ( n2565 , n1919 , n856 );
nor ( n2566 , n2564 , n2565 );
xnor ( n2567 , n2566 , n930 );
xor ( n2568 , n2563 , n2567 );
and ( n2569 , n1469 , n1107 );
and ( n2570 , n1618 , n1015 );
nor ( n2571 , n2569 , n2570 );
xnor ( n2572 , n2571 , n1113 );
xor ( n2573 , n2568 , n2572 );
and ( n2574 , n1213 , n1346 );
and ( n2575 , n1323 , n1196 );
nor ( n2576 , n2574 , n2575 );
xnor ( n2577 , n2576 , n1352 );
and ( n2578 , n1009 , n1588 );
and ( n2579 , n1123 , n1446 );
nor ( n2580 , n2578 , n2579 );
xnor ( n2581 , n2580 , n1594 );
xor ( n2582 , n2577 , n2581 );
and ( n2583 , n845 , n1894 );
and ( n2584 , n939 , n1724 );
nor ( n2585 , n2583 , n2584 );
xnor ( n2586 , n2585 , n1900 );
xor ( n2587 , n2582 , n2586 );
xor ( n2588 , n2573 , n2587 );
and ( n2589 , n2403 , n2407 );
and ( n2590 , n2407 , n2412 );
and ( n2591 , n2403 , n2412 );
or ( n2592 , n2589 , n2590 , n2591 );
xor ( n2593 , n2588 , n2592 );
xor ( n2594 , n2559 , n2593 );
and ( n2595 , n2427 , n2441 );
and ( n2596 , n2441 , n2453 );
and ( n2597 , n2427 , n2453 );
or ( n2598 , n2595 , n2596 , n2597 );
and ( n2599 , n772 , n2276 );
and ( n2600 , n784 , n2089 );
nor ( n2601 , n2599 , n2600 );
xnor ( n2602 , n2601 , n2247 );
and ( n2603 , n760 , n2244 );
xor ( n2604 , n2602 , n2603 );
xor ( n2605 , n2604 , n750 );
xor ( n2606 , n2598 , n2605 );
and ( n2607 , n2417 , n2421 );
and ( n2608 , n2421 , n2426 );
and ( n2609 , n2417 , n2426 );
or ( n2610 , n2607 , n2608 , n2609 );
and ( n2611 , n2431 , n2435 );
and ( n2612 , n2435 , n2440 );
and ( n2613 , n2431 , n2440 );
or ( n2614 , n2611 , n2612 , n2613 );
xor ( n2615 , n2610 , n2614 );
and ( n2616 , n2446 , n2450 );
and ( n2617 , n2450 , n2452 );
and ( n2618 , n2446 , n2452 );
or ( n2619 , n2616 , n2617 , n2618 );
xor ( n2620 , n2615 , n2619 );
xor ( n2621 , n2606 , n2620 );
xor ( n2622 , n2594 , n2621 );
and ( n2623 , n2395 , n2455 );
and ( n2624 , n2455 , n2460 );
and ( n2625 , n2395 , n2460 );
or ( n2626 , n2623 , n2624 , n2625 );
xor ( n2627 , n2622 , n2626 );
and ( n2628 , n2391 , n2461 );
and ( n2629 , n2462 , n2465 );
or ( n2630 , n2628 , n2629 );
xor ( n2631 , n2627 , n2630 );
buf ( n2632 , n2631 );
not ( n2633 , n455 );
and ( n2634 , n2633 , n2555 );
and ( n2635 , n2632 , n455 );
or ( n2636 , n2634 , n2635 );
and ( n2637 , n2508 , n2522 );
and ( n2638 , n2522 , n2538 );
and ( n2639 , n2508 , n2538 );
or ( n2640 , n2637 , n2638 , n2639 );
and ( n2641 , n2512 , n2516 );
and ( n2642 , n2516 , n2521 );
and ( n2643 , n2512 , n2521 );
or ( n2644 , n2641 , n2642 , n2643 );
and ( n2645 , n1791 , n895 );
and ( n2646 , n1970 , n828 );
nor ( n2647 , n2645 , n2646 );
xnor ( n2648 , n2647 , n885 );
and ( n2649 , n1251 , n1264 );
and ( n2650 , n1379 , n1175 );
nor ( n2651 , n2649 , n2650 );
xnor ( n2652 , n2651 , n1270 );
xor ( n2653 , n2648 , n2652 );
and ( n2654 , n703 , n2135 );
xor ( n2655 , n2653 , n2654 );
xor ( n2656 , n2644 , n2655 );
buf ( n2657 , n2527 );
and ( n2658 , n2175 , n692 );
not ( n2659 , n2658 );
xnor ( n2660 , n2659 , n700 );
not ( n2661 , n2660 );
xor ( n2662 , n2657 , n2661 );
and ( n2663 , n711 , n2138 );
and ( n2664 , n817 , n1981 );
nor ( n2665 , n2663 , n2664 );
xnor ( n2666 , n2665 , n2144 );
xor ( n2667 , n2662 , n2666 );
xor ( n2668 , n2656 , n2667 );
xnor ( n2669 , n2640 , n2668 );
and ( n2670 , n2475 , n2503 );
and ( n2671 , n2503 , n2539 );
and ( n2672 , n2475 , n2539 );
or ( n2673 , n2670 , n2671 , n2672 );
xor ( n2674 , n2669 , n2673 );
and ( n2675 , n2528 , n2532 );
and ( n2676 , n2532 , n2537 );
and ( n2677 , n2528 , n2537 );
or ( n2678 , n2675 , n2676 , n2677 );
and ( n2679 , n2480 , n2484 );
and ( n2680 , n2484 , n2486 );
and ( n2681 , n2480 , n2486 );
or ( n2682 , n2679 , n2680 , n2681 );
and ( n2683 , n2492 , n2496 );
and ( n2684 , n2496 , n2501 );
and ( n2685 , n2492 , n2501 );
or ( n2686 , n2683 , n2684 , n2685 );
xor ( n2687 , n2682 , n2686 );
and ( n2688 , n1540 , n1066 );
and ( n2689 , n1672 , n976 );
nor ( n2690 , n2688 , n2689 );
xnor ( n2691 , n2690 , n1047 );
and ( n2692 , n1038 , n1522 );
and ( n2693 , n1164 , n1411 );
nor ( n2694 , n2692 , n2693 );
xnor ( n2695 , n2694 , n1512 );
xor ( n2696 , n2691 , n2695 );
and ( n2697 , n876 , n1829 );
and ( n2698 , n965 , n1698 );
nor ( n2699 , n2697 , n2698 );
xnor ( n2700 , n2699 , n1800 );
xor ( n2701 , n2696 , n2700 );
xor ( n2702 , n2687 , n2701 );
xor ( n2703 , n2678 , n2702 );
and ( n2704 , n2479 , n2487 );
and ( n2705 , n2487 , n2502 );
and ( n2706 , n2479 , n2502 );
or ( n2707 , n2704 , n2705 , n2706 );
xor ( n2708 , n2703 , n2707 );
xor ( n2709 , n2674 , n2708 );
and ( n2710 , n2540 , n2544 );
and ( n2711 , n2544 , n2549 );
and ( n2712 , n2540 , n2549 );
or ( n2713 , n2710 , n2711 , n2712 );
xor ( n2714 , n2709 , n2713 );
or ( n2715 , n2550 , n2551 );
xor ( n2716 , n2714 , n2715 );
and ( n2717 , n2552 , n2553 );
xor ( n2718 , n2716 , n2717 );
buf ( n2719 , n2718 );
and ( n2720 , n2610 , n2614 );
and ( n2721 , n2614 , n2619 );
and ( n2722 , n2610 , n2619 );
or ( n2723 , n2720 , n2721 , n2722 );
and ( n2724 , n2563 , n2567 );
and ( n2725 , n2567 , n2572 );
and ( n2726 , n2563 , n2572 );
or ( n2727 , n2724 , n2725 , n2726 );
and ( n2728 , n2577 , n2581 );
and ( n2729 , n2581 , n2586 );
and ( n2730 , n2577 , n2586 );
or ( n2731 , n2728 , n2729 , n2730 );
xor ( n2732 , n2727 , n2731 );
and ( n2733 , n1919 , n924 );
and ( n2734 , n2083 , n856 );
nor ( n2735 , n2733 , n2734 );
xnor ( n2736 , n2735 , n930 );
and ( n2737 , n1618 , n1107 );
and ( n2738 , n1732 , n1015 );
nor ( n2739 , n2737 , n2738 );
xnor ( n2740 , n2739 , n1113 );
xor ( n2741 , n2736 , n2740 );
and ( n2742 , n1323 , n1346 );
and ( n2743 , n1469 , n1196 );
nor ( n2744 , n2742 , n2743 );
xnor ( n2745 , n2744 , n1352 );
xor ( n2746 , n2741 , n2745 );
xor ( n2747 , n2732 , n2746 );
xor ( n2748 , n2723 , n2747 );
and ( n2749 , n2573 , n2587 );
and ( n2750 , n2587 , n2592 );
and ( n2751 , n2573 , n2592 );
or ( n2752 , n2749 , n2750 , n2751 );
xor ( n2753 , n2748 , n2752 );
and ( n2754 , n2598 , n2605 );
and ( n2755 , n2605 , n2620 );
and ( n2756 , n2598 , n2620 );
or ( n2757 , n2754 , n2755 , n2756 );
and ( n2758 , n1123 , n1588 );
and ( n2759 , n1213 , n1446 );
nor ( n2760 , n2758 , n2759 );
xnor ( n2761 , n2760 , n1594 );
and ( n2762 , n939 , n1894 );
and ( n2763 , n1009 , n1724 );
nor ( n2764 , n2762 , n2763 );
xnor ( n2765 , n2764 , n1900 );
xor ( n2766 , n2761 , n2765 );
and ( n2767 , n772 , n2244 );
xor ( n2768 , n2766 , n2767 );
not ( n2769 , n750 );
buf ( n2770 , n2769 );
and ( n2771 , n2219 , n753 );
not ( n2772 , n2771 );
xnor ( n2773 , n2772 , n765 );
not ( n2774 , n2773 );
xor ( n2775 , n2770 , n2774 );
and ( n2776 , n784 , n2276 );
and ( n2777 , n845 , n2089 );
nor ( n2778 , n2776 , n2777 );
xnor ( n2779 , n2778 , n2247 );
xor ( n2780 , n2775 , n2779 );
xor ( n2781 , n2768 , n2780 );
and ( n2782 , n2602 , n2603 );
and ( n2783 , n2603 , n750 );
and ( n2784 , n2602 , n750 );
or ( n2785 , n2782 , n2783 , n2784 );
xor ( n2786 , n2781 , n2785 );
xor ( n2787 , n2757 , n2786 );
and ( n2788 , n2559 , n2593 );
and ( n2789 , n2593 , n2621 );
and ( n2790 , n2559 , n2621 );
or ( n2791 , n2788 , n2789 , n2790 );
xor ( n2792 , n2787 , n2791 );
xor ( n2793 , n2753 , n2792 );
and ( n2794 , n2622 , n2626 );
and ( n2795 , n2627 , n2630 );
or ( n2796 , n2794 , n2795 );
xor ( n2797 , n2793 , n2796 );
buf ( n2798 , n2797 );
not ( n2799 , n455 );
and ( n2800 , n2799 , n2719 );
and ( n2801 , n2798 , n455 );
or ( n2802 , n2800 , n2801 );
and ( n2803 , n2678 , n2702 );
and ( n2804 , n2702 , n2707 );
and ( n2805 , n2678 , n2707 );
or ( n2806 , n2803 , n2804 , n2805 );
and ( n2807 , n2669 , n2673 );
and ( n2808 , n2673 , n2708 );
and ( n2809 , n2669 , n2708 );
or ( n2810 , n2807 , n2808 , n2809 );
xor ( n2811 , n2806 , n2810 );
and ( n2812 , n2657 , n2661 );
and ( n2813 , n2661 , n2666 );
and ( n2814 , n2657 , n2666 );
or ( n2815 , n2812 , n2813 , n2814 );
and ( n2816 , n1672 , n1066 );
and ( n2817 , n1791 , n976 );
nor ( n2818 , n2816 , n2817 );
xnor ( n2819 , n2818 , n1047 );
and ( n2820 , n1164 , n1522 );
and ( n2821 , n1251 , n1411 );
nor ( n2822 , n2820 , n2821 );
xnor ( n2823 , n2822 , n1512 );
xor ( n2824 , n2819 , n2823 );
and ( n2825 , n711 , n2135 );
xor ( n2826 , n2824 , n2825 );
xor ( n2827 , n2815 , n2826 );
buf ( n2828 , n2660 );
and ( n2829 , n965 , n1829 );
and ( n2830 , n1038 , n1698 );
nor ( n2831 , n2829 , n2830 );
xnor ( n2832 , n2831 , n1800 );
xor ( n2833 , n2828 , n2832 );
and ( n2834 , n817 , n2138 );
and ( n2835 , n876 , n1981 );
nor ( n2836 , n2834 , n2835 );
xnor ( n2837 , n2836 , n2144 );
xor ( n2838 , n2833 , n2837 );
xor ( n2839 , n2827 , n2838 );
and ( n2840 , n2682 , n2686 );
and ( n2841 , n2686 , n2701 );
and ( n2842 , n2682 , n2701 );
or ( n2843 , n2840 , n2841 , n2842 );
and ( n2844 , n2644 , n2655 );
and ( n2845 , n2655 , n2667 );
and ( n2846 , n2644 , n2667 );
or ( n2847 , n2844 , n2845 , n2846 );
xor ( n2848 , n2843 , n2847 );
and ( n2849 , n2648 , n2652 );
and ( n2850 , n2652 , n2654 );
and ( n2851 , n2648 , n2654 );
or ( n2852 , n2849 , n2850 , n2851 );
and ( n2853 , n2691 , n2695 );
and ( n2854 , n2695 , n2700 );
and ( n2855 , n2691 , n2700 );
or ( n2856 , n2853 , n2854 , n2855 );
xor ( n2857 , n2852 , n2856 );
not ( n2858 , n700 );
and ( n2859 , n1970 , n895 );
and ( n2860 , n2175 , n828 );
nor ( n2861 , n2859 , n2860 );
xnor ( n2862 , n2861 , n885 );
xor ( n2863 , n2858 , n2862 );
and ( n2864 , n1379 , n1264 );
and ( n2865 , n1540 , n1175 );
nor ( n2866 , n2864 , n2865 );
xnor ( n2867 , n2866 , n1270 );
xor ( n2868 , n2863 , n2867 );
xor ( n2869 , n2857 , n2868 );
xor ( n2870 , n2848 , n2869 );
xor ( n2871 , n2839 , n2870 );
or ( n2872 , n2640 , n2668 );
xor ( n2873 , n2871 , n2872 );
xor ( n2874 , n2811 , n2873 );
and ( n2875 , n2709 , n2713 );
and ( n2876 , n2713 , n2715 );
and ( n2877 , n2709 , n2715 );
or ( n2878 , n2875 , n2876 , n2877 );
xnor ( n2879 , n2874 , n2878 );
and ( n2880 , n2716 , n2717 );
xor ( n2881 , n2879 , n2880 );
buf ( n2882 , n2881 );
and ( n2883 , n2757 , n2786 );
and ( n2884 , n2786 , n2791 );
and ( n2885 , n2757 , n2791 );
or ( n2886 , n2883 , n2884 , n2885 );
and ( n2887 , n2770 , n2774 );
and ( n2888 , n2774 , n2779 );
and ( n2889 , n2770 , n2779 );
or ( n2890 , n2887 , n2888 , n2889 );
and ( n2891 , n1732 , n1107 );
and ( n2892 , n1919 , n1015 );
nor ( n2893 , n2891 , n2892 );
xnor ( n2894 , n2893 , n1113 );
and ( n2895 , n1213 , n1588 );
and ( n2896 , n1323 , n1446 );
nor ( n2897 , n2895 , n2896 );
xnor ( n2898 , n2897 , n1594 );
xor ( n2899 , n2894 , n2898 );
and ( n2900 , n784 , n2244 );
xor ( n2901 , n2899 , n2900 );
xor ( n2902 , n2890 , n2901 );
buf ( n2903 , n2773 );
and ( n2904 , n1009 , n1894 );
and ( n2905 , n1123 , n1724 );
nor ( n2906 , n2904 , n2905 );
xnor ( n2907 , n2906 , n1900 );
xor ( n2908 , n2903 , n2907 );
and ( n2909 , n845 , n2276 );
and ( n2910 , n939 , n2089 );
nor ( n2911 , n2909 , n2910 );
xnor ( n2912 , n2911 , n2247 );
xor ( n2913 , n2908 , n2912 );
xor ( n2914 , n2902 , n2913 );
and ( n2915 , n2723 , n2747 );
and ( n2916 , n2747 , n2752 );
and ( n2917 , n2723 , n2752 );
or ( n2918 , n2915 , n2916 , n2917 );
xor ( n2919 , n2914 , n2918 );
and ( n2920 , n2727 , n2731 );
and ( n2921 , n2731 , n2746 );
and ( n2922 , n2727 , n2746 );
or ( n2923 , n2920 , n2921 , n2922 );
not ( n2924 , n765 );
and ( n2925 , n2083 , n924 );
and ( n2926 , n2219 , n856 );
nor ( n2927 , n2925 , n2926 );
xnor ( n2928 , n2927 , n930 );
xor ( n2929 , n2924 , n2928 );
and ( n2930 , n1469 , n1346 );
and ( n2931 , n1618 , n1196 );
nor ( n2932 , n2930 , n2931 );
xnor ( n2933 , n2932 , n1352 );
xor ( n2934 , n2929 , n2933 );
and ( n2935 , n2736 , n2740 );
and ( n2936 , n2740 , n2745 );
and ( n2937 , n2736 , n2745 );
or ( n2938 , n2935 , n2936 , n2937 );
xor ( n2939 , n2934 , n2938 );
and ( n2940 , n2761 , n2765 );
and ( n2941 , n2765 , n2767 );
and ( n2942 , n2761 , n2767 );
or ( n2943 , n2940 , n2941 , n2942 );
xor ( n2944 , n2939 , n2943 );
xor ( n2945 , n2923 , n2944 );
and ( n2946 , n2768 , n2780 );
and ( n2947 , n2780 , n2785 );
and ( n2948 , n2768 , n2785 );
or ( n2949 , n2946 , n2947 , n2948 );
xor ( n2950 , n2945 , n2949 );
xor ( n2951 , n2919 , n2950 );
xor ( n2952 , n2886 , n2951 );
and ( n2953 , n2753 , n2792 );
and ( n2954 , n2793 , n2796 );
or ( n2955 , n2953 , n2954 );
xor ( n2956 , n2952 , n2955 );
buf ( n2957 , n2956 );
not ( n2958 , n455 );
and ( n2959 , n2958 , n2882 );
and ( n2960 , n2957 , n455 );
or ( n2961 , n2959 , n2960 );
and ( n2962 , n2839 , n2870 );
and ( n2963 , n2870 , n2872 );
and ( n2964 , n2839 , n2872 );
or ( n2965 , n2962 , n2963 , n2964 );
and ( n2966 , n2815 , n2826 );
and ( n2967 , n2826 , n2838 );
and ( n2968 , n2815 , n2838 );
or ( n2969 , n2966 , n2967 , n2968 );
and ( n2970 , n2843 , n2847 );
and ( n2971 , n2847 , n2869 );
and ( n2972 , n2843 , n2869 );
or ( n2973 , n2970 , n2971 , n2972 );
xor ( n2974 , n2969 , n2973 );
and ( n2975 , n2852 , n2856 );
and ( n2976 , n2856 , n2868 );
and ( n2977 , n2852 , n2868 );
or ( n2978 , n2975 , n2976 , n2977 );
and ( n2979 , n2819 , n2823 );
and ( n2980 , n2823 , n2825 );
and ( n2981 , n2819 , n2825 );
or ( n2982 , n2979 , n2980 , n2981 );
and ( n2983 , n2858 , n2862 );
and ( n2984 , n2862 , n2867 );
and ( n2985 , n2858 , n2867 );
or ( n2986 , n2983 , n2984 , n2985 );
xor ( n2987 , n2982 , n2986 );
and ( n2988 , n2175 , n895 );
not ( n2989 , n2988 );
xnor ( n2990 , n2989 , n885 );
not ( n2991 , n2990 );
xor ( n2992 , n2987 , n2991 );
xor ( n2993 , n2978 , n2992 );
and ( n2994 , n2828 , n2832 );
and ( n2995 , n2832 , n2837 );
and ( n2996 , n2828 , n2837 );
or ( n2997 , n2994 , n2995 , n2996 );
and ( n2998 , n1540 , n1264 );
and ( n2999 , n1672 , n1175 );
nor ( n3000 , n2998 , n2999 );
xnor ( n3001 , n3000 , n1270 );
and ( n3002 , n876 , n2138 );
and ( n3003 , n965 , n1981 );
nor ( n3004 , n3002 , n3003 );
xnor ( n3005 , n3004 , n2144 );
xor ( n3006 , n3001 , n3005 );
and ( n3007 , n817 , n2135 );
xor ( n3008 , n3006 , n3007 );
xor ( n3009 , n2997 , n3008 );
and ( n3010 , n1791 , n1066 );
and ( n3011 , n1970 , n976 );
nor ( n3012 , n3010 , n3011 );
xnor ( n3013 , n3012 , n1047 );
and ( n3014 , n1251 , n1522 );
and ( n3015 , n1379 , n1411 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n1512 );
xor ( n3018 , n3013 , n3017 );
and ( n3019 , n1038 , n1829 );
and ( n3020 , n1164 , n1698 );
nor ( n3021 , n3019 , n3020 );
xnor ( n3022 , n3021 , n1800 );
xor ( n3023 , n3018 , n3022 );
xor ( n3024 , n3009 , n3023 );
xor ( n3025 , n2993 , n3024 );
xor ( n3026 , n2974 , n3025 );
xor ( n3027 , n2965 , n3026 );
and ( n3028 , n2806 , n2810 );
and ( n3029 , n2810 , n2873 );
and ( n3030 , n2806 , n2873 );
or ( n3031 , n3028 , n3029 , n3030 );
xor ( n3032 , n3027 , n3031 );
or ( n3033 , n2874 , n2878 );
xnor ( n3034 , n3032 , n3033 );
and ( n3035 , n2879 , n2880 );
xor ( n3036 , n3034 , n3035 );
buf ( n3037 , n3036 );
and ( n3038 , n2924 , n2928 );
and ( n3039 , n2928 , n2933 );
and ( n3040 , n2924 , n2933 );
or ( n3041 , n3038 , n3039 , n3040 );
and ( n3042 , n2894 , n2898 );
and ( n3043 , n2898 , n2900 );
and ( n3044 , n2894 , n2900 );
or ( n3045 , n3042 , n3043 , n3044 );
xor ( n3046 , n3041 , n3045 );
and ( n3047 , n2219 , n924 );
not ( n3048 , n3047 );
xnor ( n3049 , n3048 , n930 );
not ( n3050 , n3049 );
xor ( n3051 , n3046 , n3050 );
and ( n3052 , n2934 , n2938 );
and ( n3053 , n2938 , n2943 );
and ( n3054 , n2934 , n2943 );
or ( n3055 , n3052 , n3053 , n3054 );
xor ( n3056 , n3051 , n3055 );
and ( n3057 , n2903 , n2907 );
and ( n3058 , n2907 , n2912 );
and ( n3059 , n2903 , n2912 );
or ( n3060 , n3057 , n3058 , n3059 );
and ( n3061 , n1618 , n1346 );
and ( n3062 , n1732 , n1196 );
nor ( n3063 , n3061 , n3062 );
xnor ( n3064 , n3063 , n1352 );
and ( n3065 , n939 , n2276 );
and ( n3066 , n1009 , n2089 );
nor ( n3067 , n3065 , n3066 );
xnor ( n3068 , n3067 , n2247 );
xor ( n3069 , n3064 , n3068 );
and ( n3070 , n845 , n2244 );
xor ( n3071 , n3069 , n3070 );
xor ( n3072 , n3060 , n3071 );
and ( n3073 , n1919 , n1107 );
and ( n3074 , n2083 , n1015 );
nor ( n3075 , n3073 , n3074 );
xnor ( n3076 , n3075 , n1113 );
and ( n3077 , n1323 , n1588 );
and ( n3078 , n1469 , n1446 );
nor ( n3079 , n3077 , n3078 );
xnor ( n3080 , n3079 , n1594 );
xor ( n3081 , n3076 , n3080 );
and ( n3082 , n1123 , n1894 );
and ( n3083 , n1213 , n1724 );
nor ( n3084 , n3082 , n3083 );
xnor ( n3085 , n3084 , n1900 );
xor ( n3086 , n3081 , n3085 );
xor ( n3087 , n3072 , n3086 );
xor ( n3088 , n3056 , n3087 );
and ( n3089 , n2890 , n2901 );
and ( n3090 , n2901 , n2913 );
and ( n3091 , n2890 , n2913 );
or ( n3092 , n3089 , n3090 , n3091 );
and ( n3093 , n2923 , n2944 );
and ( n3094 , n2944 , n2949 );
and ( n3095 , n2923 , n2949 );
or ( n3096 , n3093 , n3094 , n3095 );
xor ( n3097 , n3092 , n3096 );
and ( n3098 , n2914 , n2918 );
and ( n3099 , n2918 , n2950 );
and ( n3100 , n2914 , n2950 );
or ( n3101 , n3098 , n3099 , n3100 );
xor ( n3102 , n3097 , n3101 );
xor ( n3103 , n3088 , n3102 );
and ( n3104 , n2886 , n2951 );
and ( n3105 , n2952 , n2955 );
or ( n3106 , n3104 , n3105 );
xor ( n3107 , n3103 , n3106 );
buf ( n3108 , n3107 );
not ( n3109 , n455 );
and ( n3110 , n3109 , n3037 );
and ( n3111 , n3108 , n455 );
or ( n3112 , n3110 , n3111 );
and ( n3113 , n2978 , n2992 );
and ( n3114 , n2992 , n3024 );
and ( n3115 , n2978 , n3024 );
or ( n3116 , n3113 , n3114 , n3115 );
and ( n3117 , n3001 , n3005 );
and ( n3118 , n3005 , n3007 );
and ( n3119 , n3001 , n3007 );
or ( n3120 , n3117 , n3118 , n3119 );
and ( n3121 , n1672 , n1264 );
and ( n3122 , n1791 , n1175 );
nor ( n3123 , n3121 , n3122 );
xnor ( n3124 , n3123 , n1270 );
and ( n3125 , n1164 , n1829 );
and ( n3126 , n1251 , n1698 );
nor ( n3127 , n3125 , n3126 );
xnor ( n3128 , n3127 , n1800 );
xor ( n3129 , n3124 , n3128 );
and ( n3130 , n965 , n2138 );
and ( n3131 , n1038 , n1981 );
nor ( n3132 , n3130 , n3131 );
xnor ( n3133 , n3132 , n2144 );
xor ( n3134 , n3129 , n3133 );
xor ( n3135 , n3120 , n3134 );
not ( n3136 , n885 );
and ( n3137 , n1970 , n1066 );
and ( n3138 , n2175 , n976 );
nor ( n3139 , n3137 , n3138 );
xnor ( n3140 , n3139 , n1047 );
xor ( n3141 , n3136 , n3140 );
and ( n3142 , n1379 , n1522 );
and ( n3143 , n1540 , n1411 );
nor ( n3144 , n3142 , n3143 );
xnor ( n3145 , n3144 , n1512 );
xor ( n3146 , n3141 , n3145 );
xor ( n3147 , n3135 , n3146 );
xor ( n3148 , n3116 , n3147 );
and ( n3149 , n2982 , n2986 );
and ( n3150 , n2986 , n2991 );
and ( n3151 , n2982 , n2991 );
or ( n3152 , n3149 , n3150 , n3151 );
and ( n3153 , n2997 , n3008 );
and ( n3154 , n3008 , n3023 );
and ( n3155 , n2997 , n3023 );
or ( n3156 , n3153 , n3154 , n3155 );
xor ( n3157 , n3152 , n3156 );
and ( n3158 , n3013 , n3017 );
and ( n3159 , n3017 , n3022 );
and ( n3160 , n3013 , n3022 );
or ( n3161 , n3158 , n3159 , n3160 );
buf ( n3162 , n2990 );
xor ( n3163 , n3161 , n3162 );
and ( n3164 , n876 , n2135 );
xor ( n3165 , n3163 , n3164 );
xor ( n3166 , n3157 , n3165 );
xor ( n3167 , n3148 , n3166 );
and ( n3168 , n2969 , n2973 );
and ( n3169 , n2973 , n3025 );
and ( n3170 , n2969 , n3025 );
or ( n3171 , n3168 , n3169 , n3170 );
xor ( n3172 , n3167 , n3171 );
and ( n3173 , n2965 , n3026 );
and ( n3174 , n3026 , n3031 );
and ( n3175 , n2965 , n3031 );
or ( n3176 , n3173 , n3174 , n3175 );
xor ( n3177 , n3172 , n3176 );
or ( n3178 , n3032 , n3033 );
xnor ( n3179 , n3177 , n3178 );
and ( n3180 , n3034 , n3035 );
xor ( n3181 , n3179 , n3180 );
buf ( n3182 , n3181 );
and ( n3183 , n3051 , n3055 );
and ( n3184 , n3055 , n3087 );
and ( n3185 , n3051 , n3087 );
or ( n3186 , n3183 , n3184 , n3185 );
and ( n3187 , n3092 , n3096 );
and ( n3188 , n3096 , n3101 );
and ( n3189 , n3092 , n3101 );
or ( n3190 , n3187 , n3188 , n3189 );
xor ( n3191 , n3186 , n3190 );
and ( n3192 , n3064 , n3068 );
and ( n3193 , n3068 , n3070 );
and ( n3194 , n3064 , n3070 );
or ( n3195 , n3192 , n3193 , n3194 );
and ( n3196 , n1009 , n2276 );
and ( n3197 , n1123 , n2089 );
nor ( n3198 , n3196 , n3197 );
xnor ( n3199 , n3198 , n2247 );
not ( n3200 , n930 );
and ( n3201 , n2083 , n1107 );
and ( n3202 , n2219 , n1015 );
nor ( n3203 , n3201 , n3202 );
xnor ( n3204 , n3203 , n1113 );
xor ( n3205 , n3200 , n3204 );
and ( n3206 , n1469 , n1588 );
and ( n3207 , n1618 , n1446 );
nor ( n3208 , n3206 , n3207 );
xnor ( n3209 , n3208 , n1594 );
xor ( n3210 , n3205 , n3209 );
xor ( n3211 , n3199 , n3210 );
and ( n3212 , n1732 , n1346 );
and ( n3213 , n1919 , n1196 );
nor ( n3214 , n3212 , n3213 );
xnor ( n3215 , n3214 , n1352 );
and ( n3216 , n1213 , n1894 );
and ( n3217 , n1323 , n1724 );
nor ( n3218 , n3216 , n3217 );
xnor ( n3219 , n3218 , n1900 );
xor ( n3220 , n3215 , n3219 );
xor ( n3221 , n3211 , n3220 );
xor ( n3222 , n3195 , n3221 );
and ( n3223 , n3041 , n3045 );
and ( n3224 , n3045 , n3050 );
and ( n3225 , n3041 , n3050 );
or ( n3226 , n3223 , n3224 , n3225 );
and ( n3227 , n3060 , n3071 );
and ( n3228 , n3071 , n3086 );
and ( n3229 , n3060 , n3086 );
or ( n3230 , n3227 , n3228 , n3229 );
xor ( n3231 , n3226 , n3230 );
and ( n3232 , n3076 , n3080 );
and ( n3233 , n3080 , n3085 );
and ( n3234 , n3076 , n3085 );
or ( n3235 , n3232 , n3233 , n3234 );
buf ( n3236 , n3049 );
xor ( n3237 , n3235 , n3236 );
and ( n3238 , n939 , n2244 );
xor ( n3239 , n3237 , n3238 );
xor ( n3240 , n3231 , n3239 );
xor ( n3241 , n3222 , n3240 );
xor ( n3242 , n3191 , n3241 );
and ( n3243 , n3088 , n3102 );
and ( n3244 , n3103 , n3106 );
or ( n3245 , n3243 , n3244 );
xor ( n3246 , n3242 , n3245 );
buf ( n3247 , n3246 );
not ( n3248 , n455 );
and ( n3249 , n3248 , n3182 );
and ( n3250 , n3247 , n455 );
or ( n3251 , n3249 , n3250 );
and ( n3252 , n3152 , n3156 );
and ( n3253 , n3156 , n3165 );
and ( n3254 , n3152 , n3165 );
or ( n3255 , n3252 , n3253 , n3254 );
and ( n3256 , n3124 , n3128 );
and ( n3257 , n3128 , n3133 );
and ( n3258 , n3124 , n3133 );
or ( n3259 , n3256 , n3257 , n3258 );
and ( n3260 , n3136 , n3140 );
and ( n3261 , n3140 , n3145 );
and ( n3262 , n3136 , n3145 );
or ( n3263 , n3260 , n3261 , n3262 );
xor ( n3264 , n3259 , n3263 );
and ( n3265 , n2175 , n1066 );
not ( n3266 , n3265 );
xnor ( n3267 , n3266 , n1047 );
and ( n3268 , n1251 , n1829 );
and ( n3269 , n1379 , n1698 );
nor ( n3270 , n3268 , n3269 );
xnor ( n3271 , n3270 , n1800 );
xor ( n3272 , n3267 , n3271 );
and ( n3273 , n1038 , n2138 );
and ( n3274 , n1164 , n1981 );
nor ( n3275 , n3273 , n3274 );
xnor ( n3276 , n3275 , n2144 );
xor ( n3277 , n3272 , n3276 );
xor ( n3278 , n3264 , n3277 );
xor ( n3279 , n3255 , n3278 );
and ( n3280 , n3161 , n3162 );
and ( n3281 , n3162 , n3164 );
and ( n3282 , n3161 , n3164 );
or ( n3283 , n3280 , n3281 , n3282 );
and ( n3284 , n3120 , n3134 );
and ( n3285 , n3134 , n3146 );
and ( n3286 , n3120 , n3146 );
or ( n3287 , n3284 , n3285 , n3286 );
xor ( n3288 , n3283 , n3287 );
and ( n3289 , n1791 , n1264 );
and ( n3290 , n1970 , n1175 );
nor ( n3291 , n3289 , n3290 );
xnor ( n3292 , n3291 , n1270 );
not ( n3293 , n3292 );
and ( n3294 , n1540 , n1522 );
and ( n3295 , n1672 , n1411 );
nor ( n3296 , n3294 , n3295 );
xnor ( n3297 , n3296 , n1512 );
xor ( n3298 , n3293 , n3297 );
and ( n3299 , n965 , n2135 );
xor ( n3300 , n3298 , n3299 );
xor ( n3301 , n3288 , n3300 );
xor ( n3302 , n3279 , n3301 );
and ( n3303 , n3116 , n3147 );
and ( n3304 , n3147 , n3166 );
and ( n3305 , n3116 , n3166 );
or ( n3306 , n3303 , n3304 , n3305 );
xor ( n3307 , n3302 , n3306 );
and ( n3308 , n3167 , n3171 );
and ( n3309 , n3171 , n3176 );
and ( n3310 , n3167 , n3176 );
or ( n3311 , n3308 , n3309 , n3310 );
xor ( n3312 , n3307 , n3311 );
or ( n3313 , n3177 , n3178 );
xnor ( n3314 , n3312 , n3313 );
and ( n3315 , n3179 , n3180 );
xor ( n3316 , n3314 , n3315 );
buf ( n3317 , n3316 );
and ( n3318 , n3186 , n3190 );
and ( n3319 , n3190 , n3241 );
and ( n3320 , n3186 , n3241 );
or ( n3321 , n3318 , n3319 , n3320 );
and ( n3322 , n3226 , n3230 );
and ( n3323 , n3230 , n3239 );
and ( n3324 , n3226 , n3239 );
or ( n3325 , n3322 , n3323 , n3324 );
and ( n3326 , n3199 , n3210 );
and ( n3327 , n3210 , n3220 );
and ( n3328 , n3199 , n3220 );
or ( n3329 , n3326 , n3327 , n3328 );
and ( n3330 , n3200 , n3204 );
and ( n3331 , n3204 , n3209 );
and ( n3332 , n3200 , n3209 );
or ( n3333 , n3330 , n3331 , n3332 );
and ( n3334 , n3215 , n3219 );
xor ( n3335 , n3333 , n3334 );
and ( n3336 , n2219 , n1107 );
not ( n3337 , n3336 );
xnor ( n3338 , n3337 , n1113 );
and ( n3339 , n1323 , n1894 );
and ( n3340 , n1469 , n1724 );
nor ( n3341 , n3339 , n3340 );
xnor ( n3342 , n3341 , n1900 );
xor ( n3343 , n3338 , n3342 );
and ( n3344 , n1123 , n2276 );
and ( n3345 , n1213 , n2089 );
nor ( n3346 , n3344 , n3345 );
xnor ( n3347 , n3346 , n2247 );
xor ( n3348 , n3343 , n3347 );
xor ( n3349 , n3335 , n3348 );
xor ( n3350 , n3329 , n3349 );
and ( n3351 , n3235 , n3236 );
and ( n3352 , n3236 , n3238 );
and ( n3353 , n3235 , n3238 );
or ( n3354 , n3351 , n3352 , n3353 );
and ( n3355 , n1919 , n1346 );
and ( n3356 , n2083 , n1196 );
nor ( n3357 , n3355 , n3356 );
xnor ( n3358 , n3357 , n1352 );
not ( n3359 , n3358 );
and ( n3360 , n1618 , n1588 );
and ( n3361 , n1732 , n1446 );
nor ( n3362 , n3360 , n3361 );
xnor ( n3363 , n3362 , n1594 );
xor ( n3364 , n3359 , n3363 );
and ( n3365 , n1009 , n2244 );
xor ( n3366 , n3364 , n3365 );
xor ( n3367 , n3354 , n3366 );
xor ( n3368 , n3350 , n3367 );
xor ( n3369 , n3325 , n3368 );
and ( n3370 , n3195 , n3221 );
and ( n3371 , n3221 , n3240 );
and ( n3372 , n3195 , n3240 );
or ( n3373 , n3370 , n3371 , n3372 );
xor ( n3374 , n3369 , n3373 );
xor ( n3375 , n3321 , n3374 );
and ( n3376 , n3242 , n3245 );
xor ( n3377 , n3375 , n3376 );
buf ( n3378 , n3377 );
not ( n3379 , n455 );
and ( n3380 , n3379 , n3317 );
and ( n3381 , n3378 , n455 );
or ( n3382 , n3380 , n3381 );
and ( n3383 , n3259 , n3263 );
and ( n3384 , n3263 , n3277 );
and ( n3385 , n3259 , n3277 );
or ( n3386 , n3383 , n3384 , n3385 );
and ( n3387 , n3283 , n3287 );
and ( n3388 , n3287 , n3300 );
and ( n3389 , n3283 , n3300 );
or ( n3390 , n3387 , n3388 , n3389 );
xor ( n3391 , n3386 , n3390 );
and ( n3392 , n3293 , n3297 );
and ( n3393 , n3297 , n3299 );
and ( n3394 , n3293 , n3299 );
or ( n3395 , n3392 , n3393 , n3394 );
not ( n3396 , n1047 );
and ( n3397 , n1970 , n1264 );
and ( n3398 , n2175 , n1175 );
nor ( n3399 , n3397 , n3398 );
xnor ( n3400 , n3399 , n1270 );
xor ( n3401 , n3396 , n3400 );
and ( n3402 , n1379 , n1829 );
and ( n3403 , n1540 , n1698 );
nor ( n3404 , n3402 , n3403 );
xnor ( n3405 , n3404 , n1800 );
xor ( n3406 , n3401 , n3405 );
xor ( n3407 , n3395 , n3406 );
and ( n3408 , n3267 , n3271 );
and ( n3409 , n3271 , n3276 );
and ( n3410 , n3267 , n3276 );
or ( n3411 , n3408 , n3409 , n3410 );
buf ( n3412 , n3292 );
xor ( n3413 , n3411 , n3412 );
and ( n3414 , n1672 , n1522 );
and ( n3415 , n1791 , n1411 );
nor ( n3416 , n3414 , n3415 );
xnor ( n3417 , n3416 , n1512 );
and ( n3418 , n1164 , n2138 );
and ( n3419 , n1251 , n1981 );
nor ( n3420 , n3418 , n3419 );
xnor ( n3421 , n3420 , n2144 );
xor ( n3422 , n3417 , n3421 );
and ( n3423 , n1038 , n2135 );
xor ( n3424 , n3422 , n3423 );
xor ( n3425 , n3413 , n3424 );
xor ( n3426 , n3407 , n3425 );
xor ( n3427 , n3391 , n3426 );
and ( n3428 , n3255 , n3278 );
and ( n3429 , n3278 , n3301 );
and ( n3430 , n3255 , n3301 );
or ( n3431 , n3428 , n3429 , n3430 );
xor ( n3432 , n3427 , n3431 );
and ( n3433 , n3302 , n3306 );
and ( n3434 , n3306 , n3311 );
and ( n3435 , n3302 , n3311 );
or ( n3436 , n3433 , n3434 , n3435 );
xor ( n3437 , n3432 , n3436 );
or ( n3438 , n3312 , n3313 );
xnor ( n3439 , n3437 , n3438 );
and ( n3440 , n3314 , n3315 );
xor ( n3441 , n3439 , n3440 );
buf ( n3442 , n3441 );
and ( n3443 , n3359 , n3363 );
and ( n3444 , n3363 , n3365 );
and ( n3445 , n3359 , n3365 );
or ( n3446 , n3443 , n3444 , n3445 );
not ( n3447 , n1113 );
and ( n3448 , n2083 , n1346 );
and ( n3449 , n2219 , n1196 );
nor ( n3450 , n3448 , n3449 );
xnor ( n3451 , n3450 , n1352 );
xor ( n3452 , n3447 , n3451 );
and ( n3453 , n1469 , n1894 );
and ( n3454 , n1618 , n1724 );
nor ( n3455 , n3453 , n3454 );
xnor ( n3456 , n3455 , n1900 );
xor ( n3457 , n3452 , n3456 );
xor ( n3458 , n3446 , n3457 );
and ( n3459 , n3333 , n3334 );
and ( n3460 , n3334 , n3348 );
and ( n3461 , n3333 , n3348 );
or ( n3462 , n3459 , n3460 , n3461 );
xor ( n3463 , n3458 , n3462 );
and ( n3464 , n1732 , n1588 );
and ( n3465 , n1919 , n1446 );
nor ( n3466 , n3464 , n3465 );
xnor ( n3467 , n3466 , n1594 );
and ( n3468 , n1213 , n2276 );
and ( n3469 , n1323 , n2089 );
nor ( n3470 , n3468 , n3469 );
xnor ( n3471 , n3470 , n2247 );
xor ( n3472 , n3467 , n3471 );
and ( n3473 , n1123 , n2244 );
xor ( n3474 , n3472 , n3473 );
buf ( n3475 , n3358 );
xor ( n3476 , n3474 , n3475 );
and ( n3477 , n3338 , n3342 );
and ( n3478 , n3342 , n3347 );
and ( n3479 , n3338 , n3347 );
or ( n3480 , n3477 , n3478 , n3479 );
xor ( n3481 , n3476 , n3480 );
xor ( n3482 , n3463 , n3481 );
and ( n3483 , n3354 , n3366 );
xor ( n3484 , n3482 , n3483 );
and ( n3485 , n3329 , n3349 );
and ( n3486 , n3349 , n3367 );
and ( n3487 , n3329 , n3367 );
or ( n3488 , n3485 , n3486 , n3487 );
xor ( n3489 , n3484 , n3488 );
and ( n3490 , n3325 , n3368 );
and ( n3491 , n3368 , n3373 );
and ( n3492 , n3325 , n3373 );
or ( n3493 , n3490 , n3491 , n3492 );
xor ( n3494 , n3489 , n3493 );
and ( n3495 , n3321 , n3374 );
and ( n3496 , n3375 , n3376 );
or ( n3497 , n3495 , n3496 );
xor ( n3498 , n3494 , n3497 );
buf ( n3499 , n3498 );
not ( n3500 , n455 );
and ( n3501 , n3500 , n3442 );
and ( n3502 , n3499 , n455 );
or ( n3503 , n3501 , n3502 );
and ( n3504 , n3411 , n3412 );
and ( n3505 , n3412 , n3424 );
and ( n3506 , n3411 , n3424 );
or ( n3507 , n3504 , n3505 , n3506 );
and ( n3508 , n3395 , n3406 );
and ( n3509 , n3406 , n3425 );
and ( n3510 , n3395 , n3425 );
or ( n3511 , n3508 , n3509 , n3510 );
xor ( n3512 , n3507 , n3511 );
and ( n3513 , n3396 , n3400 );
and ( n3514 , n3400 , n3405 );
and ( n3515 , n3396 , n3405 );
or ( n3516 , n3513 , n3514 , n3515 );
and ( n3517 , n2175 , n1264 );
not ( n3518 , n3517 );
xnor ( n3519 , n3518 , n1270 );
and ( n3520 , n1251 , n2138 );
and ( n3521 , n1379 , n1981 );
nor ( n3522 , n3520 , n3521 );
xnor ( n3523 , n3522 , n2144 );
xor ( n3524 , n3519 , n3523 );
and ( n3525 , n1164 , n2135 );
xor ( n3526 , n3524 , n3525 );
xor ( n3527 , n3516 , n3526 );
and ( n3528 , n3417 , n3421 );
and ( n3529 , n3421 , n3423 );
and ( n3530 , n3417 , n3423 );
or ( n3531 , n3528 , n3529 , n3530 );
and ( n3532 , n1791 , n1522 );
and ( n3533 , n1970 , n1411 );
nor ( n3534 , n3532 , n3533 );
xnor ( n3535 , n3534 , n1512 );
not ( n3536 , n3535 );
xor ( n3537 , n3531 , n3536 );
and ( n3538 , n1540 , n1829 );
and ( n3539 , n1672 , n1698 );
nor ( n3540 , n3538 , n3539 );
xnor ( n3541 , n3540 , n1800 );
xor ( n3542 , n3537 , n3541 );
xor ( n3543 , n3527 , n3542 );
xor ( n3544 , n3512 , n3543 );
and ( n3545 , n3386 , n3390 );
and ( n3546 , n3390 , n3426 );
and ( n3547 , n3386 , n3426 );
or ( n3548 , n3545 , n3546 , n3547 );
xor ( n3549 , n3544 , n3548 );
and ( n3550 , n3427 , n3431 );
and ( n3551 , n3431 , n3436 );
and ( n3552 , n3427 , n3436 );
or ( n3553 , n3550 , n3551 , n3552 );
xor ( n3554 , n3549 , n3553 );
or ( n3555 , n3437 , n3438 );
xnor ( n3556 , n3554 , n3555 );
and ( n3557 , n3439 , n3440 );
xor ( n3558 , n3556 , n3557 );
buf ( n3559 , n3558 );
and ( n3560 , n3458 , n3462 );
and ( n3561 , n3462 , n3481 );
and ( n3562 , n3458 , n3481 );
or ( n3563 , n3560 , n3561 , n3562 );
and ( n3564 , n3446 , n3457 );
and ( n3565 , n3474 , n3475 );
and ( n3566 , n3475 , n3480 );
and ( n3567 , n3474 , n3480 );
or ( n3568 , n3565 , n3566 , n3567 );
xor ( n3569 , n3564 , n3568 );
and ( n3570 , n3447 , n3451 );
and ( n3571 , n3451 , n3456 );
and ( n3572 , n3447 , n3456 );
or ( n3573 , n3570 , n3571 , n3572 );
and ( n3574 , n2219 , n1346 );
not ( n3575 , n3574 );
xnor ( n3576 , n3575 , n1352 );
and ( n3577 , n1323 , n2276 );
and ( n3578 , n1469 , n2089 );
nor ( n3579 , n3577 , n3578 );
xnor ( n3580 , n3579 , n2247 );
xor ( n3581 , n3576 , n3580 );
and ( n3582 , n1213 , n2244 );
xor ( n3583 , n3581 , n3582 );
xor ( n3584 , n3573 , n3583 );
and ( n3585 , n3467 , n3471 );
and ( n3586 , n3471 , n3473 );
and ( n3587 , n3467 , n3473 );
or ( n3588 , n3585 , n3586 , n3587 );
and ( n3589 , n1919 , n1588 );
and ( n3590 , n2083 , n1446 );
nor ( n3591 , n3589 , n3590 );
xnor ( n3592 , n3591 , n1594 );
not ( n3593 , n3592 );
xor ( n3594 , n3588 , n3593 );
and ( n3595 , n1618 , n1894 );
and ( n3596 , n1732 , n1724 );
nor ( n3597 , n3595 , n3596 );
xnor ( n3598 , n3597 , n1900 );
xor ( n3599 , n3594 , n3598 );
xor ( n3600 , n3584 , n3599 );
xor ( n3601 , n3569 , n3600 );
xor ( n3602 , n3563 , n3601 );
and ( n3603 , n3482 , n3483 );
and ( n3604 , n3483 , n3488 );
and ( n3605 , n3482 , n3488 );
or ( n3606 , n3603 , n3604 , n3605 );
xor ( n3607 , n3602 , n3606 );
and ( n3608 , n3489 , n3493 );
and ( n3609 , n3494 , n3497 );
or ( n3610 , n3608 , n3609 );
xor ( n3611 , n3607 , n3610 );
buf ( n3612 , n3611 );
not ( n3613 , n455 );
and ( n3614 , n3613 , n3559 );
and ( n3615 , n3612 , n455 );
or ( n3616 , n3614 , n3615 );
and ( n3617 , n3507 , n3511 );
and ( n3618 , n3511 , n3543 );
and ( n3619 , n3507 , n3543 );
or ( n3620 , n3617 , n3618 , n3619 );
and ( n3621 , n3531 , n3536 );
and ( n3622 , n3536 , n3541 );
and ( n3623 , n3531 , n3541 );
or ( n3624 , n3621 , n3622 , n3623 );
and ( n3625 , n3516 , n3526 );
and ( n3626 , n3526 , n3542 );
and ( n3627 , n3516 , n3542 );
or ( n3628 , n3625 , n3626 , n3627 );
xor ( n3629 , n3624 , n3628 );
and ( n3630 , n3519 , n3523 );
and ( n3631 , n3523 , n3525 );
and ( n3632 , n3519 , n3525 );
or ( n3633 , n3630 , n3631 , n3632 );
not ( n3634 , n1270 );
and ( n3635 , n1970 , n1522 );
and ( n3636 , n2175 , n1411 );
nor ( n3637 , n3635 , n3636 );
xnor ( n3638 , n3637 , n1512 );
xor ( n3639 , n3634 , n3638 );
and ( n3640 , n1379 , n2138 );
and ( n3641 , n1540 , n1981 );
nor ( n3642 , n3640 , n3641 );
xnor ( n3643 , n3642 , n2144 );
xor ( n3644 , n3639 , n3643 );
xor ( n3645 , n3633 , n3644 );
buf ( n3646 , n3535 );
and ( n3647 , n1672 , n1829 );
and ( n3648 , n1791 , n1698 );
nor ( n3649 , n3647 , n3648 );
xnor ( n3650 , n3649 , n1800 );
xor ( n3651 , n3646 , n3650 );
and ( n3652 , n1251 , n2135 );
xor ( n3653 , n3651 , n3652 );
xor ( n3654 , n3645 , n3653 );
xor ( n3655 , n3629 , n3654 );
xor ( n3656 , n3620 , n3655 );
and ( n3657 , n3544 , n3548 );
and ( n3658 , n3548 , n3553 );
and ( n3659 , n3544 , n3553 );
or ( n3660 , n3657 , n3658 , n3659 );
xor ( n3661 , n3656 , n3660 );
or ( n3662 , n3554 , n3555 );
xnor ( n3663 , n3661 , n3662 );
and ( n3664 , n3556 , n3557 );
xor ( n3665 , n3663 , n3664 );
buf ( n3666 , n3665 );
and ( n3667 , n3564 , n3568 );
and ( n3668 , n3568 , n3600 );
and ( n3669 , n3564 , n3600 );
or ( n3670 , n3667 , n3668 , n3669 );
and ( n3671 , n3588 , n3593 );
and ( n3672 , n3593 , n3598 );
and ( n3673 , n3588 , n3598 );
or ( n3674 , n3671 , n3672 , n3673 );
and ( n3675 , n3573 , n3583 );
and ( n3676 , n3583 , n3599 );
and ( n3677 , n3573 , n3599 );
or ( n3678 , n3675 , n3676 , n3677 );
xor ( n3679 , n3674 , n3678 );
and ( n3680 , n3576 , n3580 );
and ( n3681 , n3580 , n3582 );
and ( n3682 , n3576 , n3582 );
or ( n3683 , n3680 , n3681 , n3682 );
not ( n3684 , n1352 );
and ( n3685 , n2083 , n1588 );
and ( n3686 , n2219 , n1446 );
nor ( n3687 , n3685 , n3686 );
xnor ( n3688 , n3687 , n1594 );
xor ( n3689 , n3684 , n3688 );
and ( n3690 , n1469 , n2276 );
and ( n3691 , n1618 , n2089 );
nor ( n3692 , n3690 , n3691 );
xnor ( n3693 , n3692 , n2247 );
xor ( n3694 , n3689 , n3693 );
xor ( n3695 , n3683 , n3694 );
buf ( n3696 , n3592 );
and ( n3697 , n1732 , n1894 );
and ( n3698 , n1919 , n1724 );
nor ( n3699 , n3697 , n3698 );
xnor ( n3700 , n3699 , n1900 );
xor ( n3701 , n3696 , n3700 );
and ( n3702 , n1323 , n2244 );
xor ( n3703 , n3701 , n3702 );
xor ( n3704 , n3695 , n3703 );
xor ( n3705 , n3679 , n3704 );
xor ( n3706 , n3670 , n3705 );
and ( n3707 , n3563 , n3601 );
and ( n3708 , n3601 , n3606 );
and ( n3709 , n3563 , n3606 );
or ( n3710 , n3707 , n3708 , n3709 );
xor ( n3711 , n3706 , n3710 );
and ( n3712 , n3607 , n3610 );
xor ( n3713 , n3711 , n3712 );
buf ( n3714 , n3713 );
not ( n3715 , n455 );
and ( n3716 , n3715 , n3666 );
and ( n3717 , n3714 , n455 );
or ( n3718 , n3716 , n3717 );
and ( n3719 , n3646 , n3650 );
and ( n3720 , n3650 , n3652 );
and ( n3721 , n3646 , n3652 );
or ( n3722 , n3719 , n3720 , n3721 );
and ( n3723 , n3633 , n3644 );
and ( n3724 , n3644 , n3653 );
and ( n3725 , n3633 , n3653 );
or ( n3726 , n3723 , n3724 , n3725 );
xor ( n3727 , n3722 , n3726 );
and ( n3728 , n3634 , n3638 );
and ( n3729 , n3638 , n3643 );
and ( n3730 , n3634 , n3643 );
or ( n3731 , n3728 , n3729 , n3730 );
and ( n3732 , n2175 , n1522 );
not ( n3733 , n3732 );
xnor ( n3734 , n3733 , n1512 );
not ( n3735 , n3734 );
xor ( n3736 , n3731 , n3735 );
and ( n3737 , n1791 , n1829 );
and ( n3738 , n1970 , n1698 );
nor ( n3739 , n3737 , n3738 );
xnor ( n3740 , n3739 , n1800 );
and ( n3741 , n1540 , n2138 );
and ( n3742 , n1672 , n1981 );
nor ( n3743 , n3741 , n3742 );
xnor ( n3744 , n3743 , n2144 );
xor ( n3745 , n3740 , n3744 );
and ( n3746 , n1379 , n2135 );
xor ( n3747 , n3745 , n3746 );
xor ( n3748 , n3736 , n3747 );
xor ( n3749 , n3727 , n3748 );
and ( n3750 , n3624 , n3628 );
and ( n3751 , n3628 , n3654 );
and ( n3752 , n3624 , n3654 );
or ( n3753 , n3750 , n3751 , n3752 );
xor ( n3754 , n3749 , n3753 );
and ( n3755 , n3620 , n3655 );
and ( n3756 , n3655 , n3660 );
and ( n3757 , n3620 , n3660 );
or ( n3758 , n3755 , n3756 , n3757 );
xor ( n3759 , n3754 , n3758 );
or ( n3760 , n3661 , n3662 );
xnor ( n3761 , n3759 , n3760 );
and ( n3762 , n3663 , n3664 );
xor ( n3763 , n3761 , n3762 );
buf ( n3764 , n3763 );
and ( n3765 , n3696 , n3700 );
and ( n3766 , n3700 , n3702 );
and ( n3767 , n3696 , n3702 );
or ( n3768 , n3765 , n3766 , n3767 );
and ( n3769 , n3683 , n3694 );
and ( n3770 , n3694 , n3703 );
and ( n3771 , n3683 , n3703 );
or ( n3772 , n3769 , n3770 , n3771 );
xor ( n3773 , n3768 , n3772 );
and ( n3774 , n3684 , n3688 );
and ( n3775 , n3688 , n3693 );
and ( n3776 , n3684 , n3693 );
or ( n3777 , n3774 , n3775 , n3776 );
and ( n3778 , n2219 , n1588 );
not ( n3779 , n3778 );
xnor ( n3780 , n3779 , n1594 );
not ( n3781 , n3780 );
xor ( n3782 , n3777 , n3781 );
and ( n3783 , n1919 , n1894 );
and ( n3784 , n2083 , n1724 );
nor ( n3785 , n3783 , n3784 );
xnor ( n3786 , n3785 , n1900 );
and ( n3787 , n1618 , n2276 );
and ( n3788 , n1732 , n2089 );
nor ( n3789 , n3787 , n3788 );
xnor ( n3790 , n3789 , n2247 );
xor ( n3791 , n3786 , n3790 );
and ( n3792 , n1469 , n2244 );
xor ( n3793 , n3791 , n3792 );
xor ( n3794 , n3782 , n3793 );
xor ( n3795 , n3773 , n3794 );
and ( n3796 , n3674 , n3678 );
and ( n3797 , n3678 , n3704 );
and ( n3798 , n3674 , n3704 );
or ( n3799 , n3796 , n3797 , n3798 );
xor ( n3800 , n3795 , n3799 );
and ( n3801 , n3670 , n3705 );
and ( n3802 , n3705 , n3710 );
and ( n3803 , n3670 , n3710 );
or ( n3804 , n3801 , n3802 , n3803 );
xor ( n3805 , n3800 , n3804 );
and ( n3806 , n3711 , n3712 );
xor ( n3807 , n3805 , n3806 );
buf ( n3808 , n3807 );
not ( n3809 , n455 );
and ( n3810 , n3809 , n3764 );
and ( n3811 , n3808 , n455 );
or ( n3812 , n3810 , n3811 );
and ( n3813 , n3731 , n3735 );
and ( n3814 , n3735 , n3747 );
and ( n3815 , n3731 , n3747 );
or ( n3816 , n3813 , n3814 , n3815 );
not ( n3817 , n1512 );
and ( n3818 , n1970 , n1829 );
and ( n3819 , n2175 , n1698 );
nor ( n3820 , n3818 , n3819 );
xnor ( n3821 , n3820 , n1800 );
xor ( n3822 , n3817 , n3821 );
and ( n3823 , n1540 , n2135 );
xor ( n3824 , n3822 , n3823 );
xor ( n3825 , n3816 , n3824 );
and ( n3826 , n3740 , n3744 );
and ( n3827 , n3744 , n3746 );
and ( n3828 , n3740 , n3746 );
or ( n3829 , n3826 , n3827 , n3828 );
buf ( n3830 , n3734 );
xor ( n3831 , n3829 , n3830 );
and ( n3832 , n1672 , n2138 );
and ( n3833 , n1791 , n1981 );
nor ( n3834 , n3832 , n3833 );
xnor ( n3835 , n3834 , n2144 );
xor ( n3836 , n3831 , n3835 );
xor ( n3837 , n3825 , n3836 );
and ( n3838 , n3722 , n3726 );
and ( n3839 , n3726 , n3748 );
and ( n3840 , n3722 , n3748 );
or ( n3841 , n3838 , n3839 , n3840 );
xor ( n3842 , n3837 , n3841 );
and ( n3843 , n3749 , n3753 );
and ( n3844 , n3753 , n3758 );
and ( n3845 , n3749 , n3758 );
or ( n3846 , n3843 , n3844 , n3845 );
xor ( n3847 , n3842 , n3846 );
or ( n3848 , n3759 , n3760 );
xnor ( n3849 , n3847 , n3848 );
and ( n3850 , n3761 , n3762 );
xor ( n3851 , n3849 , n3850 );
buf ( n3852 , n3851 );
and ( n3853 , n3777 , n3781 );
and ( n3854 , n3781 , n3793 );
and ( n3855 , n3777 , n3793 );
or ( n3856 , n3853 , n3854 , n3855 );
not ( n3857 , n1594 );
and ( n3858 , n2083 , n1894 );
and ( n3859 , n2219 , n1724 );
nor ( n3860 , n3858 , n3859 );
xnor ( n3861 , n3860 , n1900 );
xor ( n3862 , n3857 , n3861 );
and ( n3863 , n1618 , n2244 );
xor ( n3864 , n3862 , n3863 );
xor ( n3865 , n3856 , n3864 );
and ( n3866 , n3786 , n3790 );
and ( n3867 , n3790 , n3792 );
and ( n3868 , n3786 , n3792 );
or ( n3869 , n3866 , n3867 , n3868 );
buf ( n3870 , n3780 );
xor ( n3871 , n3869 , n3870 );
and ( n3872 , n1732 , n2276 );
and ( n3873 , n1919 , n2089 );
nor ( n3874 , n3872 , n3873 );
xnor ( n3875 , n3874 , n2247 );
xor ( n3876 , n3871 , n3875 );
xor ( n3877 , n3865 , n3876 );
and ( n3878 , n3768 , n3772 );
and ( n3879 , n3772 , n3794 );
and ( n3880 , n3768 , n3794 );
or ( n3881 , n3878 , n3879 , n3880 );
xor ( n3882 , n3877 , n3881 );
and ( n3883 , n3795 , n3799 );
and ( n3884 , n3799 , n3804 );
and ( n3885 , n3795 , n3804 );
or ( n3886 , n3883 , n3884 , n3885 );
xor ( n3887 , n3882 , n3886 );
and ( n3888 , n3805 , n3806 );
xor ( n3889 , n3887 , n3888 );
buf ( n3890 , n3889 );
not ( n3891 , n455 );
and ( n3892 , n3891 , n3852 );
and ( n3893 , n3890 , n455 );
or ( n3894 , n3892 , n3893 );
and ( n3895 , n3817 , n3821 );
and ( n3896 , n3821 , n3823 );
and ( n3897 , n3817 , n3823 );
or ( n3898 , n3895 , n3896 , n3897 );
and ( n3899 , n3829 , n3830 );
and ( n3900 , n3830 , n3835 );
and ( n3901 , n3829 , n3835 );
or ( n3902 , n3899 , n3900 , n3901 );
xor ( n3903 , n3898 , n3902 );
and ( n3904 , n2175 , n1829 );
not ( n3905 , n3904 );
xnor ( n3906 , n3905 , n1800 );
not ( n3907 , n3906 );
and ( n3908 , n1791 , n2138 );
and ( n3909 , n1970 , n1981 );
nor ( n3910 , n3908 , n3909 );
xnor ( n3911 , n3910 , n2144 );
xor ( n3912 , n3907 , n3911 );
and ( n3913 , n1672 , n2135 );
xor ( n3914 , n3912 , n3913 );
xor ( n3915 , n3903 , n3914 );
and ( n3916 , n3816 , n3824 );
and ( n3917 , n3824 , n3836 );
and ( n3918 , n3816 , n3836 );
or ( n3919 , n3916 , n3917 , n3918 );
xor ( n3920 , n3915 , n3919 );
and ( n3921 , n3837 , n3841 );
and ( n3922 , n3841 , n3846 );
and ( n3923 , n3837 , n3846 );
or ( n3924 , n3921 , n3922 , n3923 );
xor ( n3925 , n3920 , n3924 );
or ( n3926 , n3847 , n3848 );
xnor ( n3927 , n3925 , n3926 );
and ( n3928 , n3849 , n3850 );
xor ( n3929 , n3927 , n3928 );
buf ( n3930 , n3929 );
and ( n3931 , n3857 , n3861 );
and ( n3932 , n3861 , n3863 );
and ( n3933 , n3857 , n3863 );
or ( n3934 , n3931 , n3932 , n3933 );
and ( n3935 , n3869 , n3870 );
and ( n3936 , n3870 , n3875 );
and ( n3937 , n3869 , n3875 );
or ( n3938 , n3935 , n3936 , n3937 );
xor ( n3939 , n3934 , n3938 );
and ( n3940 , n2219 , n1894 );
not ( n3941 , n3940 );
xnor ( n3942 , n3941 , n1900 );
not ( n3943 , n3942 );
and ( n3944 , n1919 , n2276 );
and ( n3945 , n2083 , n2089 );
nor ( n3946 , n3944 , n3945 );
xnor ( n3947 , n3946 , n2247 );
xor ( n3948 , n3943 , n3947 );
and ( n3949 , n1732 , n2244 );
xor ( n3950 , n3948 , n3949 );
xor ( n3951 , n3939 , n3950 );
and ( n3952 , n3856 , n3864 );
and ( n3953 , n3864 , n3876 );
and ( n3954 , n3856 , n3876 );
or ( n3955 , n3952 , n3953 , n3954 );
xor ( n3956 , n3951 , n3955 );
and ( n3957 , n3877 , n3881 );
and ( n3958 , n3881 , n3886 );
and ( n3959 , n3877 , n3886 );
or ( n3960 , n3957 , n3958 , n3959 );
xor ( n3961 , n3956 , n3960 );
and ( n3962 , n3887 , n3888 );
xor ( n3963 , n3961 , n3962 );
buf ( n3964 , n3963 );
not ( n3965 , n455 );
and ( n3966 , n3965 , n3930 );
and ( n3967 , n3964 , n455 );
or ( n3968 , n3966 , n3967 );
and ( n3969 , n3907 , n3911 );
and ( n3970 , n3911 , n3913 );
and ( n3971 , n3907 , n3913 );
or ( n3972 , n3969 , n3970 , n3971 );
buf ( n3973 , n3906 );
xor ( n3974 , n3972 , n3973 );
not ( n3975 , n1800 );
and ( n3976 , n1970 , n2138 );
and ( n3977 , n2175 , n1981 );
nor ( n3978 , n3976 , n3977 );
xnor ( n3979 , n3978 , n2144 );
xor ( n3980 , n3975 , n3979 );
and ( n3981 , n1791 , n2135 );
xor ( n3982 , n3980 , n3981 );
xor ( n3983 , n3974 , n3982 );
and ( n3984 , n3898 , n3902 );
and ( n3985 , n3902 , n3914 );
and ( n3986 , n3898 , n3914 );
or ( n3987 , n3984 , n3985 , n3986 );
xor ( n3988 , n3983 , n3987 );
and ( n3989 , n3915 , n3919 );
and ( n3990 , n3919 , n3924 );
and ( n3991 , n3915 , n3924 );
or ( n3992 , n3989 , n3990 , n3991 );
xor ( n3993 , n3988 , n3992 );
or ( n3994 , n3925 , n3926 );
xnor ( n3995 , n3993 , n3994 );
and ( n3996 , n3927 , n3928 );
xor ( n3997 , n3995 , n3996 );
buf ( n3998 , n3997 );
and ( n3999 , n3943 , n3947 );
and ( n4000 , n3947 , n3949 );
and ( n4001 , n3943 , n3949 );
or ( n4002 , n3999 , n4000 , n4001 );
buf ( n4003 , n3942 );
xor ( n4004 , n4002 , n4003 );
not ( n4005 , n1900 );
and ( n4006 , n2083 , n2276 );
and ( n4007 , n2219 , n2089 );
nor ( n4008 , n4006 , n4007 );
xnor ( n4009 , n4008 , n2247 );
xor ( n4010 , n4005 , n4009 );
and ( n4011 , n1919 , n2244 );
xor ( n4012 , n4010 , n4011 );
xor ( n4013 , n4004 , n4012 );
and ( n4014 , n3934 , n3938 );
and ( n4015 , n3938 , n3950 );
and ( n4016 , n3934 , n3950 );
or ( n4017 , n4014 , n4015 , n4016 );
xor ( n4018 , n4013 , n4017 );
and ( n4019 , n3951 , n3955 );
and ( n4020 , n3955 , n3960 );
and ( n4021 , n3951 , n3960 );
or ( n4022 , n4019 , n4020 , n4021 );
xor ( n4023 , n4018 , n4022 );
and ( n4024 , n3961 , n3962 );
xor ( n4025 , n4023 , n4024 );
buf ( n4026 , n4025 );
not ( n4027 , n455 );
and ( n4028 , n4027 , n3998 );
and ( n4029 , n4026 , n455 );
or ( n4030 , n4028 , n4029 );
and ( n4031 , n3975 , n3979 );
and ( n4032 , n3979 , n3981 );
and ( n4033 , n3975 , n3981 );
or ( n4034 , n4031 , n4032 , n4033 );
and ( n4035 , n2175 , n2138 );
not ( n4036 , n4035 );
xnor ( n4037 , n4036 , n2144 );
xor ( n4038 , n4034 , n4037 );
and ( n4039 , n1970 , n2135 );
not ( n4040 , n4039 );
xor ( n4041 , n4038 , n4040 );
and ( n4042 , n3972 , n3973 );
and ( n4043 , n3973 , n3982 );
and ( n4044 , n3972 , n3982 );
or ( n4045 , n4042 , n4043 , n4044 );
xor ( n4046 , n4041 , n4045 );
and ( n4047 , n3983 , n3987 );
and ( n4048 , n3987 , n3992 );
and ( n4049 , n3983 , n3992 );
or ( n4050 , n4047 , n4048 , n4049 );
xor ( n4051 , n4046 , n4050 );
or ( n4052 , n3993 , n3994 );
xnor ( n4053 , n4051 , n4052 );
and ( n4054 , n3995 , n3996 );
xor ( n4055 , n4053 , n4054 );
buf ( n4056 , n4055 );
and ( n4057 , n4005 , n4009 );
and ( n4058 , n4009 , n4011 );
and ( n4059 , n4005 , n4011 );
or ( n4060 , n4057 , n4058 , n4059 );
and ( n4061 , n2219 , n2276 );
not ( n4062 , n4061 );
xnor ( n4063 , n4062 , n2247 );
xor ( n4064 , n4060 , n4063 );
and ( n4065 , n2083 , n2244 );
not ( n4066 , n4065 );
xor ( n4067 , n4064 , n4066 );
and ( n4068 , n4002 , n4003 );
and ( n4069 , n4003 , n4012 );
and ( n4070 , n4002 , n4012 );
or ( n4071 , n4068 , n4069 , n4070 );
xor ( n4072 , n4067 , n4071 );
and ( n4073 , n4013 , n4017 );
and ( n4074 , n4017 , n4022 );
and ( n4075 , n4013 , n4022 );
or ( n4076 , n4073 , n4074 , n4075 );
xor ( n4077 , n4072 , n4076 );
and ( n4078 , n4023 , n4024 );
xor ( n4079 , n4077 , n4078 );
buf ( n4080 , n4079 );
not ( n4081 , n455 );
and ( n4082 , n4081 , n4056 );
and ( n4083 , n4080 , n455 );
or ( n4084 , n4082 , n4083 );
and ( n4085 , n4034 , n4037 );
and ( n4086 , n4037 , n4040 );
and ( n4087 , n4034 , n4040 );
or ( n4088 , n4085 , n4086 , n4087 );
buf ( n4089 , n4039 );
not ( n4090 , n2144 );
xor ( n4091 , n4089 , n4090 );
and ( n4092 , n2175 , n2135 );
xor ( n4093 , n4091 , n4092 );
xor ( n4094 , n4088 , n4093 );
and ( n4095 , n4041 , n4045 );
and ( n4096 , n4045 , n4050 );
and ( n4097 , n4041 , n4050 );
or ( n4098 , n4095 , n4096 , n4097 );
xor ( n4099 , n4094 , n4098 );
or ( n4100 , n4051 , n4052 );
xnor ( n4101 , n4099 , n4100 );
and ( n4102 , n4053 , n4054 );
xor ( n4103 , n4101 , n4102 );
buf ( n4104 , n4103 );
and ( n4105 , n4060 , n4063 );
and ( n4106 , n4063 , n4066 );
and ( n4107 , n4060 , n4066 );
or ( n4108 , n4105 , n4106 , n4107 );
buf ( n4109 , n4065 );
not ( n4110 , n2247 );
xor ( n4111 , n4109 , n4110 );
and ( n4112 , n2219 , n2244 );
xor ( n4113 , n4111 , n4112 );
xor ( n4114 , n4108 , n4113 );
and ( n4115 , n4067 , n4071 );
and ( n4116 , n4071 , n4076 );
and ( n4117 , n4067 , n4076 );
or ( n4118 , n4115 , n4116 , n4117 );
xor ( n4119 , n4114 , n4118 );
and ( n4120 , n4077 , n4078 );
xor ( n4121 , n4119 , n4120 );
buf ( n4122 , n4121 );
not ( n4123 , n455 );
and ( n4124 , n4123 , n4104 );
and ( n4125 , n4122 , n455 );
or ( n4126 , n4124 , n4125 );
buf ( n4127 , n504 );
buf ( n4128 , n520 );
xor ( n4129 , n4127 , n4128 );
buf ( n4130 , n4129 );
buf ( n4131 , n4130 );
buf ( n4132 , n4131 );
buf ( n4133 , n770 );
buf ( n4134 , n4133 );
and ( n4135 , n4132 , n4134 );
buf ( n4136 , n4135 );
buf ( n4137 , n4136 );
buf ( n4138 , n4137 );
buf ( n4139 , n4138 );
buf ( n4140 , n536 );
buf ( n4141 , n552 );
xor ( n4142 , n4140 , n4141 );
buf ( n4143 , n4142 );
buf ( n4144 , n4143 );
buf ( n4145 , n4144 );
and ( n4146 , n4139 , n4145 );
buf ( n4147 , n4146 );
buf ( n4148 , n4147 );
buf ( n4149 , n533 );
buf ( n4150 , n4149 );
buf ( n4151 , n471 );
buf ( n4152 , n4151 );
buf ( n4153 , n472 );
buf ( n4154 , n4153 );
xor ( n4155 , n4152 , n4154 );
not ( n4156 , n4154 );
and ( n4157 , n4155 , n4156 );
and ( n4158 , n4150 , n4157 );
buf ( n4159 , n532 );
buf ( n4160 , n4159 );
and ( n4161 , n4160 , n4154 );
nor ( n4162 , n4158 , n4161 );
xnor ( n4163 , n4162 , n4152 );
buf ( n4164 , n535 );
buf ( n4165 , n4164 );
buf ( n4166 , n469 );
buf ( n4167 , n4166 );
buf ( n4168 , n470 );
buf ( n4169 , n4168 );
xor ( n4170 , n4167 , n4169 );
xor ( n4171 , n4169 , n4152 );
not ( n4172 , n4171 );
and ( n4173 , n4170 , n4172 );
and ( n4174 , n4165 , n4173 );
buf ( n4175 , n534 );
buf ( n4176 , n4175 );
and ( n4177 , n4176 , n4171 );
nor ( n4178 , n4174 , n4177 );
and ( n4179 , n4169 , n4152 );
not ( n4180 , n4179 );
and ( n4181 , n4167 , n4180 );
xnor ( n4182 , n4178 , n4181 );
xor ( n4183 , n4163 , n4182 );
buf ( n4184 , n536 );
buf ( n4185 , n4184 );
buf ( n4186 , n468 );
buf ( n4187 , n4186 );
xor ( n4188 , n4187 , n4167 );
and ( n4189 , n4185 , n4188 );
xor ( n4190 , n4183 , n4189 );
and ( n4191 , n4176 , n4157 );
and ( n4192 , n4150 , n4154 );
nor ( n4193 , n4191 , n4192 );
xnor ( n4194 , n4193 , n4152 );
and ( n4195 , n4185 , n4171 );
not ( n4196 , n4195 );
and ( n4197 , n4196 , n4181 );
and ( n4198 , n4194 , n4197 );
xor ( n4199 , n4190 , n4198 );
and ( n4200 , n4185 , n4173 );
and ( n4201 , n4165 , n4171 );
nor ( n4202 , n4200 , n4201 );
xnor ( n4203 , n4202 , n4181 );
xor ( n4204 , n4194 , n4197 );
and ( n4205 , n4203 , n4204 );
xor ( n4206 , n4203 , n4204 );
and ( n4207 , n4165 , n4157 );
and ( n4208 , n4176 , n4154 );
nor ( n4209 , n4207 , n4208 );
xnor ( n4210 , n4209 , n4152 );
and ( n4211 , n4210 , n4195 );
xor ( n4212 , n4210 , n4195 );
and ( n4213 , n4185 , n4157 );
and ( n4214 , n4165 , n4154 );
nor ( n4215 , n4213 , n4214 );
xnor ( n4216 , n4215 , n4152 );
and ( n4217 , n4185 , n4154 );
not ( n4218 , n4217 );
and ( n4219 , n4218 , n4152 );
and ( n4220 , n4216 , n4219 );
and ( n4221 , n4212 , n4220 );
or ( n4222 , n4211 , n4221 );
and ( n4223 , n4206 , n4222 );
or ( n4224 , n4205 , n4223 );
xor ( n4225 , n4199 , n4224 );
buf ( n4226 , n4225 );
buf ( n4227 , n4226 );
buf ( n4228 , n4227 );
buf ( n4229 , n503 );
buf ( n4230 , n4229 );
buf ( n4231 , n504 );
buf ( n4232 , n4231 );
xor ( n4233 , n4230 , n4232 );
not ( n4234 , n4232 );
and ( n4235 , n4233 , n4234 );
and ( n4236 , n4228 , n4235 );
and ( n4237 , n4163 , n4182 );
and ( n4238 , n4182 , n4189 );
and ( n4239 , n4163 , n4189 );
or ( n4240 , n4237 , n4238 , n4239 );
and ( n4241 , n4160 , n4157 );
buf ( n4242 , n531 );
buf ( n4243 , n4242 );
and ( n4244 , n4243 , n4154 );
nor ( n4245 , n4241 , n4244 );
xnor ( n4246 , n4245 , n4152 );
not ( n4247 , n4189 );
buf ( n4248 , n467 );
buf ( n4249 , n4248 );
and ( n4250 , n4187 , n4167 );
not ( n4251 , n4250 );
and ( n4252 , n4249 , n4251 );
and ( n4253 , n4247 , n4252 );
xor ( n4254 , n4246 , n4253 );
and ( n4255 , n4176 , n4173 );
and ( n4256 , n4150 , n4171 );
nor ( n4257 , n4255 , n4256 );
xnor ( n4258 , n4257 , n4181 );
xor ( n4259 , n4254 , n4258 );
xor ( n4260 , n4249 , n4187 );
not ( n4261 , n4188 );
and ( n4262 , n4260 , n4261 );
and ( n4263 , n4185 , n4262 );
and ( n4264 , n4165 , n4188 );
nor ( n4265 , n4263 , n4264 );
xnor ( n4266 , n4265 , n4252 );
xor ( n4267 , n4259 , n4266 );
xor ( n4268 , n4240 , n4267 );
and ( n4269 , n4190 , n4198 );
and ( n4270 , n4199 , n4224 );
or ( n4271 , n4269 , n4270 );
xor ( n4272 , n4268 , n4271 );
buf ( n4273 , n4272 );
buf ( n4274 , n4273 );
buf ( n4275 , n4274 );
and ( n4276 , n4275 , n4232 );
nor ( n4277 , n4236 , n4276 );
xnor ( n4278 , n4277 , n4230 );
buf ( n4279 , n4217 );
buf ( n4280 , n4279 );
buf ( n4281 , n4280 );
buf ( n4282 , n4281 );
buf ( n4283 , n500 );
buf ( n4284 , n4283 );
buf ( n4285 , n501 );
buf ( n4286 , n4285 );
xor ( n4287 , n4284 , n4286 );
and ( n4288 , n4282 , n4287 );
not ( n4289 , n4288 );
buf ( n4290 , n499 );
buf ( n4291 , n4290 );
and ( n4292 , n4284 , n4286 );
not ( n4293 , n4292 );
and ( n4294 , n4291 , n4293 );
and ( n4295 , n4289 , n4294 );
xor ( n4296 , n4291 , n4284 );
not ( n4297 , n4287 );
and ( n4298 , n4296 , n4297 );
and ( n4299 , n4282 , n4298 );
xor ( n4300 , n4216 , n4219 );
buf ( n4301 , n4300 );
buf ( n4302 , n4301 );
buf ( n4303 , n4302 );
and ( n4304 , n4303 , n4287 );
nor ( n4305 , n4299 , n4304 );
xnor ( n4306 , n4305 , n4294 );
xor ( n4307 , n4295 , n4306 );
buf ( n4308 , n502 );
buf ( n4309 , n4308 );
xor ( n4310 , n4309 , n4230 );
and ( n4311 , n4282 , n4310 );
not ( n4312 , n4311 );
and ( n4313 , n4309 , n4230 );
not ( n4314 , n4313 );
and ( n4315 , n4286 , n4314 );
and ( n4316 , n4312 , n4315 );
xor ( n4317 , n4286 , n4309 );
not ( n4318 , n4310 );
and ( n4319 , n4317 , n4318 );
and ( n4320 , n4282 , n4319 );
and ( n4321 , n4303 , n4310 );
nor ( n4322 , n4320 , n4321 );
xnor ( n4323 , n4322 , n4315 );
and ( n4324 , n4316 , n4323 );
and ( n4325 , n4303 , n4319 );
xor ( n4326 , n4212 , n4220 );
buf ( n4327 , n4326 );
buf ( n4328 , n4327 );
buf ( n4329 , n4328 );
and ( n4330 , n4329 , n4310 );
nor ( n4331 , n4325 , n4330 );
xnor ( n4332 , n4331 , n4315 );
and ( n4333 , n4324 , n4332 );
and ( n4334 , n4332 , n4288 );
and ( n4335 , n4324 , n4288 );
or ( n4336 , n4333 , n4334 , n4335 );
xor ( n4337 , n4307 , n4336 );
and ( n4338 , n4329 , n4319 );
xor ( n4339 , n4206 , n4222 );
buf ( n4340 , n4339 );
buf ( n4341 , n4340 );
buf ( n4342 , n4341 );
and ( n4343 , n4342 , n4310 );
nor ( n4344 , n4338 , n4343 );
xnor ( n4345 , n4344 , n4315 );
xor ( n4346 , n4337 , n4345 );
xor ( n4347 , n4278 , n4346 );
and ( n4348 , n4342 , n4235 );
and ( n4349 , n4228 , n4232 );
nor ( n4350 , n4348 , n4349 );
xnor ( n4351 , n4350 , n4230 );
xor ( n4352 , n4324 , n4332 );
xor ( n4353 , n4352 , n4288 );
and ( n4354 , n4351 , n4353 );
xor ( n4355 , n4351 , n4353 );
and ( n4356 , n4329 , n4235 );
and ( n4357 , n4342 , n4232 );
nor ( n4358 , n4356 , n4357 );
xnor ( n4359 , n4358 , n4230 );
xor ( n4360 , n4316 , n4323 );
and ( n4361 , n4359 , n4360 );
xor ( n4362 , n4359 , n4360 );
and ( n4363 , n4303 , n4235 );
and ( n4364 , n4329 , n4232 );
nor ( n4365 , n4363 , n4364 );
xnor ( n4366 , n4365 , n4230 );
and ( n4367 , n4366 , n4311 );
xor ( n4368 , n4366 , n4311 );
and ( n4369 , n4282 , n4235 );
and ( n4370 , n4303 , n4232 );
nor ( n4371 , n4369 , n4370 );
xnor ( n4372 , n4371 , n4230 );
and ( n4373 , n4282 , n4232 );
not ( n4374 , n4373 );
and ( n4375 , n4374 , n4230 );
and ( n4376 , n4372 , n4375 );
and ( n4377 , n4368 , n4376 );
or ( n4378 , n4367 , n4377 );
and ( n4379 , n4362 , n4378 );
or ( n4380 , n4361 , n4379 );
and ( n4381 , n4355 , n4380 );
or ( n4382 , n4354 , n4381 );
xor ( n4383 , n4347 , n4382 );
buf ( n4384 , n4383 );
buf ( n4385 , n814 );
buf ( n4386 , n4385 );
buf ( n4387 , n548 );
buf ( n4388 , n4387 );
buf ( n4389 , n549 );
buf ( n4390 , n4389 );
xor ( n4391 , n4388 , n4390 );
and ( n4392 , n4386 , n4391 );
not ( n4393 , n4392 );
buf ( n4394 , n547 );
buf ( n4395 , n4394 );
and ( n4396 , n4388 , n4390 );
not ( n4397 , n4396 );
and ( n4398 , n4395 , n4397 );
and ( n4399 , n4393 , n4398 );
xor ( n4400 , n4395 , n4388 );
not ( n4401 , n4391 );
and ( n4402 , n4400 , n4401 );
and ( n4403 , n4386 , n4402 );
buf ( n4404 , n869 );
buf ( n4405 , n4404 );
and ( n4406 , n4405 , n4391 );
nor ( n4407 , n4403 , n4406 );
xnor ( n4408 , n4407 , n4398 );
xor ( n4409 , n4399 , n4408 );
buf ( n4410 , n1141 );
buf ( n4411 , n4410 );
buf ( n4412 , n551 );
buf ( n4413 , n4412 );
buf ( n4414 , n552 );
buf ( n4415 , n4414 );
xor ( n4416 , n4413 , n4415 );
not ( n4417 , n4415 );
and ( n4418 , n4416 , n4417 );
and ( n4419 , n4411 , n4418 );
buf ( n4420 , n1242 );
buf ( n4421 , n4420 );
and ( n4422 , n4421 , n4415 );
nor ( n4423 , n4419 , n4422 );
xnor ( n4424 , n4423 , n4413 );
xor ( n4425 , n4409 , n4424 );
buf ( n4426 , n956 );
buf ( n4427 , n4426 );
buf ( n4428 , n550 );
buf ( n4429 , n4428 );
xor ( n4430 , n4390 , n4429 );
xor ( n4431 , n4429 , n4413 );
not ( n4432 , n4431 );
and ( n4433 , n4430 , n4432 );
and ( n4434 , n4427 , n4433 );
buf ( n4435 , n1035 );
buf ( n4436 , n4435 );
and ( n4437 , n4436 , n4431 );
nor ( n4438 , n4434 , n4437 );
and ( n4439 , n4429 , n4413 );
not ( n4440 , n4439 );
and ( n4441 , n4390 , n4440 );
xnor ( n4442 , n4438 , n4441 );
xor ( n4443 , n4425 , n4442 );
and ( n4444 , n4386 , n4431 );
not ( n4445 , n4444 );
and ( n4446 , n4445 , n4441 );
and ( n4447 , n4386 , n4433 );
and ( n4448 , n4405 , n4431 );
nor ( n4449 , n4447 , n4448 );
xnor ( n4450 , n4449 , n4441 );
and ( n4451 , n4446 , n4450 );
and ( n4452 , n4405 , n4433 );
and ( n4453 , n4427 , n4431 );
nor ( n4454 , n4452 , n4453 );
xnor ( n4455 , n4454 , n4441 );
and ( n4456 , n4451 , n4455 );
and ( n4457 , n4455 , n4392 );
and ( n4458 , n4451 , n4392 );
or ( n4459 , n4456 , n4457 , n4458 );
xor ( n4460 , n4443 , n4459 );
and ( n4461 , n4436 , n4418 );
and ( n4462 , n4411 , n4415 );
nor ( n4463 , n4461 , n4462 );
xnor ( n4464 , n4463 , n4413 );
xor ( n4465 , n4451 , n4455 );
xor ( n4466 , n4465 , n4392 );
and ( n4467 , n4464 , n4466 );
xor ( n4468 , n4464 , n4466 );
and ( n4469 , n4427 , n4418 );
and ( n4470 , n4436 , n4415 );
nor ( n4471 , n4469 , n4470 );
xnor ( n4472 , n4471 , n4413 );
xor ( n4473 , n4446 , n4450 );
and ( n4474 , n4472 , n4473 );
xor ( n4475 , n4472 , n4473 );
and ( n4476 , n4405 , n4418 );
and ( n4477 , n4427 , n4415 );
nor ( n4478 , n4476 , n4477 );
xnor ( n4479 , n4478 , n4413 );
and ( n4480 , n4479 , n4444 );
xor ( n4481 , n4479 , n4444 );
and ( n4482 , n4386 , n4418 );
and ( n4483 , n4405 , n4415 );
nor ( n4484 , n4482 , n4483 );
xnor ( n4485 , n4484 , n4413 );
and ( n4486 , n4386 , n4415 );
not ( n4487 , n4486 );
and ( n4488 , n4487 , n4413 );
and ( n4489 , n4485 , n4488 );
and ( n4490 , n4481 , n4489 );
or ( n4491 , n4480 , n4490 );
and ( n4492 , n4475 , n4491 );
or ( n4493 , n4474 , n4492 );
and ( n4494 , n4468 , n4493 );
or ( n4495 , n4467 , n4494 );
xor ( n4496 , n4460 , n4495 );
buf ( n4497 , n4496 );
not ( n4498 , n454 );
and ( n4499 , n4498 , n4384 );
and ( n4500 , n4497 , n454 );
or ( n4501 , n4499 , n4500 );
buf ( n4502 , n4501 );
buf ( n4503 , n4502 );
buf ( n4504 , n472 );
buf ( n4505 , n4504 );
and ( n4506 , n4503 , n4505 );
buf ( n4507 , n4506 );
or ( n4508 , n456 , n455 );
and ( n4509 , n4508 , n454 );
not ( n4510 , n4509 );
and ( n4511 , n4510 , n4148 );
and ( n4512 , n4507 , n4509 );
or ( n4513 , n4511 , n4512 );
buf ( n4514 , n535 );
buf ( n4515 , n551 );
xor ( n4516 , n4514 , n4515 );
and ( n4517 , n4140 , n4141 );
xor ( n4518 , n4516 , n4517 );
buf ( n4519 , n4518 );
buf ( n4520 , n4519 );
buf ( n4521 , n4520 );
xor ( n4522 , n4521 , n4145 );
not ( n4523 , n4145 );
and ( n4524 , n4522 , n4523 );
and ( n4525 , n4139 , n4524 );
buf ( n4526 , n782 );
buf ( n4527 , n4526 );
xor ( n4528 , n4527 , n4134 );
not ( n4529 , n4134 );
and ( n4530 , n4528 , n4529 );
and ( n4531 , n4132 , n4530 );
buf ( n4532 , n503 );
buf ( n4533 , n519 );
xor ( n4534 , n4532 , n4533 );
and ( n4535 , n4127 , n4128 );
xor ( n4536 , n4534 , n4535 );
buf ( n4537 , n4536 );
buf ( n4538 , n4537 );
buf ( n4539 , n4538 );
and ( n4540 , n4539 , n4134 );
nor ( n4541 , n4531 , n4540 );
xnor ( n4542 , n4541 , n4527 );
not ( n4543 , n4135 );
and ( n4544 , n4543 , n4527 );
xor ( n4545 , n4542 , n4544 );
buf ( n4546 , n4545 );
buf ( n4547 , n4546 );
buf ( n4548 , n4547 );
and ( n4549 , n4548 , n4145 );
nor ( n4550 , n4525 , n4549 );
xnor ( n4551 , n4550 , n4521 );
not ( n4552 , n4146 );
and ( n4553 , n4552 , n4521 );
xor ( n4554 , n4551 , n4553 );
buf ( n4555 , n4554 );
buf ( n4556 , n471 );
buf ( n4557 , n4556 );
and ( n4558 , n4503 , n4557 );
and ( n4559 , n4275 , n4235 );
and ( n4560 , n4246 , n4253 );
and ( n4561 , n4165 , n4262 );
and ( n4562 , n4176 , n4188 );
nor ( n4563 , n4561 , n4562 );
xnor ( n4564 , n4563 , n4252 );
xor ( n4565 , n4560 , n4564 );
and ( n4566 , n4243 , n4157 );
buf ( n4567 , n530 );
buf ( n4568 , n4567 );
and ( n4569 , n4568 , n4154 );
nor ( n4570 , n4566 , n4569 );
xnor ( n4571 , n4570 , n4152 );
and ( n4572 , n4150 , n4173 );
and ( n4573 , n4160 , n4171 );
nor ( n4574 , n4572 , n4573 );
xnor ( n4575 , n4574 , n4181 );
xor ( n4576 , n4571 , n4575 );
buf ( n4577 , n466 );
buf ( n4578 , n4577 );
xor ( n4579 , n4578 , n4249 );
and ( n4580 , n4185 , n4579 );
xor ( n4581 , n4576 , n4580 );
xor ( n4582 , n4565 , n4581 );
and ( n4583 , n4254 , n4258 );
and ( n4584 , n4258 , n4266 );
and ( n4585 , n4254 , n4266 );
or ( n4586 , n4583 , n4584 , n4585 );
xor ( n4587 , n4582 , n4586 );
and ( n4588 , n4240 , n4267 );
and ( n4589 , n4268 , n4271 );
or ( n4590 , n4588 , n4589 );
xor ( n4591 , n4587 , n4590 );
buf ( n4592 , n4591 );
buf ( n4593 , n4592 );
buf ( n4594 , n4593 );
and ( n4595 , n4594 , n4232 );
nor ( n4596 , n4559 , n4595 );
xnor ( n4597 , n4596 , n4230 );
and ( n4598 , n4342 , n4319 );
and ( n4599 , n4228 , n4310 );
nor ( n4600 , n4598 , n4599 );
xnor ( n4601 , n4600 , n4315 );
xor ( n4602 , n4597 , n4601 );
and ( n4603 , n4295 , n4306 );
and ( n4604 , n4303 , n4298 );
and ( n4605 , n4329 , n4287 );
nor ( n4606 , n4604 , n4605 );
xnor ( n4607 , n4606 , n4294 );
xor ( n4608 , n4603 , n4607 );
buf ( n4609 , n498 );
buf ( n4610 , n4609 );
xor ( n4611 , n4610 , n4291 );
and ( n4612 , n4282 , n4611 );
xor ( n4613 , n4608 , n4612 );
xor ( n4614 , n4602 , n4613 );
and ( n4615 , n4307 , n4336 );
and ( n4616 , n4336 , n4345 );
and ( n4617 , n4307 , n4345 );
or ( n4618 , n4615 , n4616 , n4617 );
xor ( n4619 , n4614 , n4618 );
and ( n4620 , n4278 , n4346 );
and ( n4621 , n4347 , n4382 );
or ( n4622 , n4620 , n4621 );
xor ( n4623 , n4619 , n4622 );
buf ( n4624 , n4623 );
and ( n4625 , n4409 , n4424 );
and ( n4626 , n4424 , n4442 );
and ( n4627 , n4409 , n4442 );
or ( n4628 , n4625 , n4626 , n4627 );
and ( n4629 , n4421 , n4418 );
buf ( n4630 , n1372 );
buf ( n4631 , n4630 );
and ( n4632 , n4631 , n4415 );
nor ( n4633 , n4629 , n4632 );
xnor ( n4634 , n4633 , n4413 );
and ( n4635 , n4436 , n4433 );
and ( n4636 , n4411 , n4431 );
nor ( n4637 , n4635 , n4636 );
xnor ( n4638 , n4637 , n4441 );
xor ( n4639 , n4634 , n4638 );
and ( n4640 , n4399 , n4408 );
and ( n4641 , n4405 , n4402 );
and ( n4642 , n4427 , n4391 );
nor ( n4643 , n4641 , n4642 );
xnor ( n4644 , n4643 , n4398 );
xor ( n4645 , n4640 , n4644 );
buf ( n4646 , n546 );
buf ( n4647 , n4646 );
xor ( n4648 , n4647 , n4395 );
and ( n4649 , n4386 , n4648 );
xor ( n4650 , n4645 , n4649 );
xor ( n4651 , n4639 , n4650 );
xor ( n4652 , n4628 , n4651 );
and ( n4653 , n4443 , n4459 );
and ( n4654 , n4460 , n4495 );
or ( n4655 , n4653 , n4654 );
xor ( n4656 , n4652 , n4655 );
buf ( n4657 , n4656 );
not ( n4658 , n454 );
and ( n4659 , n4658 , n4624 );
and ( n4660 , n4657 , n454 );
or ( n4661 , n4659 , n4660 );
buf ( n4662 , n4661 );
buf ( n4663 , n4662 );
and ( n4664 , n4663 , n4505 );
xor ( n4665 , n4558 , n4664 );
buf ( n4666 , n4665 );
not ( n4667 , n4509 );
and ( n4668 , n4667 , n4555 );
and ( n4669 , n4666 , n4509 );
or ( n4670 , n4668 , n4669 );
and ( n4671 , n4548 , n4524 );
and ( n4672 , n4539 , n4530 );
buf ( n4673 , n502 );
buf ( n4674 , n518 );
xor ( n4675 , n4673 , n4674 );
and ( n4676 , n4532 , n4533 );
and ( n4677 , n4533 , n4535 );
and ( n4678 , n4532 , n4535 );
or ( n4679 , n4676 , n4677 , n4678 );
xor ( n4680 , n4675 , n4679 );
buf ( n4681 , n4680 );
buf ( n4682 , n4681 );
buf ( n4683 , n4682 );
and ( n4684 , n4683 , n4134 );
nor ( n4685 , n4672 , n4684 );
xnor ( n4686 , n4685 , n4527 );
buf ( n4687 , n843 );
buf ( n4688 , n4687 );
xor ( n4689 , n4688 , n4527 );
and ( n4690 , n4132 , n4689 );
xor ( n4691 , n4686 , n4690 );
and ( n4692 , n4542 , n4544 );
xor ( n4693 , n4691 , n4692 );
buf ( n4694 , n4693 );
buf ( n4695 , n4694 );
buf ( n4696 , n4695 );
and ( n4697 , n4696 , n4145 );
nor ( n4698 , n4671 , n4697 );
xnor ( n4699 , n4698 , n4521 );
buf ( n4700 , n534 );
buf ( n4701 , n550 );
xor ( n4702 , n4700 , n4701 );
and ( n4703 , n4514 , n4515 );
and ( n4704 , n4515 , n4517 );
and ( n4705 , n4514 , n4517 );
or ( n4706 , n4703 , n4704 , n4705 );
xor ( n4707 , n4702 , n4706 );
buf ( n4708 , n4707 );
buf ( n4709 , n4708 );
buf ( n4710 , n4709 );
xor ( n4711 , n4710 , n4521 );
and ( n4712 , n4139 , n4711 );
xor ( n4713 , n4699 , n4712 );
and ( n4714 , n4551 , n4553 );
xor ( n4715 , n4713 , n4714 );
buf ( n4716 , n4715 );
and ( n4717 , n4597 , n4601 );
and ( n4718 , n4601 , n4613 );
and ( n4719 , n4597 , n4613 );
or ( n4720 , n4717 , n4718 , n4719 );
and ( n4721 , n4594 , n4235 );
and ( n4722 , n4568 , n4157 );
buf ( n4723 , n529 );
buf ( n4724 , n4723 );
and ( n4725 , n4724 , n4154 );
nor ( n4726 , n4722 , n4725 );
xnor ( n4727 , n4726 , n4152 );
not ( n4728 , n4580 );
buf ( n4729 , n465 );
buf ( n4730 , n4729 );
and ( n4731 , n4578 , n4249 );
not ( n4732 , n4731 );
and ( n4733 , n4730 , n4732 );
and ( n4734 , n4728 , n4733 );
xor ( n4735 , n4727 , n4734 );
and ( n4736 , n4571 , n4575 );
and ( n4737 , n4575 , n4580 );
and ( n4738 , n4571 , n4580 );
or ( n4739 , n4736 , n4737 , n4738 );
xor ( n4740 , n4735 , n4739 );
and ( n4741 , n4160 , n4173 );
and ( n4742 , n4243 , n4171 );
nor ( n4743 , n4741 , n4742 );
xnor ( n4744 , n4743 , n4181 );
and ( n4745 , n4176 , n4262 );
and ( n4746 , n4150 , n4188 );
nor ( n4747 , n4745 , n4746 );
xnor ( n4748 , n4747 , n4252 );
xor ( n4749 , n4744 , n4748 );
xor ( n4750 , n4730 , n4578 );
not ( n4751 , n4579 );
and ( n4752 , n4750 , n4751 );
and ( n4753 , n4185 , n4752 );
and ( n4754 , n4165 , n4579 );
nor ( n4755 , n4753 , n4754 );
xnor ( n4756 , n4755 , n4733 );
xor ( n4757 , n4749 , n4756 );
xor ( n4758 , n4740 , n4757 );
and ( n4759 , n4560 , n4564 );
and ( n4760 , n4564 , n4581 );
and ( n4761 , n4560 , n4581 );
or ( n4762 , n4759 , n4760 , n4761 );
xor ( n4763 , n4758 , n4762 );
and ( n4764 , n4582 , n4586 );
and ( n4765 , n4587 , n4590 );
or ( n4766 , n4764 , n4765 );
xor ( n4767 , n4763 , n4766 );
buf ( n4768 , n4767 );
buf ( n4769 , n4768 );
buf ( n4770 , n4769 );
and ( n4771 , n4770 , n4232 );
nor ( n4772 , n4721 , n4771 );
xnor ( n4773 , n4772 , n4230 );
and ( n4774 , n4228 , n4319 );
and ( n4775 , n4275 , n4310 );
nor ( n4776 , n4774 , n4775 );
xnor ( n4777 , n4776 , n4315 );
xor ( n4778 , n4773 , n4777 );
not ( n4779 , n4612 );
buf ( n4780 , n497 );
buf ( n4781 , n4780 );
and ( n4782 , n4610 , n4291 );
not ( n4783 , n4782 );
and ( n4784 , n4781 , n4783 );
and ( n4785 , n4779 , n4784 );
xor ( n4786 , n4781 , n4610 );
not ( n4787 , n4611 );
and ( n4788 , n4786 , n4787 );
and ( n4789 , n4282 , n4788 );
and ( n4790 , n4303 , n4611 );
nor ( n4791 , n4789 , n4790 );
xnor ( n4792 , n4791 , n4784 );
xor ( n4793 , n4785 , n4792 );
and ( n4794 , n4603 , n4607 );
and ( n4795 , n4607 , n4612 );
and ( n4796 , n4603 , n4612 );
or ( n4797 , n4794 , n4795 , n4796 );
xor ( n4798 , n4793 , n4797 );
and ( n4799 , n4329 , n4298 );
and ( n4800 , n4342 , n4287 );
nor ( n4801 , n4799 , n4800 );
xnor ( n4802 , n4801 , n4294 );
xor ( n4803 , n4798 , n4802 );
xor ( n4804 , n4778 , n4803 );
xor ( n4805 , n4720 , n4804 );
and ( n4806 , n4614 , n4618 );
and ( n4807 , n4619 , n4622 );
or ( n4808 , n4806 , n4807 );
xor ( n4809 , n4805 , n4808 );
buf ( n4810 , n4809 );
and ( n4811 , n4634 , n4638 );
and ( n4812 , n4638 , n4650 );
and ( n4813 , n4634 , n4650 );
or ( n4814 , n4811 , n4812 , n4813 );
and ( n4815 , n4631 , n4418 );
buf ( n4816 , n1498 );
buf ( n4817 , n4816 );
and ( n4818 , n4817 , n4415 );
nor ( n4819 , n4815 , n4818 );
xnor ( n4820 , n4819 , n4413 );
and ( n4821 , n4411 , n4433 );
and ( n4822 , n4421 , n4431 );
nor ( n4823 , n4821 , n4822 );
xnor ( n4824 , n4823 , n4441 );
xor ( n4825 , n4820 , n4824 );
not ( n4826 , n4649 );
buf ( n4827 , n545 );
buf ( n4828 , n4827 );
and ( n4829 , n4647 , n4395 );
not ( n4830 , n4829 );
and ( n4831 , n4828 , n4830 );
and ( n4832 , n4826 , n4831 );
xor ( n4833 , n4828 , n4647 );
not ( n4834 , n4648 );
and ( n4835 , n4833 , n4834 );
and ( n4836 , n4386 , n4835 );
and ( n4837 , n4405 , n4648 );
nor ( n4838 , n4836 , n4837 );
xnor ( n4839 , n4838 , n4831 );
xor ( n4840 , n4832 , n4839 );
and ( n4841 , n4640 , n4644 );
and ( n4842 , n4644 , n4649 );
and ( n4843 , n4640 , n4649 );
or ( n4844 , n4841 , n4842 , n4843 );
xor ( n4845 , n4840 , n4844 );
and ( n4846 , n4427 , n4402 );
and ( n4847 , n4436 , n4391 );
nor ( n4848 , n4846 , n4847 );
xnor ( n4849 , n4848 , n4398 );
xor ( n4850 , n4845 , n4849 );
xor ( n4851 , n4825 , n4850 );
xor ( n4852 , n4814 , n4851 );
and ( n4853 , n4628 , n4651 );
and ( n4854 , n4652 , n4655 );
or ( n4855 , n4853 , n4854 );
xor ( n4856 , n4852 , n4855 );
buf ( n4857 , n4856 );
not ( n4858 , n454 );
and ( n4859 , n4858 , n4810 );
and ( n4860 , n4857 , n454 );
or ( n4861 , n4859 , n4860 );
buf ( n4862 , n4861 );
buf ( n4863 , n4862 );
and ( n4864 , n4863 , n4505 );
buf ( n4865 , n470 );
buf ( n4866 , n4865 );
and ( n4867 , n4503 , n4866 );
and ( n4868 , n4663 , n4557 );
xor ( n4869 , n4867 , n4868 );
xor ( n4870 , n4864 , n4869 );
and ( n4871 , n4558 , n4664 );
xor ( n4872 , n4870 , n4871 );
buf ( n4873 , n4872 );
not ( n4874 , n4509 );
and ( n4875 , n4874 , n4716 );
and ( n4876 , n4873 , n4509 );
or ( n4877 , n4875 , n4876 );
and ( n4878 , n4696 , n4524 );
and ( n4879 , n4683 , n4530 );
buf ( n4880 , n501 );
buf ( n4881 , n517 );
xor ( n4882 , n4880 , n4881 );
and ( n4883 , n4673 , n4674 );
and ( n4884 , n4674 , n4679 );
and ( n4885 , n4673 , n4679 );
or ( n4886 , n4883 , n4884 , n4885 );
xor ( n4887 , n4882 , n4886 );
buf ( n4888 , n4887 );
buf ( n4889 , n4888 );
buf ( n4890 , n4889 );
and ( n4891 , n4890 , n4134 );
nor ( n4892 , n4879 , n4891 );
xnor ( n4893 , n4892 , n4527 );
buf ( n4894 , n937 );
buf ( n4895 , n4894 );
xor ( n4896 , n4895 , n4688 );
not ( n4897 , n4689 );
and ( n4898 , n4896 , n4897 );
and ( n4899 , n4132 , n4898 );
and ( n4900 , n4539 , n4689 );
nor ( n4901 , n4899 , n4900 );
and ( n4902 , n4688 , n4527 );
not ( n4903 , n4902 );
and ( n4904 , n4895 , n4903 );
xnor ( n4905 , n4901 , n4904 );
xor ( n4906 , n4893 , n4905 );
not ( n4907 , n4690 );
and ( n4908 , n4907 , n4904 );
xor ( n4909 , n4906 , n4908 );
and ( n4910 , n4686 , n4690 );
and ( n4911 , n4691 , n4692 );
or ( n4912 , n4910 , n4911 );
xor ( n4913 , n4909 , n4912 );
buf ( n4914 , n4913 );
buf ( n4915 , n4914 );
buf ( n4916 , n4915 );
and ( n4917 , n4916 , n4145 );
nor ( n4918 , n4878 , n4917 );
xnor ( n4919 , n4918 , n4521 );
not ( n4920 , n4712 );
buf ( n4921 , n533 );
buf ( n4922 , n549 );
xor ( n4923 , n4921 , n4922 );
and ( n4924 , n4700 , n4701 );
and ( n4925 , n4701 , n4706 );
and ( n4926 , n4700 , n4706 );
or ( n4927 , n4924 , n4925 , n4926 );
xor ( n4928 , n4923 , n4927 );
buf ( n4929 , n4928 );
buf ( n4930 , n4929 );
buf ( n4931 , n4930 );
and ( n4932 , n4710 , n4521 );
not ( n4933 , n4932 );
and ( n4934 , n4931 , n4933 );
and ( n4935 , n4920 , n4934 );
xor ( n4936 , n4931 , n4710 );
not ( n4937 , n4711 );
and ( n4938 , n4936 , n4937 );
and ( n4939 , n4139 , n4938 );
and ( n4940 , n4548 , n4711 );
nor ( n4941 , n4939 , n4940 );
xnor ( n4942 , n4941 , n4934 );
xor ( n4943 , n4935 , n4942 );
xor ( n4944 , n4919 , n4943 );
and ( n4945 , n4699 , n4712 );
and ( n4946 , n4713 , n4714 );
or ( n4947 , n4945 , n4946 );
xor ( n4948 , n4944 , n4947 );
buf ( n4949 , n4948 );
and ( n4950 , n4793 , n4797 );
and ( n4951 , n4797 , n4802 );
and ( n4952 , n4793 , n4802 );
or ( n4953 , n4950 , n4951 , n4952 );
and ( n4954 , n4770 , n4235 );
and ( n4955 , n4735 , n4739 );
and ( n4956 , n4739 , n4757 );
and ( n4957 , n4735 , n4757 );
or ( n4958 , n4955 , n4956 , n4957 );
and ( n4959 , n4744 , n4748 );
and ( n4960 , n4748 , n4756 );
and ( n4961 , n4744 , n4756 );
or ( n4962 , n4959 , n4960 , n4961 );
and ( n4963 , n4724 , n4157 );
buf ( n4964 , n528 );
buf ( n4965 , n4964 );
and ( n4966 , n4965 , n4154 );
nor ( n4967 , n4963 , n4966 );
xnor ( n4968 , n4967 , n4152 );
and ( n4969 , n4165 , n4752 );
and ( n4970 , n4176 , n4579 );
nor ( n4971 , n4969 , n4970 );
xnor ( n4972 , n4971 , n4733 );
xor ( n4973 , n4968 , n4972 );
buf ( n4974 , n464 );
buf ( n4975 , n4974 );
xor ( n4976 , n4975 , n4730 );
and ( n4977 , n4185 , n4976 );
xor ( n4978 , n4973 , n4977 );
xor ( n4979 , n4962 , n4978 );
and ( n4980 , n4727 , n4734 );
and ( n4981 , n4243 , n4173 );
and ( n4982 , n4568 , n4171 );
nor ( n4983 , n4981 , n4982 );
xnor ( n4984 , n4983 , n4181 );
xor ( n4985 , n4980 , n4984 );
and ( n4986 , n4150 , n4262 );
and ( n4987 , n4160 , n4188 );
nor ( n4988 , n4986 , n4987 );
xnor ( n4989 , n4988 , n4252 );
xor ( n4990 , n4985 , n4989 );
xor ( n4991 , n4979 , n4990 );
xor ( n4992 , n4958 , n4991 );
and ( n4993 , n4758 , n4762 );
and ( n4994 , n4763 , n4766 );
or ( n4995 , n4993 , n4994 );
xor ( n4996 , n4992 , n4995 );
buf ( n4997 , n4996 );
buf ( n4998 , n4997 );
buf ( n4999 , n4998 );
and ( n5000 , n4999 , n4232 );
nor ( n5001 , n4954 , n5000 );
xnor ( n5002 , n5001 , n4230 );
xor ( n5003 , n4953 , n5002 );
and ( n5004 , n4275 , n4319 );
and ( n5005 , n4594 , n4310 );
nor ( n5006 , n5004 , n5005 );
xnor ( n5007 , n5006 , n4315 );
and ( n5008 , n4342 , n4298 );
and ( n5009 , n4228 , n4287 );
nor ( n5010 , n5008 , n5009 );
xnor ( n5011 , n5010 , n4294 );
xor ( n5012 , n5007 , n5011 );
and ( n5013 , n4785 , n4792 );
and ( n5014 , n4303 , n4788 );
and ( n5015 , n4329 , n4611 );
nor ( n5016 , n5014 , n5015 );
xnor ( n5017 , n5016 , n4784 );
xor ( n5018 , n5013 , n5017 );
buf ( n5019 , n496 );
buf ( n5020 , n5019 );
xor ( n5021 , n5020 , n4781 );
and ( n5022 , n4282 , n5021 );
xor ( n5023 , n5018 , n5022 );
xor ( n5024 , n5012 , n5023 );
xor ( n5025 , n5003 , n5024 );
and ( n5026 , n4773 , n4777 );
and ( n5027 , n4777 , n4803 );
and ( n5028 , n4773 , n4803 );
or ( n5029 , n5026 , n5027 , n5028 );
xor ( n5030 , n5025 , n5029 );
and ( n5031 , n4720 , n4804 );
and ( n5032 , n4805 , n4808 );
or ( n5033 , n5031 , n5032 );
xor ( n5034 , n5030 , n5033 );
buf ( n5035 , n5034 );
and ( n5036 , n4840 , n4844 );
and ( n5037 , n4844 , n4849 );
and ( n5038 , n4840 , n4849 );
or ( n5039 , n5036 , n5037 , n5038 );
and ( n5040 , n4817 , n4418 );
buf ( n5041 , n1645 );
buf ( n5042 , n5041 );
and ( n5043 , n5042 , n4415 );
nor ( n5044 , n5040 , n5043 );
xnor ( n5045 , n5044 , n4413 );
xor ( n5046 , n5039 , n5045 );
and ( n5047 , n4421 , n4433 );
and ( n5048 , n4631 , n4431 );
nor ( n5049 , n5047 , n5048 );
xnor ( n5050 , n5049 , n4441 );
and ( n5051 , n4436 , n4402 );
and ( n5052 , n4411 , n4391 );
nor ( n5053 , n5051 , n5052 );
xnor ( n5054 , n5053 , n4398 );
xor ( n5055 , n5050 , n5054 );
and ( n5056 , n4832 , n4839 );
and ( n5057 , n4405 , n4835 );
and ( n5058 , n4427 , n4648 );
nor ( n5059 , n5057 , n5058 );
xnor ( n5060 , n5059 , n4831 );
xor ( n5061 , n5056 , n5060 );
buf ( n5062 , n544 );
buf ( n5063 , n5062 );
xor ( n5064 , n5063 , n4828 );
and ( n5065 , n4386 , n5064 );
xor ( n5066 , n5061 , n5065 );
xor ( n5067 , n5055 , n5066 );
xor ( n5068 , n5046 , n5067 );
and ( n5069 , n4820 , n4824 );
and ( n5070 , n4824 , n4850 );
and ( n5071 , n4820 , n4850 );
or ( n5072 , n5069 , n5070 , n5071 );
xor ( n5073 , n5068 , n5072 );
and ( n5074 , n4814 , n4851 );
and ( n5075 , n4852 , n4855 );
or ( n5076 , n5074 , n5075 );
xor ( n5077 , n5073 , n5076 );
buf ( n5078 , n5077 );
not ( n5079 , n454 );
and ( n5080 , n5079 , n5035 );
and ( n5081 , n5078 , n454 );
or ( n5082 , n5080 , n5081 );
buf ( n5083 , n5082 );
buf ( n5084 , n5083 );
and ( n5085 , n5084 , n4505 );
and ( n5086 , n4867 , n4868 );
xor ( n5087 , n5085 , n5086 );
buf ( n5088 , n469 );
buf ( n5089 , n5088 );
and ( n5090 , n4503 , n5089 );
and ( n5091 , n4663 , n4866 );
xor ( n5092 , n5090 , n5091 );
and ( n5093 , n4863 , n4557 );
xor ( n5094 , n5092 , n5093 );
xor ( n5095 , n5087 , n5094 );
and ( n5096 , n4864 , n4869 );
and ( n5097 , n4870 , n4871 );
or ( n5098 , n5096 , n5097 );
xor ( n5099 , n5095 , n5098 );
buf ( n5100 , n5099 );
not ( n5101 , n4509 );
and ( n5102 , n5101 , n4949 );
and ( n5103 , n5100 , n4509 );
or ( n5104 , n5102 , n5103 );
and ( n5105 , n4916 , n4524 );
and ( n5106 , n4893 , n4905 );
and ( n5107 , n4905 , n4908 );
and ( n5108 , n4893 , n4908 );
or ( n5109 , n5106 , n5107 , n5108 );
and ( n5110 , n4890 , n4530 );
buf ( n5111 , n500 );
buf ( n5112 , n516 );
xor ( n5113 , n5111 , n5112 );
and ( n5114 , n4880 , n4881 );
and ( n5115 , n4881 , n4886 );
and ( n5116 , n4880 , n4886 );
or ( n5117 , n5114 , n5115 , n5116 );
xor ( n5118 , n5113 , n5117 );
buf ( n5119 , n5118 );
buf ( n5120 , n5119 );
buf ( n5121 , n5120 );
and ( n5122 , n5121 , n4134 );
nor ( n5123 , n5110 , n5122 );
xnor ( n5124 , n5123 , n4527 );
and ( n5125 , n4539 , n4898 );
and ( n5126 , n4683 , n4689 );
nor ( n5127 , n5125 , n5126 );
xnor ( n5128 , n5127 , n4904 );
xor ( n5129 , n5124 , n5128 );
buf ( n5130 , n1007 );
buf ( n5131 , n5130 );
xor ( n5132 , n5131 , n4895 );
and ( n5133 , n4132 , n5132 );
xor ( n5134 , n5129 , n5133 );
xor ( n5135 , n5109 , n5134 );
and ( n5136 , n4909 , n4912 );
xor ( n5137 , n5135 , n5136 );
buf ( n5138 , n5137 );
buf ( n5139 , n5138 );
buf ( n5140 , n5139 );
and ( n5141 , n5140 , n4145 );
nor ( n5142 , n5105 , n5141 );
xnor ( n5143 , n5142 , n4521 );
and ( n5144 , n4935 , n4942 );
and ( n5145 , n4548 , n4938 );
and ( n5146 , n4696 , n4711 );
nor ( n5147 , n5145 , n5146 );
xnor ( n5148 , n5147 , n4934 );
xor ( n5149 , n5144 , n5148 );
buf ( n5150 , n532 );
buf ( n5151 , n548 );
xor ( n5152 , n5150 , n5151 );
and ( n5153 , n4921 , n4922 );
and ( n5154 , n4922 , n4927 );
and ( n5155 , n4921 , n4927 );
or ( n5156 , n5153 , n5154 , n5155 );
xor ( n5157 , n5152 , n5156 );
buf ( n5158 , n5157 );
buf ( n5159 , n5158 );
buf ( n5160 , n5159 );
xor ( n5161 , n5160 , n4931 );
and ( n5162 , n4139 , n5161 );
xor ( n5163 , n5149 , n5162 );
xor ( n5164 , n5143 , n5163 );
and ( n5165 , n4919 , n4943 );
and ( n5166 , n4944 , n4947 );
or ( n5167 , n5165 , n5166 );
xor ( n5168 , n5164 , n5167 );
buf ( n5169 , n5168 );
and ( n5170 , n5090 , n5091 );
and ( n5171 , n5091 , n5093 );
and ( n5172 , n5090 , n5093 );
or ( n5173 , n5170 , n5171 , n5172 );
and ( n5174 , n5085 , n5086 );
and ( n5175 , n5086 , n5094 );
and ( n5176 , n5085 , n5094 );
or ( n5177 , n5174 , n5175 , n5176 );
xor ( n5178 , n5173 , n5177 );
and ( n5179 , n5084 , n4557 );
and ( n5180 , n4953 , n5002 );
and ( n5181 , n5002 , n5024 );
and ( n5182 , n4953 , n5024 );
or ( n5183 , n5180 , n5181 , n5182 );
and ( n5184 , n5007 , n5011 );
and ( n5185 , n5011 , n5023 );
and ( n5186 , n5007 , n5023 );
or ( n5187 , n5184 , n5185 , n5186 );
and ( n5188 , n4999 , n4235 );
and ( n5189 , n4980 , n4984 );
and ( n5190 , n4984 , n4989 );
and ( n5191 , n4980 , n4989 );
or ( n5192 , n5189 , n5190 , n5191 );
and ( n5193 , n4965 , n4157 );
buf ( n5194 , n527 );
buf ( n5195 , n5194 );
and ( n5196 , n5195 , n4154 );
nor ( n5197 , n5193 , n5196 );
xnor ( n5198 , n5197 , n4152 );
and ( n5199 , n4176 , n4752 );
and ( n5200 , n4150 , n4579 );
nor ( n5201 , n5199 , n5200 );
xnor ( n5202 , n5201 , n4733 );
xor ( n5203 , n5198 , n5202 );
buf ( n5204 , n463 );
buf ( n5205 , n5204 );
xor ( n5206 , n5205 , n4975 );
not ( n5207 , n4976 );
and ( n5208 , n5206 , n5207 );
and ( n5209 , n4185 , n5208 );
and ( n5210 , n4165 , n4976 );
nor ( n5211 , n5209 , n5210 );
and ( n5212 , n4975 , n4730 );
not ( n5213 , n5212 );
and ( n5214 , n5205 , n5213 );
xnor ( n5215 , n5211 , n5214 );
xor ( n5216 , n5203 , n5215 );
xor ( n5217 , n5192 , n5216 );
and ( n5218 , n4568 , n4173 );
and ( n5219 , n4724 , n4171 );
nor ( n5220 , n5218 , n5219 );
xnor ( n5221 , n5220 , n4181 );
not ( n5222 , n4977 );
and ( n5223 , n5222 , n5214 );
xor ( n5224 , n5221 , n5223 );
and ( n5225 , n4968 , n4972 );
and ( n5226 , n4972 , n4977 );
and ( n5227 , n4968 , n4977 );
or ( n5228 , n5225 , n5226 , n5227 );
xor ( n5229 , n5224 , n5228 );
and ( n5230 , n4160 , n4262 );
and ( n5231 , n4243 , n4188 );
nor ( n5232 , n5230 , n5231 );
xnor ( n5233 , n5232 , n4252 );
xor ( n5234 , n5229 , n5233 );
xor ( n5235 , n5217 , n5234 );
and ( n5236 , n4962 , n4978 );
and ( n5237 , n4978 , n4990 );
and ( n5238 , n4962 , n4990 );
or ( n5239 , n5236 , n5237 , n5238 );
xor ( n5240 , n5235 , n5239 );
and ( n5241 , n4958 , n4991 );
and ( n5242 , n4992 , n4995 );
or ( n5243 , n5241 , n5242 );
xor ( n5244 , n5240 , n5243 );
buf ( n5245 , n5244 );
buf ( n5246 , n5245 );
buf ( n5247 , n5246 );
and ( n5248 , n5247 , n4232 );
nor ( n5249 , n5188 , n5248 );
xnor ( n5250 , n5249 , n4230 );
xor ( n5251 , n5187 , n5250 );
and ( n5252 , n4594 , n4319 );
and ( n5253 , n4770 , n4310 );
nor ( n5254 , n5252 , n5253 );
xnor ( n5255 , n5254 , n4315 );
and ( n5256 , n4228 , n4298 );
and ( n5257 , n4275 , n4287 );
nor ( n5258 , n5256 , n5257 );
xnor ( n5259 , n5258 , n4294 );
xor ( n5260 , n5255 , n5259 );
not ( n5261 , n5022 );
buf ( n5262 , n495 );
buf ( n5263 , n5262 );
and ( n5264 , n5020 , n4781 );
not ( n5265 , n5264 );
and ( n5266 , n5263 , n5265 );
and ( n5267 , n5261 , n5266 );
xor ( n5268 , n5263 , n5020 );
not ( n5269 , n5021 );
and ( n5270 , n5268 , n5269 );
and ( n5271 , n4282 , n5270 );
and ( n5272 , n4303 , n5021 );
nor ( n5273 , n5271 , n5272 );
xnor ( n5274 , n5273 , n5266 );
xor ( n5275 , n5267 , n5274 );
and ( n5276 , n5013 , n5017 );
and ( n5277 , n5017 , n5022 );
and ( n5278 , n5013 , n5022 );
or ( n5279 , n5276 , n5277 , n5278 );
xor ( n5280 , n5275 , n5279 );
and ( n5281 , n4329 , n4788 );
and ( n5282 , n4342 , n4611 );
nor ( n5283 , n5281 , n5282 );
xnor ( n5284 , n5283 , n4784 );
xor ( n5285 , n5280 , n5284 );
xor ( n5286 , n5260 , n5285 );
xor ( n5287 , n5251 , n5286 );
xor ( n5288 , n5183 , n5287 );
and ( n5289 , n5025 , n5029 );
and ( n5290 , n5030 , n5033 );
or ( n5291 , n5289 , n5290 );
xor ( n5292 , n5288 , n5291 );
buf ( n5293 , n5292 );
and ( n5294 , n5050 , n5054 );
and ( n5295 , n5054 , n5066 );
and ( n5296 , n5050 , n5066 );
or ( n5297 , n5294 , n5295 , n5296 );
and ( n5298 , n5042 , n4418 );
buf ( n5299 , n1784 );
buf ( n5300 , n5299 );
and ( n5301 , n5300 , n4415 );
nor ( n5302 , n5298 , n5301 );
xnor ( n5303 , n5302 , n4413 );
xor ( n5304 , n5297 , n5303 );
and ( n5305 , n5056 , n5060 );
and ( n5306 , n5060 , n5065 );
and ( n5307 , n5056 , n5065 );
or ( n5308 , n5305 , n5306 , n5307 );
and ( n5309 , n4631 , n4433 );
and ( n5310 , n4817 , n4431 );
nor ( n5311 , n5309 , n5310 );
xnor ( n5312 , n5311 , n4441 );
xor ( n5313 , n5308 , n5312 );
not ( n5314 , n5065 );
buf ( n5315 , n543 );
buf ( n5316 , n5315 );
and ( n5317 , n5063 , n4828 );
not ( n5318 , n5317 );
and ( n5319 , n5316 , n5318 );
and ( n5320 , n5314 , n5319 );
xor ( n5321 , n5316 , n5063 );
not ( n5322 , n5064 );
and ( n5323 , n5321 , n5322 );
and ( n5324 , n4386 , n5323 );
and ( n5325 , n4405 , n5064 );
nor ( n5326 , n5324 , n5325 );
xnor ( n5327 , n5326 , n5319 );
xor ( n5328 , n5320 , n5327 );
and ( n5329 , n4411 , n4402 );
and ( n5330 , n4421 , n4391 );
nor ( n5331 , n5329 , n5330 );
xnor ( n5332 , n5331 , n4398 );
xor ( n5333 , n5328 , n5332 );
and ( n5334 , n4427 , n4835 );
and ( n5335 , n4436 , n4648 );
nor ( n5336 , n5334 , n5335 );
xnor ( n5337 , n5336 , n4831 );
xor ( n5338 , n5333 , n5337 );
xor ( n5339 , n5313 , n5338 );
xor ( n5340 , n5304 , n5339 );
and ( n5341 , n5039 , n5045 );
and ( n5342 , n5045 , n5067 );
and ( n5343 , n5039 , n5067 );
or ( n5344 , n5341 , n5342 , n5343 );
xor ( n5345 , n5340 , n5344 );
and ( n5346 , n5068 , n5072 );
and ( n5347 , n5073 , n5076 );
or ( n5348 , n5346 , n5347 );
xor ( n5349 , n5345 , n5348 );
buf ( n5350 , n5349 );
not ( n5351 , n454 );
and ( n5352 , n5351 , n5293 );
and ( n5353 , n5350 , n454 );
or ( n5354 , n5352 , n5353 );
buf ( n5355 , n5354 );
buf ( n5356 , n5355 );
and ( n5357 , n5356 , n4505 );
xor ( n5358 , n5179 , n5357 );
and ( n5359 , n4663 , n5089 );
and ( n5360 , n4863 , n4866 );
xor ( n5361 , n5359 , n5360 );
xor ( n5362 , n5358 , n5361 );
xor ( n5363 , n5178 , n5362 );
and ( n5364 , n5095 , n5098 );
xor ( n5365 , n5363 , n5364 );
buf ( n5366 , n5365 );
not ( n5367 , n4509 );
and ( n5368 , n5367 , n5169 );
and ( n5369 , n5366 , n4509 );
or ( n5370 , n5368 , n5369 );
and ( n5371 , n5140 , n4524 );
and ( n5372 , n5124 , n5128 );
and ( n5373 , n5128 , n5133 );
and ( n5374 , n5124 , n5133 );
or ( n5375 , n5372 , n5373 , n5374 );
and ( n5376 , n5121 , n4530 );
buf ( n5377 , n499 );
buf ( n5378 , n515 );
xor ( n5379 , n5377 , n5378 );
and ( n5380 , n5111 , n5112 );
and ( n5381 , n5112 , n5117 );
and ( n5382 , n5111 , n5117 );
or ( n5383 , n5380 , n5381 , n5382 );
xor ( n5384 , n5379 , n5383 );
buf ( n5385 , n5384 );
buf ( n5386 , n5385 );
buf ( n5387 , n5386 );
and ( n5388 , n5387 , n4134 );
nor ( n5389 , n5376 , n5388 );
xnor ( n5390 , n5389 , n4527 );
and ( n5391 , n4683 , n4898 );
and ( n5392 , n4890 , n4689 );
nor ( n5393 , n5391 , n5392 );
xnor ( n5394 , n5393 , n4904 );
xor ( n5395 , n5390 , n5394 );
not ( n5396 , n5133 );
buf ( n5397 , n1121 );
buf ( n5398 , n5397 );
and ( n5399 , n5131 , n4895 );
not ( n5400 , n5399 );
and ( n5401 , n5398 , n5400 );
and ( n5402 , n5396 , n5401 );
xor ( n5403 , n5398 , n5131 );
not ( n5404 , n5132 );
and ( n5405 , n5403 , n5404 );
and ( n5406 , n4132 , n5405 );
and ( n5407 , n4539 , n5132 );
nor ( n5408 , n5406 , n5407 );
xnor ( n5409 , n5408 , n5401 );
xor ( n5410 , n5402 , n5409 );
xor ( n5411 , n5395 , n5410 );
xor ( n5412 , n5375 , n5411 );
and ( n5413 , n5109 , n5134 );
and ( n5414 , n5135 , n5136 );
or ( n5415 , n5413 , n5414 );
xor ( n5416 , n5412 , n5415 );
buf ( n5417 , n5416 );
buf ( n5418 , n5417 );
buf ( n5419 , n5418 );
and ( n5420 , n5419 , n4145 );
nor ( n5421 , n5371 , n5420 );
xnor ( n5422 , n5421 , n4521 );
not ( n5423 , n5162 );
buf ( n5424 , n531 );
buf ( n5425 , n547 );
xor ( n5426 , n5424 , n5425 );
and ( n5427 , n5150 , n5151 );
and ( n5428 , n5151 , n5156 );
and ( n5429 , n5150 , n5156 );
or ( n5430 , n5427 , n5428 , n5429 );
xor ( n5431 , n5426 , n5430 );
buf ( n5432 , n5431 );
buf ( n5433 , n5432 );
buf ( n5434 , n5433 );
and ( n5435 , n5160 , n4931 );
not ( n5436 , n5435 );
and ( n5437 , n5434 , n5436 );
and ( n5438 , n5423 , n5437 );
xor ( n5439 , n5434 , n5160 );
not ( n5440 , n5161 );
and ( n5441 , n5439 , n5440 );
and ( n5442 , n4139 , n5441 );
and ( n5443 , n4548 , n5161 );
nor ( n5444 , n5442 , n5443 );
xnor ( n5445 , n5444 , n5437 );
xor ( n5446 , n5438 , n5445 );
and ( n5447 , n5144 , n5148 );
and ( n5448 , n5148 , n5162 );
and ( n5449 , n5144 , n5162 );
or ( n5450 , n5447 , n5448 , n5449 );
xor ( n5451 , n5446 , n5450 );
and ( n5452 , n4696 , n4938 );
and ( n5453 , n4916 , n4711 );
nor ( n5454 , n5452 , n5453 );
xnor ( n5455 , n5454 , n4934 );
xor ( n5456 , n5451 , n5455 );
xor ( n5457 , n5422 , n5456 );
and ( n5458 , n5143 , n5163 );
and ( n5459 , n5164 , n5167 );
or ( n5460 , n5458 , n5459 );
xor ( n5461 , n5457 , n5460 );
buf ( n5462 , n5461 );
and ( n5463 , n5179 , n5357 );
and ( n5464 , n5357 , n5361 );
and ( n5465 , n5179 , n5361 );
or ( n5466 , n5463 , n5464 , n5465 );
and ( n5467 , n4863 , n5089 );
and ( n5468 , n5084 , n4866 );
xor ( n5469 , n5467 , n5468 );
and ( n5470 , n5356 , n4557 );
xor ( n5471 , n5469 , n5470 );
and ( n5472 , n5187 , n5250 );
and ( n5473 , n5250 , n5286 );
and ( n5474 , n5187 , n5286 );
or ( n5475 , n5472 , n5473 , n5474 );
and ( n5476 , n5255 , n5259 );
and ( n5477 , n5259 , n5285 );
and ( n5478 , n5255 , n5285 );
or ( n5479 , n5476 , n5477 , n5478 );
and ( n5480 , n5247 , n4235 );
and ( n5481 , n5224 , n5228 );
and ( n5482 , n5228 , n5233 );
and ( n5483 , n5224 , n5233 );
or ( n5484 , n5481 , n5482 , n5483 );
and ( n5485 , n5195 , n4157 );
buf ( n5486 , n526 );
buf ( n5487 , n5486 );
and ( n5488 , n5487 , n4154 );
nor ( n5489 , n5485 , n5488 );
xnor ( n5490 , n5489 , n4152 );
and ( n5491 , n4243 , n4262 );
and ( n5492 , n4568 , n4188 );
nor ( n5493 , n5491 , n5492 );
xnor ( n5494 , n5493 , n4252 );
xor ( n5495 , n5490 , n5494 );
and ( n5496 , n4165 , n5208 );
and ( n5497 , n4176 , n4976 );
nor ( n5498 , n5496 , n5497 );
xnor ( n5499 , n5498 , n5214 );
xor ( n5500 , n5495 , n5499 );
xor ( n5501 , n5484 , n5500 );
and ( n5502 , n5198 , n5202 );
and ( n5503 , n5202 , n5215 );
and ( n5504 , n5198 , n5215 );
or ( n5505 , n5502 , n5503 , n5504 );
and ( n5506 , n5221 , n5223 );
xor ( n5507 , n5505 , n5506 );
and ( n5508 , n4724 , n4173 );
and ( n5509 , n4965 , n4171 );
nor ( n5510 , n5508 , n5509 );
xnor ( n5511 , n5510 , n4181 );
and ( n5512 , n4150 , n4752 );
and ( n5513 , n4160 , n4579 );
nor ( n5514 , n5512 , n5513 );
xnor ( n5515 , n5514 , n4733 );
xor ( n5516 , n5511 , n5515 );
buf ( n5517 , n462 );
buf ( n5518 , n5517 );
xor ( n5519 , n5518 , n5205 );
and ( n5520 , n4185 , n5519 );
xor ( n5521 , n5516 , n5520 );
xor ( n5522 , n5507 , n5521 );
xor ( n5523 , n5501 , n5522 );
and ( n5524 , n5192 , n5216 );
and ( n5525 , n5216 , n5234 );
and ( n5526 , n5192 , n5234 );
or ( n5527 , n5524 , n5525 , n5526 );
xor ( n5528 , n5523 , n5527 );
and ( n5529 , n5235 , n5239 );
and ( n5530 , n5240 , n5243 );
or ( n5531 , n5529 , n5530 );
xor ( n5532 , n5528 , n5531 );
buf ( n5533 , n5532 );
buf ( n5534 , n5533 );
buf ( n5535 , n5534 );
and ( n5536 , n5535 , n4232 );
nor ( n5537 , n5480 , n5536 );
xnor ( n5538 , n5537 , n4230 );
xor ( n5539 , n5479 , n5538 );
and ( n5540 , n4770 , n4319 );
and ( n5541 , n4999 , n4310 );
nor ( n5542 , n5540 , n5541 );
xnor ( n5543 , n5542 , n4315 );
and ( n5544 , n4275 , n4298 );
and ( n5545 , n4594 , n4287 );
nor ( n5546 , n5544 , n5545 );
xnor ( n5547 , n5546 , n4294 );
xor ( n5548 , n5543 , n5547 );
and ( n5549 , n5275 , n5279 );
and ( n5550 , n5279 , n5284 );
and ( n5551 , n5275 , n5284 );
or ( n5552 , n5549 , n5550 , n5551 );
and ( n5553 , n4342 , n4788 );
and ( n5554 , n4228 , n4611 );
nor ( n5555 , n5553 , n5554 );
xnor ( n5556 , n5555 , n4784 );
xor ( n5557 , n5552 , n5556 );
and ( n5558 , n5267 , n5274 );
and ( n5559 , n4303 , n5270 );
and ( n5560 , n4329 , n5021 );
nor ( n5561 , n5559 , n5560 );
xnor ( n5562 , n5561 , n5266 );
xor ( n5563 , n5558 , n5562 );
buf ( n5564 , n494 );
buf ( n5565 , n5564 );
xor ( n5566 , n5565 , n5263 );
and ( n5567 , n4282 , n5566 );
xor ( n5568 , n5563 , n5567 );
xor ( n5569 , n5557 , n5568 );
xor ( n5570 , n5548 , n5569 );
xor ( n5571 , n5539 , n5570 );
xor ( n5572 , n5475 , n5571 );
and ( n5573 , n5183 , n5287 );
and ( n5574 , n5288 , n5291 );
or ( n5575 , n5573 , n5574 );
xor ( n5576 , n5572 , n5575 );
buf ( n5577 , n5576 );
and ( n5578 , n5308 , n5312 );
and ( n5579 , n5312 , n5338 );
and ( n5580 , n5308 , n5338 );
or ( n5581 , n5578 , n5579 , n5580 );
and ( n5582 , n5328 , n5332 );
and ( n5583 , n5332 , n5337 );
and ( n5584 , n5328 , n5337 );
or ( n5585 , n5582 , n5583 , n5584 );
and ( n5586 , n5300 , n4418 );
buf ( n5587 , n1954 );
buf ( n5588 , n5587 );
and ( n5589 , n5588 , n4415 );
nor ( n5590 , n5586 , n5589 );
xnor ( n5591 , n5590 , n4413 );
xor ( n5592 , n5585 , n5591 );
and ( n5593 , n4817 , n4433 );
and ( n5594 , n5042 , n4431 );
nor ( n5595 , n5593 , n5594 );
xnor ( n5596 , n5595 , n4441 );
xor ( n5597 , n5592 , n5596 );
xor ( n5598 , n5581 , n5597 );
and ( n5599 , n4421 , n4402 );
and ( n5600 , n4631 , n4391 );
nor ( n5601 , n5599 , n5600 );
xnor ( n5602 , n5601 , n4398 );
and ( n5603 , n4436 , n4835 );
and ( n5604 , n4411 , n4648 );
nor ( n5605 , n5603 , n5604 );
xnor ( n5606 , n5605 , n4831 );
xor ( n5607 , n5602 , n5606 );
and ( n5608 , n5320 , n5327 );
and ( n5609 , n4405 , n5323 );
and ( n5610 , n4427 , n5064 );
nor ( n5611 , n5609 , n5610 );
xnor ( n5612 , n5611 , n5319 );
xor ( n5613 , n5608 , n5612 );
buf ( n5614 , n542 );
buf ( n5615 , n5614 );
xor ( n5616 , n5615 , n5316 );
and ( n5617 , n4386 , n5616 );
xor ( n5618 , n5613 , n5617 );
xor ( n5619 , n5607 , n5618 );
xor ( n5620 , n5598 , n5619 );
and ( n5621 , n5297 , n5303 );
and ( n5622 , n5303 , n5339 );
and ( n5623 , n5297 , n5339 );
or ( n5624 , n5621 , n5622 , n5623 );
xor ( n5625 , n5620 , n5624 );
and ( n5626 , n5340 , n5344 );
and ( n5627 , n5345 , n5348 );
or ( n5628 , n5626 , n5627 );
xor ( n5629 , n5625 , n5628 );
buf ( n5630 , n5629 );
not ( n5631 , n454 );
and ( n5632 , n5631 , n5577 );
and ( n5633 , n5630 , n454 );
or ( n5634 , n5632 , n5633 );
buf ( n5635 , n5634 );
buf ( n5636 , n5635 );
and ( n5637 , n5636 , n4505 );
not ( n5638 , n5637 );
xor ( n5639 , n5471 , n5638 );
and ( n5640 , n5359 , n5360 );
xor ( n5641 , n5639 , n5640 );
xor ( n5642 , n5466 , n5641 );
and ( n5643 , n5173 , n5177 );
and ( n5644 , n5177 , n5362 );
and ( n5645 , n5173 , n5362 );
or ( n5646 , n5643 , n5644 , n5645 );
xor ( n5647 , n5642 , n5646 );
not ( n5648 , n5647 );
and ( n5649 , n5363 , n5364 );
xor ( n5650 , n5648 , n5649 );
buf ( n5651 , n5650 );
not ( n5652 , n4509 );
and ( n5653 , n5652 , n5462 );
and ( n5654 , n5651 , n4509 );
or ( n5655 , n5653 , n5654 );
and ( n5656 , n5419 , n4524 );
and ( n5657 , n5390 , n5394 );
and ( n5658 , n5394 , n5410 );
and ( n5659 , n5390 , n5410 );
or ( n5660 , n5657 , n5658 , n5659 );
and ( n5661 , n5387 , n4530 );
buf ( n5662 , n498 );
buf ( n5663 , n514 );
xor ( n5664 , n5662 , n5663 );
and ( n5665 , n5377 , n5378 );
and ( n5666 , n5378 , n5383 );
and ( n5667 , n5377 , n5383 );
or ( n5668 , n5665 , n5666 , n5667 );
xor ( n5669 , n5664 , n5668 );
buf ( n5670 , n5669 );
buf ( n5671 , n5670 );
buf ( n5672 , n5671 );
and ( n5673 , n5672 , n4134 );
nor ( n5674 , n5661 , n5673 );
xnor ( n5675 , n5674 , n4527 );
and ( n5676 , n4890 , n4898 );
and ( n5677 , n5121 , n4689 );
nor ( n5678 , n5676 , n5677 );
xnor ( n5679 , n5678 , n4904 );
xor ( n5680 , n5675 , n5679 );
and ( n5681 , n5402 , n5409 );
and ( n5682 , n4539 , n5405 );
and ( n5683 , n4683 , n5132 );
nor ( n5684 , n5682 , n5683 );
xnor ( n5685 , n5684 , n5401 );
xor ( n5686 , n5681 , n5685 );
buf ( n5687 , n1211 );
buf ( n5688 , n5687 );
xor ( n5689 , n5688 , n5398 );
and ( n5690 , n4132 , n5689 );
xor ( n5691 , n5686 , n5690 );
xor ( n5692 , n5680 , n5691 );
xor ( n5693 , n5660 , n5692 );
and ( n5694 , n5375 , n5411 );
and ( n5695 , n5412 , n5415 );
or ( n5696 , n5694 , n5695 );
xor ( n5697 , n5693 , n5696 );
buf ( n5698 , n5697 );
buf ( n5699 , n5698 );
buf ( n5700 , n5699 );
and ( n5701 , n5700 , n4145 );
nor ( n5702 , n5656 , n5701 );
xnor ( n5703 , n5702 , n4521 );
and ( n5704 , n5446 , n5450 );
and ( n5705 , n5450 , n5455 );
and ( n5706 , n5446 , n5455 );
or ( n5707 , n5704 , n5705 , n5706 );
and ( n5708 , n4916 , n4938 );
and ( n5709 , n5140 , n4711 );
nor ( n5710 , n5708 , n5709 );
xnor ( n5711 , n5710 , n4934 );
xor ( n5712 , n5707 , n5711 );
and ( n5713 , n5438 , n5445 );
and ( n5714 , n4548 , n5441 );
and ( n5715 , n4696 , n5161 );
nor ( n5716 , n5714 , n5715 );
xnor ( n5717 , n5716 , n5437 );
xor ( n5718 , n5713 , n5717 );
buf ( n5719 , n530 );
buf ( n5720 , n546 );
xor ( n5721 , n5719 , n5720 );
and ( n5722 , n5424 , n5425 );
and ( n5723 , n5425 , n5430 );
and ( n5724 , n5424 , n5430 );
or ( n5725 , n5722 , n5723 , n5724 );
xor ( n5726 , n5721 , n5725 );
buf ( n5727 , n5726 );
buf ( n5728 , n5727 );
buf ( n5729 , n5728 );
xor ( n5730 , n5729 , n5434 );
and ( n5731 , n4139 , n5730 );
xor ( n5732 , n5718 , n5731 );
xor ( n5733 , n5712 , n5732 );
xor ( n5734 , n5703 , n5733 );
and ( n5735 , n5422 , n5456 );
and ( n5736 , n5457 , n5460 );
or ( n5737 , n5735 , n5736 );
xor ( n5738 , n5734 , n5737 );
buf ( n5739 , n5738 );
buf ( n5740 , n5637 );
and ( n5741 , n5467 , n5468 );
and ( n5742 , n5468 , n5470 );
and ( n5743 , n5467 , n5470 );
or ( n5744 , n5741 , n5742 , n5743 );
and ( n5745 , n5543 , n5547 );
and ( n5746 , n5547 , n5569 );
and ( n5747 , n5543 , n5569 );
or ( n5748 , n5745 , n5746 , n5747 );
and ( n5749 , n5535 , n4235 );
and ( n5750 , n5505 , n5506 );
and ( n5751 , n5506 , n5521 );
and ( n5752 , n5505 , n5521 );
or ( n5753 , n5750 , n5751 , n5752 );
and ( n5754 , n4965 , n4173 );
and ( n5755 , n5195 , n4171 );
nor ( n5756 , n5754 , n5755 );
xnor ( n5757 , n5756 , n4181 );
not ( n5758 , n5520 );
buf ( n5759 , n461 );
buf ( n5760 , n5759 );
and ( n5761 , n5518 , n5205 );
not ( n5762 , n5761 );
and ( n5763 , n5760 , n5762 );
and ( n5764 , n5758 , n5763 );
xor ( n5765 , n5757 , n5764 );
and ( n5766 , n4568 , n4262 );
and ( n5767 , n4724 , n4188 );
nor ( n5768 , n5766 , n5767 );
xnor ( n5769 , n5768 , n4252 );
xor ( n5770 , n5765 , n5769 );
xor ( n5771 , n5760 , n5518 );
not ( n5772 , n5519 );
and ( n5773 , n5771 , n5772 );
and ( n5774 , n4185 , n5773 );
and ( n5775 , n4165 , n5519 );
nor ( n5776 , n5774 , n5775 );
xnor ( n5777 , n5776 , n5763 );
xor ( n5778 , n5770 , n5777 );
xor ( n5779 , n5753 , n5778 );
and ( n5780 , n5490 , n5494 );
and ( n5781 , n5494 , n5499 );
and ( n5782 , n5490 , n5499 );
or ( n5783 , n5780 , n5781 , n5782 );
and ( n5784 , n5511 , n5515 );
and ( n5785 , n5515 , n5520 );
and ( n5786 , n5511 , n5520 );
or ( n5787 , n5784 , n5785 , n5786 );
xor ( n5788 , n5783 , n5787 );
and ( n5789 , n5487 , n4157 );
buf ( n5790 , n525 );
buf ( n5791 , n5790 );
and ( n5792 , n5791 , n4154 );
nor ( n5793 , n5789 , n5792 );
xnor ( n5794 , n5793 , n4152 );
and ( n5795 , n4160 , n4752 );
and ( n5796 , n4243 , n4579 );
nor ( n5797 , n5795 , n5796 );
xnor ( n5798 , n5797 , n4733 );
xor ( n5799 , n5794 , n5798 );
and ( n5800 , n4176 , n5208 );
and ( n5801 , n4150 , n4976 );
nor ( n5802 , n5800 , n5801 );
xnor ( n5803 , n5802 , n5214 );
xor ( n5804 , n5799 , n5803 );
xor ( n5805 , n5788 , n5804 );
xor ( n5806 , n5779 , n5805 );
and ( n5807 , n5484 , n5500 );
and ( n5808 , n5500 , n5522 );
and ( n5809 , n5484 , n5522 );
or ( n5810 , n5807 , n5808 , n5809 );
xor ( n5811 , n5806 , n5810 );
and ( n5812 , n5523 , n5527 );
and ( n5813 , n5528 , n5531 );
or ( n5814 , n5812 , n5813 );
xor ( n5815 , n5811 , n5814 );
buf ( n5816 , n5815 );
buf ( n5817 , n5816 );
buf ( n5818 , n5817 );
and ( n5819 , n5818 , n4232 );
nor ( n5820 , n5749 , n5819 );
xnor ( n5821 , n5820 , n4230 );
xor ( n5822 , n5748 , n5821 );
and ( n5823 , n5552 , n5556 );
and ( n5824 , n5556 , n5568 );
and ( n5825 , n5552 , n5568 );
or ( n5826 , n5823 , n5824 , n5825 );
and ( n5827 , n4999 , n4319 );
and ( n5828 , n5247 , n4310 );
nor ( n5829 , n5827 , n5828 );
xnor ( n5830 , n5829 , n4315 );
xor ( n5831 , n5826 , n5830 );
and ( n5832 , n4594 , n4298 );
and ( n5833 , n4770 , n4287 );
nor ( n5834 , n5832 , n5833 );
xnor ( n5835 , n5834 , n4294 );
and ( n5836 , n4228 , n4788 );
and ( n5837 , n4275 , n4611 );
nor ( n5838 , n5836 , n5837 );
xnor ( n5839 , n5838 , n4784 );
xor ( n5840 , n5835 , n5839 );
not ( n5841 , n5567 );
buf ( n5842 , n493 );
buf ( n5843 , n5842 );
and ( n5844 , n5565 , n5263 );
not ( n5845 , n5844 );
and ( n5846 , n5843 , n5845 );
and ( n5847 , n5841 , n5846 );
xor ( n5848 , n5843 , n5565 );
not ( n5849 , n5566 );
and ( n5850 , n5848 , n5849 );
and ( n5851 , n4282 , n5850 );
and ( n5852 , n4303 , n5566 );
nor ( n5853 , n5851 , n5852 );
xnor ( n5854 , n5853 , n5846 );
xor ( n5855 , n5847 , n5854 );
and ( n5856 , n5558 , n5562 );
and ( n5857 , n5562 , n5567 );
and ( n5858 , n5558 , n5567 );
or ( n5859 , n5856 , n5857 , n5858 );
xor ( n5860 , n5855 , n5859 );
and ( n5861 , n4329 , n5270 );
and ( n5862 , n4342 , n5021 );
nor ( n5863 , n5861 , n5862 );
xnor ( n5864 , n5863 , n5266 );
xor ( n5865 , n5860 , n5864 );
xor ( n5866 , n5840 , n5865 );
xor ( n5867 , n5831 , n5866 );
xor ( n5868 , n5822 , n5867 );
and ( n5869 , n5479 , n5538 );
and ( n5870 , n5538 , n5570 );
and ( n5871 , n5479 , n5570 );
or ( n5872 , n5869 , n5870 , n5871 );
xor ( n5873 , n5868 , n5872 );
and ( n5874 , n5475 , n5571 );
and ( n5875 , n5572 , n5575 );
or ( n5876 , n5874 , n5875 );
xor ( n5877 , n5873 , n5876 );
buf ( n5878 , n5877 );
and ( n5879 , n5581 , n5597 );
and ( n5880 , n5597 , n5619 );
and ( n5881 , n5581 , n5619 );
or ( n5882 , n5879 , n5880 , n5881 );
and ( n5883 , n5585 , n5591 );
and ( n5884 , n5591 , n5596 );
and ( n5885 , n5585 , n5596 );
or ( n5886 , n5883 , n5884 , n5885 );
and ( n5887 , n5602 , n5606 );
and ( n5888 , n5606 , n5618 );
and ( n5889 , n5602 , n5618 );
or ( n5890 , n5887 , n5888 , n5889 );
and ( n5891 , n5588 , n4418 );
buf ( n5892 , n2116 );
buf ( n5893 , n5892 );
and ( n5894 , n5893 , n4415 );
nor ( n5895 , n5891 , n5894 );
xnor ( n5896 , n5895 , n4413 );
xor ( n5897 , n5890 , n5896 );
and ( n5898 , n5042 , n4433 );
and ( n5899 , n5300 , n4431 );
nor ( n5900 , n5898 , n5899 );
xnor ( n5901 , n5900 , n4441 );
xor ( n5902 , n5897 , n5901 );
xor ( n5903 , n5886 , n5902 );
and ( n5904 , n4631 , n4402 );
and ( n5905 , n4817 , n4391 );
nor ( n5906 , n5904 , n5905 );
xnor ( n5907 , n5906 , n4398 );
and ( n5908 , n4411 , n4835 );
and ( n5909 , n4421 , n4648 );
nor ( n5910 , n5908 , n5909 );
xnor ( n5911 , n5910 , n4831 );
xor ( n5912 , n5907 , n5911 );
not ( n5913 , n5617 );
buf ( n5914 , n541 );
buf ( n5915 , n5914 );
and ( n5916 , n5615 , n5316 );
not ( n5917 , n5916 );
and ( n5918 , n5915 , n5917 );
and ( n5919 , n5913 , n5918 );
xor ( n5920 , n5915 , n5615 );
not ( n5921 , n5616 );
and ( n5922 , n5920 , n5921 );
and ( n5923 , n4386 , n5922 );
and ( n5924 , n4405 , n5616 );
nor ( n5925 , n5923 , n5924 );
xnor ( n5926 , n5925 , n5918 );
xor ( n5927 , n5919 , n5926 );
and ( n5928 , n5608 , n5612 );
and ( n5929 , n5612 , n5617 );
and ( n5930 , n5608 , n5617 );
or ( n5931 , n5928 , n5929 , n5930 );
xor ( n5932 , n5927 , n5931 );
and ( n5933 , n4427 , n5323 );
and ( n5934 , n4436 , n5064 );
nor ( n5935 , n5933 , n5934 );
xnor ( n5936 , n5935 , n5319 );
xor ( n5937 , n5932 , n5936 );
xor ( n5938 , n5912 , n5937 );
xor ( n5939 , n5903 , n5938 );
xor ( n5940 , n5882 , n5939 );
and ( n5941 , n5620 , n5624 );
and ( n5942 , n5625 , n5628 );
or ( n5943 , n5941 , n5942 );
xor ( n5944 , n5940 , n5943 );
buf ( n5945 , n5944 );
not ( n5946 , n454 );
and ( n5947 , n5946 , n5878 );
and ( n5948 , n5945 , n454 );
or ( n5949 , n5947 , n5948 );
buf ( n5950 , n5949 );
buf ( n5951 , n5950 );
and ( n5952 , n5951 , n4505 );
xor ( n5953 , n5744 , n5952 );
and ( n5954 , n5084 , n5089 );
and ( n5955 , n5356 , n4866 );
xor ( n5956 , n5954 , n5955 );
and ( n5957 , n5636 , n4557 );
xor ( n5958 , n5956 , n5957 );
xor ( n5959 , n5953 , n5958 );
xor ( n5960 , n5740 , n5959 );
and ( n5961 , n5471 , n5638 );
and ( n5962 , n5638 , n5640 );
and ( n5963 , n5471 , n5640 );
or ( n5964 , n5961 , n5962 , n5963 );
xor ( n5965 , n5960 , n5964 );
and ( n5966 , n5466 , n5641 );
and ( n5967 , n5641 , n5646 );
and ( n5968 , n5466 , n5646 );
or ( n5969 , n5966 , n5967 , n5968 );
xnor ( n5970 , n5965 , n5969 );
and ( n5971 , n5648 , n5649 );
or ( n5972 , n5647 , n5971 );
xor ( n5973 , n5970 , n5972 );
buf ( n5974 , n5973 );
not ( n5975 , n4509 );
and ( n5976 , n5975 , n5739 );
and ( n5977 , n5974 , n4509 );
or ( n5978 , n5976 , n5977 );
and ( n5979 , n5700 , n4524 );
and ( n5980 , n5675 , n5679 );
and ( n5981 , n5679 , n5691 );
and ( n5982 , n5675 , n5691 );
or ( n5983 , n5980 , n5981 , n5982 );
and ( n5984 , n5672 , n4530 );
buf ( n5985 , n497 );
buf ( n5986 , n513 );
xor ( n5987 , n5985 , n5986 );
and ( n5988 , n5662 , n5663 );
and ( n5989 , n5663 , n5668 );
and ( n5990 , n5662 , n5668 );
or ( n5991 , n5988 , n5989 , n5990 );
xor ( n5992 , n5987 , n5991 );
buf ( n5993 , n5992 );
buf ( n5994 , n5993 );
buf ( n5995 , n5994 );
and ( n5996 , n5995 , n4134 );
nor ( n5997 , n5984 , n5996 );
xnor ( n5998 , n5997 , n4527 );
not ( n5999 , n5690 );
buf ( n6000 , n1321 );
buf ( n6001 , n6000 );
and ( n6002 , n5688 , n5398 );
not ( n6003 , n6002 );
and ( n6004 , n6001 , n6003 );
and ( n6005 , n5999 , n6004 );
xor ( n6006 , n6001 , n5688 );
not ( n6007 , n5689 );
and ( n6008 , n6006 , n6007 );
and ( n6009 , n4132 , n6008 );
and ( n6010 , n4539 , n5689 );
nor ( n6011 , n6009 , n6010 );
xnor ( n6012 , n6011 , n6004 );
xor ( n6013 , n6005 , n6012 );
and ( n6014 , n5121 , n4898 );
and ( n6015 , n5387 , n4689 );
nor ( n6016 , n6014 , n6015 );
xnor ( n6017 , n6016 , n4904 );
xor ( n6018 , n6013 , n6017 );
and ( n6019 , n4683 , n5405 );
and ( n6020 , n4890 , n5132 );
nor ( n6021 , n6019 , n6020 );
xnor ( n6022 , n6021 , n5401 );
xor ( n6023 , n6018 , n6022 );
xor ( n6024 , n5998 , n6023 );
and ( n6025 , n5681 , n5685 );
and ( n6026 , n5685 , n5690 );
and ( n6027 , n5681 , n5690 );
or ( n6028 , n6025 , n6026 , n6027 );
xor ( n6029 , n6024 , n6028 );
xor ( n6030 , n5983 , n6029 );
and ( n6031 , n5660 , n5692 );
and ( n6032 , n5693 , n5696 );
or ( n6033 , n6031 , n6032 );
xor ( n6034 , n6030 , n6033 );
buf ( n6035 , n6034 );
buf ( n6036 , n6035 );
buf ( n6037 , n6036 );
and ( n6038 , n6037 , n4145 );
nor ( n6039 , n5979 , n6038 );
xnor ( n6040 , n6039 , n4521 );
and ( n6041 , n5707 , n5711 );
and ( n6042 , n5711 , n5732 );
and ( n6043 , n5707 , n5732 );
or ( n6044 , n6041 , n6042 , n6043 );
and ( n6045 , n5140 , n4938 );
and ( n6046 , n5419 , n4711 );
nor ( n6047 , n6045 , n6046 );
xnor ( n6048 , n6047 , n4934 );
xor ( n6049 , n6044 , n6048 );
not ( n6050 , n5731 );
buf ( n6051 , n529 );
buf ( n6052 , n545 );
xor ( n6053 , n6051 , n6052 );
and ( n6054 , n5719 , n5720 );
and ( n6055 , n5720 , n5725 );
and ( n6056 , n5719 , n5725 );
or ( n6057 , n6054 , n6055 , n6056 );
xor ( n6058 , n6053 , n6057 );
buf ( n6059 , n6058 );
buf ( n6060 , n6059 );
buf ( n6061 , n6060 );
and ( n6062 , n5729 , n5434 );
not ( n6063 , n6062 );
and ( n6064 , n6061 , n6063 );
and ( n6065 , n6050 , n6064 );
xor ( n6066 , n6061 , n5729 );
not ( n6067 , n5730 );
and ( n6068 , n6066 , n6067 );
and ( n6069 , n4139 , n6068 );
and ( n6070 , n4548 , n5730 );
nor ( n6071 , n6069 , n6070 );
xnor ( n6072 , n6071 , n6064 );
xor ( n6073 , n6065 , n6072 );
and ( n6074 , n5713 , n5717 );
and ( n6075 , n5717 , n5731 );
and ( n6076 , n5713 , n5731 );
or ( n6077 , n6074 , n6075 , n6076 );
xor ( n6078 , n6073 , n6077 );
and ( n6079 , n4696 , n5441 );
and ( n6080 , n4916 , n5161 );
nor ( n6081 , n6079 , n6080 );
xnor ( n6082 , n6081 , n5437 );
xor ( n6083 , n6078 , n6082 );
xor ( n6084 , n6049 , n6083 );
xor ( n6085 , n6040 , n6084 );
and ( n6086 , n5703 , n5733 );
and ( n6087 , n5734 , n5737 );
or ( n6088 , n6086 , n6087 );
xor ( n6089 , n6085 , n6088 );
buf ( n6090 , n6089 );
and ( n6091 , n5954 , n5955 );
and ( n6092 , n5955 , n5957 );
and ( n6093 , n5954 , n5957 );
or ( n6094 , n6091 , n6092 , n6093 );
and ( n6095 , n5826 , n5830 );
and ( n6096 , n5830 , n5866 );
and ( n6097 , n5826 , n5866 );
or ( n6098 , n6095 , n6096 , n6097 );
and ( n6099 , n5835 , n5839 );
and ( n6100 , n5839 , n5865 );
and ( n6101 , n5835 , n5865 );
or ( n6102 , n6099 , n6100 , n6101 );
and ( n6103 , n5818 , n4235 );
and ( n6104 , n5195 , n4173 );
and ( n6105 , n5487 , n4171 );
nor ( n6106 , n6104 , n6105 );
xnor ( n6107 , n6106 , n4181 );
and ( n6108 , n4243 , n4752 );
and ( n6109 , n4568 , n4579 );
nor ( n6110 , n6108 , n6109 );
xnor ( n6111 , n6110 , n4733 );
xor ( n6112 , n6107 , n6111 );
buf ( n6113 , n460 );
buf ( n6114 , n6113 );
xor ( n6115 , n6114 , n5760 );
and ( n6116 , n4185 , n6115 );
xor ( n6117 , n6112 , n6116 );
and ( n6118 , n5791 , n4157 );
buf ( n6119 , n524 );
buf ( n6120 , n6119 );
and ( n6121 , n6120 , n4154 );
nor ( n6122 , n6118 , n6121 );
xnor ( n6123 , n6122 , n4152 );
and ( n6124 , n4150 , n5208 );
and ( n6125 , n4160 , n4976 );
nor ( n6126 , n6124 , n6125 );
xnor ( n6127 , n6126 , n5214 );
xor ( n6128 , n6123 , n6127 );
and ( n6129 , n4165 , n5773 );
and ( n6130 , n4176 , n5519 );
nor ( n6131 , n6129 , n6130 );
xnor ( n6132 , n6131 , n5763 );
xor ( n6133 , n6128 , n6132 );
xor ( n6134 , n6117 , n6133 );
and ( n6135 , n5794 , n5798 );
and ( n6136 , n5798 , n5803 );
and ( n6137 , n5794 , n5803 );
or ( n6138 , n6135 , n6136 , n6137 );
and ( n6139 , n5757 , n5764 );
xor ( n6140 , n6138 , n6139 );
and ( n6141 , n4724 , n4262 );
and ( n6142 , n4965 , n4188 );
nor ( n6143 , n6141 , n6142 );
xnor ( n6144 , n6143 , n4252 );
xor ( n6145 , n6140 , n6144 );
xor ( n6146 , n6134 , n6145 );
and ( n6147 , n5765 , n5769 );
and ( n6148 , n5769 , n5777 );
and ( n6149 , n5765 , n5777 );
or ( n6150 , n6147 , n6148 , n6149 );
and ( n6151 , n5783 , n5787 );
and ( n6152 , n5787 , n5804 );
and ( n6153 , n5783 , n5804 );
or ( n6154 , n6151 , n6152 , n6153 );
xor ( n6155 , n6150 , n6154 );
and ( n6156 , n5753 , n5778 );
and ( n6157 , n5778 , n5805 );
and ( n6158 , n5753 , n5805 );
or ( n6159 , n6156 , n6157 , n6158 );
xor ( n6160 , n6155 , n6159 );
xor ( n6161 , n6146 , n6160 );
and ( n6162 , n5806 , n5810 );
and ( n6163 , n5811 , n5814 );
or ( n6164 , n6162 , n6163 );
xor ( n6165 , n6161 , n6164 );
buf ( n6166 , n6165 );
buf ( n6167 , n6166 );
buf ( n6168 , n6167 );
and ( n6169 , n6168 , n4232 );
nor ( n6170 , n6103 , n6169 );
xnor ( n6171 , n6170 , n4230 );
xor ( n6172 , n6102 , n6171 );
and ( n6173 , n5247 , n4319 );
and ( n6174 , n5535 , n4310 );
nor ( n6175 , n6173 , n6174 );
xnor ( n6176 , n6175 , n4315 );
xor ( n6177 , n6172 , n6176 );
xor ( n6178 , n6098 , n6177 );
and ( n6179 , n4770 , n4298 );
and ( n6180 , n4999 , n4287 );
nor ( n6181 , n6179 , n6180 );
xnor ( n6182 , n6181 , n4294 );
and ( n6183 , n4275 , n4788 );
and ( n6184 , n4594 , n4611 );
nor ( n6185 , n6183 , n6184 );
xnor ( n6186 , n6185 , n4784 );
xor ( n6187 , n6182 , n6186 );
and ( n6188 , n5855 , n5859 );
and ( n6189 , n5859 , n5864 );
and ( n6190 , n5855 , n5864 );
or ( n6191 , n6188 , n6189 , n6190 );
and ( n6192 , n4342 , n5270 );
and ( n6193 , n4228 , n5021 );
nor ( n6194 , n6192 , n6193 );
xnor ( n6195 , n6194 , n5266 );
xor ( n6196 , n6191 , n6195 );
and ( n6197 , n5847 , n5854 );
and ( n6198 , n4303 , n5850 );
and ( n6199 , n4329 , n5566 );
nor ( n6200 , n6198 , n6199 );
xnor ( n6201 , n6200 , n5846 );
xor ( n6202 , n6197 , n6201 );
buf ( n6203 , n492 );
buf ( n6204 , n6203 );
xor ( n6205 , n6204 , n5843 );
and ( n6206 , n4282 , n6205 );
xor ( n6207 , n6202 , n6206 );
xor ( n6208 , n6196 , n6207 );
xor ( n6209 , n6187 , n6208 );
xor ( n6210 , n6178 , n6209 );
and ( n6211 , n5748 , n5821 );
and ( n6212 , n5821 , n5867 );
and ( n6213 , n5748 , n5867 );
or ( n6214 , n6211 , n6212 , n6213 );
xor ( n6215 , n6210 , n6214 );
and ( n6216 , n5868 , n5872 );
and ( n6217 , n5873 , n5876 );
or ( n6218 , n6216 , n6217 );
xor ( n6219 , n6215 , n6218 );
buf ( n6220 , n6219 );
and ( n6221 , n5886 , n5902 );
and ( n6222 , n5902 , n5938 );
and ( n6223 , n5886 , n5938 );
or ( n6224 , n6221 , n6222 , n6223 );
and ( n6225 , n5890 , n5896 );
and ( n6226 , n5896 , n5901 );
and ( n6227 , n5890 , n5901 );
or ( n6228 , n6225 , n6226 , n6227 );
and ( n6229 , n5907 , n5911 );
and ( n6230 , n5911 , n5937 );
and ( n6231 , n5907 , n5937 );
or ( n6232 , n6229 , n6230 , n6231 );
and ( n6233 , n5893 , n4418 );
buf ( n6234 , n2305 );
buf ( n6235 , n6234 );
and ( n6236 , n6235 , n4415 );
nor ( n6237 , n6233 , n6236 );
xnor ( n6238 , n6237 , n4413 );
xor ( n6239 , n6232 , n6238 );
and ( n6240 , n5300 , n4433 );
and ( n6241 , n5588 , n4431 );
nor ( n6242 , n6240 , n6241 );
xnor ( n6243 , n6242 , n4441 );
xor ( n6244 , n6239 , n6243 );
xor ( n6245 , n6228 , n6244 );
and ( n6246 , n5927 , n5931 );
and ( n6247 , n5931 , n5936 );
and ( n6248 , n5927 , n5936 );
or ( n6249 , n6246 , n6247 , n6248 );
and ( n6250 , n4817 , n4402 );
and ( n6251 , n5042 , n4391 );
nor ( n6252 , n6250 , n6251 );
xnor ( n6253 , n6252 , n4398 );
xor ( n6254 , n6249 , n6253 );
and ( n6255 , n4421 , n4835 );
and ( n6256 , n4631 , n4648 );
nor ( n6257 , n6255 , n6256 );
xnor ( n6258 , n6257 , n4831 );
and ( n6259 , n4436 , n5323 );
and ( n6260 , n4411 , n5064 );
nor ( n6261 , n6259 , n6260 );
xnor ( n6262 , n6261 , n5319 );
xor ( n6263 , n6258 , n6262 );
and ( n6264 , n5919 , n5926 );
and ( n6265 , n4405 , n5922 );
and ( n6266 , n4427 , n5616 );
nor ( n6267 , n6265 , n6266 );
xnor ( n6268 , n6267 , n5918 );
xor ( n6269 , n6264 , n6268 );
buf ( n6270 , n540 );
buf ( n6271 , n6270 );
xor ( n6272 , n6271 , n5915 );
and ( n6273 , n4386 , n6272 );
xor ( n6274 , n6269 , n6273 );
xor ( n6275 , n6263 , n6274 );
xor ( n6276 , n6254 , n6275 );
xor ( n6277 , n6245 , n6276 );
xor ( n6278 , n6224 , n6277 );
and ( n6279 , n5882 , n5939 );
and ( n6280 , n5940 , n5943 );
or ( n6281 , n6279 , n6280 );
xor ( n6282 , n6278 , n6281 );
buf ( n6283 , n6282 );
not ( n6284 , n454 );
and ( n6285 , n6284 , n6220 );
and ( n6286 , n6283 , n454 );
or ( n6287 , n6285 , n6286 );
buf ( n6288 , n6287 );
buf ( n6289 , n6288 );
and ( n6290 , n6289 , n4505 );
xor ( n6291 , n6094 , n6290 );
and ( n6292 , n5356 , n5089 );
and ( n6293 , n5636 , n4866 );
xor ( n6294 , n6292 , n6293 );
and ( n6295 , n5951 , n4557 );
xor ( n6296 , n6294 , n6295 );
xor ( n6297 , n6291 , n6296 );
and ( n6298 , n5744 , n5952 );
and ( n6299 , n5952 , n5958 );
and ( n6300 , n5744 , n5958 );
or ( n6301 , n6298 , n6299 , n6300 );
xor ( n6302 , n6297 , n6301 );
and ( n6303 , n5740 , n5959 );
and ( n6304 , n5959 , n5964 );
and ( n6305 , n5740 , n5964 );
or ( n6306 , n6303 , n6304 , n6305 );
xor ( n6307 , n6302 , n6306 );
or ( n6308 , n5965 , n5969 );
xnor ( n6309 , n6307 , n6308 );
and ( n6310 , n5970 , n5972 );
xor ( n6311 , n6309 , n6310 );
buf ( n6312 , n6311 );
not ( n6313 , n4509 );
and ( n6314 , n6313 , n6090 );
and ( n6315 , n6312 , n4509 );
or ( n6316 , n6314 , n6315 );
and ( n6317 , n4548 , n6068 );
and ( n6318 , n4696 , n5730 );
nor ( n6319 , n6317 , n6318 );
xnor ( n6320 , n6319 , n6064 );
buf ( n6321 , n528 );
buf ( n6322 , n544 );
xor ( n6323 , n6321 , n6322 );
and ( n6324 , n6051 , n6052 );
and ( n6325 , n6052 , n6057 );
and ( n6326 , n6051 , n6057 );
or ( n6327 , n6324 , n6325 , n6326 );
xor ( n6328 , n6323 , n6327 );
buf ( n6329 , n6328 );
buf ( n6330 , n6329 );
buf ( n6331 , n6330 );
xor ( n6332 , n6331 , n6061 );
and ( n6333 , n4139 , n6332 );
xor ( n6334 , n6320 , n6333 );
and ( n6335 , n6065 , n6072 );
xor ( n6336 , n6334 , n6335 );
and ( n6337 , n6037 , n4524 );
and ( n6338 , n5998 , n6023 );
and ( n6339 , n6023 , n6028 );
and ( n6340 , n5998 , n6028 );
or ( n6341 , n6338 , n6339 , n6340 );
and ( n6342 , n5995 , n4530 );
buf ( n6343 , n496 );
buf ( n6344 , n512 );
xor ( n6345 , n6343 , n6344 );
and ( n6346 , n5985 , n5986 );
and ( n6347 , n5986 , n5991 );
and ( n6348 , n5985 , n5991 );
or ( n6349 , n6346 , n6347 , n6348 );
xor ( n6350 , n6345 , n6349 );
buf ( n6351 , n6350 );
buf ( n6352 , n6351 );
buf ( n6353 , n6352 );
and ( n6354 , n6353 , n4134 );
nor ( n6355 , n6342 , n6354 );
xnor ( n6356 , n6355 , n4527 );
and ( n6357 , n6005 , n6012 );
and ( n6358 , n5387 , n4898 );
and ( n6359 , n5672 , n4689 );
nor ( n6360 , n6358 , n6359 );
xnor ( n6361 , n6360 , n4904 );
xor ( n6362 , n6357 , n6361 );
xor ( n6363 , n6356 , n6362 );
and ( n6364 , n6013 , n6017 );
and ( n6365 , n6017 , n6022 );
and ( n6366 , n6013 , n6022 );
or ( n6367 , n6364 , n6365 , n6366 );
and ( n6368 , n4890 , n5405 );
and ( n6369 , n5121 , n5132 );
nor ( n6370 , n6368 , n6369 );
xnor ( n6371 , n6370 , n5401 );
and ( n6372 , n4539 , n6008 );
and ( n6373 , n4683 , n5689 );
nor ( n6374 , n6372 , n6373 );
xnor ( n6375 , n6374 , n6004 );
xor ( n6376 , n6371 , n6375 );
buf ( n6377 , n1467 );
buf ( n6378 , n6377 );
xor ( n6379 , n6378 , n6001 );
and ( n6380 , n4132 , n6379 );
xor ( n6381 , n6376 , n6380 );
xor ( n6382 , n6367 , n6381 );
xor ( n6383 , n6363 , n6382 );
xor ( n6384 , n6341 , n6383 );
and ( n6385 , n5983 , n6029 );
and ( n6386 , n6030 , n6033 );
or ( n6387 , n6385 , n6386 );
xor ( n6388 , n6384 , n6387 );
buf ( n6389 , n6388 );
buf ( n6390 , n6389 );
buf ( n6391 , n6390 );
and ( n6392 , n6391 , n4145 );
nor ( n6393 , n6337 , n6392 );
xnor ( n6394 , n6393 , n4521 );
and ( n6395 , n5419 , n4938 );
and ( n6396 , n5700 , n4711 );
nor ( n6397 , n6395 , n6396 );
xnor ( n6398 , n6397 , n4934 );
xor ( n6399 , n6394 , n6398 );
and ( n6400 , n4916 , n5441 );
and ( n6401 , n5140 , n5161 );
nor ( n6402 , n6400 , n6401 );
xnor ( n6403 , n6402 , n5437 );
xor ( n6404 , n6399 , n6403 );
xor ( n6405 , n6336 , n6404 );
and ( n6406 , n6073 , n6077 );
and ( n6407 , n6077 , n6082 );
and ( n6408 , n6073 , n6082 );
or ( n6409 , n6406 , n6407 , n6408 );
xor ( n6410 , n6405 , n6409 );
and ( n6411 , n6044 , n6048 );
and ( n6412 , n6048 , n6083 );
and ( n6413 , n6044 , n6083 );
or ( n6414 , n6411 , n6412 , n6413 );
xor ( n6415 , n6410 , n6414 );
and ( n6416 , n6040 , n6084 );
and ( n6417 , n6085 , n6088 );
or ( n6418 , n6416 , n6417 );
xor ( n6419 , n6415 , n6418 );
buf ( n6420 , n6419 );
and ( n6421 , n6292 , n6293 );
and ( n6422 , n6293 , n6295 );
and ( n6423 , n6292 , n6295 );
or ( n6424 , n6421 , n6422 , n6423 );
and ( n6425 , n6098 , n6177 );
and ( n6426 , n6177 , n6209 );
and ( n6427 , n6098 , n6209 );
or ( n6428 , n6425 , n6426 , n6427 );
and ( n6429 , n6102 , n6171 );
and ( n6430 , n6171 , n6176 );
and ( n6431 , n6102 , n6176 );
or ( n6432 , n6429 , n6430 , n6431 );
and ( n6433 , n6182 , n6186 );
and ( n6434 , n6186 , n6208 );
and ( n6435 , n6182 , n6208 );
or ( n6436 , n6433 , n6434 , n6435 );
and ( n6437 , n6168 , n4235 );
and ( n6438 , n6150 , n6154 );
and ( n6439 , n6154 , n6159 );
and ( n6440 , n6150 , n6159 );
or ( n6441 , n6438 , n6439 , n6440 );
and ( n6442 , n6120 , n4157 );
buf ( n6443 , n523 );
buf ( n6444 , n6443 );
and ( n6445 , n6444 , n4154 );
nor ( n6446 , n6442 , n6445 );
xnor ( n6447 , n6446 , n4152 );
not ( n6448 , n6116 );
buf ( n6449 , n459 );
buf ( n6450 , n6449 );
and ( n6451 , n6114 , n5760 );
not ( n6452 , n6451 );
and ( n6453 , n6450 , n6452 );
and ( n6454 , n6448 , n6453 );
xor ( n6455 , n6447 , n6454 );
and ( n6456 , n6107 , n6111 );
and ( n6457 , n6111 , n6116 );
and ( n6458 , n6107 , n6116 );
or ( n6459 , n6456 , n6457 , n6458 );
xor ( n6460 , n6455 , n6459 );
and ( n6461 , n6123 , n6127 );
and ( n6462 , n6127 , n6132 );
and ( n6463 , n6123 , n6132 );
or ( n6464 , n6461 , n6462 , n6463 );
xor ( n6465 , n6460 , n6464 );
and ( n6466 , n6138 , n6139 );
and ( n6467 , n6139 , n6144 );
and ( n6468 , n6138 , n6144 );
or ( n6469 , n6466 , n6467 , n6468 );
and ( n6470 , n5487 , n4173 );
and ( n6471 , n5791 , n4171 );
nor ( n6472 , n6470 , n6471 );
xnor ( n6473 , n6472 , n4181 );
and ( n6474 , n4568 , n4752 );
and ( n6475 , n4724 , n4579 );
nor ( n6476 , n6474 , n6475 );
xnor ( n6477 , n6476 , n4733 );
xor ( n6478 , n6473 , n6477 );
and ( n6479 , n4160 , n5208 );
and ( n6480 , n4243 , n4976 );
nor ( n6481 , n6479 , n6480 );
xnor ( n6482 , n6481 , n5214 );
xor ( n6483 , n6478 , n6482 );
xor ( n6484 , n6469 , n6483 );
and ( n6485 , n4965 , n4262 );
and ( n6486 , n5195 , n4188 );
nor ( n6487 , n6485 , n6486 );
xnor ( n6488 , n6487 , n4252 );
and ( n6489 , n4176 , n5773 );
and ( n6490 , n4150 , n5519 );
nor ( n6491 , n6489 , n6490 );
xnor ( n6492 , n6491 , n5763 );
xor ( n6493 , n6488 , n6492 );
xor ( n6494 , n6450 , n6114 );
not ( n6495 , n6115 );
and ( n6496 , n6494 , n6495 );
and ( n6497 , n4185 , n6496 );
and ( n6498 , n4165 , n6115 );
nor ( n6499 , n6497 , n6498 );
xnor ( n6500 , n6499 , n6453 );
xor ( n6501 , n6493 , n6500 );
xor ( n6502 , n6484 , n6501 );
xor ( n6503 , n6465 , n6502 );
and ( n6504 , n6117 , n6133 );
and ( n6505 , n6133 , n6145 );
and ( n6506 , n6117 , n6145 );
or ( n6507 , n6504 , n6505 , n6506 );
xor ( n6508 , n6503 , n6507 );
xor ( n6509 , n6441 , n6508 );
and ( n6510 , n6146 , n6160 );
and ( n6511 , n6161 , n6164 );
or ( n6512 , n6510 , n6511 );
xor ( n6513 , n6509 , n6512 );
buf ( n6514 , n6513 );
buf ( n6515 , n6514 );
buf ( n6516 , n6515 );
and ( n6517 , n6516 , n4232 );
nor ( n6518 , n6437 , n6517 );
xnor ( n6519 , n6518 , n4230 );
xor ( n6520 , n6436 , n6519 );
and ( n6521 , n5535 , n4319 );
and ( n6522 , n5818 , n4310 );
nor ( n6523 , n6521 , n6522 );
xnor ( n6524 , n6523 , n4315 );
xor ( n6525 , n6520 , n6524 );
xor ( n6526 , n6432 , n6525 );
and ( n6527 , n6191 , n6195 );
and ( n6528 , n6195 , n6207 );
and ( n6529 , n6191 , n6207 );
or ( n6530 , n6527 , n6528 , n6529 );
and ( n6531 , n4999 , n4298 );
and ( n6532 , n5247 , n4287 );
nor ( n6533 , n6531 , n6532 );
xnor ( n6534 , n6533 , n4294 );
xor ( n6535 , n6530 , n6534 );
and ( n6536 , n4594 , n4788 );
and ( n6537 , n4770 , n4611 );
nor ( n6538 , n6536 , n6537 );
xnor ( n6539 , n6538 , n4784 );
and ( n6540 , n4228 , n5270 );
and ( n6541 , n4275 , n5021 );
nor ( n6542 , n6540 , n6541 );
xnor ( n6543 , n6542 , n5266 );
xor ( n6544 , n6539 , n6543 );
not ( n6545 , n6206 );
buf ( n6546 , n491 );
buf ( n6547 , n6546 );
and ( n6548 , n6204 , n5843 );
not ( n6549 , n6548 );
and ( n6550 , n6547 , n6549 );
and ( n6551 , n6545 , n6550 );
xor ( n6552 , n6547 , n6204 );
not ( n6553 , n6205 );
and ( n6554 , n6552 , n6553 );
and ( n6555 , n4282 , n6554 );
and ( n6556 , n4303 , n6205 );
nor ( n6557 , n6555 , n6556 );
xnor ( n6558 , n6557 , n6550 );
xor ( n6559 , n6551 , n6558 );
and ( n6560 , n6197 , n6201 );
and ( n6561 , n6201 , n6206 );
and ( n6562 , n6197 , n6206 );
or ( n6563 , n6560 , n6561 , n6562 );
xor ( n6564 , n6559 , n6563 );
and ( n6565 , n4329 , n5850 );
and ( n6566 , n4342 , n5566 );
nor ( n6567 , n6565 , n6566 );
xnor ( n6568 , n6567 , n5846 );
xor ( n6569 , n6564 , n6568 );
xor ( n6570 , n6544 , n6569 );
xor ( n6571 , n6535 , n6570 );
xor ( n6572 , n6526 , n6571 );
xor ( n6573 , n6428 , n6572 );
and ( n6574 , n6210 , n6214 );
and ( n6575 , n6215 , n6218 );
or ( n6576 , n6574 , n6575 );
xor ( n6577 , n6573 , n6576 );
buf ( n6578 , n6577 );
and ( n6579 , n6232 , n6238 );
and ( n6580 , n6238 , n6243 );
and ( n6581 , n6232 , n6243 );
or ( n6582 , n6579 , n6580 , n6581 );
and ( n6583 , n6258 , n6262 );
and ( n6584 , n6262 , n6274 );
and ( n6585 , n6258 , n6274 );
or ( n6586 , n6583 , n6584 , n6585 );
and ( n6587 , n5588 , n4433 );
and ( n6588 , n5893 , n4431 );
nor ( n6589 , n6587 , n6588 );
xnor ( n6590 , n6589 , n4441 );
xor ( n6591 , n6586 , n6590 );
and ( n6592 , n5042 , n4402 );
and ( n6593 , n5300 , n4391 );
nor ( n6594 , n6592 , n6593 );
xnor ( n6595 , n6594 , n4398 );
xor ( n6596 , n6591 , n6595 );
xor ( n6597 , n6582 , n6596 );
and ( n6598 , n6249 , n6253 );
and ( n6599 , n6253 , n6275 );
and ( n6600 , n6249 , n6275 );
or ( n6601 , n6598 , n6599 , n6600 );
and ( n6602 , n6235 , n4418 );
buf ( n6603 , n2471 );
buf ( n6604 , n6603 );
and ( n6605 , n6604 , n4415 );
nor ( n6606 , n6602 , n6605 );
xnor ( n6607 , n6606 , n4413 );
xor ( n6608 , n6601 , n6607 );
and ( n6609 , n4631 , n4835 );
and ( n6610 , n4817 , n4648 );
nor ( n6611 , n6609 , n6610 );
xnor ( n6612 , n6611 , n4831 );
and ( n6613 , n4411 , n5323 );
and ( n6614 , n4421 , n5064 );
nor ( n6615 , n6613 , n6614 );
xnor ( n6616 , n6615 , n5319 );
xor ( n6617 , n6612 , n6616 );
not ( n6618 , n6273 );
buf ( n6619 , n539 );
buf ( n6620 , n6619 );
and ( n6621 , n6271 , n5915 );
not ( n6622 , n6621 );
and ( n6623 , n6620 , n6622 );
and ( n6624 , n6618 , n6623 );
xor ( n6625 , n6620 , n6271 );
not ( n6626 , n6272 );
and ( n6627 , n6625 , n6626 );
and ( n6628 , n4386 , n6627 );
and ( n6629 , n4405 , n6272 );
nor ( n6630 , n6628 , n6629 );
xnor ( n6631 , n6630 , n6623 );
xor ( n6632 , n6624 , n6631 );
and ( n6633 , n6264 , n6268 );
and ( n6634 , n6268 , n6273 );
and ( n6635 , n6264 , n6273 );
or ( n6636 , n6633 , n6634 , n6635 );
xor ( n6637 , n6632 , n6636 );
and ( n6638 , n4427 , n5922 );
and ( n6639 , n4436 , n5616 );
nor ( n6640 , n6638 , n6639 );
xnor ( n6641 , n6640 , n5918 );
xor ( n6642 , n6637 , n6641 );
xor ( n6643 , n6617 , n6642 );
xor ( n6644 , n6608 , n6643 );
xor ( n6645 , n6597 , n6644 );
and ( n6646 , n6228 , n6244 );
and ( n6647 , n6244 , n6276 );
and ( n6648 , n6228 , n6276 );
or ( n6649 , n6646 , n6647 , n6648 );
xor ( n6650 , n6645 , n6649 );
and ( n6651 , n6224 , n6277 );
and ( n6652 , n6278 , n6281 );
or ( n6653 , n6651 , n6652 );
xor ( n6654 , n6650 , n6653 );
buf ( n6655 , n6654 );
not ( n6656 , n454 );
and ( n6657 , n6656 , n6578 );
and ( n6658 , n6655 , n454 );
or ( n6659 , n6657 , n6658 );
buf ( n6660 , n6659 );
buf ( n6661 , n6660 );
and ( n6662 , n6661 , n4505 );
xor ( n6663 , n6424 , n6662 );
and ( n6664 , n5636 , n5089 );
and ( n6665 , n5951 , n4866 );
xor ( n6666 , n6664 , n6665 );
and ( n6667 , n6289 , n4557 );
xor ( n6668 , n6666 , n6667 );
xor ( n6669 , n6663 , n6668 );
and ( n6670 , n6094 , n6290 );
and ( n6671 , n6290 , n6296 );
and ( n6672 , n6094 , n6296 );
or ( n6673 , n6670 , n6671 , n6672 );
xor ( n6674 , n6669 , n6673 );
and ( n6675 , n6297 , n6301 );
and ( n6676 , n6301 , n6306 );
and ( n6677 , n6297 , n6306 );
or ( n6678 , n6675 , n6676 , n6677 );
xor ( n6679 , n6674 , n6678 );
or ( n6680 , n6307 , n6308 );
xnor ( n6681 , n6679 , n6680 );
and ( n6682 , n6309 , n6310 );
xor ( n6683 , n6681 , n6682 );
buf ( n6684 , n6683 );
not ( n6685 , n4509 );
and ( n6686 , n6685 , n6420 );
and ( n6687 , n6684 , n4509 );
or ( n6688 , n6686 , n6687 );
and ( n6689 , n4696 , n6068 );
and ( n6690 , n4916 , n5730 );
nor ( n6691 , n6689 , n6690 );
xnor ( n6692 , n6691 , n6064 );
not ( n6693 , n6333 );
buf ( n6694 , n527 );
buf ( n6695 , n543 );
xor ( n6696 , n6694 , n6695 );
and ( n6697 , n6321 , n6322 );
and ( n6698 , n6322 , n6327 );
and ( n6699 , n6321 , n6327 );
or ( n6700 , n6697 , n6698 , n6699 );
xor ( n6701 , n6696 , n6700 );
buf ( n6702 , n6701 );
buf ( n6703 , n6702 );
buf ( n6704 , n6703 );
and ( n6705 , n6331 , n6061 );
not ( n6706 , n6705 );
and ( n6707 , n6704 , n6706 );
and ( n6708 , n6693 , n6707 );
xor ( n6709 , n6704 , n6331 );
not ( n6710 , n6332 );
and ( n6711 , n6709 , n6710 );
and ( n6712 , n4139 , n6711 );
and ( n6713 , n4548 , n6332 );
nor ( n6714 , n6712 , n6713 );
xnor ( n6715 , n6714 , n6707 );
xor ( n6716 , n6708 , n6715 );
xor ( n6717 , n6692 , n6716 );
and ( n6718 , n6334 , n6335 );
and ( n6719 , n6335 , n6404 );
and ( n6720 , n6334 , n6404 );
or ( n6721 , n6718 , n6719 , n6720 );
xor ( n6722 , n6717 , n6721 );
and ( n6723 , n6320 , n6333 );
and ( n6724 , n6394 , n6398 );
and ( n6725 , n6398 , n6403 );
and ( n6726 , n6394 , n6403 );
or ( n6727 , n6724 , n6725 , n6726 );
xor ( n6728 , n6723 , n6727 );
and ( n6729 , n6391 , n4524 );
and ( n6730 , n6356 , n6362 );
and ( n6731 , n6362 , n6382 );
and ( n6732 , n6356 , n6382 );
or ( n6733 , n6730 , n6731 , n6732 );
and ( n6734 , n6357 , n6361 );
and ( n6735 , n6367 , n6381 );
xor ( n6736 , n6734 , n6735 );
and ( n6737 , n6353 , n4530 );
buf ( n6738 , n495 );
buf ( n6739 , n511 );
xor ( n6740 , n6738 , n6739 );
and ( n6741 , n6343 , n6344 );
and ( n6742 , n6344 , n6349 );
and ( n6743 , n6343 , n6349 );
or ( n6744 , n6741 , n6742 , n6743 );
xor ( n6745 , n6740 , n6744 );
buf ( n6746 , n6745 );
buf ( n6747 , n6746 );
buf ( n6748 , n6747 );
and ( n6749 , n6748 , n4134 );
nor ( n6750 , n6737 , n6749 );
xnor ( n6751 , n6750 , n4527 );
not ( n6752 , n6380 );
buf ( n6753 , n1616 );
buf ( n6754 , n6753 );
and ( n6755 , n6378 , n6001 );
not ( n6756 , n6755 );
and ( n6757 , n6754 , n6756 );
and ( n6758 , n6752 , n6757 );
xor ( n6759 , n6754 , n6378 );
not ( n6760 , n6379 );
and ( n6761 , n6759 , n6760 );
and ( n6762 , n4132 , n6761 );
and ( n6763 , n4539 , n6379 );
nor ( n6764 , n6762 , n6763 );
xnor ( n6765 , n6764 , n6757 );
xor ( n6766 , n6758 , n6765 );
and ( n6767 , n5672 , n4898 );
and ( n6768 , n5995 , n4689 );
nor ( n6769 , n6767 , n6768 );
xnor ( n6770 , n6769 , n4904 );
xor ( n6771 , n6766 , n6770 );
and ( n6772 , n4683 , n6008 );
and ( n6773 , n4890 , n5689 );
nor ( n6774 , n6772 , n6773 );
xnor ( n6775 , n6774 , n6004 );
xor ( n6776 , n6771 , n6775 );
xor ( n6777 , n6751 , n6776 );
and ( n6778 , n6371 , n6375 );
and ( n6779 , n6375 , n6380 );
and ( n6780 , n6371 , n6380 );
or ( n6781 , n6778 , n6779 , n6780 );
and ( n6782 , n5121 , n5405 );
and ( n6783 , n5387 , n5132 );
nor ( n6784 , n6782 , n6783 );
xnor ( n6785 , n6784 , n5401 );
xor ( n6786 , n6781 , n6785 );
xor ( n6787 , n6777 , n6786 );
xor ( n6788 , n6736 , n6787 );
xor ( n6789 , n6733 , n6788 );
and ( n6790 , n6341 , n6383 );
and ( n6791 , n6384 , n6387 );
or ( n6792 , n6790 , n6791 );
xor ( n6793 , n6789 , n6792 );
buf ( n6794 , n6793 );
buf ( n6795 , n6794 );
buf ( n6796 , n6795 );
and ( n6797 , n6796 , n4145 );
nor ( n6798 , n6729 , n6797 );
xnor ( n6799 , n6798 , n4521 );
and ( n6800 , n5700 , n4938 );
and ( n6801 , n6037 , n4711 );
nor ( n6802 , n6800 , n6801 );
xnor ( n6803 , n6802 , n4934 );
xor ( n6804 , n6799 , n6803 );
and ( n6805 , n5140 , n5441 );
and ( n6806 , n5419 , n5161 );
nor ( n6807 , n6805 , n6806 );
xnor ( n6808 , n6807 , n5437 );
xor ( n6809 , n6804 , n6808 );
xor ( n6810 , n6728 , n6809 );
xor ( n6811 , n6722 , n6810 );
and ( n6812 , n6405 , n6409 );
and ( n6813 , n6409 , n6414 );
and ( n6814 , n6405 , n6414 );
or ( n6815 , n6812 , n6813 , n6814 );
xor ( n6816 , n6811 , n6815 );
and ( n6817 , n6415 , n6418 );
xor ( n6818 , n6816 , n6817 );
buf ( n6819 , n6818 );
and ( n6820 , n6664 , n6665 );
and ( n6821 , n6665 , n6667 );
and ( n6822 , n6664 , n6667 );
or ( n6823 , n6820 , n6821 , n6822 );
and ( n6824 , n6436 , n6519 );
and ( n6825 , n6519 , n6524 );
and ( n6826 , n6436 , n6524 );
or ( n6827 , n6824 , n6825 , n6826 );
and ( n6828 , n6530 , n6534 );
and ( n6829 , n6534 , n6570 );
and ( n6830 , n6530 , n6570 );
or ( n6831 , n6828 , n6829 , n6830 );
and ( n6832 , n6516 , n4235 );
and ( n6833 , n6469 , n6483 );
and ( n6834 , n6483 , n6501 );
and ( n6835 , n6469 , n6501 );
or ( n6836 , n6833 , n6834 , n6835 );
and ( n6837 , n6465 , n6502 );
and ( n6838 , n6502 , n6507 );
and ( n6839 , n6465 , n6507 );
or ( n6840 , n6837 , n6838 , n6839 );
xor ( n6841 , n6836 , n6840 );
and ( n6842 , n6473 , n6477 );
and ( n6843 , n6477 , n6482 );
and ( n6844 , n6473 , n6482 );
or ( n6845 , n6842 , n6843 , n6844 );
and ( n6846 , n6488 , n6492 );
and ( n6847 , n6492 , n6500 );
and ( n6848 , n6488 , n6500 );
or ( n6849 , n6846 , n6847 , n6848 );
xor ( n6850 , n6845 , n6849 );
and ( n6851 , n6444 , n4157 );
buf ( n6852 , n522 );
buf ( n6853 , n6852 );
and ( n6854 , n6853 , n4154 );
nor ( n6855 , n6851 , n6854 );
xnor ( n6856 , n6855 , n4152 );
and ( n6857 , n5791 , n4173 );
and ( n6858 , n6120 , n4171 );
nor ( n6859 , n6857 , n6858 );
xnor ( n6860 , n6859 , n4181 );
xor ( n6861 , n6856 , n6860 );
buf ( n6862 , n458 );
buf ( n6863 , n6862 );
xor ( n6864 , n6863 , n6450 );
and ( n6865 , n4185 , n6864 );
xor ( n6866 , n6861 , n6865 );
xor ( n6867 , n6850 , n6866 );
and ( n6868 , n6455 , n6459 );
and ( n6869 , n6459 , n6464 );
and ( n6870 , n6455 , n6464 );
or ( n6871 , n6868 , n6869 , n6870 );
xor ( n6872 , n6867 , n6871 );
and ( n6873 , n5195 , n4262 );
and ( n6874 , n5487 , n4188 );
nor ( n6875 , n6873 , n6874 );
xnor ( n6876 , n6875 , n4252 );
and ( n6877 , n4724 , n4752 );
and ( n6878 , n4965 , n4579 );
nor ( n6879 , n6877 , n6878 );
xnor ( n6880 , n6879 , n4733 );
xor ( n6881 , n6876 , n6880 );
and ( n6882 , n4243 , n5208 );
and ( n6883 , n4568 , n4976 );
nor ( n6884 , n6882 , n6883 );
xnor ( n6885 , n6884 , n5214 );
xor ( n6886 , n6881 , n6885 );
and ( n6887 , n6447 , n6454 );
and ( n6888 , n4150 , n5773 );
and ( n6889 , n4160 , n5519 );
nor ( n6890 , n6888 , n6889 );
xnor ( n6891 , n6890 , n5763 );
xor ( n6892 , n6887 , n6891 );
and ( n6893 , n4165 , n6496 );
and ( n6894 , n4176 , n6115 );
nor ( n6895 , n6893 , n6894 );
xnor ( n6896 , n6895 , n6453 );
xor ( n6897 , n6892 , n6896 );
xor ( n6898 , n6886 , n6897 );
xor ( n6899 , n6872 , n6898 );
xor ( n6900 , n6841 , n6899 );
and ( n6901 , n6441 , n6508 );
and ( n6902 , n6509 , n6512 );
or ( n6903 , n6901 , n6902 );
xor ( n6904 , n6900 , n6903 );
buf ( n6905 , n6904 );
buf ( n6906 , n6905 );
buf ( n6907 , n6906 );
and ( n6908 , n6907 , n4232 );
nor ( n6909 , n6832 , n6908 );
xnor ( n6910 , n6909 , n4230 );
xor ( n6911 , n6831 , n6910 );
and ( n6912 , n5818 , n4319 );
and ( n6913 , n6168 , n4310 );
nor ( n6914 , n6912 , n6913 );
xnor ( n6915 , n6914 , n4315 );
xor ( n6916 , n6911 , n6915 );
xor ( n6917 , n6827 , n6916 );
and ( n6918 , n6539 , n6543 );
and ( n6919 , n6543 , n6569 );
and ( n6920 , n6539 , n6569 );
or ( n6921 , n6918 , n6919 , n6920 );
and ( n6922 , n5247 , n4298 );
and ( n6923 , n5535 , n4287 );
nor ( n6924 , n6922 , n6923 );
xnor ( n6925 , n6924 , n4294 );
xor ( n6926 , n6921 , n6925 );
and ( n6927 , n4770 , n4788 );
and ( n6928 , n4999 , n4611 );
nor ( n6929 , n6927 , n6928 );
xnor ( n6930 , n6929 , n4784 );
and ( n6931 , n4275 , n5270 );
and ( n6932 , n4594 , n5021 );
nor ( n6933 , n6931 , n6932 );
xnor ( n6934 , n6933 , n5266 );
xor ( n6935 , n6930 , n6934 );
and ( n6936 , n6559 , n6563 );
and ( n6937 , n6563 , n6568 );
and ( n6938 , n6559 , n6568 );
or ( n6939 , n6936 , n6937 , n6938 );
and ( n6940 , n4342 , n5850 );
and ( n6941 , n4228 , n5566 );
nor ( n6942 , n6940 , n6941 );
xnor ( n6943 , n6942 , n5846 );
xor ( n6944 , n6939 , n6943 );
and ( n6945 , n6551 , n6558 );
and ( n6946 , n4303 , n6554 );
and ( n6947 , n4329 , n6205 );
nor ( n6948 , n6946 , n6947 );
xnor ( n6949 , n6948 , n6550 );
xor ( n6950 , n6945 , n6949 );
buf ( n6951 , n490 );
buf ( n6952 , n6951 );
xor ( n6953 , n6952 , n6547 );
and ( n6954 , n4282 , n6953 );
xor ( n6955 , n6950 , n6954 );
xor ( n6956 , n6944 , n6955 );
xor ( n6957 , n6935 , n6956 );
xor ( n6958 , n6926 , n6957 );
xor ( n6959 , n6917 , n6958 );
and ( n6960 , n6432 , n6525 );
and ( n6961 , n6525 , n6571 );
and ( n6962 , n6432 , n6571 );
or ( n6963 , n6960 , n6961 , n6962 );
xor ( n6964 , n6959 , n6963 );
and ( n6965 , n6428 , n6572 );
and ( n6966 , n6573 , n6576 );
or ( n6967 , n6965 , n6966 );
xor ( n6968 , n6964 , n6967 );
buf ( n6969 , n6968 );
and ( n6970 , n6601 , n6607 );
and ( n6971 , n6607 , n6643 );
and ( n6972 , n6601 , n6643 );
or ( n6973 , n6970 , n6971 , n6972 );
and ( n6974 , n6612 , n6616 );
and ( n6975 , n6616 , n6642 );
and ( n6976 , n6612 , n6642 );
or ( n6977 , n6974 , n6975 , n6976 );
and ( n6978 , n5893 , n4433 );
and ( n6979 , n6235 , n4431 );
nor ( n6980 , n6978 , n6979 );
xnor ( n6981 , n6980 , n4441 );
xor ( n6982 , n6977 , n6981 );
and ( n6983 , n5300 , n4402 );
and ( n6984 , n5588 , n4391 );
nor ( n6985 , n6983 , n6984 );
xnor ( n6986 , n6985 , n4398 );
xor ( n6987 , n6982 , n6986 );
xor ( n6988 , n6973 , n6987 );
and ( n6989 , n6586 , n6590 );
and ( n6990 , n6590 , n6595 );
and ( n6991 , n6586 , n6595 );
or ( n6992 , n6989 , n6990 , n6991 );
and ( n6993 , n6604 , n4418 );
buf ( n6994 , n2636 );
buf ( n6995 , n6994 );
and ( n6996 , n6995 , n4415 );
nor ( n6997 , n6993 , n6996 );
xnor ( n6998 , n6997 , n4413 );
xor ( n6999 , n6992 , n6998 );
and ( n7000 , n6632 , n6636 );
and ( n7001 , n6636 , n6641 );
and ( n7002 , n6632 , n6641 );
or ( n7003 , n7000 , n7001 , n7002 );
and ( n7004 , n4817 , n4835 );
and ( n7005 , n5042 , n4648 );
nor ( n7006 , n7004 , n7005 );
xnor ( n7007 , n7006 , n4831 );
xor ( n7008 , n7003 , n7007 );
and ( n7009 , n4421 , n5323 );
and ( n7010 , n4631 , n5064 );
nor ( n7011 , n7009 , n7010 );
xnor ( n7012 , n7011 , n5319 );
and ( n7013 , n4436 , n5922 );
and ( n7014 , n4411 , n5616 );
nor ( n7015 , n7013 , n7014 );
xnor ( n7016 , n7015 , n5918 );
xor ( n7017 , n7012 , n7016 );
and ( n7018 , n6624 , n6631 );
and ( n7019 , n4405 , n6627 );
and ( n7020 , n4427 , n6272 );
nor ( n7021 , n7019 , n7020 );
xnor ( n7022 , n7021 , n6623 );
xor ( n7023 , n7018 , n7022 );
buf ( n7024 , n538 );
buf ( n7025 , n7024 );
xor ( n7026 , n7025 , n6620 );
and ( n7027 , n4386 , n7026 );
xor ( n7028 , n7023 , n7027 );
xor ( n7029 , n7017 , n7028 );
xor ( n7030 , n7008 , n7029 );
xor ( n7031 , n6999 , n7030 );
xor ( n7032 , n6988 , n7031 );
and ( n7033 , n6582 , n6596 );
and ( n7034 , n6596 , n6644 );
and ( n7035 , n6582 , n6644 );
or ( n7036 , n7033 , n7034 , n7035 );
xor ( n7037 , n7032 , n7036 );
and ( n7038 , n6645 , n6649 );
and ( n7039 , n6650 , n6653 );
or ( n7040 , n7038 , n7039 );
xor ( n7041 , n7037 , n7040 );
buf ( n7042 , n7041 );
not ( n7043 , n454 );
and ( n7044 , n7043 , n6969 );
and ( n7045 , n7042 , n454 );
or ( n7046 , n7044 , n7045 );
buf ( n7047 , n7046 );
buf ( n7048 , n7047 );
and ( n7049 , n7048 , n4505 );
xor ( n7050 , n6823 , n7049 );
and ( n7051 , n5951 , n5089 );
and ( n7052 , n6289 , n4866 );
xor ( n7053 , n7051 , n7052 );
and ( n7054 , n6661 , n4557 );
xor ( n7055 , n7053 , n7054 );
xor ( n7056 , n7050 , n7055 );
and ( n7057 , n6424 , n6662 );
and ( n7058 , n6662 , n6668 );
and ( n7059 , n6424 , n6668 );
or ( n7060 , n7057 , n7058 , n7059 );
xor ( n7061 , n7056 , n7060 );
and ( n7062 , n6669 , n6673 );
and ( n7063 , n6673 , n6678 );
and ( n7064 , n6669 , n6678 );
or ( n7065 , n7062 , n7063 , n7064 );
xor ( n7066 , n7061 , n7065 );
or ( n7067 , n6679 , n6680 );
xnor ( n7068 , n7066 , n7067 );
and ( n7069 , n6681 , n6682 );
xor ( n7070 , n7068 , n7069 );
buf ( n7071 , n7070 );
not ( n7072 , n4509 );
and ( n7073 , n7072 , n6819 );
and ( n7074 , n7071 , n4509 );
or ( n7075 , n7073 , n7074 );
and ( n7076 , n6799 , n6803 );
and ( n7077 , n6803 , n6808 );
and ( n7078 , n6799 , n6808 );
or ( n7079 , n7076 , n7077 , n7078 );
and ( n7080 , n6796 , n4524 );
and ( n7081 , n6748 , n4530 );
buf ( n7082 , n494 );
buf ( n7083 , n510 );
xor ( n7084 , n7082 , n7083 );
and ( n7085 , n6738 , n6739 );
and ( n7086 , n6739 , n6744 );
and ( n7087 , n6738 , n6744 );
or ( n7088 , n7085 , n7086 , n7087 );
xor ( n7089 , n7084 , n7088 );
buf ( n7090 , n7089 );
buf ( n7091 , n7090 );
buf ( n7092 , n7091 );
and ( n7093 , n7092 , n4134 );
nor ( n7094 , n7081 , n7093 );
xnor ( n7095 , n7094 , n4527 );
and ( n7096 , n4890 , n6008 );
and ( n7097 , n5121 , n5689 );
nor ( n7098 , n7096 , n7097 );
xnor ( n7099 , n7098 , n6004 );
and ( n7100 , n4539 , n6761 );
and ( n7101 , n4683 , n6379 );
nor ( n7102 , n7100 , n7101 );
xnor ( n7103 , n7102 , n6757 );
xor ( n7104 , n7099 , n7103 );
buf ( n7105 , n1730 );
buf ( n7106 , n7105 );
xor ( n7107 , n7106 , n6754 );
and ( n7108 , n4132 , n7107 );
xor ( n7109 , n7104 , n7108 );
xor ( n7110 , n7095 , n7109 );
and ( n7111 , n6758 , n6765 );
and ( n7112 , n5995 , n4898 );
and ( n7113 , n6353 , n4689 );
nor ( n7114 , n7112 , n7113 );
xnor ( n7115 , n7114 , n4904 );
xor ( n7116 , n7111 , n7115 );
and ( n7117 , n5387 , n5405 );
and ( n7118 , n5672 , n5132 );
nor ( n7119 , n7117 , n7118 );
xnor ( n7120 , n7119 , n5401 );
xor ( n7121 , n7116 , n7120 );
xor ( n7122 , n7110 , n7121 );
and ( n7123 , n6734 , n6735 );
and ( n7124 , n6735 , n6787 );
and ( n7125 , n6734 , n6787 );
or ( n7126 , n7123 , n7124 , n7125 );
xor ( n7127 , n7122 , n7126 );
and ( n7128 , n6766 , n6770 );
and ( n7129 , n6770 , n6775 );
and ( n7130 , n6766 , n6775 );
or ( n7131 , n7128 , n7129 , n7130 );
and ( n7132 , n6781 , n6785 );
xor ( n7133 , n7131 , n7132 );
and ( n7134 , n6751 , n6776 );
and ( n7135 , n6776 , n6786 );
and ( n7136 , n6751 , n6786 );
or ( n7137 , n7134 , n7135 , n7136 );
xor ( n7138 , n7133 , n7137 );
xor ( n7139 , n7127 , n7138 );
and ( n7140 , n6733 , n6788 );
and ( n7141 , n6789 , n6792 );
or ( n7142 , n7140 , n7141 );
xor ( n7143 , n7139 , n7142 );
buf ( n7144 , n7143 );
buf ( n7145 , n7144 );
buf ( n7146 , n7145 );
and ( n7147 , n7146 , n4145 );
nor ( n7148 , n7080 , n7147 );
xnor ( n7149 , n7148 , n4521 );
and ( n7150 , n6037 , n4938 );
and ( n7151 , n6391 , n4711 );
nor ( n7152 , n7150 , n7151 );
xnor ( n7153 , n7152 , n4934 );
xor ( n7154 , n7149 , n7153 );
and ( n7155 , n5419 , n5441 );
and ( n7156 , n5700 , n5161 );
nor ( n7157 , n7155 , n7156 );
xnor ( n7158 , n7157 , n5437 );
xor ( n7159 , n7154 , n7158 );
xor ( n7160 , n7079 , n7159 );
and ( n7161 , n6692 , n6716 );
xor ( n7162 , n7160 , n7161 );
and ( n7163 , n6723 , n6727 );
and ( n7164 , n6727 , n6809 );
and ( n7165 , n6723 , n6809 );
or ( n7166 , n7163 , n7164 , n7165 );
and ( n7167 , n4916 , n6068 );
and ( n7168 , n5140 , n5730 );
nor ( n7169 , n7167 , n7168 );
xnor ( n7170 , n7169 , n6064 );
and ( n7171 , n6708 , n6715 );
and ( n7172 , n4548 , n6711 );
and ( n7173 , n4696 , n6332 );
nor ( n7174 , n7172 , n7173 );
xnor ( n7175 , n7174 , n6707 );
xor ( n7176 , n7171 , n7175 );
buf ( n7177 , n526 );
buf ( n7178 , n542 );
xor ( n7179 , n7177 , n7178 );
and ( n7180 , n6694 , n6695 );
and ( n7181 , n6695 , n6700 );
and ( n7182 , n6694 , n6700 );
or ( n7183 , n7180 , n7181 , n7182 );
xor ( n7184 , n7179 , n7183 );
buf ( n7185 , n7184 );
buf ( n7186 , n7185 );
buf ( n7187 , n7186 );
xor ( n7188 , n7187 , n6704 );
and ( n7189 , n4139 , n7188 );
xor ( n7190 , n7176 , n7189 );
xor ( n7191 , n7170 , n7190 );
xor ( n7192 , n7166 , n7191 );
and ( n7193 , n6717 , n6721 );
and ( n7194 , n6721 , n6810 );
and ( n7195 , n6717 , n6810 );
or ( n7196 , n7193 , n7194 , n7195 );
xor ( n7197 , n7192 , n7196 );
xor ( n7198 , n7162 , n7197 );
and ( n7199 , n6811 , n6815 );
and ( n7200 , n6816 , n6817 );
or ( n7201 , n7199 , n7200 );
xor ( n7202 , n7198 , n7201 );
buf ( n7203 , n7202 );
and ( n7204 , n7051 , n7052 );
and ( n7205 , n7052 , n7054 );
and ( n7206 , n7051 , n7054 );
or ( n7207 , n7204 , n7205 , n7206 );
and ( n7208 , n6827 , n6916 );
and ( n7209 , n6916 , n6958 );
and ( n7210 , n6827 , n6958 );
or ( n7211 , n7208 , n7209 , n7210 );
and ( n7212 , n6831 , n6910 );
and ( n7213 , n6910 , n6915 );
and ( n7214 , n6831 , n6915 );
or ( n7215 , n7212 , n7213 , n7214 );
and ( n7216 , n6930 , n6934 );
and ( n7217 , n6934 , n6956 );
and ( n7218 , n6930 , n6956 );
or ( n7219 , n7216 , n7217 , n7218 );
and ( n7220 , n6168 , n4319 );
and ( n7221 , n6516 , n4310 );
nor ( n7222 , n7220 , n7221 );
xnor ( n7223 , n7222 , n4315 );
xor ( n7224 , n7219 , n7223 );
and ( n7225 , n5535 , n4298 );
and ( n7226 , n5818 , n4287 );
nor ( n7227 , n7225 , n7226 );
xnor ( n7228 , n7227 , n4294 );
xor ( n7229 , n7224 , n7228 );
xor ( n7230 , n7215 , n7229 );
and ( n7231 , n6921 , n6925 );
and ( n7232 , n6925 , n6957 );
and ( n7233 , n6921 , n6957 );
or ( n7234 , n7231 , n7232 , n7233 );
and ( n7235 , n6907 , n4235 );
and ( n7236 , n6836 , n6840 );
and ( n7237 , n6840 , n6899 );
and ( n7238 , n6836 , n6899 );
or ( n7239 , n7236 , n7237 , n7238 );
and ( n7240 , n6886 , n6897 );
and ( n7241 , n6867 , n6871 );
and ( n7242 , n6871 , n6898 );
and ( n7243 , n6867 , n6898 );
or ( n7244 , n7241 , n7242 , n7243 );
xor ( n7245 , n7240 , n7244 );
and ( n7246 , n6876 , n6880 );
and ( n7247 , n6880 , n6885 );
and ( n7248 , n6876 , n6885 );
or ( n7249 , n7246 , n7247 , n7248 );
and ( n7250 , n4965 , n4752 );
and ( n7251 , n5195 , n4579 );
nor ( n7252 , n7250 , n7251 );
xnor ( n7253 , n7252 , n4733 );
and ( n7254 , n5487 , n4262 );
and ( n7255 , n5791 , n4188 );
nor ( n7256 , n7254 , n7255 );
xnor ( n7257 , n7256 , n4252 );
and ( n7258 , n4568 , n5208 );
and ( n7259 , n4724 , n4976 );
nor ( n7260 , n7258 , n7259 );
xnor ( n7261 , n7260 , n5214 );
xor ( n7262 , n7257 , n7261 );
and ( n7263 , n4160 , n5773 );
and ( n7264 , n4243 , n5519 );
nor ( n7265 , n7263 , n7264 );
xnor ( n7266 , n7265 , n5763 );
xor ( n7267 , n7262 , n7266 );
xor ( n7268 , n7253 , n7267 );
and ( n7269 , n6120 , n4173 );
and ( n7270 , n6444 , n4171 );
nor ( n7271 , n7269 , n7270 );
xnor ( n7272 , n7271 , n4181 );
buf ( n7273 , n457 );
buf ( n7274 , n7273 );
xor ( n7275 , n7274 , n6863 );
not ( n7276 , n6864 );
and ( n7277 , n7275 , n7276 );
and ( n7278 , n4185 , n7277 );
and ( n7279 , n4165 , n6864 );
nor ( n7280 , n7278 , n7279 );
and ( n7281 , n6863 , n6450 );
not ( n7282 , n7281 );
and ( n7283 , n7274 , n7282 );
xnor ( n7284 , n7280 , n7283 );
xor ( n7285 , n7272 , n7284 );
xor ( n7286 , n7268 , n7285 );
xor ( n7287 , n7249 , n7286 );
and ( n7288 , n6887 , n6891 );
and ( n7289 , n6891 , n6896 );
and ( n7290 , n6887 , n6896 );
or ( n7291 , n7288 , n7289 , n7290 );
and ( n7292 , n6845 , n6849 );
and ( n7293 , n6849 , n6866 );
and ( n7294 , n6845 , n6866 );
or ( n7295 , n7292 , n7293 , n7294 );
xor ( n7296 , n7291 , n7295 );
and ( n7297 , n6853 , n4157 );
buf ( n7298 , n521 );
buf ( n7299 , n7298 );
and ( n7300 , n7299 , n4154 );
nor ( n7301 , n7297 , n7300 );
xnor ( n7302 , n7301 , n4152 );
not ( n7303 , n6865 );
and ( n7304 , n7303 , n7283 );
xor ( n7305 , n7302 , n7304 );
and ( n7306 , n6856 , n6860 );
and ( n7307 , n6860 , n6865 );
and ( n7308 , n6856 , n6865 );
or ( n7309 , n7306 , n7307 , n7308 );
xor ( n7310 , n7305 , n7309 );
and ( n7311 , n4176 , n6496 );
and ( n7312 , n4150 , n6115 );
nor ( n7313 , n7311 , n7312 );
xnor ( n7314 , n7313 , n6453 );
xor ( n7315 , n7310 , n7314 );
xor ( n7316 , n7296 , n7315 );
xor ( n7317 , n7287 , n7316 );
xor ( n7318 , n7245 , n7317 );
xor ( n7319 , n7239 , n7318 );
and ( n7320 , n6900 , n6903 );
xor ( n7321 , n7319 , n7320 );
buf ( n7322 , n7321 );
buf ( n7323 , n7322 );
buf ( n7324 , n7323 );
and ( n7325 , n7324 , n4232 );
nor ( n7326 , n7235 , n7325 );
xnor ( n7327 , n7326 , n4230 );
xor ( n7328 , n7234 , n7327 );
and ( n7329 , n6939 , n6943 );
and ( n7330 , n6943 , n6955 );
and ( n7331 , n6939 , n6955 );
or ( n7332 , n7329 , n7330 , n7331 );
and ( n7333 , n4999 , n4788 );
and ( n7334 , n5247 , n4611 );
nor ( n7335 , n7333 , n7334 );
xnor ( n7336 , n7335 , n4784 );
xor ( n7337 , n7332 , n7336 );
and ( n7338 , n4594 , n5270 );
and ( n7339 , n4770 , n5021 );
nor ( n7340 , n7338 , n7339 );
xnor ( n7341 , n7340 , n5266 );
and ( n7342 , n4228 , n5850 );
and ( n7343 , n4275 , n5566 );
nor ( n7344 , n7342 , n7343 );
xnor ( n7345 , n7344 , n5846 );
xor ( n7346 , n7341 , n7345 );
not ( n7347 , n6954 );
buf ( n7348 , n489 );
buf ( n7349 , n7348 );
and ( n7350 , n6952 , n6547 );
not ( n7351 , n7350 );
and ( n7352 , n7349 , n7351 );
and ( n7353 , n7347 , n7352 );
xor ( n7354 , n7349 , n6952 );
not ( n7355 , n6953 );
and ( n7356 , n7354 , n7355 );
and ( n7357 , n4282 , n7356 );
and ( n7358 , n4303 , n6953 );
nor ( n7359 , n7357 , n7358 );
xnor ( n7360 , n7359 , n7352 );
xor ( n7361 , n7353 , n7360 );
and ( n7362 , n6945 , n6949 );
and ( n7363 , n6949 , n6954 );
and ( n7364 , n6945 , n6954 );
or ( n7365 , n7362 , n7363 , n7364 );
xor ( n7366 , n7361 , n7365 );
and ( n7367 , n4329 , n6554 );
and ( n7368 , n4342 , n6205 );
nor ( n7369 , n7367 , n7368 );
xnor ( n7370 , n7369 , n6550 );
xor ( n7371 , n7366 , n7370 );
xor ( n7372 , n7346 , n7371 );
xor ( n7373 , n7337 , n7372 );
xor ( n7374 , n7328 , n7373 );
xor ( n7375 , n7230 , n7374 );
xor ( n7376 , n7211 , n7375 );
and ( n7377 , n6959 , n6963 );
and ( n7378 , n6964 , n6967 );
or ( n7379 , n7377 , n7378 );
xor ( n7380 , n7376 , n7379 );
buf ( n7381 , n7380 );
and ( n7382 , n6973 , n6987 );
and ( n7383 , n6987 , n7031 );
and ( n7384 , n6973 , n7031 );
or ( n7385 , n7382 , n7383 , n7384 );
and ( n7386 , n6992 , n6998 );
and ( n7387 , n6998 , n7030 );
and ( n7388 , n6992 , n7030 );
or ( n7389 , n7386 , n7387 , n7388 );
and ( n7390 , n6977 , n6981 );
and ( n7391 , n6981 , n6986 );
and ( n7392 , n6977 , n6986 );
or ( n7393 , n7390 , n7391 , n7392 );
and ( n7394 , n7003 , n7007 );
and ( n7395 , n7007 , n7029 );
and ( n7396 , n7003 , n7029 );
or ( n7397 , n7394 , n7395 , n7396 );
xor ( n7398 , n7393 , n7397 );
and ( n7399 , n7012 , n7016 );
and ( n7400 , n7016 , n7028 );
and ( n7401 , n7012 , n7028 );
or ( n7402 , n7399 , n7400 , n7401 );
and ( n7403 , n5588 , n4402 );
and ( n7404 , n5893 , n4391 );
nor ( n7405 , n7403 , n7404 );
xnor ( n7406 , n7405 , n4398 );
xor ( n7407 , n7402 , n7406 );
and ( n7408 , n5042 , n4835 );
and ( n7409 , n5300 , n4648 );
nor ( n7410 , n7408 , n7409 );
xnor ( n7411 , n7410 , n4831 );
xor ( n7412 , n7407 , n7411 );
xor ( n7413 , n7398 , n7412 );
xor ( n7414 , n7389 , n7413 );
and ( n7415 , n6995 , n4418 );
buf ( n7416 , n2802 );
buf ( n7417 , n7416 );
and ( n7418 , n7417 , n4415 );
nor ( n7419 , n7415 , n7418 );
xnor ( n7420 , n7419 , n4413 );
and ( n7421 , n6235 , n4433 );
and ( n7422 , n6604 , n4431 );
nor ( n7423 , n7421 , n7422 );
xnor ( n7424 , n7423 , n4441 );
xor ( n7425 , n7420 , n7424 );
and ( n7426 , n4631 , n5323 );
and ( n7427 , n4817 , n5064 );
nor ( n7428 , n7426 , n7427 );
xnor ( n7429 , n7428 , n5319 );
and ( n7430 , n4411 , n5922 );
and ( n7431 , n4421 , n5616 );
nor ( n7432 , n7430 , n7431 );
xnor ( n7433 , n7432 , n5918 );
xor ( n7434 , n7429 , n7433 );
not ( n7435 , n7027 );
buf ( n7436 , n537 );
buf ( n7437 , n7436 );
and ( n7438 , n7025 , n6620 );
not ( n7439 , n7438 );
and ( n7440 , n7437 , n7439 );
and ( n7441 , n7435 , n7440 );
xor ( n7442 , n7437 , n7025 );
not ( n7443 , n7026 );
and ( n7444 , n7442 , n7443 );
and ( n7445 , n4386 , n7444 );
and ( n7446 , n4405 , n7026 );
nor ( n7447 , n7445 , n7446 );
xnor ( n7448 , n7447 , n7440 );
xor ( n7449 , n7441 , n7448 );
and ( n7450 , n7018 , n7022 );
and ( n7451 , n7022 , n7027 );
and ( n7452 , n7018 , n7027 );
or ( n7453 , n7450 , n7451 , n7452 );
xor ( n7454 , n7449 , n7453 );
and ( n7455 , n4427 , n6627 );
and ( n7456 , n4436 , n6272 );
nor ( n7457 , n7455 , n7456 );
xnor ( n7458 , n7457 , n6623 );
xor ( n7459 , n7454 , n7458 );
xor ( n7460 , n7434 , n7459 );
xor ( n7461 , n7425 , n7460 );
xor ( n7462 , n7414 , n7461 );
xor ( n7463 , n7385 , n7462 );
and ( n7464 , n7032 , n7036 );
and ( n7465 , n7037 , n7040 );
or ( n7466 , n7464 , n7465 );
xor ( n7467 , n7463 , n7466 );
buf ( n7468 , n7467 );
not ( n7469 , n454 );
and ( n7470 , n7469 , n7381 );
and ( n7471 , n7468 , n454 );
or ( n7472 , n7470 , n7471 );
buf ( n7473 , n7472 );
buf ( n7474 , n7473 );
and ( n7475 , n7474 , n4505 );
xor ( n7476 , n7207 , n7475 );
and ( n7477 , n6289 , n5089 );
and ( n7478 , n6661 , n4866 );
xor ( n7479 , n7477 , n7478 );
and ( n7480 , n7048 , n4557 );
xor ( n7481 , n7479 , n7480 );
xor ( n7482 , n7476 , n7481 );
and ( n7483 , n6823 , n7049 );
and ( n7484 , n7049 , n7055 );
and ( n7485 , n6823 , n7055 );
or ( n7486 , n7483 , n7484 , n7485 );
xor ( n7487 , n7482 , n7486 );
and ( n7488 , n7056 , n7060 );
and ( n7489 , n7060 , n7065 );
and ( n7490 , n7056 , n7065 );
or ( n7491 , n7488 , n7489 , n7490 );
xor ( n7492 , n7487 , n7491 );
or ( n7493 , n7066 , n7067 );
xnor ( n7494 , n7492 , n7493 );
and ( n7495 , n7068 , n7069 );
xor ( n7496 , n7494 , n7495 );
buf ( n7497 , n7496 );
not ( n7498 , n4509 );
and ( n7499 , n7498 , n7203 );
and ( n7500 , n7497 , n4509 );
or ( n7501 , n7499 , n7500 );
and ( n7502 , n7149 , n7153 );
and ( n7503 , n7153 , n7158 );
and ( n7504 , n7149 , n7158 );
or ( n7505 , n7502 , n7503 , n7504 );
and ( n7506 , n7146 , n4524 );
and ( n7507 , n7131 , n7132 );
and ( n7508 , n7132 , n7137 );
and ( n7509 , n7131 , n7137 );
or ( n7510 , n7507 , n7508 , n7509 );
and ( n7511 , n7111 , n7115 );
and ( n7512 , n7115 , n7120 );
and ( n7513 , n7111 , n7120 );
or ( n7514 , n7511 , n7512 , n7513 );
and ( n7515 , n7095 , n7109 );
and ( n7516 , n7109 , n7121 );
and ( n7517 , n7095 , n7121 );
or ( n7518 , n7515 , n7516 , n7517 );
xor ( n7519 , n7514 , n7518 );
and ( n7520 , n7092 , n4530 );
buf ( n7521 , n493 );
buf ( n7522 , n509 );
xor ( n7523 , n7521 , n7522 );
and ( n7524 , n7082 , n7083 );
and ( n7525 , n7083 , n7088 );
and ( n7526 , n7082 , n7088 );
or ( n7527 , n7524 , n7525 , n7526 );
xor ( n7528 , n7523 , n7527 );
buf ( n7529 , n7528 );
buf ( n7530 , n7529 );
buf ( n7531 , n7530 );
and ( n7532 , n7531 , n4134 );
nor ( n7533 , n7520 , n7532 );
xnor ( n7534 , n7533 , n4527 );
and ( n7535 , n7099 , n7103 );
and ( n7536 , n7103 , n7108 );
and ( n7537 , n7099 , n7108 );
or ( n7538 , n7535 , n7536 , n7537 );
and ( n7539 , n6353 , n4898 );
and ( n7540 , n6748 , n4689 );
nor ( n7541 , n7539 , n7540 );
xnor ( n7542 , n7541 , n4904 );
xor ( n7543 , n7538 , n7542 );
and ( n7544 , n5672 , n5405 );
and ( n7545 , n5995 , n5132 );
nor ( n7546 , n7544 , n7545 );
xnor ( n7547 , n7546 , n5401 );
xor ( n7548 , n7543 , n7547 );
xor ( n7549 , n7534 , n7548 );
not ( n7550 , n7108 );
buf ( n7551 , n1917 );
buf ( n7552 , n7551 );
and ( n7553 , n7106 , n6754 );
not ( n7554 , n7553 );
and ( n7555 , n7552 , n7554 );
and ( n7556 , n7550 , n7555 );
xor ( n7557 , n7552 , n7106 );
not ( n7558 , n7107 );
and ( n7559 , n7557 , n7558 );
and ( n7560 , n4132 , n7559 );
and ( n7561 , n4539 , n7107 );
nor ( n7562 , n7560 , n7561 );
xnor ( n7563 , n7562 , n7555 );
xor ( n7564 , n7556 , n7563 );
and ( n7565 , n5121 , n6008 );
and ( n7566 , n5387 , n5689 );
nor ( n7567 , n7565 , n7566 );
xnor ( n7568 , n7567 , n6004 );
xor ( n7569 , n7564 , n7568 );
and ( n7570 , n4683 , n6761 );
and ( n7571 , n4890 , n6379 );
nor ( n7572 , n7570 , n7571 );
xnor ( n7573 , n7572 , n6757 );
xor ( n7574 , n7569 , n7573 );
xor ( n7575 , n7549 , n7574 );
xor ( n7576 , n7519 , n7575 );
xor ( n7577 , n7510 , n7576 );
and ( n7578 , n7122 , n7126 );
and ( n7579 , n7126 , n7138 );
and ( n7580 , n7122 , n7138 );
or ( n7581 , n7578 , n7579 , n7580 );
xor ( n7582 , n7577 , n7581 );
and ( n7583 , n7139 , n7142 );
xor ( n7584 , n7582 , n7583 );
buf ( n7585 , n7584 );
buf ( n7586 , n7585 );
buf ( n7587 , n7586 );
and ( n7588 , n7587 , n4145 );
nor ( n7589 , n7506 , n7588 );
xnor ( n7590 , n7589 , n4521 );
and ( n7591 , n6391 , n4938 );
and ( n7592 , n6796 , n4711 );
nor ( n7593 , n7591 , n7592 );
xnor ( n7594 , n7593 , n4934 );
xor ( n7595 , n7590 , n7594 );
and ( n7596 , n5700 , n5441 );
and ( n7597 , n6037 , n5161 );
nor ( n7598 , n7596 , n7597 );
xnor ( n7599 , n7598 , n5437 );
xor ( n7600 , n7595 , n7599 );
xor ( n7601 , n7505 , n7600 );
and ( n7602 , n7170 , n7190 );
xor ( n7603 , n7601 , n7602 );
and ( n7604 , n7079 , n7159 );
and ( n7605 , n7159 , n7161 );
and ( n7606 , n7079 , n7161 );
or ( n7607 , n7604 , n7605 , n7606 );
and ( n7608 , n5140 , n6068 );
and ( n7609 , n5419 , n5730 );
nor ( n7610 , n7608 , n7609 );
xnor ( n7611 , n7610 , n6064 );
not ( n7612 , n7189 );
buf ( n7613 , n525 );
buf ( n7614 , n541 );
xor ( n7615 , n7613 , n7614 );
and ( n7616 , n7177 , n7178 );
and ( n7617 , n7178 , n7183 );
and ( n7618 , n7177 , n7183 );
or ( n7619 , n7616 , n7617 , n7618 );
xor ( n7620 , n7615 , n7619 );
buf ( n7621 , n7620 );
buf ( n7622 , n7621 );
buf ( n7623 , n7622 );
and ( n7624 , n7187 , n6704 );
not ( n7625 , n7624 );
and ( n7626 , n7623 , n7625 );
and ( n7627 , n7612 , n7626 );
xor ( n7628 , n7623 , n7187 );
not ( n7629 , n7188 );
and ( n7630 , n7628 , n7629 );
and ( n7631 , n4139 , n7630 );
and ( n7632 , n4548 , n7188 );
nor ( n7633 , n7631 , n7632 );
xnor ( n7634 , n7633 , n7626 );
xor ( n7635 , n7627 , n7634 );
and ( n7636 , n7171 , n7175 );
and ( n7637 , n7175 , n7189 );
and ( n7638 , n7171 , n7189 );
or ( n7639 , n7636 , n7637 , n7638 );
xor ( n7640 , n7635 , n7639 );
and ( n7641 , n4696 , n6711 );
and ( n7642 , n4916 , n6332 );
nor ( n7643 , n7641 , n7642 );
xnor ( n7644 , n7643 , n6707 );
xor ( n7645 , n7640 , n7644 );
xor ( n7646 , n7611 , n7645 );
xor ( n7647 , n7607 , n7646 );
and ( n7648 , n7166 , n7191 );
and ( n7649 , n7191 , n7196 );
and ( n7650 , n7166 , n7196 );
or ( n7651 , n7648 , n7649 , n7650 );
xor ( n7652 , n7647 , n7651 );
xor ( n7653 , n7603 , n7652 );
and ( n7654 , n7162 , n7197 );
and ( n7655 , n7198 , n7201 );
or ( n7656 , n7654 , n7655 );
xor ( n7657 , n7653 , n7656 );
buf ( n7658 , n7657 );
and ( n7659 , n7477 , n7478 );
and ( n7660 , n7478 , n7480 );
and ( n7661 , n7477 , n7480 );
or ( n7662 , n7659 , n7660 , n7661 );
and ( n7663 , n7234 , n7327 );
and ( n7664 , n7327 , n7373 );
and ( n7665 , n7234 , n7373 );
or ( n7666 , n7663 , n7664 , n7665 );
and ( n7667 , n7219 , n7223 );
and ( n7668 , n7223 , n7228 );
and ( n7669 , n7219 , n7228 );
or ( n7670 , n7667 , n7668 , n7669 );
and ( n7671 , n7324 , n4235 );
and ( n7672 , n7240 , n7244 );
and ( n7673 , n7244 , n7317 );
and ( n7674 , n7240 , n7317 );
or ( n7675 , n7672 , n7673 , n7674 );
and ( n7676 , n7305 , n7309 );
and ( n7677 , n7309 , n7314 );
and ( n7678 , n7305 , n7314 );
or ( n7679 , n7676 , n7677 , n7678 );
and ( n7680 , n7253 , n7267 );
and ( n7681 , n7267 , n7285 );
and ( n7682 , n7253 , n7285 );
or ( n7683 , n7680 , n7681 , n7682 );
xor ( n7684 , n7679 , n7683 );
and ( n7685 , n7257 , n7261 );
and ( n7686 , n7261 , n7266 );
and ( n7687 , n7257 , n7266 );
or ( n7688 , n7685 , n7686 , n7687 );
and ( n7689 , n7302 , n7304 );
xor ( n7690 , n7688 , n7689 );
and ( n7691 , n7272 , n7284 );
xor ( n7692 , n7690 , n7691 );
xor ( n7693 , n7684 , n7692 );
and ( n7694 , n7291 , n7295 );
and ( n7695 , n7295 , n7315 );
and ( n7696 , n7291 , n7315 );
or ( n7697 , n7694 , n7695 , n7696 );
and ( n7698 , n7299 , n4157 );
not ( n7699 , n7698 );
xnor ( n7700 , n7699 , n4152 );
and ( n7701 , n6444 , n4173 );
and ( n7702 , n6853 , n4171 );
nor ( n7703 , n7701 , n7702 );
xnor ( n7704 , n7703 , n4181 );
xor ( n7705 , n7700 , n7704 );
and ( n7706 , n4185 , n7274 );
xor ( n7707 , n7705 , n7706 );
and ( n7708 , n5195 , n4752 );
and ( n7709 , n5487 , n4579 );
nor ( n7710 , n7708 , n7709 );
xnor ( n7711 , n7710 , n4733 );
and ( n7712 , n4724 , n5208 );
and ( n7713 , n4965 , n4976 );
nor ( n7714 , n7712 , n7713 );
xnor ( n7715 , n7714 , n5214 );
xor ( n7716 , n7711 , n7715 );
and ( n7717 , n4165 , n7277 );
and ( n7718 , n4176 , n6864 );
nor ( n7719 , n7717 , n7718 );
xnor ( n7720 , n7719 , n7283 );
xor ( n7721 , n7716 , n7720 );
xor ( n7722 , n7707 , n7721 );
and ( n7723 , n5791 , n4262 );
and ( n7724 , n6120 , n4188 );
nor ( n7725 , n7723 , n7724 );
xnor ( n7726 , n7725 , n4252 );
and ( n7727 , n4243 , n5773 );
and ( n7728 , n4568 , n5519 );
nor ( n7729 , n7727 , n7728 );
xnor ( n7730 , n7729 , n5763 );
xor ( n7731 , n7726 , n7730 );
and ( n7732 , n4150 , n6496 );
and ( n7733 , n4160 , n6115 );
nor ( n7734 , n7732 , n7733 );
xnor ( n7735 , n7734 , n6453 );
xor ( n7736 , n7731 , n7735 );
xor ( n7737 , n7722 , n7736 );
xor ( n7738 , n7697 , n7737 );
xor ( n7739 , n7693 , n7738 );
and ( n7740 , n7249 , n7286 );
and ( n7741 , n7286 , n7316 );
and ( n7742 , n7249 , n7316 );
or ( n7743 , n7740 , n7741 , n7742 );
xor ( n7744 , n7739 , n7743 );
xor ( n7745 , n7675 , n7744 );
and ( n7746 , n7239 , n7318 );
and ( n7747 , n7319 , n7320 );
or ( n7748 , n7746 , n7747 );
xor ( n7749 , n7745 , n7748 );
buf ( n7750 , n7749 );
buf ( n7751 , n7750 );
buf ( n7752 , n7751 );
and ( n7753 , n7752 , n4232 );
nor ( n7754 , n7671 , n7753 );
xnor ( n7755 , n7754 , n4230 );
xor ( n7756 , n7670 , n7755 );
and ( n7757 , n7341 , n7345 );
and ( n7758 , n7345 , n7371 );
and ( n7759 , n7341 , n7371 );
or ( n7760 , n7757 , n7758 , n7759 );
and ( n7761 , n5818 , n4298 );
and ( n7762 , n6168 , n4287 );
nor ( n7763 , n7761 , n7762 );
xnor ( n7764 , n7763 , n4294 );
xor ( n7765 , n7760 , n7764 );
and ( n7766 , n5247 , n4788 );
and ( n7767 , n5535 , n4611 );
nor ( n7768 , n7766 , n7767 );
xnor ( n7769 , n7768 , n4784 );
xor ( n7770 , n7765 , n7769 );
xor ( n7771 , n7756 , n7770 );
xor ( n7772 , n7666 , n7771 );
and ( n7773 , n7332 , n7336 );
and ( n7774 , n7336 , n7372 );
and ( n7775 , n7332 , n7372 );
or ( n7776 , n7773 , n7774 , n7775 );
and ( n7777 , n6516 , n4319 );
and ( n7778 , n6907 , n4310 );
nor ( n7779 , n7777 , n7778 );
xnor ( n7780 , n7779 , n4315 );
xor ( n7781 , n7776 , n7780 );
and ( n7782 , n4770 , n5270 );
and ( n7783 , n4999 , n5021 );
nor ( n7784 , n7782 , n7783 );
xnor ( n7785 , n7784 , n5266 );
and ( n7786 , n4275 , n5850 );
and ( n7787 , n4594 , n5566 );
nor ( n7788 , n7786 , n7787 );
xnor ( n7789 , n7788 , n5846 );
xor ( n7790 , n7785 , n7789 );
and ( n7791 , n7361 , n7365 );
and ( n7792 , n7365 , n7370 );
and ( n7793 , n7361 , n7370 );
or ( n7794 , n7791 , n7792 , n7793 );
and ( n7795 , n4342 , n6554 );
and ( n7796 , n4228 , n6205 );
nor ( n7797 , n7795 , n7796 );
xnor ( n7798 , n7797 , n6550 );
xor ( n7799 , n7794 , n7798 );
and ( n7800 , n7353 , n7360 );
and ( n7801 , n4303 , n7356 );
and ( n7802 , n4329 , n6953 );
nor ( n7803 , n7801 , n7802 );
xnor ( n7804 , n7803 , n7352 );
xor ( n7805 , n7800 , n7804 );
and ( n7806 , n4282 , n7349 );
xor ( n7807 , n7805 , n7806 );
xor ( n7808 , n7799 , n7807 );
xor ( n7809 , n7790 , n7808 );
xor ( n7810 , n7781 , n7809 );
xor ( n7811 , n7772 , n7810 );
and ( n7812 , n7215 , n7229 );
and ( n7813 , n7229 , n7374 );
and ( n7814 , n7215 , n7374 );
or ( n7815 , n7812 , n7813 , n7814 );
xor ( n7816 , n7811 , n7815 );
and ( n7817 , n7211 , n7375 );
and ( n7818 , n7376 , n7379 );
or ( n7819 , n7817 , n7818 );
xor ( n7820 , n7816 , n7819 );
buf ( n7821 , n7820 );
and ( n7822 , n7393 , n7397 );
and ( n7823 , n7397 , n7412 );
and ( n7824 , n7393 , n7412 );
or ( n7825 , n7822 , n7823 , n7824 );
and ( n7826 , n7402 , n7406 );
and ( n7827 , n7406 , n7411 );
and ( n7828 , n7402 , n7411 );
or ( n7829 , n7826 , n7827 , n7828 );
and ( n7830 , n6604 , n4433 );
and ( n7831 , n6995 , n4431 );
nor ( n7832 , n7830 , n7831 );
xnor ( n7833 , n7832 , n4441 );
xor ( n7834 , n7829 , n7833 );
and ( n7835 , n7449 , n7453 );
and ( n7836 , n7453 , n7458 );
and ( n7837 , n7449 , n7458 );
or ( n7838 , n7835 , n7836 , n7837 );
and ( n7839 , n5300 , n4835 );
and ( n7840 , n5588 , n4648 );
nor ( n7841 , n7839 , n7840 );
xnor ( n7842 , n7841 , n4831 );
xor ( n7843 , n7838 , n7842 );
and ( n7844 , n4817 , n5323 );
and ( n7845 , n5042 , n5064 );
nor ( n7846 , n7844 , n7845 );
xnor ( n7847 , n7846 , n5319 );
xor ( n7848 , n7843 , n7847 );
xor ( n7849 , n7834 , n7848 );
xor ( n7850 , n7825 , n7849 );
and ( n7851 , n7420 , n7424 );
and ( n7852 , n7424 , n7460 );
and ( n7853 , n7420 , n7460 );
or ( n7854 , n7851 , n7852 , n7853 );
and ( n7855 , n7417 , n4418 );
buf ( n7856 , n2961 );
buf ( n7857 , n7856 );
and ( n7858 , n7857 , n4415 );
nor ( n7859 , n7855 , n7858 );
xnor ( n7860 , n7859 , n4413 );
xor ( n7861 , n7854 , n7860 );
and ( n7862 , n7429 , n7433 );
and ( n7863 , n7433 , n7459 );
and ( n7864 , n7429 , n7459 );
or ( n7865 , n7862 , n7863 , n7864 );
and ( n7866 , n5893 , n4402 );
and ( n7867 , n6235 , n4391 );
nor ( n7868 , n7866 , n7867 );
xnor ( n7869 , n7868 , n4398 );
xor ( n7870 , n7865 , n7869 );
and ( n7871 , n4421 , n5922 );
and ( n7872 , n4631 , n5616 );
nor ( n7873 , n7871 , n7872 );
xnor ( n7874 , n7873 , n5918 );
and ( n7875 , n4436 , n6627 );
and ( n7876 , n4411 , n6272 );
nor ( n7877 , n7875 , n7876 );
xnor ( n7878 , n7877 , n6623 );
xor ( n7879 , n7874 , n7878 );
and ( n7880 , n7441 , n7448 );
and ( n7881 , n4405 , n7444 );
and ( n7882 , n4427 , n7026 );
nor ( n7883 , n7881 , n7882 );
xnor ( n7884 , n7883 , n7440 );
xor ( n7885 , n7880 , n7884 );
and ( n7886 , n4386 , n7437 );
xor ( n7887 , n7885 , n7886 );
xor ( n7888 , n7879 , n7887 );
xor ( n7889 , n7870 , n7888 );
xor ( n7890 , n7861 , n7889 );
xor ( n7891 , n7850 , n7890 );
and ( n7892 , n7389 , n7413 );
and ( n7893 , n7413 , n7461 );
and ( n7894 , n7389 , n7461 );
or ( n7895 , n7892 , n7893 , n7894 );
xor ( n7896 , n7891 , n7895 );
and ( n7897 , n7385 , n7462 );
and ( n7898 , n7463 , n7466 );
or ( n7899 , n7897 , n7898 );
xor ( n7900 , n7896 , n7899 );
buf ( n7901 , n7900 );
not ( n7902 , n454 );
and ( n7903 , n7902 , n7821 );
and ( n7904 , n7901 , n454 );
or ( n7905 , n7903 , n7904 );
buf ( n7906 , n7905 );
buf ( n7907 , n7906 );
and ( n7908 , n7907 , n4505 );
xor ( n7909 , n7662 , n7908 );
and ( n7910 , n6661 , n5089 );
and ( n7911 , n7048 , n4866 );
xor ( n7912 , n7910 , n7911 );
and ( n7913 , n7474 , n4557 );
xor ( n7914 , n7912 , n7913 );
xor ( n7915 , n7909 , n7914 );
and ( n7916 , n7207 , n7475 );
and ( n7917 , n7475 , n7481 );
and ( n7918 , n7207 , n7481 );
or ( n7919 , n7916 , n7917 , n7918 );
xor ( n7920 , n7915 , n7919 );
and ( n7921 , n7482 , n7486 );
and ( n7922 , n7486 , n7491 );
and ( n7923 , n7482 , n7491 );
or ( n7924 , n7921 , n7922 , n7923 );
xor ( n7925 , n7920 , n7924 );
or ( n7926 , n7492 , n7493 );
xnor ( n7927 , n7925 , n7926 );
and ( n7928 , n7494 , n7495 );
xor ( n7929 , n7927 , n7928 );
buf ( n7930 , n7929 );
not ( n7931 , n4509 );
and ( n7932 , n7931 , n7658 );
and ( n7933 , n7930 , n4509 );
or ( n7934 , n7932 , n7933 );
and ( n7935 , n6037 , n5441 );
and ( n7936 , n6391 , n5161 );
nor ( n7937 , n7935 , n7936 );
xnor ( n7938 , n7937 , n5437 );
and ( n7939 , n5419 , n6068 );
and ( n7940 , n5700 , n5730 );
nor ( n7941 , n7939 , n7940 );
xnor ( n7942 , n7941 , n6064 );
xor ( n7943 , n7938 , n7942 );
and ( n7944 , n7635 , n7639 );
and ( n7945 , n7639 , n7644 );
and ( n7946 , n7635 , n7644 );
or ( n7947 , n7944 , n7945 , n7946 );
and ( n7948 , n4916 , n6711 );
and ( n7949 , n5140 , n6332 );
nor ( n7950 , n7948 , n7949 );
xnor ( n7951 , n7950 , n6707 );
xor ( n7952 , n7947 , n7951 );
and ( n7953 , n7627 , n7634 );
and ( n7954 , n4548 , n7630 );
and ( n7955 , n4696 , n7188 );
nor ( n7956 , n7954 , n7955 );
xnor ( n7957 , n7956 , n7626 );
xor ( n7958 , n7953 , n7957 );
buf ( n7959 , n524 );
buf ( n7960 , n540 );
xor ( n7961 , n7959 , n7960 );
and ( n7962 , n7613 , n7614 );
and ( n7963 , n7614 , n7619 );
and ( n7964 , n7613 , n7619 );
or ( n7965 , n7962 , n7963 , n7964 );
xor ( n7966 , n7961 , n7965 );
buf ( n7967 , n7966 );
buf ( n7968 , n7967 );
buf ( n7969 , n7968 );
xor ( n7970 , n7969 , n7623 );
and ( n7971 , n4139 , n7970 );
xor ( n7972 , n7958 , n7971 );
xor ( n7973 , n7952 , n7972 );
xor ( n7974 , n7943 , n7973 );
and ( n7975 , n7607 , n7646 );
and ( n7976 , n7646 , n7651 );
and ( n7977 , n7607 , n7651 );
or ( n7978 , n7975 , n7976 , n7977 );
xor ( n7979 , n7974 , n7978 );
and ( n7980 , n7587 , n4524 );
and ( n7981 , n7534 , n7548 );
and ( n7982 , n7548 , n7574 );
and ( n7983 , n7534 , n7574 );
or ( n7984 , n7981 , n7982 , n7983 );
and ( n7985 , n7514 , n7518 );
and ( n7986 , n7518 , n7575 );
and ( n7987 , n7514 , n7575 );
or ( n7988 , n7985 , n7986 , n7987 );
xor ( n7989 , n7984 , n7988 );
and ( n7990 , n7531 , n4530 );
buf ( n7991 , n492 );
buf ( n7992 , n508 );
xor ( n7993 , n7991 , n7992 );
and ( n7994 , n7521 , n7522 );
and ( n7995 , n7522 , n7527 );
and ( n7996 , n7521 , n7527 );
or ( n7997 , n7994 , n7995 , n7996 );
xor ( n7998 , n7993 , n7997 );
buf ( n7999 , n7998 );
buf ( n8000 , n7999 );
buf ( n8001 , n8000 );
and ( n8002 , n8001 , n4134 );
nor ( n8003 , n7990 , n8002 );
xnor ( n8004 , n8003 , n4527 );
and ( n8005 , n7538 , n7542 );
and ( n8006 , n7542 , n7547 );
and ( n8007 , n7538 , n7547 );
or ( n8008 , n8005 , n8006 , n8007 );
and ( n8009 , n7564 , n7568 );
and ( n8010 , n7568 , n7573 );
and ( n8011 , n7564 , n7573 );
or ( n8012 , n8009 , n8010 , n8011 );
xor ( n8013 , n8008 , n8012 );
and ( n8014 , n5995 , n5405 );
and ( n8015 , n6353 , n5132 );
nor ( n8016 , n8014 , n8015 );
xnor ( n8017 , n8016 , n5401 );
and ( n8018 , n5387 , n6008 );
and ( n8019 , n5672 , n5689 );
nor ( n8020 , n8018 , n8019 );
xnor ( n8021 , n8020 , n6004 );
xor ( n8022 , n8017 , n8021 );
and ( n8023 , n4890 , n6761 );
and ( n8024 , n5121 , n6379 );
nor ( n8025 , n8023 , n8024 );
xnor ( n8026 , n8025 , n6757 );
xor ( n8027 , n8022 , n8026 );
xor ( n8028 , n8013 , n8027 );
xor ( n8029 , n8004 , n8028 );
and ( n8030 , n6748 , n4898 );
and ( n8031 , n7092 , n4689 );
nor ( n8032 , n8030 , n8031 );
xnor ( n8033 , n8032 , n4904 );
and ( n8034 , n7556 , n7563 );
and ( n8035 , n4539 , n7559 );
and ( n8036 , n4683 , n7107 );
nor ( n8037 , n8035 , n8036 );
xnor ( n8038 , n8037 , n7555 );
xor ( n8039 , n8034 , n8038 );
buf ( n8040 , n2081 );
buf ( n8041 , n8040 );
xor ( n8042 , n8041 , n7552 );
and ( n8043 , n4132 , n8042 );
xor ( n8044 , n8039 , n8043 );
xor ( n8045 , n8033 , n8044 );
xor ( n8046 , n8029 , n8045 );
xor ( n8047 , n7989 , n8046 );
and ( n8048 , n7510 , n7576 );
and ( n8049 , n7576 , n7581 );
and ( n8050 , n7510 , n7581 );
or ( n8051 , n8048 , n8049 , n8050 );
xor ( n8052 , n8047 , n8051 );
and ( n8053 , n7582 , n7583 );
xor ( n8054 , n8052 , n8053 );
buf ( n8055 , n8054 );
buf ( n8056 , n8055 );
buf ( n8057 , n8056 );
and ( n8058 , n8057 , n4145 );
nor ( n8059 , n7980 , n8058 );
xnor ( n8060 , n8059 , n4521 );
and ( n8061 , n6796 , n4938 );
and ( n8062 , n7146 , n4711 );
nor ( n8063 , n8061 , n8062 );
xnor ( n8064 , n8063 , n4934 );
xor ( n8065 , n8060 , n8064 );
and ( n8066 , n7590 , n7594 );
and ( n8067 , n7594 , n7599 );
and ( n8068 , n7590 , n7599 );
or ( n8069 , n8066 , n8067 , n8068 );
xor ( n8070 , n8065 , n8069 );
and ( n8071 , n7611 , n7645 );
xor ( n8072 , n8070 , n8071 );
and ( n8073 , n7505 , n7600 );
and ( n8074 , n7600 , n7602 );
and ( n8075 , n7505 , n7602 );
or ( n8076 , n8073 , n8074 , n8075 );
xor ( n8077 , n8072 , n8076 );
xor ( n8078 , n7979 , n8077 );
and ( n8079 , n7603 , n7652 );
and ( n8080 , n7653 , n7656 );
or ( n8081 , n8079 , n8080 );
xor ( n8082 , n8078 , n8081 );
buf ( n8083 , n8082 );
and ( n8084 , n7910 , n7911 );
and ( n8085 , n7911 , n7913 );
and ( n8086 , n7910 , n7913 );
or ( n8087 , n8084 , n8085 , n8086 );
and ( n8088 , n7670 , n7755 );
and ( n8089 , n7755 , n7770 );
and ( n8090 , n7670 , n7770 );
or ( n8091 , n8088 , n8089 , n8090 );
and ( n8092 , n7776 , n7780 );
and ( n8093 , n7780 , n7809 );
and ( n8094 , n7776 , n7809 );
or ( n8095 , n8092 , n8093 , n8094 );
and ( n8096 , n7752 , n4235 );
and ( n8097 , n7693 , n7738 );
and ( n8098 , n7738 , n7743 );
and ( n8099 , n7693 , n7743 );
or ( n8100 , n8097 , n8098 , n8099 );
and ( n8101 , n7679 , n7683 );
and ( n8102 , n7683 , n7692 );
and ( n8103 , n7679 , n7692 );
or ( n8104 , n8101 , n8102 , n8103 );
and ( n8105 , n7697 , n7737 );
xor ( n8106 , n8104 , n8105 );
and ( n8107 , n6853 , n4173 );
and ( n8108 , n7299 , n4171 );
nor ( n8109 , n8107 , n8108 );
xnor ( n8110 , n8109 , n4181 );
and ( n8111 , n6120 , n4262 );
and ( n8112 , n6444 , n4188 );
nor ( n8113 , n8111 , n8112 );
xnor ( n8114 , n8113 , n4252 );
xor ( n8115 , n8110 , n8114 );
and ( n8116 , n4965 , n5208 );
and ( n8117 , n5195 , n4976 );
nor ( n8118 , n8116 , n8117 );
xnor ( n8119 , n8118 , n5214 );
xor ( n8120 , n8115 , n8119 );
not ( n8121 , n4152 );
and ( n8122 , n4176 , n7277 );
and ( n8123 , n4150 , n6864 );
nor ( n8124 , n8122 , n8123 );
xnor ( n8125 , n8124 , n7283 );
xor ( n8126 , n8121 , n8125 );
and ( n8127 , n4165 , n7274 );
xor ( n8128 , n8126 , n8127 );
xor ( n8129 , n8120 , n8128 );
and ( n8130 , n7688 , n7689 );
and ( n8131 , n7689 , n7691 );
and ( n8132 , n7688 , n7691 );
or ( n8133 , n8130 , n8131 , n8132 );
xor ( n8134 , n8129 , n8133 );
and ( n8135 , n7707 , n7721 );
and ( n8136 , n7721 , n7736 );
and ( n8137 , n7707 , n7736 );
or ( n8138 , n8135 , n8136 , n8137 );
and ( n8139 , n7700 , n7704 );
and ( n8140 , n7704 , n7706 );
and ( n8141 , n7700 , n7706 );
or ( n8142 , n8139 , n8140 , n8141 );
and ( n8143 , n7711 , n7715 );
and ( n8144 , n7715 , n7720 );
and ( n8145 , n7711 , n7720 );
or ( n8146 , n8143 , n8144 , n8145 );
xor ( n8147 , n8142 , n8146 );
and ( n8148 , n7726 , n7730 );
and ( n8149 , n7730 , n7735 );
and ( n8150 , n7726 , n7735 );
or ( n8151 , n8148 , n8149 , n8150 );
xor ( n8152 , n8147 , n8151 );
xor ( n8153 , n8138 , n8152 );
and ( n8154 , n5487 , n4752 );
and ( n8155 , n5791 , n4579 );
nor ( n8156 , n8154 , n8155 );
xnor ( n8157 , n8156 , n4733 );
not ( n8158 , n8157 );
and ( n8159 , n4568 , n5773 );
and ( n8160 , n4724 , n5519 );
nor ( n8161 , n8159 , n8160 );
xnor ( n8162 , n8161 , n5763 );
xor ( n8163 , n8158 , n8162 );
and ( n8164 , n4160 , n6496 );
and ( n8165 , n4243 , n6115 );
nor ( n8166 , n8164 , n8165 );
xnor ( n8167 , n8166 , n6453 );
xor ( n8168 , n8163 , n8167 );
xor ( n8169 , n8153 , n8168 );
xor ( n8170 , n8134 , n8169 );
xor ( n8171 , n8106 , n8170 );
xor ( n8172 , n8100 , n8171 );
and ( n8173 , n7675 , n7744 );
and ( n8174 , n7745 , n7748 );
or ( n8175 , n8173 , n8174 );
xor ( n8176 , n8172 , n8175 );
buf ( n8177 , n8176 );
buf ( n8178 , n8177 );
buf ( n8179 , n8178 );
and ( n8180 , n8179 , n4232 );
nor ( n8181 , n8096 , n8180 );
xnor ( n8182 , n8181 , n4230 );
xor ( n8183 , n8095 , n8182 );
and ( n8184 , n7785 , n7789 );
and ( n8185 , n7789 , n7808 );
and ( n8186 , n7785 , n7808 );
or ( n8187 , n8184 , n8185 , n8186 );
and ( n8188 , n6168 , n4298 );
and ( n8189 , n6516 , n4287 );
nor ( n8190 , n8188 , n8189 );
xnor ( n8191 , n8190 , n4294 );
xor ( n8192 , n8187 , n8191 );
and ( n8193 , n5535 , n4788 );
and ( n8194 , n5818 , n4611 );
nor ( n8195 , n8193 , n8194 );
xnor ( n8196 , n8195 , n4784 );
xor ( n8197 , n8192 , n8196 );
xor ( n8198 , n8183 , n8197 );
xor ( n8199 , n8091 , n8198 );
and ( n8200 , n7760 , n7764 );
and ( n8201 , n7764 , n7769 );
and ( n8202 , n7760 , n7769 );
or ( n8203 , n8200 , n8201 , n8202 );
and ( n8204 , n6907 , n4319 );
and ( n8205 , n7324 , n4310 );
nor ( n8206 , n8204 , n8205 );
xnor ( n8207 , n8206 , n4315 );
xor ( n8208 , n8203 , n8207 );
and ( n8209 , n7794 , n7798 );
and ( n8210 , n7798 , n7807 );
and ( n8211 , n7794 , n7807 );
or ( n8212 , n8209 , n8210 , n8211 );
and ( n8213 , n4999 , n5270 );
and ( n8214 , n5247 , n5021 );
nor ( n8215 , n8213 , n8214 );
xnor ( n8216 , n8215 , n5266 );
xor ( n8217 , n8212 , n8216 );
and ( n8218 , n4594 , n5850 );
and ( n8219 , n4770 , n5566 );
nor ( n8220 , n8218 , n8219 );
xnor ( n8221 , n8220 , n5846 );
and ( n8222 , n4228 , n6554 );
and ( n8223 , n4275 , n6205 );
nor ( n8224 , n8222 , n8223 );
xnor ( n8225 , n8224 , n6550 );
xor ( n8226 , n8221 , n8225 );
and ( n8227 , n7800 , n7804 );
and ( n8228 , n7804 , n7806 );
and ( n8229 , n7800 , n7806 );
or ( n8230 , n8227 , n8228 , n8229 );
and ( n8231 , n4329 , n7356 );
and ( n8232 , n4342 , n6953 );
nor ( n8233 , n8231 , n8232 );
xnor ( n8234 , n8233 , n7352 );
xor ( n8235 , n8230 , n8234 );
and ( n8236 , n4303 , n7349 );
xor ( n8237 , n8235 , n8236 );
xor ( n8238 , n8226 , n8237 );
xor ( n8239 , n8217 , n8238 );
xor ( n8240 , n8208 , n8239 );
xor ( n8241 , n8199 , n8240 );
and ( n8242 , n7666 , n7771 );
and ( n8243 , n7771 , n7810 );
and ( n8244 , n7666 , n7810 );
or ( n8245 , n8242 , n8243 , n8244 );
xor ( n8246 , n8241 , n8245 );
and ( n8247 , n7811 , n7815 );
and ( n8248 , n7816 , n7819 );
or ( n8249 , n8247 , n8248 );
xor ( n8250 , n8246 , n8249 );
buf ( n8251 , n8250 );
and ( n8252 , n4411 , n6627 );
and ( n8253 , n4421 , n6272 );
nor ( n8254 , n8252 , n8253 );
xnor ( n8255 , n8254 , n6623 );
and ( n8256 , n4427 , n7444 );
and ( n8257 , n4436 , n7026 );
nor ( n8258 , n8256 , n8257 );
xnor ( n8259 , n8258 , n7440 );
xor ( n8260 , n8255 , n8259 );
and ( n8261 , n4405 , n7437 );
xor ( n8262 , n8260 , n8261 );
and ( n8263 , n6995 , n4433 );
and ( n8264 , n7417 , n4431 );
nor ( n8265 , n8263 , n8264 );
xnor ( n8266 , n8265 , n4441 );
and ( n8267 , n6235 , n4402 );
and ( n8268 , n6604 , n4391 );
nor ( n8269 , n8267 , n8268 );
xnor ( n8270 , n8269 , n4398 );
xor ( n8271 , n8266 , n8270 );
and ( n8272 , n4631 , n5922 );
and ( n8273 , n4817 , n5616 );
nor ( n8274 , n8272 , n8273 );
xnor ( n8275 , n8274 , n5918 );
xor ( n8276 , n8271 , n8275 );
xor ( n8277 , n8262 , n8276 );
and ( n8278 , n7880 , n7884 );
and ( n8279 , n7884 , n7886 );
and ( n8280 , n7880 , n7886 );
or ( n8281 , n8278 , n8279 , n8280 );
xor ( n8282 , n8277 , n8281 );
and ( n8283 , n7829 , n7833 );
and ( n8284 , n7833 , n7848 );
and ( n8285 , n7829 , n7848 );
or ( n8286 , n8283 , n8284 , n8285 );
xor ( n8287 , n8282 , n8286 );
and ( n8288 , n7865 , n7869 );
and ( n8289 , n7869 , n7888 );
and ( n8290 , n7865 , n7888 );
or ( n8291 , n8288 , n8289 , n8290 );
xor ( n8292 , n8287 , n8291 );
and ( n8293 , n7854 , n7860 );
and ( n8294 , n7860 , n7889 );
and ( n8295 , n7854 , n7889 );
or ( n8296 , n8293 , n8294 , n8295 );
and ( n8297 , n7838 , n7842 );
and ( n8298 , n7842 , n7847 );
and ( n8299 , n7838 , n7847 );
or ( n8300 , n8297 , n8298 , n8299 );
and ( n8301 , n7857 , n4418 );
buf ( n8302 , n3112 );
buf ( n8303 , n8302 );
and ( n8304 , n8303 , n4415 );
nor ( n8305 , n8301 , n8304 );
xnor ( n8306 , n8305 , n4413 );
xor ( n8307 , n8300 , n8306 );
and ( n8308 , n7874 , n7878 );
and ( n8309 , n7878 , n7887 );
and ( n8310 , n7874 , n7887 );
or ( n8311 , n8308 , n8309 , n8310 );
and ( n8312 , n5588 , n4835 );
and ( n8313 , n5893 , n4648 );
nor ( n8314 , n8312 , n8313 );
xnor ( n8315 , n8314 , n4831 );
xor ( n8316 , n8311 , n8315 );
and ( n8317 , n5042 , n5323 );
and ( n8318 , n5300 , n5064 );
nor ( n8319 , n8317 , n8318 );
xnor ( n8320 , n8319 , n5319 );
xor ( n8321 , n8316 , n8320 );
xor ( n8322 , n8307 , n8321 );
xor ( n8323 , n8296 , n8322 );
xor ( n8324 , n8292 , n8323 );
and ( n8325 , n7825 , n7849 );
and ( n8326 , n7849 , n7890 );
and ( n8327 , n7825 , n7890 );
or ( n8328 , n8325 , n8326 , n8327 );
xor ( n8329 , n8324 , n8328 );
and ( n8330 , n7891 , n7895 );
and ( n8331 , n7896 , n7899 );
or ( n8332 , n8330 , n8331 );
xor ( n8333 , n8329 , n8332 );
buf ( n8334 , n8333 );
not ( n8335 , n454 );
and ( n8336 , n8335 , n8251 );
and ( n8337 , n8334 , n454 );
or ( n8338 , n8336 , n8337 );
buf ( n8339 , n8338 );
buf ( n8340 , n8339 );
and ( n8341 , n8340 , n4505 );
xor ( n8342 , n8087 , n8341 );
and ( n8343 , n7048 , n5089 );
and ( n8344 , n7474 , n4866 );
xor ( n8345 , n8343 , n8344 );
and ( n8346 , n7907 , n4557 );
xor ( n8347 , n8345 , n8346 );
xor ( n8348 , n8342 , n8347 );
and ( n8349 , n7662 , n7908 );
and ( n8350 , n7908 , n7914 );
and ( n8351 , n7662 , n7914 );
or ( n8352 , n8349 , n8350 , n8351 );
xor ( n8353 , n8348 , n8352 );
and ( n8354 , n7915 , n7919 );
and ( n8355 , n7919 , n7924 );
and ( n8356 , n7915 , n7924 );
or ( n8357 , n8354 , n8355 , n8356 );
xor ( n8358 , n8353 , n8357 );
or ( n8359 , n7925 , n7926 );
xnor ( n8360 , n8358 , n8359 );
and ( n8361 , n7927 , n7928 );
xor ( n8362 , n8360 , n8361 );
buf ( n8363 , n8362 );
not ( n8364 , n4509 );
and ( n8365 , n8364 , n8083 );
and ( n8366 , n8363 , n4509 );
or ( n8367 , n8365 , n8366 );
and ( n8368 , n7974 , n7978 );
and ( n8369 , n7978 , n8077 );
and ( n8370 , n7974 , n8077 );
or ( n8371 , n8368 , n8369 , n8370 );
and ( n8372 , n8057 , n4524 );
not ( n8373 , n8043 );
buf ( n8374 , n2217 );
buf ( n8375 , n8374 );
and ( n8376 , n8041 , n7552 );
not ( n8377 , n8376 );
and ( n8378 , n8375 , n8377 );
and ( n8379 , n8373 , n8378 );
xor ( n8380 , n8375 , n8041 );
not ( n8381 , n8042 );
and ( n8382 , n8380 , n8381 );
and ( n8383 , n4132 , n8382 );
and ( n8384 , n4539 , n8042 );
nor ( n8385 , n8383 , n8384 );
xnor ( n8386 , n8385 , n8378 );
xor ( n8387 , n8379 , n8386 );
and ( n8388 , n5121 , n6761 );
and ( n8389 , n5387 , n6379 );
nor ( n8390 , n8388 , n8389 );
xnor ( n8391 , n8390 , n6757 );
xor ( n8392 , n8387 , n8391 );
and ( n8393 , n4683 , n7559 );
and ( n8394 , n4890 , n7107 );
nor ( n8395 , n8393 , n8394 );
xnor ( n8396 , n8395 , n7555 );
xor ( n8397 , n8392 , n8396 );
and ( n8398 , n8001 , n4530 );
buf ( n8399 , n491 );
buf ( n8400 , n507 );
xor ( n8401 , n8399 , n8400 );
and ( n8402 , n7991 , n7992 );
and ( n8403 , n7992 , n7997 );
and ( n8404 , n7991 , n7997 );
or ( n8405 , n8402 , n8403 , n8404 );
xor ( n8406 , n8401 , n8405 );
buf ( n8407 , n8406 );
buf ( n8408 , n8407 );
buf ( n8409 , n8408 );
and ( n8410 , n8409 , n4134 );
nor ( n8411 , n8398 , n8410 );
xnor ( n8412 , n8411 , n4527 );
and ( n8413 , n6353 , n5405 );
and ( n8414 , n6748 , n5132 );
nor ( n8415 , n8413 , n8414 );
xnor ( n8416 , n8415 , n5401 );
xor ( n8417 , n8412 , n8416 );
and ( n8418 , n8017 , n8021 );
and ( n8419 , n8021 , n8026 );
and ( n8420 , n8017 , n8026 );
or ( n8421 , n8418 , n8419 , n8420 );
xor ( n8422 , n8417 , n8421 );
xor ( n8423 , n8397 , n8422 );
and ( n8424 , n8034 , n8038 );
and ( n8425 , n8038 , n8043 );
and ( n8426 , n8034 , n8043 );
or ( n8427 , n8424 , n8425 , n8426 );
and ( n8428 , n7092 , n4898 );
and ( n8429 , n7531 , n4689 );
nor ( n8430 , n8428 , n8429 );
xnor ( n8431 , n8430 , n4904 );
xor ( n8432 , n8427 , n8431 );
and ( n8433 , n5672 , n6008 );
and ( n8434 , n5995 , n5689 );
nor ( n8435 , n8433 , n8434 );
xnor ( n8436 , n8435 , n6004 );
xor ( n8437 , n8432 , n8436 );
xor ( n8438 , n8423 , n8437 );
and ( n8439 , n7984 , n7988 );
and ( n8440 , n7988 , n8046 );
and ( n8441 , n7984 , n8046 );
or ( n8442 , n8439 , n8440 , n8441 );
xor ( n8443 , n8438 , n8442 );
and ( n8444 , n8008 , n8012 );
and ( n8445 , n8012 , n8027 );
and ( n8446 , n8008 , n8027 );
or ( n8447 , n8444 , n8445 , n8446 );
and ( n8448 , n8033 , n8044 );
xor ( n8449 , n8447 , n8448 );
and ( n8450 , n8004 , n8028 );
and ( n8451 , n8028 , n8045 );
and ( n8452 , n8004 , n8045 );
or ( n8453 , n8450 , n8451 , n8452 );
xor ( n8454 , n8449 , n8453 );
xor ( n8455 , n8443 , n8454 );
and ( n8456 , n8047 , n8051 );
and ( n8457 , n8052 , n8053 );
or ( n8458 , n8456 , n8457 );
xor ( n8459 , n8455 , n8458 );
buf ( n8460 , n8459 );
buf ( n8461 , n8460 );
buf ( n8462 , n8461 );
and ( n8463 , n8462 , n4145 );
nor ( n8464 , n8372 , n8463 );
xnor ( n8465 , n8464 , n4521 );
and ( n8466 , n6391 , n5441 );
and ( n8467 , n6796 , n5161 );
nor ( n8468 , n8466 , n8467 );
xnor ( n8469 , n8468 , n5437 );
and ( n8470 , n5700 , n6068 );
and ( n8471 , n6037 , n5730 );
nor ( n8472 , n8470 , n8471 );
xnor ( n8473 , n8472 , n6064 );
xor ( n8474 , n8469 , n8473 );
and ( n8475 , n7947 , n7951 );
and ( n8476 , n7951 , n7972 );
and ( n8477 , n7947 , n7972 );
or ( n8478 , n8475 , n8476 , n8477 );
and ( n8479 , n5140 , n6711 );
and ( n8480 , n5419 , n6332 );
nor ( n8481 , n8479 , n8480 );
xnor ( n8482 , n8481 , n6707 );
xor ( n8483 , n8478 , n8482 );
not ( n8484 , n7971 );
buf ( n8485 , n523 );
buf ( n8486 , n539 );
xor ( n8487 , n8485 , n8486 );
and ( n8488 , n7959 , n7960 );
and ( n8489 , n7960 , n7965 );
and ( n8490 , n7959 , n7965 );
or ( n8491 , n8488 , n8489 , n8490 );
xor ( n8492 , n8487 , n8491 );
buf ( n8493 , n8492 );
buf ( n8494 , n8493 );
buf ( n8495 , n8494 );
and ( n8496 , n7969 , n7623 );
not ( n8497 , n8496 );
and ( n8498 , n8495 , n8497 );
and ( n8499 , n8484 , n8498 );
xor ( n8500 , n8495 , n7969 );
not ( n8501 , n7970 );
and ( n8502 , n8500 , n8501 );
and ( n8503 , n4139 , n8502 );
and ( n8504 , n4548 , n7970 );
nor ( n8505 , n8503 , n8504 );
xnor ( n8506 , n8505 , n8498 );
xor ( n8507 , n8499 , n8506 );
and ( n8508 , n7953 , n7957 );
and ( n8509 , n7957 , n7971 );
and ( n8510 , n7953 , n7971 );
or ( n8511 , n8508 , n8509 , n8510 );
xor ( n8512 , n8507 , n8511 );
and ( n8513 , n4696 , n7630 );
and ( n8514 , n4916 , n7188 );
nor ( n8515 , n8513 , n8514 );
xnor ( n8516 , n8515 , n7626 );
xor ( n8517 , n8512 , n8516 );
xor ( n8518 , n8483 , n8517 );
xor ( n8519 , n8474 , n8518 );
xor ( n8520 , n8465 , n8519 );
xor ( n8521 , n8371 , n8520 );
and ( n8522 , n8060 , n8064 );
and ( n8523 , n8064 , n8069 );
and ( n8524 , n8060 , n8069 );
or ( n8525 , n8522 , n8523 , n8524 );
and ( n8526 , n8070 , n8071 );
and ( n8527 , n8071 , n8076 );
and ( n8528 , n8070 , n8076 );
or ( n8529 , n8526 , n8527 , n8528 );
xor ( n8530 , n8525 , n8529 );
and ( n8531 , n7938 , n7942 );
and ( n8532 , n7942 , n7973 );
and ( n8533 , n7938 , n7973 );
or ( n8534 , n8531 , n8532 , n8533 );
and ( n8535 , n7146 , n4938 );
and ( n8536 , n7587 , n4711 );
nor ( n8537 , n8535 , n8536 );
xnor ( n8538 , n8537 , n4934 );
xor ( n8539 , n8534 , n8538 );
xor ( n8540 , n8530 , n8539 );
xor ( n8541 , n8521 , n8540 );
and ( n8542 , n8078 , n8081 );
xor ( n8543 , n8541 , n8542 );
buf ( n8544 , n8543 );
and ( n8545 , n8343 , n8344 );
and ( n8546 , n8344 , n8346 );
and ( n8547 , n8343 , n8346 );
or ( n8548 , n8545 , n8546 , n8547 );
and ( n8549 , n8340 , n4557 );
xor ( n8550 , n8548 , n8549 );
and ( n8551 , n7474 , n5089 );
and ( n8552 , n7907 , n4866 );
xor ( n8553 , n8551 , n8552 );
and ( n8554 , n8095 , n8182 );
and ( n8555 , n8182 , n8197 );
and ( n8556 , n8095 , n8197 );
or ( n8557 , n8554 , n8555 , n8556 );
and ( n8558 , n8179 , n4235 );
and ( n8559 , n8104 , n8105 );
and ( n8560 , n8105 , n8170 );
and ( n8561 , n8104 , n8170 );
or ( n8562 , n8559 , n8560 , n8561 );
and ( n8563 , n8138 , n8152 );
and ( n8564 , n8152 , n8168 );
and ( n8565 , n8138 , n8168 );
or ( n8566 , n8563 , n8564 , n8565 );
and ( n8567 , n8129 , n8133 );
and ( n8568 , n8133 , n8169 );
and ( n8569 , n8129 , n8169 );
or ( n8570 , n8567 , n8568 , n8569 );
xor ( n8571 , n8566 , n8570 );
and ( n8572 , n8120 , n8128 );
and ( n8573 , n8142 , n8146 );
and ( n8574 , n8146 , n8151 );
and ( n8575 , n8142 , n8151 );
or ( n8576 , n8573 , n8574 , n8575 );
and ( n8577 , n6444 , n4262 );
and ( n8578 , n6853 , n4188 );
nor ( n8579 , n8577 , n8578 );
xnor ( n8580 , n8579 , n4252 );
and ( n8581 , n5195 , n5208 );
and ( n8582 , n5487 , n4976 );
nor ( n8583 , n8581 , n8582 );
xnor ( n8584 , n8583 , n5214 );
xor ( n8585 , n8580 , n8584 );
and ( n8586 , n4176 , n7274 );
xor ( n8587 , n8585 , n8586 );
xor ( n8588 , n8576 , n8587 );
buf ( n8589 , n8157 );
and ( n8590 , n7299 , n4173 );
not ( n8591 , n8590 );
xnor ( n8592 , n8591 , n4181 );
not ( n8593 , n8592 );
xor ( n8594 , n8589 , n8593 );
and ( n8595 , n4150 , n7277 );
and ( n8596 , n4160 , n6864 );
nor ( n8597 , n8595 , n8596 );
xnor ( n8598 , n8597 , n7283 );
xor ( n8599 , n8594 , n8598 );
xor ( n8600 , n8588 , n8599 );
xor ( n8601 , n8572 , n8600 );
and ( n8602 , n8158 , n8162 );
and ( n8603 , n8162 , n8167 );
and ( n8604 , n8158 , n8167 );
or ( n8605 , n8602 , n8603 , n8604 );
and ( n8606 , n8110 , n8114 );
and ( n8607 , n8114 , n8119 );
and ( n8608 , n8110 , n8119 );
or ( n8609 , n8606 , n8607 , n8608 );
and ( n8610 , n8121 , n8125 );
and ( n8611 , n8125 , n8127 );
and ( n8612 , n8121 , n8127 );
or ( n8613 , n8610 , n8611 , n8612 );
xor ( n8614 , n8609 , n8613 );
and ( n8615 , n5791 , n4752 );
and ( n8616 , n6120 , n4579 );
nor ( n8617 , n8615 , n8616 );
xnor ( n8618 , n8617 , n4733 );
and ( n8619 , n4724 , n5773 );
and ( n8620 , n4965 , n5519 );
nor ( n8621 , n8619 , n8620 );
xnor ( n8622 , n8621 , n5763 );
xor ( n8623 , n8618 , n8622 );
and ( n8624 , n4243 , n6496 );
and ( n8625 , n4568 , n6115 );
nor ( n8626 , n8624 , n8625 );
xnor ( n8627 , n8626 , n6453 );
xor ( n8628 , n8623 , n8627 );
xor ( n8629 , n8614 , n8628 );
xor ( n8630 , n8605 , n8629 );
xor ( n8631 , n8601 , n8630 );
xor ( n8632 , n8571 , n8631 );
xor ( n8633 , n8562 , n8632 );
and ( n8634 , n8100 , n8171 );
and ( n8635 , n8172 , n8175 );
or ( n8636 , n8634 , n8635 );
xor ( n8637 , n8633 , n8636 );
buf ( n8638 , n8637 );
buf ( n8639 , n8638 );
buf ( n8640 , n8639 );
and ( n8641 , n8640 , n4232 );
nor ( n8642 , n8558 , n8641 );
xnor ( n8643 , n8642 , n4230 );
and ( n8644 , n7324 , n4319 );
and ( n8645 , n7752 , n4310 );
nor ( n8646 , n8644 , n8645 );
xnor ( n8647 , n8646 , n4315 );
xor ( n8648 , n8643 , n8647 );
and ( n8649 , n8221 , n8225 );
and ( n8650 , n8225 , n8237 );
and ( n8651 , n8221 , n8237 );
or ( n8652 , n8649 , n8650 , n8651 );
and ( n8653 , n5818 , n4788 );
and ( n8654 , n6168 , n4611 );
nor ( n8655 , n8653 , n8654 );
xnor ( n8656 , n8655 , n4784 );
xor ( n8657 , n8652 , n8656 );
and ( n8658 , n5247 , n5270 );
and ( n8659 , n5535 , n5021 );
nor ( n8660 , n8658 , n8659 );
xnor ( n8661 , n8660 , n5266 );
xor ( n8662 , n8657 , n8661 );
xor ( n8663 , n8648 , n8662 );
xor ( n8664 , n8557 , n8663 );
and ( n8665 , n8187 , n8191 );
and ( n8666 , n8191 , n8196 );
and ( n8667 , n8187 , n8196 );
or ( n8668 , n8665 , n8666 , n8667 );
and ( n8669 , n8203 , n8207 );
and ( n8670 , n8207 , n8239 );
and ( n8671 , n8203 , n8239 );
or ( n8672 , n8669 , n8670 , n8671 );
xor ( n8673 , n8668 , n8672 );
and ( n8674 , n8212 , n8216 );
and ( n8675 , n8216 , n8238 );
and ( n8676 , n8212 , n8238 );
or ( n8677 , n8674 , n8675 , n8676 );
and ( n8678 , n6516 , n4298 );
and ( n8679 , n6907 , n4287 );
nor ( n8680 , n8678 , n8679 );
xnor ( n8681 , n8680 , n4294 );
xor ( n8682 , n8677 , n8681 );
and ( n8683 , n8230 , n8234 );
and ( n8684 , n8234 , n8236 );
and ( n8685 , n8230 , n8236 );
or ( n8686 , n8683 , n8684 , n8685 );
and ( n8687 , n4770 , n5850 );
and ( n8688 , n4999 , n5566 );
nor ( n8689 , n8687 , n8688 );
xnor ( n8690 , n8689 , n5846 );
xor ( n8691 , n8686 , n8690 );
and ( n8692 , n4275 , n6554 );
and ( n8693 , n4594 , n6205 );
nor ( n8694 , n8692 , n8693 );
xnor ( n8695 , n8694 , n6550 );
and ( n8696 , n4342 , n7356 );
and ( n8697 , n4228 , n6953 );
nor ( n8698 , n8696 , n8697 );
xnor ( n8699 , n8698 , n7352 );
xor ( n8700 , n8695 , n8699 );
and ( n8701 , n4329 , n7349 );
xor ( n8702 , n8700 , n8701 );
xor ( n8703 , n8691 , n8702 );
xor ( n8704 , n8682 , n8703 );
xor ( n8705 , n8673 , n8704 );
xor ( n8706 , n8664 , n8705 );
and ( n8707 , n8091 , n8198 );
and ( n8708 , n8198 , n8240 );
and ( n8709 , n8091 , n8240 );
or ( n8710 , n8707 , n8708 , n8709 );
xor ( n8711 , n8706 , n8710 );
and ( n8712 , n8241 , n8245 );
and ( n8713 , n8246 , n8249 );
or ( n8714 , n8712 , n8713 );
xor ( n8715 , n8711 , n8714 );
buf ( n8716 , n8715 );
and ( n8717 , n8296 , n8322 );
and ( n8718 , n8300 , n8306 );
and ( n8719 , n8306 , n8321 );
and ( n8720 , n8300 , n8321 );
or ( n8721 , n8718 , n8719 , n8720 );
and ( n8722 , n8262 , n8276 );
and ( n8723 , n8276 , n8281 );
and ( n8724 , n8262 , n8281 );
or ( n8725 , n8722 , n8723 , n8724 );
and ( n8726 , n8303 , n4418 );
buf ( n8727 , n3251 );
buf ( n8728 , n8727 );
and ( n8729 , n8728 , n4415 );
nor ( n8730 , n8726 , n8729 );
xnor ( n8731 , n8730 , n4413 );
and ( n8732 , n7417 , n4433 );
and ( n8733 , n7857 , n4431 );
nor ( n8734 , n8732 , n8733 );
xnor ( n8735 , n8734 , n4441 );
xor ( n8736 , n8731 , n8735 );
and ( n8737 , n6604 , n4402 );
and ( n8738 , n6995 , n4391 );
nor ( n8739 , n8737 , n8738 );
xnor ( n8740 , n8739 , n4398 );
xor ( n8741 , n8736 , n8740 );
and ( n8742 , n5893 , n4835 );
and ( n8743 , n6235 , n4648 );
nor ( n8744 , n8742 , n8743 );
xnor ( n8745 , n8744 , n4831 );
and ( n8746 , n5300 , n5323 );
and ( n8747 , n5588 , n5064 );
nor ( n8748 , n8746 , n8747 );
xnor ( n8749 , n8748 , n5319 );
xor ( n8750 , n8745 , n8749 );
and ( n8751 , n4817 , n5922 );
and ( n8752 , n5042 , n5616 );
nor ( n8753 , n8751 , n8752 );
xnor ( n8754 , n8753 , n5918 );
xor ( n8755 , n8750 , n8754 );
xor ( n8756 , n8741 , n8755 );
and ( n8757 , n4421 , n6627 );
and ( n8758 , n4631 , n6272 );
nor ( n8759 , n8757 , n8758 );
xnor ( n8760 , n8759 , n6623 );
and ( n8761 , n4436 , n7444 );
and ( n8762 , n4411 , n7026 );
nor ( n8763 , n8761 , n8762 );
xnor ( n8764 , n8763 , n7440 );
xor ( n8765 , n8760 , n8764 );
and ( n8766 , n4427 , n7437 );
xor ( n8767 , n8765 , n8766 );
and ( n8768 , n8255 , n8259 );
and ( n8769 , n8259 , n8261 );
and ( n8770 , n8255 , n8261 );
or ( n8771 , n8768 , n8769 , n8770 );
xor ( n8772 , n8767 , n8771 );
and ( n8773 , n8266 , n8270 );
and ( n8774 , n8270 , n8275 );
and ( n8775 , n8266 , n8275 );
or ( n8776 , n8773 , n8774 , n8775 );
xor ( n8777 , n8772 , n8776 );
xor ( n8778 , n8756 , n8777 );
xor ( n8779 , n8725 , n8778 );
and ( n8780 , n8311 , n8315 );
and ( n8781 , n8315 , n8320 );
and ( n8782 , n8311 , n8320 );
or ( n8783 , n8780 , n8781 , n8782 );
xor ( n8784 , n8779 , n8783 );
xor ( n8785 , n8721 , n8784 );
and ( n8786 , n8282 , n8286 );
and ( n8787 , n8286 , n8291 );
and ( n8788 , n8282 , n8291 );
or ( n8789 , n8786 , n8787 , n8788 );
xor ( n8790 , n8785 , n8789 );
xor ( n8791 , n8717 , n8790 );
and ( n8792 , n8292 , n8323 );
and ( n8793 , n8323 , n8328 );
and ( n8794 , n8292 , n8328 );
or ( n8795 , n8792 , n8793 , n8794 );
xor ( n8796 , n8791 , n8795 );
and ( n8797 , n8329 , n8332 );
xor ( n8798 , n8796 , n8797 );
buf ( n8799 , n8798 );
not ( n8800 , n454 );
and ( n8801 , n8800 , n8716 );
and ( n8802 , n8799 , n454 );
or ( n8803 , n8801 , n8802 );
buf ( n8804 , n8803 );
buf ( n8805 , n8804 );
and ( n8806 , n8805 , n4505 );
xor ( n8807 , n8553 , n8806 );
xor ( n8808 , n8550 , n8807 );
and ( n8809 , n8087 , n8341 );
and ( n8810 , n8341 , n8347 );
and ( n8811 , n8087 , n8347 );
or ( n8812 , n8809 , n8810 , n8811 );
xor ( n8813 , n8808 , n8812 );
and ( n8814 , n8348 , n8352 );
and ( n8815 , n8352 , n8357 );
and ( n8816 , n8348 , n8357 );
or ( n8817 , n8814 , n8815 , n8816 );
xor ( n8818 , n8813 , n8817 );
or ( n8819 , n8358 , n8359 );
xnor ( n8820 , n8818 , n8819 );
and ( n8821 , n8360 , n8361 );
xor ( n8822 , n8820 , n8821 );
buf ( n8823 , n8822 );
not ( n8824 , n4509 );
and ( n8825 , n8824 , n8544 );
and ( n8826 , n8823 , n4509 );
or ( n8827 , n8825 , n8826 );
and ( n8828 , n8478 , n8482 );
and ( n8829 , n8482 , n8517 );
and ( n8830 , n8478 , n8517 );
or ( n8831 , n8828 , n8829 , n8830 );
and ( n8832 , n6796 , n5441 );
and ( n8833 , n7146 , n5161 );
nor ( n8834 , n8832 , n8833 );
xnor ( n8835 , n8834 , n5437 );
xor ( n8836 , n8831 , n8835 );
and ( n8837 , n6037 , n6068 );
and ( n8838 , n6391 , n5730 );
nor ( n8839 , n8837 , n8838 );
xnor ( n8840 , n8839 , n6064 );
and ( n8841 , n5419 , n6711 );
and ( n8842 , n5700 , n6332 );
nor ( n8843 , n8841 , n8842 );
xnor ( n8844 , n8843 , n6707 );
xor ( n8845 , n8840 , n8844 );
and ( n8846 , n8507 , n8511 );
and ( n8847 , n8511 , n8516 );
and ( n8848 , n8507 , n8516 );
or ( n8849 , n8846 , n8847 , n8848 );
and ( n8850 , n4916 , n7630 );
and ( n8851 , n5140 , n7188 );
nor ( n8852 , n8850 , n8851 );
xnor ( n8853 , n8852 , n7626 );
xor ( n8854 , n8849 , n8853 );
and ( n8855 , n8499 , n8506 );
and ( n8856 , n4548 , n8502 );
and ( n8857 , n4696 , n7970 );
nor ( n8858 , n8856 , n8857 );
xnor ( n8859 , n8858 , n8498 );
xor ( n8860 , n8855 , n8859 );
buf ( n8861 , n522 );
buf ( n8862 , n538 );
xor ( n8863 , n8861 , n8862 );
and ( n8864 , n8485 , n8486 );
and ( n8865 , n8486 , n8491 );
and ( n8866 , n8485 , n8491 );
or ( n8867 , n8864 , n8865 , n8866 );
xor ( n8868 , n8863 , n8867 );
buf ( n8869 , n8868 );
buf ( n8870 , n8869 );
buf ( n8871 , n8870 );
xor ( n8872 , n8871 , n8495 );
and ( n8873 , n4139 , n8872 );
xor ( n8874 , n8860 , n8873 );
xor ( n8875 , n8854 , n8874 );
xor ( n8876 , n8845 , n8875 );
xor ( n8877 , n8836 , n8876 );
and ( n8878 , n8534 , n8538 );
xor ( n8879 , n8877 , n8878 );
and ( n8880 , n8469 , n8473 );
and ( n8881 , n8473 , n8518 );
and ( n8882 , n8469 , n8518 );
or ( n8883 , n8880 , n8881 , n8882 );
and ( n8884 , n8462 , n4524 );
and ( n8885 , n8438 , n8442 );
and ( n8886 , n8442 , n8454 );
and ( n8887 , n8438 , n8454 );
or ( n8888 , n8885 , n8886 , n8887 );
and ( n8889 , n8409 , n4530 );
buf ( n8890 , n490 );
buf ( n8891 , n506 );
xor ( n8892 , n8890 , n8891 );
and ( n8893 , n8399 , n8400 );
and ( n8894 , n8400 , n8405 );
and ( n8895 , n8399 , n8405 );
or ( n8896 , n8893 , n8894 , n8895 );
xor ( n8897 , n8892 , n8896 );
buf ( n8898 , n8897 );
buf ( n8899 , n8898 );
buf ( n8900 , n8899 );
and ( n8901 , n8900 , n4134 );
nor ( n8902 , n8889 , n8901 );
xnor ( n8903 , n8902 , n4527 );
and ( n8904 , n8412 , n8416 );
and ( n8905 , n8416 , n8421 );
and ( n8906 , n8412 , n8421 );
or ( n8907 , n8904 , n8905 , n8906 );
xor ( n8908 , n8903 , n8907 );
and ( n8909 , n8387 , n8391 );
and ( n8910 , n8391 , n8396 );
and ( n8911 , n8387 , n8396 );
or ( n8912 , n8909 , n8910 , n8911 );
and ( n8913 , n6748 , n5405 );
and ( n8914 , n7092 , n5132 );
nor ( n8915 , n8913 , n8914 );
xnor ( n8916 , n8915 , n5401 );
xor ( n8917 , n8912 , n8916 );
and ( n8918 , n5995 , n6008 );
and ( n8919 , n6353 , n5689 );
nor ( n8920 , n8918 , n8919 );
xnor ( n8921 , n8920 , n6004 );
and ( n8922 , n5387 , n6761 );
and ( n8923 , n5672 , n6379 );
nor ( n8924 , n8922 , n8923 );
xnor ( n8925 , n8924 , n6757 );
xor ( n8926 , n8921 , n8925 );
and ( n8927 , n4890 , n7559 );
and ( n8928 , n5121 , n7107 );
nor ( n8929 , n8927 , n8928 );
xnor ( n8930 , n8929 , n7555 );
xor ( n8931 , n8926 , n8930 );
xor ( n8932 , n8917 , n8931 );
xor ( n8933 , n8908 , n8932 );
and ( n8934 , n8447 , n8448 );
and ( n8935 , n8448 , n8453 );
and ( n8936 , n8447 , n8453 );
or ( n8937 , n8934 , n8935 , n8936 );
xor ( n8938 , n8933 , n8937 );
and ( n8939 , n7531 , n4898 );
and ( n8940 , n8001 , n4689 );
nor ( n8941 , n8939 , n8940 );
xnor ( n8942 , n8941 , n4904 );
and ( n8943 , n8379 , n8386 );
and ( n8944 , n4539 , n8382 );
and ( n8945 , n4683 , n8042 );
nor ( n8946 , n8944 , n8945 );
xnor ( n8947 , n8946 , n8378 );
xor ( n8948 , n8943 , n8947 );
and ( n8949 , n4132 , n8375 );
xor ( n8950 , n8948 , n8949 );
xor ( n8951 , n8942 , n8950 );
and ( n8952 , n8427 , n8431 );
and ( n8953 , n8431 , n8436 );
and ( n8954 , n8427 , n8436 );
or ( n8955 , n8952 , n8953 , n8954 );
xor ( n8956 , n8951 , n8955 );
and ( n8957 , n8397 , n8422 );
and ( n8958 , n8422 , n8437 );
and ( n8959 , n8397 , n8437 );
or ( n8960 , n8957 , n8958 , n8959 );
xor ( n8961 , n8956 , n8960 );
xor ( n8962 , n8938 , n8961 );
xor ( n8963 , n8888 , n8962 );
and ( n8964 , n8455 , n8458 );
xor ( n8965 , n8963 , n8964 );
buf ( n8966 , n8965 );
buf ( n8967 , n8966 );
buf ( n8968 , n8967 );
and ( n8969 , n8968 , n4145 );
nor ( n8970 , n8884 , n8969 );
xnor ( n8971 , n8970 , n4521 );
xor ( n8972 , n8883 , n8971 );
and ( n8973 , n7587 , n4938 );
and ( n8974 , n8057 , n4711 );
nor ( n8975 , n8973 , n8974 );
xnor ( n8976 , n8975 , n4934 );
xor ( n8977 , n8972 , n8976 );
xor ( n8978 , n8879 , n8977 );
and ( n8979 , n8465 , n8519 );
and ( n8980 , n8525 , n8529 );
and ( n8981 , n8529 , n8539 );
and ( n8982 , n8525 , n8539 );
or ( n8983 , n8980 , n8981 , n8982 );
xor ( n8984 , n8979 , n8983 );
and ( n8985 , n8371 , n8520 );
and ( n8986 , n8520 , n8540 );
and ( n8987 , n8371 , n8540 );
or ( n8988 , n8985 , n8986 , n8987 );
xor ( n8989 , n8984 , n8988 );
xor ( n8990 , n8978 , n8989 );
and ( n8991 , n8541 , n8542 );
xor ( n8992 , n8990 , n8991 );
buf ( n8993 , n8992 );
and ( n8994 , n8551 , n8552 );
and ( n8995 , n8552 , n8806 );
and ( n8996 , n8551 , n8806 );
or ( n8997 , n8994 , n8995 , n8996 );
and ( n8998 , n8668 , n8672 );
and ( n8999 , n8672 , n8704 );
and ( n9000 , n8668 , n8704 );
or ( n9001 , n8998 , n8999 , n9000 );
and ( n9002 , n8677 , n8681 );
and ( n9003 , n8681 , n8703 );
and ( n9004 , n8677 , n8703 );
or ( n9005 , n9002 , n9003 , n9004 );
and ( n9006 , n7752 , n4319 );
and ( n9007 , n8179 , n4310 );
nor ( n9008 , n9006 , n9007 );
xnor ( n9009 , n9008 , n4315 );
xor ( n9010 , n9005 , n9009 );
and ( n9011 , n8686 , n8690 );
and ( n9012 , n8690 , n8702 );
and ( n9013 , n8686 , n8702 );
or ( n9014 , n9011 , n9012 , n9013 );
and ( n9015 , n6168 , n4788 );
and ( n9016 , n6516 , n4611 );
nor ( n9017 , n9015 , n9016 );
xnor ( n9018 , n9017 , n4784 );
xor ( n9019 , n9014 , n9018 );
and ( n9020 , n5535 , n5270 );
and ( n9021 , n5818 , n5021 );
nor ( n9022 , n9020 , n9021 );
xnor ( n9023 , n9022 , n5266 );
xor ( n9024 , n9019 , n9023 );
xor ( n9025 , n9010 , n9024 );
xor ( n9026 , n9001 , n9025 );
and ( n9027 , n8643 , n8647 );
and ( n9028 , n8647 , n8662 );
and ( n9029 , n8643 , n8662 );
or ( n9030 , n9027 , n9028 , n9029 );
and ( n9031 , n8640 , n4235 );
and ( n9032 , n8566 , n8570 );
and ( n9033 , n8570 , n8631 );
and ( n9034 , n8566 , n8631 );
or ( n9035 , n9032 , n9033 , n9034 );
and ( n9036 , n8605 , n8629 );
and ( n9037 , n8572 , n8600 );
and ( n9038 , n8600 , n8630 );
and ( n9039 , n8572 , n8630 );
or ( n9040 , n9037 , n9038 , n9039 );
xor ( n9041 , n9036 , n9040 );
and ( n9042 , n8589 , n8593 );
and ( n9043 , n8593 , n8598 );
and ( n9044 , n8589 , n8598 );
or ( n9045 , n9042 , n9043 , n9044 );
and ( n9046 , n6120 , n4752 );
and ( n9047 , n6444 , n4579 );
nor ( n9048 , n9046 , n9047 );
xnor ( n9049 , n9048 , n4733 );
and ( n9050 , n4965 , n5773 );
and ( n9051 , n5195 , n5519 );
nor ( n9052 , n9050 , n9051 );
xnor ( n9053 , n9052 , n5763 );
xor ( n9054 , n9049 , n9053 );
and ( n9055 , n4150 , n7274 );
xor ( n9056 , n9054 , n9055 );
xor ( n9057 , n9045 , n9056 );
buf ( n9058 , n8592 );
and ( n9059 , n4568 , n6496 );
and ( n9060 , n4724 , n6115 );
nor ( n9061 , n9059 , n9060 );
xnor ( n9062 , n9061 , n6453 );
xor ( n9063 , n9058 , n9062 );
and ( n9064 , n4160 , n7277 );
and ( n9065 , n4243 , n6864 );
nor ( n9066 , n9064 , n9065 );
xnor ( n9067 , n9066 , n7283 );
xor ( n9068 , n9063 , n9067 );
xor ( n9069 , n9057 , n9068 );
and ( n9070 , n8609 , n8613 );
and ( n9071 , n8613 , n8628 );
and ( n9072 , n8609 , n8628 );
or ( n9073 , n9070 , n9071 , n9072 );
and ( n9074 , n8576 , n8587 );
and ( n9075 , n8587 , n8599 );
and ( n9076 , n8576 , n8599 );
or ( n9077 , n9074 , n9075 , n9076 );
xor ( n9078 , n9073 , n9077 );
and ( n9079 , n8618 , n8622 );
and ( n9080 , n8622 , n8627 );
and ( n9081 , n8618 , n8627 );
or ( n9082 , n9079 , n9080 , n9081 );
and ( n9083 , n8580 , n8584 );
and ( n9084 , n8584 , n8586 );
and ( n9085 , n8580 , n8586 );
or ( n9086 , n9083 , n9084 , n9085 );
xor ( n9087 , n9082 , n9086 );
not ( n9088 , n4181 );
and ( n9089 , n6853 , n4262 );
and ( n9090 , n7299 , n4188 );
nor ( n9091 , n9089 , n9090 );
xnor ( n9092 , n9091 , n4252 );
xor ( n9093 , n9088 , n9092 );
and ( n9094 , n5487 , n5208 );
and ( n9095 , n5791 , n4976 );
nor ( n9096 , n9094 , n9095 );
xnor ( n9097 , n9096 , n5214 );
xor ( n9098 , n9093 , n9097 );
xor ( n9099 , n9087 , n9098 );
xor ( n9100 , n9078 , n9099 );
xor ( n9101 , n9069 , n9100 );
xor ( n9102 , n9041 , n9101 );
xor ( n9103 , n9035 , n9102 );
and ( n9104 , n8562 , n8632 );
and ( n9105 , n8633 , n8636 );
or ( n9106 , n9104 , n9105 );
xor ( n9107 , n9103 , n9106 );
buf ( n9108 , n9107 );
buf ( n9109 , n9108 );
buf ( n9110 , n9109 );
and ( n9111 , n9110 , n4232 );
nor ( n9112 , n9031 , n9111 );
xnor ( n9113 , n9112 , n4230 );
xor ( n9114 , n9030 , n9113 );
and ( n9115 , n8652 , n8656 );
and ( n9116 , n8656 , n8661 );
and ( n9117 , n8652 , n8661 );
or ( n9118 , n9115 , n9116 , n9117 );
and ( n9119 , n6907 , n4298 );
and ( n9120 , n7324 , n4287 );
nor ( n9121 , n9119 , n9120 );
xnor ( n9122 , n9121 , n4294 );
xor ( n9123 , n9118 , n9122 );
and ( n9124 , n8695 , n8699 );
and ( n9125 , n8699 , n8701 );
and ( n9126 , n8695 , n8701 );
or ( n9127 , n9124 , n9125 , n9126 );
and ( n9128 , n4999 , n5850 );
and ( n9129 , n5247 , n5566 );
nor ( n9130 , n9128 , n9129 );
xnor ( n9131 , n9130 , n5846 );
xor ( n9132 , n9127 , n9131 );
and ( n9133 , n4594 , n6554 );
and ( n9134 , n4770 , n6205 );
nor ( n9135 , n9133 , n9134 );
xnor ( n9136 , n9135 , n6550 );
and ( n9137 , n4228 , n7356 );
and ( n9138 , n4275 , n6953 );
nor ( n9139 , n9137 , n9138 );
xnor ( n9140 , n9139 , n7352 );
xor ( n9141 , n9136 , n9140 );
and ( n9142 , n4342 , n7349 );
xor ( n9143 , n9141 , n9142 );
xor ( n9144 , n9132 , n9143 );
xor ( n9145 , n9123 , n9144 );
xor ( n9146 , n9114 , n9145 );
xor ( n9147 , n9026 , n9146 );
and ( n9148 , n8557 , n8663 );
and ( n9149 , n8663 , n8705 );
and ( n9150 , n8557 , n8705 );
or ( n9151 , n9148 , n9149 , n9150 );
xor ( n9152 , n9147 , n9151 );
and ( n9153 , n8706 , n8710 );
and ( n9154 , n8711 , n8714 );
or ( n9155 , n9153 , n9154 );
xor ( n9156 , n9152 , n9155 );
buf ( n9157 , n9156 );
and ( n9158 , n8745 , n8749 );
and ( n9159 , n8749 , n8754 );
and ( n9160 , n8745 , n8754 );
or ( n9161 , n9158 , n9159 , n9160 );
and ( n9162 , n8728 , n4418 );
buf ( n9163 , n3382 );
buf ( n9164 , n9163 );
and ( n9165 , n9164 , n4415 );
nor ( n9166 , n9162 , n9165 );
xnor ( n9167 , n9166 , n4413 );
and ( n9168 , n7857 , n4433 );
and ( n9169 , n8303 , n4431 );
nor ( n9170 , n9168 , n9169 );
xnor ( n9171 , n9170 , n4441 );
xor ( n9172 , n9167 , n9171 );
and ( n9173 , n5588 , n5323 );
and ( n9174 , n5893 , n5064 );
nor ( n9175 , n9173 , n9174 );
xnor ( n9176 , n9175 , n5319 );
xor ( n9177 , n9172 , n9176 );
xor ( n9178 , n9161 , n9177 );
and ( n9179 , n6995 , n4402 );
and ( n9180 , n7417 , n4391 );
nor ( n9181 , n9179 , n9180 );
xnor ( n9182 , n9181 , n4398 );
and ( n9183 , n6235 , n4835 );
and ( n9184 , n6604 , n4648 );
nor ( n9185 , n9183 , n9184 );
xnor ( n9186 , n9185 , n4831 );
xor ( n9187 , n9182 , n9186 );
and ( n9188 , n4631 , n6627 );
and ( n9189 , n4817 , n6272 );
nor ( n9190 , n9188 , n9189 );
xnor ( n9191 , n9190 , n6623 );
and ( n9192 , n4411 , n7444 );
and ( n9193 , n4421 , n7026 );
nor ( n9194 , n9192 , n9193 );
xnor ( n9195 , n9194 , n7440 );
xor ( n9196 , n9191 , n9195 );
and ( n9197 , n4436 , n7437 );
xor ( n9198 , n9196 , n9197 );
xor ( n9199 , n9187 , n9198 );
xor ( n9200 , n9178 , n9199 );
and ( n9201 , n8767 , n8771 );
and ( n9202 , n8771 , n8776 );
and ( n9203 , n8767 , n8776 );
or ( n9204 , n9201 , n9202 , n9203 );
and ( n9205 , n5042 , n5922 );
and ( n9206 , n5300 , n5616 );
nor ( n9207 , n9205 , n9206 );
xnor ( n9208 , n9207 , n5918 );
and ( n9209 , n8760 , n8764 );
and ( n9210 , n8764 , n8766 );
and ( n9211 , n8760 , n8766 );
or ( n9212 , n9209 , n9210 , n9211 );
xor ( n9213 , n9208 , n9212 );
and ( n9214 , n8731 , n8735 );
and ( n9215 , n8735 , n8740 );
and ( n9216 , n8731 , n8740 );
or ( n9217 , n9214 , n9215 , n9216 );
xor ( n9218 , n9213 , n9217 );
xor ( n9219 , n9204 , n9218 );
and ( n9220 , n8741 , n8755 );
and ( n9221 , n8755 , n8777 );
and ( n9222 , n8741 , n8777 );
or ( n9223 , n9220 , n9221 , n9222 );
xor ( n9224 , n9219 , n9223 );
xor ( n9225 , n9200 , n9224 );
and ( n9226 , n8725 , n8778 );
and ( n9227 , n8778 , n8783 );
and ( n9228 , n8725 , n8783 );
or ( n9229 , n9226 , n9227 , n9228 );
xor ( n9230 , n9225 , n9229 );
and ( n9231 , n8721 , n8784 );
and ( n9232 , n8784 , n8789 );
and ( n9233 , n8721 , n8789 );
or ( n9234 , n9231 , n9232 , n9233 );
xor ( n9235 , n9230 , n9234 );
and ( n9236 , n8717 , n8790 );
and ( n9237 , n8790 , n8795 );
and ( n9238 , n8717 , n8795 );
or ( n9239 , n9236 , n9237 , n9238 );
xor ( n9240 , n9235 , n9239 );
and ( n9241 , n8796 , n8797 );
xor ( n9242 , n9240 , n9241 );
buf ( n9243 , n9242 );
not ( n9244 , n454 );
and ( n9245 , n9244 , n9157 );
and ( n9246 , n9243 , n454 );
or ( n9247 , n9245 , n9246 );
buf ( n9248 , n9247 );
buf ( n9249 , n9248 );
and ( n9250 , n9249 , n4505 );
xor ( n9251 , n8997 , n9250 );
and ( n9252 , n7907 , n5089 );
and ( n9253 , n8340 , n4866 );
xor ( n9254 , n9252 , n9253 );
and ( n9255 , n8805 , n4557 );
xor ( n9256 , n9254 , n9255 );
xor ( n9257 , n9251 , n9256 );
and ( n9258 , n8548 , n8549 );
and ( n9259 , n8549 , n8807 );
and ( n9260 , n8548 , n8807 );
or ( n9261 , n9258 , n9259 , n9260 );
xor ( n9262 , n9257 , n9261 );
and ( n9263 , n8808 , n8812 );
and ( n9264 , n8812 , n8817 );
and ( n9265 , n8808 , n8817 );
or ( n9266 , n9263 , n9264 , n9265 );
xor ( n9267 , n9262 , n9266 );
or ( n9268 , n8818 , n8819 );
xnor ( n9269 , n9267 , n9268 );
and ( n9270 , n8820 , n8821 );
xor ( n9271 , n9269 , n9270 );
buf ( n9272 , n9271 );
not ( n9273 , n4509 );
and ( n9274 , n9273 , n8993 );
and ( n9275 , n9272 , n4509 );
or ( n9276 , n9274 , n9275 );
and ( n9277 , n8979 , n8983 );
and ( n9278 , n8983 , n8988 );
and ( n9279 , n8979 , n8988 );
or ( n9280 , n9277 , n9278 , n9279 );
and ( n9281 , n8968 , n4524 );
and ( n9282 , n8951 , n8955 );
and ( n9283 , n8955 , n8960 );
and ( n9284 , n8951 , n8960 );
or ( n9285 , n9282 , n9283 , n9284 );
and ( n9286 , n8900 , n4530 );
buf ( n9287 , n489 );
buf ( n9288 , n505 );
xor ( n9289 , n9287 , n9288 );
and ( n9290 , n8890 , n8891 );
and ( n9291 , n8891 , n8896 );
and ( n9292 , n8890 , n8896 );
or ( n9293 , n9290 , n9291 , n9292 );
xor ( n9294 , n9289 , n9293 );
buf ( n9295 , n9294 );
buf ( n9296 , n9295 );
buf ( n9297 , n9296 );
and ( n9298 , n9297 , n4134 );
nor ( n9299 , n9286 , n9298 );
xnor ( n9300 , n9299 , n4527 );
and ( n9301 , n6353 , n6008 );
and ( n9302 , n6748 , n5689 );
nor ( n9303 , n9301 , n9302 );
xnor ( n9304 , n9303 , n6004 );
and ( n9305 , n5672 , n6761 );
and ( n9306 , n5995 , n6379 );
nor ( n9307 , n9305 , n9306 );
xnor ( n9308 , n9307 , n6757 );
xor ( n9309 , n9304 , n9308 );
xor ( n9310 , n9300 , n9309 );
and ( n9311 , n8921 , n8925 );
and ( n9312 , n8925 , n8930 );
and ( n9313 , n8921 , n8930 );
or ( n9314 , n9311 , n9312 , n9313 );
and ( n9315 , n5121 , n7559 );
and ( n9316 , n5387 , n7107 );
nor ( n9317 , n9315 , n9316 );
xnor ( n9318 , n9317 , n7555 );
and ( n9319 , n4683 , n8382 );
and ( n9320 , n4890 , n8042 );
nor ( n9321 , n9319 , n9320 );
xnor ( n9322 , n9321 , n8378 );
xor ( n9323 , n9318 , n9322 );
and ( n9324 , n4539 , n8375 );
xor ( n9325 , n9323 , n9324 );
xor ( n9326 , n9314 , n9325 );
xor ( n9327 , n9310 , n9326 );
and ( n9328 , n8903 , n8907 );
and ( n9329 , n8907 , n8932 );
and ( n9330 , n8903 , n8932 );
or ( n9331 , n9328 , n9329 , n9330 );
xor ( n9332 , n9327 , n9331 );
and ( n9333 , n8943 , n8947 );
and ( n9334 , n8947 , n8949 );
and ( n9335 , n8943 , n8949 );
or ( n9336 , n9333 , n9334 , n9335 );
and ( n9337 , n8001 , n4898 );
and ( n9338 , n8409 , n4689 );
nor ( n9339 , n9337 , n9338 );
xnor ( n9340 , n9339 , n4904 );
xor ( n9341 , n9336 , n9340 );
and ( n9342 , n7092 , n5405 );
and ( n9343 , n7531 , n5132 );
nor ( n9344 , n9342 , n9343 );
xnor ( n9345 , n9344 , n5401 );
xor ( n9346 , n9341 , n9345 );
and ( n9347 , n8912 , n8916 );
and ( n9348 , n8916 , n8931 );
and ( n9349 , n8912 , n8931 );
or ( n9350 , n9347 , n9348 , n9349 );
xor ( n9351 , n9346 , n9350 );
and ( n9352 , n8942 , n8950 );
xor ( n9353 , n9351 , n9352 );
xor ( n9354 , n9332 , n9353 );
xor ( n9355 , n9285 , n9354 );
and ( n9356 , n8933 , n8937 );
and ( n9357 , n8937 , n8961 );
and ( n9358 , n8933 , n8961 );
or ( n9359 , n9356 , n9357 , n9358 );
xor ( n9360 , n9355 , n9359 );
and ( n9361 , n8888 , n8962 );
and ( n9362 , n8963 , n8964 );
or ( n9363 , n9361 , n9362 );
xor ( n9364 , n9360 , n9363 );
buf ( n9365 , n9364 );
buf ( n9366 , n9365 );
buf ( n9367 , n9366 );
and ( n9368 , n9367 , n4145 );
nor ( n9369 , n9281 , n9368 );
xnor ( n9370 , n9369 , n4521 );
and ( n9371 , n6391 , n6068 );
and ( n9372 , n6796 , n5730 );
nor ( n9373 , n9371 , n9372 );
xnor ( n9374 , n9373 , n6064 );
and ( n9375 , n5700 , n6711 );
and ( n9376 , n6037 , n6332 );
nor ( n9377 , n9375 , n9376 );
xnor ( n9378 , n9377 , n6707 );
xor ( n9379 , n9374 , n9378 );
and ( n9380 , n8849 , n8853 );
and ( n9381 , n8853 , n8874 );
and ( n9382 , n8849 , n8874 );
or ( n9383 , n9380 , n9381 , n9382 );
and ( n9384 , n5140 , n7630 );
and ( n9385 , n5419 , n7188 );
nor ( n9386 , n9384 , n9385 );
xnor ( n9387 , n9386 , n7626 );
xor ( n9388 , n9383 , n9387 );
not ( n9389 , n8873 );
buf ( n9390 , n521 );
buf ( n9391 , n537 );
xor ( n9392 , n9390 , n9391 );
and ( n9393 , n8861 , n8862 );
and ( n9394 , n8862 , n8867 );
and ( n9395 , n8861 , n8867 );
or ( n9396 , n9393 , n9394 , n9395 );
xor ( n9397 , n9392 , n9396 );
buf ( n9398 , n9397 );
buf ( n9399 , n9398 );
buf ( n9400 , n9399 );
and ( n9401 , n8871 , n8495 );
not ( n9402 , n9401 );
and ( n9403 , n9400 , n9402 );
and ( n9404 , n9389 , n9403 );
xor ( n9405 , n9400 , n8871 );
not ( n9406 , n8872 );
and ( n9407 , n9405 , n9406 );
and ( n9408 , n4139 , n9407 );
and ( n9409 , n4548 , n8872 );
nor ( n9410 , n9408 , n9409 );
xnor ( n9411 , n9410 , n9403 );
xor ( n9412 , n9404 , n9411 );
and ( n9413 , n8855 , n8859 );
and ( n9414 , n8859 , n8873 );
and ( n9415 , n8855 , n8873 );
or ( n9416 , n9413 , n9414 , n9415 );
xor ( n9417 , n9412 , n9416 );
and ( n9418 , n4696 , n8502 );
and ( n9419 , n4916 , n7970 );
nor ( n9420 , n9418 , n9419 );
xnor ( n9421 , n9420 , n8498 );
xor ( n9422 , n9417 , n9421 );
xor ( n9423 , n9388 , n9422 );
xor ( n9424 , n9379 , n9423 );
xor ( n9425 , n9370 , n9424 );
and ( n9426 , n8831 , n8835 );
and ( n9427 , n8835 , n8876 );
and ( n9428 , n8831 , n8876 );
or ( n9429 , n9426 , n9427 , n9428 );
xor ( n9430 , n9425 , n9429 );
and ( n9431 , n8883 , n8971 );
and ( n9432 , n8971 , n8976 );
and ( n9433 , n8883 , n8976 );
or ( n9434 , n9431 , n9432 , n9433 );
and ( n9435 , n8840 , n8844 );
and ( n9436 , n8844 , n8875 );
and ( n9437 , n8840 , n8875 );
or ( n9438 , n9435 , n9436 , n9437 );
and ( n9439 , n8057 , n4938 );
and ( n9440 , n8462 , n4711 );
nor ( n9441 , n9439 , n9440 );
xnor ( n9442 , n9441 , n4934 );
xor ( n9443 , n9438 , n9442 );
and ( n9444 , n7146 , n5441 );
and ( n9445 , n7587 , n5161 );
nor ( n9446 , n9444 , n9445 );
xnor ( n9447 , n9446 , n5437 );
xor ( n9448 , n9443 , n9447 );
xor ( n9449 , n9434 , n9448 );
xor ( n9450 , n9430 , n9449 );
and ( n9451 , n8877 , n8878 );
and ( n9452 , n8878 , n8977 );
and ( n9453 , n8877 , n8977 );
or ( n9454 , n9451 , n9452 , n9453 );
xor ( n9455 , n9450 , n9454 );
xor ( n9456 , n9280 , n9455 );
and ( n9457 , n8978 , n8989 );
and ( n9458 , n8990 , n8991 );
or ( n9459 , n9457 , n9458 );
xor ( n9460 , n9456 , n9459 );
buf ( n9461 , n9460 );
and ( n9462 , n9252 , n9253 );
and ( n9463 , n9253 , n9255 );
and ( n9464 , n9252 , n9255 );
or ( n9465 , n9462 , n9463 , n9464 );
and ( n9466 , n9249 , n4557 );
xor ( n9467 , n9465 , n9466 );
and ( n9468 , n8340 , n5089 );
and ( n9469 , n8805 , n4866 );
xor ( n9470 , n9468 , n9469 );
and ( n9471 , n9001 , n9025 );
and ( n9472 , n9025 , n9146 );
and ( n9473 , n9001 , n9146 );
or ( n9474 , n9471 , n9472 , n9473 );
and ( n9475 , n9030 , n9113 );
and ( n9476 , n9113 , n9145 );
and ( n9477 , n9030 , n9145 );
or ( n9478 , n9475 , n9476 , n9477 );
and ( n9479 , n9014 , n9018 );
and ( n9480 , n9018 , n9023 );
and ( n9481 , n9014 , n9023 );
or ( n9482 , n9479 , n9480 , n9481 );
and ( n9483 , n9118 , n9122 );
and ( n9484 , n9122 , n9144 );
and ( n9485 , n9118 , n9144 );
or ( n9486 , n9483 , n9484 , n9485 );
xor ( n9487 , n9482 , n9486 );
and ( n9488 , n9127 , n9131 );
and ( n9489 , n9131 , n9143 );
and ( n9490 , n9127 , n9143 );
or ( n9491 , n9488 , n9489 , n9490 );
and ( n9492 , n6516 , n4788 );
and ( n9493 , n6907 , n4611 );
nor ( n9494 , n9492 , n9493 );
xnor ( n9495 , n9494 , n4784 );
xor ( n9496 , n9491 , n9495 );
and ( n9497 , n5818 , n5270 );
and ( n9498 , n6168 , n5021 );
nor ( n9499 , n9497 , n9498 );
xnor ( n9500 , n9499 , n5266 );
xor ( n9501 , n9496 , n9500 );
xor ( n9502 , n9487 , n9501 );
xor ( n9503 , n9478 , n9502 );
and ( n9504 , n9005 , n9009 );
and ( n9505 , n9009 , n9024 );
and ( n9506 , n9005 , n9024 );
or ( n9507 , n9504 , n9505 , n9506 );
and ( n9508 , n9110 , n4235 );
and ( n9509 , n9069 , n9100 );
and ( n9510 , n9045 , n9056 );
and ( n9511 , n9056 , n9068 );
and ( n9512 , n9045 , n9068 );
or ( n9513 , n9510 , n9511 , n9512 );
and ( n9514 , n9073 , n9077 );
and ( n9515 , n9077 , n9099 );
and ( n9516 , n9073 , n9099 );
or ( n9517 , n9514 , n9515 , n9516 );
xor ( n9518 , n9513 , n9517 );
and ( n9519 , n9082 , n9086 );
and ( n9520 , n9086 , n9098 );
and ( n9521 , n9082 , n9098 );
or ( n9522 , n9519 , n9520 , n9521 );
and ( n9523 , n9088 , n9092 );
and ( n9524 , n9092 , n9097 );
and ( n9525 , n9088 , n9097 );
or ( n9526 , n9523 , n9524 , n9525 );
and ( n9527 , n9049 , n9053 );
and ( n9528 , n9053 , n9055 );
and ( n9529 , n9049 , n9055 );
or ( n9530 , n9527 , n9528 , n9529 );
xor ( n9531 , n9526 , n9530 );
and ( n9532 , n7299 , n4262 );
not ( n9533 , n9532 );
xnor ( n9534 , n9533 , n4252 );
not ( n9535 , n9534 );
xor ( n9536 , n9531 , n9535 );
xor ( n9537 , n9522 , n9536 );
and ( n9538 , n9058 , n9062 );
and ( n9539 , n9062 , n9067 );
and ( n9540 , n9058 , n9067 );
or ( n9541 , n9538 , n9539 , n9540 );
and ( n9542 , n5791 , n5208 );
and ( n9543 , n6120 , n4976 );
nor ( n9544 , n9542 , n9543 );
xnor ( n9545 , n9544 , n5214 );
and ( n9546 , n4243 , n7277 );
and ( n9547 , n4568 , n6864 );
nor ( n9548 , n9546 , n9547 );
xnor ( n9549 , n9548 , n7283 );
xor ( n9550 , n9545 , n9549 );
and ( n9551 , n4160 , n7274 );
xor ( n9552 , n9550 , n9551 );
xor ( n9553 , n9541 , n9552 );
and ( n9554 , n6444 , n4752 );
and ( n9555 , n6853 , n4579 );
nor ( n9556 , n9554 , n9555 );
xnor ( n9557 , n9556 , n4733 );
and ( n9558 , n5195 , n5773 );
and ( n9559 , n5487 , n5519 );
nor ( n9560 , n9558 , n9559 );
xnor ( n9561 , n9560 , n5763 );
xor ( n9562 , n9557 , n9561 );
and ( n9563 , n4724 , n6496 );
and ( n9564 , n4965 , n6115 );
nor ( n9565 , n9563 , n9564 );
xnor ( n9566 , n9565 , n6453 );
xor ( n9567 , n9562 , n9566 );
xor ( n9568 , n9553 , n9567 );
xor ( n9569 , n9537 , n9568 );
xor ( n9570 , n9518 , n9569 );
xor ( n9571 , n9509 , n9570 );
and ( n9572 , n9036 , n9040 );
and ( n9573 , n9040 , n9101 );
and ( n9574 , n9036 , n9101 );
or ( n9575 , n9572 , n9573 , n9574 );
xor ( n9576 , n9571 , n9575 );
and ( n9577 , n9035 , n9102 );
and ( n9578 , n9103 , n9106 );
or ( n9579 , n9577 , n9578 );
xor ( n9580 , n9576 , n9579 );
buf ( n9581 , n9580 );
buf ( n9582 , n9581 );
buf ( n9583 , n9582 );
and ( n9584 , n9583 , n4232 );
nor ( n9585 , n9508 , n9584 );
xnor ( n9586 , n9585 , n4230 );
xor ( n9587 , n9507 , n9586 );
and ( n9588 , n8179 , n4319 );
and ( n9589 , n8640 , n4310 );
nor ( n9590 , n9588 , n9589 );
xnor ( n9591 , n9590 , n4315 );
and ( n9592 , n7324 , n4298 );
and ( n9593 , n7752 , n4287 );
nor ( n9594 , n9592 , n9593 );
xnor ( n9595 , n9594 , n4294 );
xor ( n9596 , n9591 , n9595 );
and ( n9597 , n9136 , n9140 );
and ( n9598 , n9140 , n9142 );
and ( n9599 , n9136 , n9142 );
or ( n9600 , n9597 , n9598 , n9599 );
and ( n9601 , n5247 , n5850 );
and ( n9602 , n5535 , n5566 );
nor ( n9603 , n9601 , n9602 );
xnor ( n9604 , n9603 , n5846 );
xor ( n9605 , n9600 , n9604 );
and ( n9606 , n4770 , n6554 );
and ( n9607 , n4999 , n6205 );
nor ( n9608 , n9606 , n9607 );
xnor ( n9609 , n9608 , n6550 );
and ( n9610 , n4275 , n7356 );
and ( n9611 , n4594 , n6953 );
nor ( n9612 , n9610 , n9611 );
xnor ( n9613 , n9612 , n7352 );
xor ( n9614 , n9609 , n9613 );
and ( n9615 , n4228 , n7349 );
xor ( n9616 , n9614 , n9615 );
xor ( n9617 , n9605 , n9616 );
xor ( n9618 , n9596 , n9617 );
xor ( n9619 , n9587 , n9618 );
xor ( n9620 , n9503 , n9619 );
xor ( n9621 , n9474 , n9620 );
and ( n9622 , n9147 , n9151 );
and ( n9623 , n9152 , n9155 );
or ( n9624 , n9622 , n9623 );
xor ( n9625 , n9621 , n9624 );
buf ( n9626 , n9625 );
and ( n9627 , n9164 , n4418 );
buf ( n9628 , n3503 );
buf ( n9629 , n9628 );
and ( n9630 , n9629 , n4415 );
nor ( n9631 , n9627 , n9630 );
xnor ( n9632 , n9631 , n4413 );
and ( n9633 , n9182 , n9186 );
and ( n9634 , n9186 , n9198 );
and ( n9635 , n9182 , n9198 );
or ( n9636 , n9633 , n9634 , n9635 );
and ( n9637 , n7417 , n4402 );
and ( n9638 , n7857 , n4391 );
nor ( n9639 , n9637 , n9638 );
xnor ( n9640 , n9639 , n4398 );
xor ( n9641 , n9636 , n9640 );
and ( n9642 , n9191 , n9195 );
and ( n9643 , n9195 , n9197 );
and ( n9644 , n9191 , n9197 );
or ( n9645 , n9642 , n9643 , n9644 );
and ( n9646 , n5893 , n5323 );
and ( n9647 , n6235 , n5064 );
nor ( n9648 , n9646 , n9647 );
xnor ( n9649 , n9648 , n5319 );
xor ( n9650 , n9645 , n9649 );
and ( n9651 , n5300 , n5922 );
and ( n9652 , n5588 , n5616 );
nor ( n9653 , n9651 , n9652 );
xnor ( n9654 , n9653 , n5918 );
xor ( n9655 , n9650 , n9654 );
xor ( n9656 , n9641 , n9655 );
xor ( n9657 , n9632 , n9656 );
and ( n9658 , n9204 , n9218 );
and ( n9659 , n9218 , n9223 );
and ( n9660 , n9204 , n9223 );
or ( n9661 , n9658 , n9659 , n9660 );
xor ( n9662 , n9657 , n9661 );
and ( n9663 , n9208 , n9212 );
and ( n9664 , n9212 , n9217 );
and ( n9665 , n9208 , n9217 );
or ( n9666 , n9663 , n9664 , n9665 );
and ( n9667 , n9161 , n9177 );
and ( n9668 , n9177 , n9199 );
and ( n9669 , n9161 , n9199 );
or ( n9670 , n9667 , n9668 , n9669 );
xor ( n9671 , n9666 , n9670 );
and ( n9672 , n8303 , n4433 );
and ( n9673 , n8728 , n4431 );
nor ( n9674 , n9672 , n9673 );
xnor ( n9675 , n9674 , n4441 );
and ( n9676 , n9167 , n9171 );
and ( n9677 , n9171 , n9176 );
and ( n9678 , n9167 , n9176 );
or ( n9679 , n9676 , n9677 , n9678 );
xor ( n9680 , n9675 , n9679 );
and ( n9681 , n6604 , n4835 );
and ( n9682 , n6995 , n4648 );
nor ( n9683 , n9681 , n9682 );
xnor ( n9684 , n9683 , n4831 );
and ( n9685 , n4817 , n6627 );
and ( n9686 , n5042 , n6272 );
nor ( n9687 , n9685 , n9686 );
xnor ( n9688 , n9687 , n6623 );
and ( n9689 , n4421 , n7444 );
and ( n9690 , n4631 , n7026 );
nor ( n9691 , n9689 , n9690 );
xnor ( n9692 , n9691 , n7440 );
xor ( n9693 , n9688 , n9692 );
and ( n9694 , n4411 , n7437 );
xor ( n9695 , n9693 , n9694 );
xor ( n9696 , n9684 , n9695 );
xor ( n9697 , n9680 , n9696 );
xor ( n9698 , n9671 , n9697 );
xor ( n9699 , n9662 , n9698 );
and ( n9700 , n9200 , n9224 );
and ( n9701 , n9224 , n9229 );
and ( n9702 , n9200 , n9229 );
or ( n9703 , n9700 , n9701 , n9702 );
xor ( n9704 , n9699 , n9703 );
and ( n9705 , n9230 , n9234 );
and ( n9706 , n9234 , n9239 );
and ( n9707 , n9230 , n9239 );
or ( n9708 , n9705 , n9706 , n9707 );
xor ( n9709 , n9704 , n9708 );
and ( n9710 , n9240 , n9241 );
xor ( n9711 , n9709 , n9710 );
buf ( n9712 , n9711 );
not ( n9713 , n454 );
and ( n9714 , n9713 , n9626 );
and ( n9715 , n9712 , n454 );
or ( n9716 , n9714 , n9715 );
buf ( n9717 , n9716 );
buf ( n9718 , n9717 );
and ( n9719 , n9718 , n4505 );
xor ( n9720 , n9470 , n9719 );
xor ( n9721 , n9467 , n9720 );
and ( n9722 , n8997 , n9250 );
and ( n9723 , n9250 , n9256 );
and ( n9724 , n8997 , n9256 );
or ( n9725 , n9722 , n9723 , n9724 );
xor ( n9726 , n9721 , n9725 );
and ( n9727 , n9257 , n9261 );
and ( n9728 , n9261 , n9266 );
and ( n9729 , n9257 , n9266 );
or ( n9730 , n9727 , n9728 , n9729 );
xor ( n9731 , n9726 , n9730 );
or ( n9732 , n9267 , n9268 );
xnor ( n9733 , n9731 , n9732 );
and ( n9734 , n9269 , n9270 );
xor ( n9735 , n9733 , n9734 );
buf ( n9736 , n9735 );
not ( n9737 , n4509 );
and ( n9738 , n9737 , n9461 );
and ( n9739 , n9736 , n4509 );
or ( n9740 , n9738 , n9739 );
and ( n9741 , n9434 , n9448 );
and ( n9742 , n9374 , n9378 );
and ( n9743 , n9378 , n9423 );
and ( n9744 , n9374 , n9423 );
or ( n9745 , n9742 , n9743 , n9744 );
and ( n9746 , n7587 , n5441 );
and ( n9747 , n8057 , n5161 );
nor ( n9748 , n9746 , n9747 );
xnor ( n9749 , n9748 , n5437 );
xor ( n9750 , n9745 , n9749 );
and ( n9751 , n9383 , n9387 );
and ( n9752 , n9387 , n9422 );
and ( n9753 , n9383 , n9422 );
or ( n9754 , n9751 , n9752 , n9753 );
and ( n9755 , n6796 , n6068 );
and ( n9756 , n7146 , n5730 );
nor ( n9757 , n9755 , n9756 );
xnor ( n9758 , n9757 , n6064 );
xor ( n9759 , n9754 , n9758 );
and ( n9760 , n6037 , n6711 );
and ( n9761 , n6391 , n6332 );
nor ( n9762 , n9760 , n9761 );
xnor ( n9763 , n9762 , n6707 );
and ( n9764 , n5419 , n7630 );
and ( n9765 , n5700 , n7188 );
nor ( n9766 , n9764 , n9765 );
xnor ( n9767 , n9766 , n7626 );
xor ( n9768 , n9763 , n9767 );
and ( n9769 , n9412 , n9416 );
and ( n9770 , n9416 , n9421 );
and ( n9771 , n9412 , n9421 );
or ( n9772 , n9769 , n9770 , n9771 );
and ( n9773 , n4916 , n8502 );
and ( n9774 , n5140 , n7970 );
nor ( n9775 , n9773 , n9774 );
xnor ( n9776 , n9775 , n8498 );
xor ( n9777 , n9772 , n9776 );
and ( n9778 , n9404 , n9411 );
and ( n9779 , n4548 , n9407 );
and ( n9780 , n4696 , n8872 );
nor ( n9781 , n9779 , n9780 );
xnor ( n9782 , n9781 , n9403 );
xor ( n9783 , n9778 , n9782 );
and ( n9784 , n9390 , n9391 );
and ( n9785 , n9391 , n9396 );
and ( n9786 , n9390 , n9396 );
or ( n9787 , n9784 , n9785 , n9786 );
buf ( n9788 , n9787 );
buf ( n9789 , n9788 );
buf ( n9790 , n9789 );
xor ( n9791 , n9790 , n9400 );
and ( n9792 , n4139 , n9791 );
xor ( n9793 , n9783 , n9792 );
xor ( n9794 , n9777 , n9793 );
xor ( n9795 , n9768 , n9794 );
xor ( n9796 , n9759 , n9795 );
xor ( n9797 , n9750 , n9796 );
and ( n9798 , n9370 , n9424 );
and ( n9799 , n9424 , n9429 );
and ( n9800 , n9370 , n9429 );
or ( n9801 , n9798 , n9799 , n9800 );
xor ( n9802 , n9797 , n9801 );
and ( n9803 , n9367 , n4524 );
and ( n9804 , n9327 , n9331 );
and ( n9805 , n9331 , n9353 );
and ( n9806 , n9327 , n9353 );
or ( n9807 , n9804 , n9805 , n9806 );
and ( n9808 , n9318 , n9322 );
and ( n9809 , n9322 , n9324 );
and ( n9810 , n9318 , n9324 );
or ( n9811 , n9808 , n9809 , n9810 );
and ( n9812 , n8409 , n4898 );
and ( n9813 , n8900 , n4689 );
nor ( n9814 , n9812 , n9813 );
xnor ( n9815 , n9814 , n4904 );
xor ( n9816 , n9811 , n9815 );
and ( n9817 , n7531 , n5405 );
and ( n9818 , n8001 , n5132 );
nor ( n9819 , n9817 , n9818 );
xnor ( n9820 , n9819 , n5401 );
xor ( n9821 , n9816 , n9820 );
and ( n9822 , n5995 , n6761 );
and ( n9823 , n6353 , n6379 );
nor ( n9824 , n9822 , n9823 );
xnor ( n9825 , n9824 , n6757 );
and ( n9826 , n4890 , n8382 );
and ( n9827 , n5121 , n8042 );
nor ( n9828 , n9826 , n9827 );
xnor ( n9829 , n9828 , n8378 );
and ( n9830 , n4683 , n8375 );
xor ( n9831 , n9829 , n9830 );
xor ( n9832 , n9825 , n9831 );
xor ( n9833 , n9821 , n9832 );
and ( n9834 , n9314 , n9325 );
xor ( n9835 , n9833 , n9834 );
and ( n9836 , n9346 , n9350 );
and ( n9837 , n9350 , n9352 );
and ( n9838 , n9346 , n9352 );
or ( n9839 , n9836 , n9837 , n9838 );
xor ( n9840 , n9835 , n9839 );
and ( n9841 , n9297 , n4530 );
and ( n9842 , n9287 , n9288 );
and ( n9843 , n9288 , n9293 );
and ( n9844 , n9287 , n9293 );
or ( n9845 , n9842 , n9843 , n9844 );
buf ( n9846 , n9845 );
buf ( n9847 , n9846 );
buf ( n9848 , n9847 );
and ( n9849 , n9848 , n4134 );
nor ( n9850 , n9841 , n9849 );
xnor ( n9851 , n9850 , n4527 );
and ( n9852 , n6748 , n6008 );
and ( n9853 , n7092 , n5689 );
nor ( n9854 , n9852 , n9853 );
xnor ( n9855 , n9854 , n6004 );
and ( n9856 , n5387 , n7559 );
and ( n9857 , n5672 , n7107 );
nor ( n9858 , n9856 , n9857 );
xnor ( n9859 , n9858 , n7555 );
xor ( n9860 , n9855 , n9859 );
xor ( n9861 , n9851 , n9860 );
and ( n9862 , n9304 , n9308 );
xor ( n9863 , n9861 , n9862 );
and ( n9864 , n9336 , n9340 );
and ( n9865 , n9340 , n9345 );
and ( n9866 , n9336 , n9345 );
or ( n9867 , n9864 , n9865 , n9866 );
xor ( n9868 , n9863 , n9867 );
and ( n9869 , n9300 , n9309 );
and ( n9870 , n9309 , n9326 );
and ( n9871 , n9300 , n9326 );
or ( n9872 , n9869 , n9870 , n9871 );
xor ( n9873 , n9868 , n9872 );
xor ( n9874 , n9840 , n9873 );
xor ( n9875 , n9807 , n9874 );
and ( n9876 , n9285 , n9354 );
and ( n9877 , n9354 , n9359 );
and ( n9878 , n9285 , n9359 );
or ( n9879 , n9876 , n9877 , n9878 );
xor ( n9880 , n9875 , n9879 );
and ( n9881 , n9360 , n9363 );
xor ( n9882 , n9880 , n9881 );
buf ( n9883 , n9882 );
buf ( n9884 , n9883 );
buf ( n9885 , n9884 );
and ( n9886 , n9885 , n4145 );
nor ( n9887 , n9803 , n9886 );
xnor ( n9888 , n9887 , n4521 );
and ( n9889 , n8462 , n4938 );
and ( n9890 , n8968 , n4711 );
nor ( n9891 , n9889 , n9890 );
xnor ( n9892 , n9891 , n4934 );
xor ( n9893 , n9888 , n9892 );
and ( n9894 , n9438 , n9442 );
and ( n9895 , n9442 , n9447 );
and ( n9896 , n9438 , n9447 );
or ( n9897 , n9894 , n9895 , n9896 );
xor ( n9898 , n9893 , n9897 );
xor ( n9899 , n9802 , n9898 );
xor ( n9900 , n9741 , n9899 );
and ( n9901 , n9430 , n9449 );
and ( n9902 , n9449 , n9454 );
and ( n9903 , n9430 , n9454 );
or ( n9904 , n9901 , n9902 , n9903 );
xor ( n9905 , n9900 , n9904 );
and ( n9906 , n9280 , n9455 );
and ( n9907 , n9456 , n9459 );
or ( n9908 , n9906 , n9907 );
xor ( n9909 , n9905 , n9908 );
buf ( n9910 , n9909 );
and ( n9911 , n9468 , n9469 );
and ( n9912 , n9469 , n9719 );
and ( n9913 , n9468 , n9719 );
or ( n9914 , n9911 , n9912 , n9913 );
and ( n9915 , n9507 , n9586 );
and ( n9916 , n9586 , n9618 );
and ( n9917 , n9507 , n9618 );
or ( n9918 , n9915 , n9916 , n9917 );
and ( n9919 , n9583 , n4235 );
and ( n9920 , n9522 , n9536 );
and ( n9921 , n9536 , n9568 );
and ( n9922 , n9522 , n9568 );
or ( n9923 , n9920 , n9921 , n9922 );
and ( n9924 , n9545 , n9549 );
and ( n9925 , n9549 , n9551 );
and ( n9926 , n9545 , n9551 );
or ( n9927 , n9924 , n9925 , n9926 );
and ( n9928 , n6120 , n5208 );
and ( n9929 , n6444 , n4976 );
nor ( n9930 , n9928 , n9929 );
xnor ( n9931 , n9930 , n5214 );
and ( n9932 , n4965 , n6496 );
and ( n9933 , n5195 , n6115 );
nor ( n9934 , n9932 , n9933 );
xnor ( n9935 , n9934 , n6453 );
xor ( n9936 , n9931 , n9935 );
and ( n9937 , n4568 , n7277 );
and ( n9938 , n4724 , n6864 );
nor ( n9939 , n9937 , n9938 );
xnor ( n9940 , n9939 , n7283 );
xor ( n9941 , n9936 , n9940 );
xor ( n9942 , n9927 , n9941 );
not ( n9943 , n4252 );
and ( n9944 , n6853 , n4752 );
and ( n9945 , n7299 , n4579 );
nor ( n9946 , n9944 , n9945 );
xnor ( n9947 , n9946 , n4733 );
xor ( n9948 , n9943 , n9947 );
and ( n9949 , n5487 , n5773 );
and ( n9950 , n5791 , n5519 );
nor ( n9951 , n9949 , n9950 );
xnor ( n9952 , n9951 , n5763 );
xor ( n9953 , n9948 , n9952 );
xor ( n9954 , n9942 , n9953 );
xor ( n9955 , n9923 , n9954 );
and ( n9956 , n9526 , n9530 );
and ( n9957 , n9530 , n9535 );
and ( n9958 , n9526 , n9535 );
or ( n9959 , n9956 , n9957 , n9958 );
and ( n9960 , n9541 , n9552 );
and ( n9961 , n9552 , n9567 );
and ( n9962 , n9541 , n9567 );
or ( n9963 , n9960 , n9961 , n9962 );
xor ( n9964 , n9959 , n9963 );
and ( n9965 , n9557 , n9561 );
and ( n9966 , n9561 , n9566 );
and ( n9967 , n9557 , n9566 );
or ( n9968 , n9965 , n9966 , n9967 );
buf ( n9969 , n9534 );
xor ( n9970 , n9968 , n9969 );
and ( n9971 , n4243 , n7274 );
xor ( n9972 , n9970 , n9971 );
xor ( n9973 , n9964 , n9972 );
xor ( n9974 , n9955 , n9973 );
and ( n9975 , n9513 , n9517 );
and ( n9976 , n9517 , n9569 );
and ( n9977 , n9513 , n9569 );
or ( n9978 , n9975 , n9976 , n9977 );
xor ( n9979 , n9974 , n9978 );
and ( n9980 , n9509 , n9570 );
and ( n9981 , n9570 , n9575 );
and ( n9982 , n9509 , n9575 );
or ( n9983 , n9980 , n9981 , n9982 );
xor ( n9984 , n9979 , n9983 );
and ( n9985 , n9576 , n9579 );
xor ( n9986 , n9984 , n9985 );
buf ( n9987 , n9986 );
buf ( n9988 , n9987 );
buf ( n9989 , n9988 );
and ( n9990 , n9989 , n4232 );
nor ( n9991 , n9919 , n9990 );
xnor ( n9992 , n9991 , n4230 );
and ( n9993 , n8640 , n4319 );
and ( n9994 , n9110 , n4310 );
nor ( n9995 , n9993 , n9994 );
xnor ( n9996 , n9995 , n4315 );
xor ( n9997 , n9992 , n9996 );
and ( n9998 , n9600 , n9604 );
and ( n9999 , n9604 , n9616 );
and ( n10000 , n9600 , n9616 );
or ( n10001 , n9998 , n9999 , n10000 );
and ( n10002 , n6907 , n4788 );
and ( n10003 , n7324 , n4611 );
nor ( n10004 , n10002 , n10003 );
xnor ( n10005 , n10004 , n4784 );
xor ( n10006 , n10001 , n10005 );
and ( n10007 , n6168 , n5270 );
and ( n10008 , n6516 , n5021 );
nor ( n10009 , n10007 , n10008 );
xnor ( n10010 , n10009 , n5266 );
xor ( n10011 , n10006 , n10010 );
xor ( n10012 , n9997 , n10011 );
xor ( n10013 , n9918 , n10012 );
and ( n10014 , n9482 , n9486 );
and ( n10015 , n9486 , n9501 );
and ( n10016 , n9482 , n9501 );
or ( n10017 , n10014 , n10015 , n10016 );
and ( n10018 , n9591 , n9595 );
and ( n10019 , n9595 , n9617 );
and ( n10020 , n9591 , n9617 );
or ( n10021 , n10018 , n10019 , n10020 );
xor ( n10022 , n10017 , n10021 );
and ( n10023 , n9491 , n9495 );
and ( n10024 , n9495 , n9500 );
and ( n10025 , n9491 , n9500 );
or ( n10026 , n10023 , n10024 , n10025 );
and ( n10027 , n7752 , n4298 );
and ( n10028 , n8179 , n4287 );
nor ( n10029 , n10027 , n10028 );
xnor ( n10030 , n10029 , n4294 );
xor ( n10031 , n10026 , n10030 );
and ( n10032 , n9609 , n9613 );
and ( n10033 , n9613 , n9615 );
and ( n10034 , n9609 , n9615 );
or ( n10035 , n10032 , n10033 , n10034 );
and ( n10036 , n5535 , n5850 );
and ( n10037 , n5818 , n5566 );
nor ( n10038 , n10036 , n10037 );
xnor ( n10039 , n10038 , n5846 );
xor ( n10040 , n10035 , n10039 );
and ( n10041 , n4999 , n6554 );
and ( n10042 , n5247 , n6205 );
nor ( n10043 , n10041 , n10042 );
xnor ( n10044 , n10043 , n6550 );
and ( n10045 , n4594 , n7356 );
and ( n10046 , n4770 , n6953 );
nor ( n10047 , n10045 , n10046 );
xnor ( n10048 , n10047 , n7352 );
xor ( n10049 , n10044 , n10048 );
and ( n10050 , n4275 , n7349 );
xor ( n10051 , n10049 , n10050 );
xor ( n10052 , n10040 , n10051 );
xor ( n10053 , n10031 , n10052 );
xor ( n10054 , n10022 , n10053 );
xor ( n10055 , n10013 , n10054 );
and ( n10056 , n9478 , n9502 );
and ( n10057 , n9502 , n9619 );
and ( n10058 , n9478 , n9619 );
or ( n10059 , n10056 , n10057 , n10058 );
xor ( n10060 , n10055 , n10059 );
and ( n10061 , n9474 , n9620 );
and ( n10062 , n9621 , n9624 );
or ( n10063 , n10061 , n10062 );
xor ( n10064 , n10060 , n10063 );
buf ( n10065 , n10064 );
and ( n10066 , n9675 , n9679 );
and ( n10067 , n9679 , n9696 );
and ( n10068 , n9675 , n9696 );
or ( n10069 , n10066 , n10067 , n10068 );
and ( n10070 , n9629 , n4418 );
buf ( n10071 , n3616 );
buf ( n10072 , n10071 );
and ( n10073 , n10072 , n4415 );
nor ( n10074 , n10070 , n10073 );
xnor ( n10075 , n10074 , n4413 );
and ( n10076 , n9688 , n9692 );
and ( n10077 , n9692 , n9694 );
and ( n10078 , n9688 , n9694 );
or ( n10079 , n10076 , n10077 , n10078 );
and ( n10080 , n6235 , n5323 );
and ( n10081 , n6604 , n5064 );
nor ( n10082 , n10080 , n10081 );
xnor ( n10083 , n10082 , n5319 );
xor ( n10084 , n10079 , n10083 );
and ( n10085 , n5588 , n5922 );
and ( n10086 , n5893 , n5616 );
nor ( n10087 , n10085 , n10086 );
xnor ( n10088 , n10087 , n5918 );
xor ( n10089 , n10084 , n10088 );
xor ( n10090 , n10075 , n10089 );
and ( n10091 , n5042 , n6627 );
and ( n10092 , n5300 , n6272 );
nor ( n10093 , n10091 , n10092 );
xnor ( n10094 , n10093 , n6623 );
and ( n10095 , n4631 , n7444 );
and ( n10096 , n4817 , n7026 );
nor ( n10097 , n10095 , n10096 );
xnor ( n10098 , n10097 , n7440 );
and ( n10099 , n4421 , n7437 );
xor ( n10100 , n10098 , n10099 );
xor ( n10101 , n10094 , n10100 );
and ( n10102 , n7857 , n4402 );
and ( n10103 , n8303 , n4391 );
nor ( n10104 , n10102 , n10103 );
xnor ( n10105 , n10104 , n4398 );
xor ( n10106 , n10101 , n10105 );
and ( n10107 , n6995 , n4835 );
and ( n10108 , n7417 , n4648 );
nor ( n10109 , n10107 , n10108 );
xnor ( n10110 , n10109 , n4831 );
xor ( n10111 , n10106 , n10110 );
xor ( n10112 , n10090 , n10111 );
xor ( n10113 , n10069 , n10112 );
and ( n10114 , n9632 , n9656 );
xor ( n10115 , n10113 , n10114 );
and ( n10116 , n9666 , n9670 );
and ( n10117 , n9670 , n9697 );
and ( n10118 , n9666 , n9697 );
or ( n10119 , n10116 , n10117 , n10118 );
and ( n10120 , n9684 , n9695 );
and ( n10121 , n9645 , n9649 );
and ( n10122 , n9649 , n9654 );
and ( n10123 , n9645 , n9654 );
or ( n10124 , n10121 , n10122 , n10123 );
and ( n10125 , n8728 , n4433 );
and ( n10126 , n9164 , n4431 );
nor ( n10127 , n10125 , n10126 );
xnor ( n10128 , n10127 , n4441 );
xor ( n10129 , n10124 , n10128 );
xor ( n10130 , n10120 , n10129 );
and ( n10131 , n9636 , n9640 );
and ( n10132 , n9640 , n9655 );
and ( n10133 , n9636 , n9655 );
or ( n10134 , n10131 , n10132 , n10133 );
xor ( n10135 , n10130 , n10134 );
xor ( n10136 , n10119 , n10135 );
and ( n10137 , n9657 , n9661 );
and ( n10138 , n9661 , n9698 );
and ( n10139 , n9657 , n9698 );
or ( n10140 , n10137 , n10138 , n10139 );
xor ( n10141 , n10136 , n10140 );
xor ( n10142 , n10115 , n10141 );
and ( n10143 , n9699 , n9703 );
and ( n10144 , n9703 , n9708 );
and ( n10145 , n9699 , n9708 );
or ( n10146 , n10143 , n10144 , n10145 );
xor ( n10147 , n10142 , n10146 );
and ( n10148 , n9709 , n9710 );
xor ( n10149 , n10147 , n10148 );
buf ( n10150 , n10149 );
not ( n10151 , n454 );
and ( n10152 , n10151 , n10065 );
and ( n10153 , n10150 , n454 );
or ( n10154 , n10152 , n10153 );
buf ( n10155 , n10154 );
buf ( n10156 , n10155 );
and ( n10157 , n10156 , n4505 );
xor ( n10158 , n9914 , n10157 );
and ( n10159 , n8805 , n5089 );
and ( n10160 , n9249 , n4866 );
xor ( n10161 , n10159 , n10160 );
and ( n10162 , n9718 , n4557 );
xor ( n10163 , n10161 , n10162 );
xor ( n10164 , n10158 , n10163 );
and ( n10165 , n9465 , n9466 );
and ( n10166 , n9466 , n9720 );
and ( n10167 , n9465 , n9720 );
or ( n10168 , n10165 , n10166 , n10167 );
xor ( n10169 , n10164 , n10168 );
and ( n10170 , n9721 , n9725 );
and ( n10171 , n9725 , n9730 );
and ( n10172 , n9721 , n9730 );
or ( n10173 , n10170 , n10171 , n10172 );
xor ( n10174 , n10169 , n10173 );
or ( n10175 , n9731 , n9732 );
xnor ( n10176 , n10174 , n10175 );
and ( n10177 , n9733 , n9734 );
xor ( n10178 , n10176 , n10177 );
buf ( n10179 , n10178 );
not ( n10180 , n4509 );
and ( n10181 , n10180 , n9910 );
and ( n10182 , n10179 , n4509 );
or ( n10183 , n10181 , n10182 );
and ( n10184 , n9797 , n9801 );
and ( n10185 , n9801 , n9898 );
and ( n10186 , n9797 , n9898 );
or ( n10187 , n10184 , n10185 , n10186 );
and ( n10188 , n9754 , n9758 );
and ( n10189 , n9758 , n9795 );
and ( n10190 , n9754 , n9795 );
or ( n10191 , n10188 , n10189 , n10190 );
and ( n10192 , n8968 , n4938 );
and ( n10193 , n9367 , n4711 );
nor ( n10194 , n10192 , n10193 );
xnor ( n10195 , n10194 , n4934 );
xor ( n10196 , n10191 , n10195 );
and ( n10197 , n8057 , n5441 );
and ( n10198 , n8462 , n5161 );
nor ( n10199 , n10197 , n10198 );
xnor ( n10200 , n10199 , n5437 );
xor ( n10201 , n10196 , n10200 );
and ( n10202 , n9888 , n9892 );
and ( n10203 , n9892 , n9897 );
and ( n10204 , n9888 , n9897 );
or ( n10205 , n10202 , n10203 , n10204 );
xor ( n10206 , n10201 , n10205 );
and ( n10207 , n9745 , n9749 );
and ( n10208 , n9749 , n9796 );
and ( n10209 , n9745 , n9796 );
or ( n10210 , n10207 , n10208 , n10209 );
and ( n10211 , n9885 , n4524 );
and ( n10212 , n9835 , n9839 );
and ( n10213 , n9839 , n9873 );
and ( n10214 , n9835 , n9873 );
or ( n10215 , n10212 , n10213 , n10214 );
and ( n10216 , n9829 , n9830 );
and ( n10217 , n5672 , n7559 );
and ( n10218 , n5995 , n7107 );
nor ( n10219 , n10217 , n10218 );
xnor ( n10220 , n10219 , n7555 );
xor ( n10221 , n10216 , n10220 );
and ( n10222 , n5121 , n8382 );
and ( n10223 , n5387 , n8042 );
nor ( n10224 , n10222 , n10223 );
xnor ( n10225 , n10224 , n8378 );
xor ( n10226 , n10221 , n10225 );
and ( n10227 , n9811 , n9815 );
and ( n10228 , n9815 , n9820 );
and ( n10229 , n9811 , n9820 );
or ( n10230 , n10227 , n10228 , n10229 );
xor ( n10231 , n10226 , n10230 );
and ( n10232 , n9825 , n9831 );
xor ( n10233 , n10231 , n10232 );
and ( n10234 , n9863 , n9867 );
and ( n10235 , n9867 , n9872 );
and ( n10236 , n9863 , n9872 );
or ( n10237 , n10234 , n10235 , n10236 );
xor ( n10238 , n10233 , n10237 );
and ( n10239 , n9851 , n9860 );
and ( n10240 , n9860 , n9862 );
and ( n10241 , n9851 , n9862 );
or ( n10242 , n10239 , n10240 , n10241 );
and ( n10243 , n8900 , n4898 );
and ( n10244 , n9297 , n4689 );
nor ( n10245 , n10243 , n10244 );
xnor ( n10246 , n10245 , n4904 );
and ( n10247 , n7092 , n6008 );
and ( n10248 , n7531 , n5689 );
nor ( n10249 , n10247 , n10248 );
xnor ( n10250 , n10249 , n6004 );
xor ( n10251 , n10246 , n10250 );
and ( n10252 , n6353 , n6761 );
and ( n10253 , n6748 , n6379 );
nor ( n10254 , n10252 , n10253 );
xnor ( n10255 , n10254 , n6757 );
xor ( n10256 , n10251 , n10255 );
and ( n10257 , n9855 , n9859 );
xor ( n10258 , n10256 , n10257 );
and ( n10259 , n9848 , n4530 );
not ( n10260 , n10259 );
xnor ( n10261 , n10260 , n4527 );
and ( n10262 , n8001 , n5405 );
and ( n10263 , n8409 , n5132 );
nor ( n10264 , n10262 , n10263 );
xnor ( n10265 , n10264 , n5401 );
xor ( n10266 , n10261 , n10265 );
and ( n10267 , n4890 , n8375 );
xor ( n10268 , n10266 , n10267 );
xor ( n10269 , n10258 , n10268 );
xor ( n10270 , n10242 , n10269 );
and ( n10271 , n9821 , n9832 );
and ( n10272 , n9832 , n9834 );
and ( n10273 , n9821 , n9834 );
or ( n10274 , n10271 , n10272 , n10273 );
xor ( n10275 , n10270 , n10274 );
xor ( n10276 , n10238 , n10275 );
xor ( n10277 , n10215 , n10276 );
and ( n10278 , n9807 , n9874 );
and ( n10279 , n9874 , n9879 );
and ( n10280 , n9807 , n9879 );
or ( n10281 , n10278 , n10279 , n10280 );
xor ( n10282 , n10277 , n10281 );
and ( n10283 , n9880 , n9881 );
xor ( n10284 , n10282 , n10283 );
buf ( n10285 , n10284 );
buf ( n10286 , n10285 );
buf ( n10287 , n10286 );
and ( n10288 , n10287 , n4145 );
nor ( n10289 , n10211 , n10288 );
xnor ( n10290 , n10289 , n4521 );
xor ( n10291 , n10210 , n10290 );
and ( n10292 , n9763 , n9767 );
and ( n10293 , n9767 , n9794 );
and ( n10294 , n9763 , n9794 );
or ( n10295 , n10292 , n10293 , n10294 );
and ( n10296 , n7146 , n6068 );
and ( n10297 , n7587 , n5730 );
nor ( n10298 , n10296 , n10297 );
xnor ( n10299 , n10298 , n6064 );
xor ( n10300 , n10295 , n10299 );
and ( n10301 , n6391 , n6711 );
and ( n10302 , n6796 , n6332 );
nor ( n10303 , n10301 , n10302 );
xnor ( n10304 , n10303 , n6707 );
and ( n10305 , n5700 , n7630 );
and ( n10306 , n6037 , n7188 );
nor ( n10307 , n10305 , n10306 );
xnor ( n10308 , n10307 , n7626 );
xor ( n10309 , n10304 , n10308 );
and ( n10310 , n9772 , n9776 );
and ( n10311 , n9776 , n9793 );
and ( n10312 , n9772 , n9793 );
or ( n10313 , n10310 , n10311 , n10312 );
and ( n10314 , n5140 , n8502 );
and ( n10315 , n5419 , n7970 );
nor ( n10316 , n10314 , n10315 );
xnor ( n10317 , n10316 , n8498 );
xor ( n10318 , n10313 , n10317 );
and ( n10319 , n9778 , n9782 );
and ( n10320 , n9782 , n9792 );
and ( n10321 , n9778 , n9792 );
or ( n10322 , n10319 , n10320 , n10321 );
and ( n10323 , n4696 , n9407 );
and ( n10324 , n4916 , n8872 );
nor ( n10325 , n10323 , n10324 );
xnor ( n10326 , n10325 , n9403 );
xor ( n10327 , n10322 , n10326 );
not ( n10328 , n9791 );
and ( n10329 , n9790 , n10328 );
and ( n10330 , n4139 , n10329 );
and ( n10331 , n4548 , n9791 );
nor ( n10332 , n10330 , n10331 );
not ( n10333 , n10332 );
xor ( n10334 , n10327 , n10333 );
xor ( n10335 , n10318 , n10334 );
xor ( n10336 , n10309 , n10335 );
xor ( n10337 , n10300 , n10336 );
xor ( n10338 , n10291 , n10337 );
xor ( n10339 , n10206 , n10338 );
xor ( n10340 , n10187 , n10339 );
and ( n10341 , n9741 , n9899 );
and ( n10342 , n9899 , n9904 );
and ( n10343 , n9741 , n9904 );
or ( n10344 , n10341 , n10342 , n10343 );
xor ( n10345 , n10340 , n10344 );
and ( n10346 , n9905 , n9908 );
xor ( n10347 , n10345 , n10346 );
buf ( n10348 , n10347 );
and ( n10349 , n10159 , n10160 );
and ( n10350 , n10160 , n10162 );
and ( n10351 , n10159 , n10162 );
or ( n10352 , n10349 , n10350 , n10351 );
and ( n10353 , n10156 , n4557 );
xor ( n10354 , n10352 , n10353 );
and ( n10355 , n9249 , n5089 );
and ( n10356 , n9718 , n4866 );
xor ( n10357 , n10355 , n10356 );
and ( n10358 , n10017 , n10021 );
and ( n10359 , n10021 , n10053 );
and ( n10360 , n10017 , n10053 );
or ( n10361 , n10358 , n10359 , n10360 );
and ( n10362 , n10001 , n10005 );
and ( n10363 , n10005 , n10010 );
and ( n10364 , n10001 , n10010 );
or ( n10365 , n10362 , n10363 , n10364 );
and ( n10366 , n10026 , n10030 );
and ( n10367 , n10030 , n10052 );
and ( n10368 , n10026 , n10052 );
or ( n10369 , n10366 , n10367 , n10368 );
xor ( n10370 , n10365 , n10369 );
and ( n10371 , n9989 , n4235 );
and ( n10372 , n9959 , n9963 );
and ( n10373 , n9963 , n9972 );
and ( n10374 , n9959 , n9972 );
or ( n10375 , n10372 , n10373 , n10374 );
and ( n10376 , n9931 , n9935 );
and ( n10377 , n9935 , n9940 );
and ( n10378 , n9931 , n9940 );
or ( n10379 , n10376 , n10377 , n10378 );
and ( n10380 , n9943 , n9947 );
and ( n10381 , n9947 , n9952 );
and ( n10382 , n9943 , n9952 );
or ( n10383 , n10380 , n10381 , n10382 );
xor ( n10384 , n10379 , n10383 );
and ( n10385 , n7299 , n4752 );
not ( n10386 , n10385 );
xnor ( n10387 , n10386 , n4733 );
and ( n10388 , n5195 , n6496 );
and ( n10389 , n5487 , n6115 );
nor ( n10390 , n10388 , n10389 );
xnor ( n10391 , n10390 , n6453 );
xor ( n10392 , n10387 , n10391 );
and ( n10393 , n4724 , n7277 );
and ( n10394 , n4965 , n6864 );
nor ( n10395 , n10393 , n10394 );
xnor ( n10396 , n10395 , n7283 );
xor ( n10397 , n10392 , n10396 );
xor ( n10398 , n10384 , n10397 );
xor ( n10399 , n10375 , n10398 );
and ( n10400 , n9968 , n9969 );
and ( n10401 , n9969 , n9971 );
and ( n10402 , n9968 , n9971 );
or ( n10403 , n10400 , n10401 , n10402 );
and ( n10404 , n9927 , n9941 );
and ( n10405 , n9941 , n9953 );
and ( n10406 , n9927 , n9953 );
or ( n10407 , n10404 , n10405 , n10406 );
xor ( n10408 , n10403 , n10407 );
and ( n10409 , n6444 , n5208 );
and ( n10410 , n6853 , n4976 );
nor ( n10411 , n10409 , n10410 );
xnor ( n10412 , n10411 , n5214 );
not ( n10413 , n10412 );
and ( n10414 , n5791 , n5773 );
and ( n10415 , n6120 , n5519 );
nor ( n10416 , n10414 , n10415 );
xnor ( n10417 , n10416 , n5763 );
xor ( n10418 , n10413 , n10417 );
and ( n10419 , n4568 , n7274 );
xor ( n10420 , n10418 , n10419 );
xor ( n10421 , n10408 , n10420 );
xor ( n10422 , n10399 , n10421 );
and ( n10423 , n9923 , n9954 );
and ( n10424 , n9954 , n9973 );
and ( n10425 , n9923 , n9973 );
or ( n10426 , n10423 , n10424 , n10425 );
xor ( n10427 , n10422 , n10426 );
and ( n10428 , n9974 , n9978 );
and ( n10429 , n9978 , n9983 );
and ( n10430 , n9974 , n9983 );
or ( n10431 , n10428 , n10429 , n10430 );
xor ( n10432 , n10427 , n10431 );
and ( n10433 , n9984 , n9985 );
xor ( n10434 , n10432 , n10433 );
buf ( n10435 , n10434 );
buf ( n10436 , n10435 );
buf ( n10437 , n10436 );
and ( n10438 , n10437 , n4232 );
nor ( n10439 , n10371 , n10438 );
xnor ( n10440 , n10439 , n4230 );
xor ( n10441 , n10370 , n10440 );
xor ( n10442 , n10361 , n10441 );
and ( n10443 , n9992 , n9996 );
and ( n10444 , n9996 , n10011 );
and ( n10445 , n9992 , n10011 );
or ( n10446 , n10443 , n10444 , n10445 );
and ( n10447 , n8179 , n4298 );
and ( n10448 , n8640 , n4287 );
nor ( n10449 , n10447 , n10448 );
xnor ( n10450 , n10449 , n4294 );
and ( n10451 , n7324 , n4788 );
and ( n10452 , n7752 , n4611 );
nor ( n10453 , n10451 , n10452 );
xnor ( n10454 , n10453 , n4784 );
xor ( n10455 , n10450 , n10454 );
and ( n10456 , n5247 , n6554 );
and ( n10457 , n5535 , n6205 );
nor ( n10458 , n10456 , n10457 );
xnor ( n10459 , n10458 , n6550 );
and ( n10460 , n4770 , n7356 );
and ( n10461 , n4999 , n6953 );
nor ( n10462 , n10460 , n10461 );
xnor ( n10463 , n10462 , n7352 );
xor ( n10464 , n10459 , n10463 );
and ( n10465 , n4594 , n7349 );
xor ( n10466 , n10464 , n10465 );
xor ( n10467 , n10455 , n10466 );
xor ( n10468 , n10446 , n10467 );
and ( n10469 , n10035 , n10039 );
and ( n10470 , n10039 , n10051 );
and ( n10471 , n10035 , n10051 );
or ( n10472 , n10469 , n10470 , n10471 );
and ( n10473 , n9110 , n4319 );
and ( n10474 , n9583 , n4310 );
nor ( n10475 , n10473 , n10474 );
xnor ( n10476 , n10475 , n4315 );
xor ( n10477 , n10472 , n10476 );
and ( n10478 , n10044 , n10048 );
and ( n10479 , n10048 , n10050 );
and ( n10480 , n10044 , n10050 );
or ( n10481 , n10478 , n10479 , n10480 );
and ( n10482 , n6516 , n5270 );
and ( n10483 , n6907 , n5021 );
nor ( n10484 , n10482 , n10483 );
xnor ( n10485 , n10484 , n5266 );
xor ( n10486 , n10481 , n10485 );
and ( n10487 , n5818 , n5850 );
and ( n10488 , n6168 , n5566 );
nor ( n10489 , n10487 , n10488 );
xnor ( n10490 , n10489 , n5846 );
xor ( n10491 , n10486 , n10490 );
xor ( n10492 , n10477 , n10491 );
xor ( n10493 , n10468 , n10492 );
xor ( n10494 , n10442 , n10493 );
and ( n10495 , n9918 , n10012 );
and ( n10496 , n10012 , n10054 );
and ( n10497 , n9918 , n10054 );
or ( n10498 , n10495 , n10496 , n10497 );
xor ( n10499 , n10494 , n10498 );
and ( n10500 , n10055 , n10059 );
and ( n10501 , n10060 , n10063 );
or ( n10502 , n10500 , n10501 );
xor ( n10503 , n10499 , n10502 );
buf ( n10504 , n10503 );
and ( n10505 , n10124 , n10128 );
and ( n10506 , n10079 , n10083 );
and ( n10507 , n10083 , n10088 );
and ( n10508 , n10079 , n10088 );
or ( n10509 , n10506 , n10507 , n10508 );
and ( n10510 , n9164 , n4433 );
and ( n10511 , n9629 , n4431 );
nor ( n10512 , n10510 , n10511 );
xnor ( n10513 , n10512 , n4441 );
xor ( n10514 , n10509 , n10513 );
and ( n10515 , n10094 , n10100 );
and ( n10516 , n6604 , n5323 );
and ( n10517 , n6995 , n5064 );
nor ( n10518 , n10516 , n10517 );
xnor ( n10519 , n10518 , n5319 );
xor ( n10520 , n10515 , n10519 );
and ( n10521 , n5893 , n5922 );
and ( n10522 , n6235 , n5616 );
nor ( n10523 , n10521 , n10522 );
xnor ( n10524 , n10523 , n5918 );
xor ( n10525 , n10520 , n10524 );
xor ( n10526 , n10514 , n10525 );
xor ( n10527 , n10505 , n10526 );
and ( n10528 , n10101 , n10105 );
and ( n10529 , n10105 , n10110 );
and ( n10530 , n10101 , n10110 );
or ( n10531 , n10528 , n10529 , n10530 );
and ( n10532 , n10072 , n4418 );
buf ( n10533 , n3718 );
buf ( n10534 , n10533 );
and ( n10535 , n10534 , n4415 );
nor ( n10536 , n10532 , n10535 );
xnor ( n10537 , n10536 , n4413 );
xor ( n10538 , n10531 , n10537 );
and ( n10539 , n8303 , n4402 );
and ( n10540 , n8728 , n4391 );
nor ( n10541 , n10539 , n10540 );
xnor ( n10542 , n10541 , n4398 );
and ( n10543 , n7417 , n4835 );
and ( n10544 , n7857 , n4648 );
nor ( n10545 , n10543 , n10544 );
xnor ( n10546 , n10545 , n4831 );
xor ( n10547 , n10542 , n10546 );
and ( n10548 , n4817 , n7444 );
and ( n10549 , n5042 , n7026 );
nor ( n10550 , n10548 , n10549 );
xnor ( n10551 , n10550 , n7440 );
and ( n10552 , n4631 , n7437 );
xor ( n10553 , n10551 , n10552 );
and ( n10554 , n10098 , n10099 );
xor ( n10555 , n10553 , n10554 );
and ( n10556 , n5300 , n6627 );
and ( n10557 , n5588 , n6272 );
nor ( n10558 , n10556 , n10557 );
xnor ( n10559 , n10558 , n6623 );
xor ( n10560 , n10555 , n10559 );
xor ( n10561 , n10547 , n10560 );
xor ( n10562 , n10538 , n10561 );
xor ( n10563 , n10527 , n10562 );
and ( n10564 , n10119 , n10135 );
and ( n10565 , n10135 , n10140 );
and ( n10566 , n10119 , n10140 );
or ( n10567 , n10564 , n10565 , n10566 );
xor ( n10568 , n10563 , n10567 );
and ( n10569 , n10075 , n10089 );
and ( n10570 , n10089 , n10111 );
and ( n10571 , n10075 , n10111 );
or ( n10572 , n10569 , n10570 , n10571 );
and ( n10573 , n10120 , n10129 );
and ( n10574 , n10129 , n10134 );
and ( n10575 , n10120 , n10134 );
or ( n10576 , n10573 , n10574 , n10575 );
xor ( n10577 , n10572 , n10576 );
and ( n10578 , n10069 , n10112 );
and ( n10579 , n10112 , n10114 );
and ( n10580 , n10069 , n10114 );
or ( n10581 , n10578 , n10579 , n10580 );
xor ( n10582 , n10577 , n10581 );
xor ( n10583 , n10568 , n10582 );
and ( n10584 , n10115 , n10141 );
and ( n10585 , n10141 , n10146 );
and ( n10586 , n10115 , n10146 );
or ( n10587 , n10584 , n10585 , n10586 );
xor ( n10588 , n10583 , n10587 );
and ( n10589 , n10147 , n10148 );
xor ( n10590 , n10588 , n10589 );
buf ( n10591 , n10590 );
not ( n10592 , n454 );
and ( n10593 , n10592 , n10504 );
and ( n10594 , n10591 , n454 );
or ( n10595 , n10593 , n10594 );
buf ( n10596 , n10595 );
buf ( n10597 , n10596 );
and ( n10598 , n10597 , n4505 );
xor ( n10599 , n10357 , n10598 );
xor ( n10600 , n10354 , n10599 );
and ( n10601 , n9914 , n10157 );
and ( n10602 , n10157 , n10163 );
and ( n10603 , n9914 , n10163 );
or ( n10604 , n10601 , n10602 , n10603 );
xor ( n10605 , n10600 , n10604 );
and ( n10606 , n10164 , n10168 );
and ( n10607 , n10168 , n10173 );
and ( n10608 , n10164 , n10173 );
or ( n10609 , n10606 , n10607 , n10608 );
xor ( n10610 , n10605 , n10609 );
or ( n10611 , n10174 , n10175 );
xnor ( n10612 , n10610 , n10611 );
and ( n10613 , n10176 , n10177 );
xor ( n10614 , n10612 , n10613 );
buf ( n10615 , n10614 );
not ( n10616 , n4509 );
and ( n10617 , n10616 , n10348 );
and ( n10618 , n10615 , n4509 );
or ( n10619 , n10617 , n10618 );
and ( n10620 , n10210 , n10290 );
and ( n10621 , n10290 , n10337 );
and ( n10622 , n10210 , n10337 );
or ( n10623 , n10620 , n10621 , n10622 );
and ( n10624 , n10191 , n10195 );
and ( n10625 , n10195 , n10200 );
and ( n10626 , n10191 , n10200 );
or ( n10627 , n10624 , n10625 , n10626 );
and ( n10628 , n10287 , n4524 );
and ( n10629 , n10233 , n10237 );
and ( n10630 , n10237 , n10275 );
and ( n10631 , n10233 , n10275 );
or ( n10632 , n10629 , n10630 , n10631 );
not ( n10633 , n4527 );
and ( n10634 , n5121 , n8375 );
xnor ( n10635 , n10633 , n10634 );
and ( n10636 , n10261 , n10265 );
and ( n10637 , n10265 , n10267 );
and ( n10638 , n10261 , n10267 );
or ( n10639 , n10636 , n10637 , n10638 );
xor ( n10640 , n10635 , n10639 );
and ( n10641 , n10246 , n10250 );
and ( n10642 , n10250 , n10255 );
and ( n10643 , n10246 , n10255 );
or ( n10644 , n10641 , n10642 , n10643 );
and ( n10645 , n7531 , n6008 );
and ( n10646 , n8001 , n5689 );
nor ( n10647 , n10645 , n10646 );
xnor ( n10648 , n10647 , n6004 );
and ( n10649 , n5995 , n7559 );
and ( n10650 , n6353 , n7107 );
nor ( n10651 , n10649 , n10650 );
xnor ( n10652 , n10651 , n7555 );
xor ( n10653 , n10648 , n10652 );
and ( n10654 , n5387 , n8382 );
and ( n10655 , n5672 , n8042 );
nor ( n10656 , n10654 , n10655 );
xnor ( n10657 , n10656 , n8378 );
xor ( n10658 , n10653 , n10657 );
xor ( n10659 , n10644 , n10658 );
and ( n10660 , n9297 , n4898 );
and ( n10661 , n9848 , n4689 );
nor ( n10662 , n10660 , n10661 );
xnor ( n10663 , n10662 , n4904 );
and ( n10664 , n8409 , n5405 );
and ( n10665 , n8900 , n5132 );
nor ( n10666 , n10664 , n10665 );
xnor ( n10667 , n10666 , n5401 );
xor ( n10668 , n10663 , n10667 );
and ( n10669 , n6748 , n6761 );
and ( n10670 , n7092 , n6379 );
nor ( n10671 , n10669 , n10670 );
xnor ( n10672 , n10671 , n6757 );
xor ( n10673 , n10668 , n10672 );
xor ( n10674 , n10659 , n10673 );
xor ( n10675 , n10640 , n10674 );
and ( n10676 , n10242 , n10269 );
and ( n10677 , n10269 , n10274 );
and ( n10678 , n10242 , n10274 );
or ( n10679 , n10676 , n10677 , n10678 );
xor ( n10680 , n10675 , n10679 );
and ( n10681 , n10216 , n10220 );
and ( n10682 , n10220 , n10225 );
and ( n10683 , n10216 , n10225 );
or ( n10684 , n10681 , n10682 , n10683 );
and ( n10685 , n10256 , n10257 );
and ( n10686 , n10257 , n10268 );
and ( n10687 , n10256 , n10268 );
or ( n10688 , n10685 , n10686 , n10687 );
xor ( n10689 , n10684 , n10688 );
and ( n10690 , n10226 , n10230 );
and ( n10691 , n10230 , n10232 );
and ( n10692 , n10226 , n10232 );
or ( n10693 , n10690 , n10691 , n10692 );
xor ( n10694 , n10689 , n10693 );
xor ( n10695 , n10680 , n10694 );
xor ( n10696 , n10632 , n10695 );
and ( n10697 , n10215 , n10276 );
and ( n10698 , n10276 , n10281 );
and ( n10699 , n10215 , n10281 );
or ( n10700 , n10697 , n10698 , n10699 );
xor ( n10701 , n10696 , n10700 );
and ( n10702 , n10282 , n10283 );
xor ( n10703 , n10701 , n10702 );
buf ( n10704 , n10703 );
buf ( n10705 , n10704 );
buf ( n10706 , n10705 );
and ( n10707 , n10706 , n4145 );
nor ( n10708 , n10628 , n10707 );
xnor ( n10709 , n10708 , n4521 );
xor ( n10710 , n10627 , n10709 );
and ( n10711 , n10304 , n10308 );
and ( n10712 , n10308 , n10335 );
and ( n10713 , n10304 , n10335 );
or ( n10714 , n10711 , n10712 , n10713 );
and ( n10715 , n8462 , n5441 );
and ( n10716 , n8968 , n5161 );
nor ( n10717 , n10715 , n10716 );
xnor ( n10718 , n10717 , n5437 );
xor ( n10719 , n10714 , n10718 );
and ( n10720 , n7587 , n6068 );
and ( n10721 , n8057 , n5730 );
nor ( n10722 , n10720 , n10721 );
xnor ( n10723 , n10722 , n6064 );
xor ( n10724 , n10719 , n10723 );
xor ( n10725 , n10710 , n10724 );
xor ( n10726 , n10623 , n10725 );
and ( n10727 , n10295 , n10299 );
and ( n10728 , n10299 , n10336 );
and ( n10729 , n10295 , n10336 );
or ( n10730 , n10727 , n10728 , n10729 );
and ( n10731 , n9367 , n4938 );
and ( n10732 , n9885 , n4711 );
nor ( n10733 , n10731 , n10732 );
xnor ( n10734 , n10733 , n4934 );
xor ( n10735 , n10730 , n10734 );
and ( n10736 , n10313 , n10317 );
and ( n10737 , n10317 , n10334 );
and ( n10738 , n10313 , n10334 );
or ( n10739 , n10736 , n10737 , n10738 );
and ( n10740 , n6796 , n6711 );
and ( n10741 , n7146 , n6332 );
nor ( n10742 , n10740 , n10741 );
xnor ( n10743 , n10742 , n6707 );
xor ( n10744 , n10739 , n10743 );
and ( n10745 , n6037 , n7630 );
and ( n10746 , n6391 , n7188 );
nor ( n10747 , n10745 , n10746 );
xnor ( n10748 , n10747 , n7626 );
and ( n10749 , n5419 , n8502 );
and ( n10750 , n5700 , n7970 );
nor ( n10751 , n10749 , n10750 );
xnor ( n10752 , n10751 , n8498 );
xor ( n10753 , n10748 , n10752 );
and ( n10754 , n10322 , n10326 );
and ( n10755 , n10326 , n10333 );
and ( n10756 , n10322 , n10333 );
or ( n10757 , n10754 , n10755 , n10756 );
and ( n10758 , n4916 , n9407 );
and ( n10759 , n5140 , n8872 );
nor ( n10760 , n10758 , n10759 );
xnor ( n10761 , n10760 , n9403 );
xor ( n10762 , n10757 , n10761 );
and ( n10763 , n4548 , n10329 );
and ( n10764 , n4696 , n9791 );
nor ( n10765 , n10763 , n10764 );
not ( n10766 , n10765 );
xor ( n10767 , n10762 , n10766 );
xor ( n10768 , n10753 , n10767 );
xor ( n10769 , n10744 , n10768 );
xor ( n10770 , n10735 , n10769 );
xor ( n10771 , n10726 , n10770 );
and ( n10772 , n10201 , n10205 );
and ( n10773 , n10205 , n10338 );
and ( n10774 , n10201 , n10338 );
or ( n10775 , n10772 , n10773 , n10774 );
xor ( n10776 , n10771 , n10775 );
and ( n10777 , n10187 , n10339 );
and ( n10778 , n10339 , n10344 );
and ( n10779 , n10187 , n10344 );
or ( n10780 , n10777 , n10778 , n10779 );
xor ( n10781 , n10776 , n10780 );
and ( n10782 , n10345 , n10346 );
xor ( n10783 , n10781 , n10782 );
buf ( n10784 , n10783 );
and ( n10785 , n10355 , n10356 );
and ( n10786 , n10356 , n10598 );
and ( n10787 , n10355 , n10598 );
or ( n10788 , n10785 , n10786 , n10787 );
and ( n10789 , n10446 , n10467 );
and ( n10790 , n10467 , n10492 );
and ( n10791 , n10446 , n10492 );
or ( n10792 , n10789 , n10790 , n10791 );
and ( n10793 , n10450 , n10454 );
and ( n10794 , n10454 , n10466 );
and ( n10795 , n10450 , n10466 );
or ( n10796 , n10793 , n10794 , n10795 );
and ( n10797 , n10437 , n4235 );
and ( n10798 , n10379 , n10383 );
and ( n10799 , n10383 , n10397 );
and ( n10800 , n10379 , n10397 );
or ( n10801 , n10798 , n10799 , n10800 );
and ( n10802 , n10403 , n10407 );
and ( n10803 , n10407 , n10420 );
and ( n10804 , n10403 , n10420 );
or ( n10805 , n10802 , n10803 , n10804 );
xor ( n10806 , n10801 , n10805 );
and ( n10807 , n10413 , n10417 );
and ( n10808 , n10417 , n10419 );
and ( n10809 , n10413 , n10419 );
or ( n10810 , n10807 , n10808 , n10809 );
not ( n10811 , n4733 );
and ( n10812 , n6853 , n5208 );
and ( n10813 , n7299 , n4976 );
nor ( n10814 , n10812 , n10813 );
xnor ( n10815 , n10814 , n5214 );
xor ( n10816 , n10811 , n10815 );
and ( n10817 , n5487 , n6496 );
and ( n10818 , n5791 , n6115 );
nor ( n10819 , n10817 , n10818 );
xnor ( n10820 , n10819 , n6453 );
xor ( n10821 , n10816 , n10820 );
xor ( n10822 , n10810 , n10821 );
and ( n10823 , n10387 , n10391 );
and ( n10824 , n10391 , n10396 );
and ( n10825 , n10387 , n10396 );
or ( n10826 , n10823 , n10824 , n10825 );
buf ( n10827 , n10412 );
xor ( n10828 , n10826 , n10827 );
and ( n10829 , n6120 , n5773 );
and ( n10830 , n6444 , n5519 );
nor ( n10831 , n10829 , n10830 );
xnor ( n10832 , n10831 , n5763 );
and ( n10833 , n4965 , n7277 );
and ( n10834 , n5195 , n6864 );
nor ( n10835 , n10833 , n10834 );
xnor ( n10836 , n10835 , n7283 );
xor ( n10837 , n10832 , n10836 );
and ( n10838 , n4724 , n7274 );
xor ( n10839 , n10837 , n10838 );
xor ( n10840 , n10828 , n10839 );
xor ( n10841 , n10822 , n10840 );
xor ( n10842 , n10806 , n10841 );
and ( n10843 , n10375 , n10398 );
and ( n10844 , n10398 , n10421 );
and ( n10845 , n10375 , n10421 );
or ( n10846 , n10843 , n10844 , n10845 );
xor ( n10847 , n10842 , n10846 );
and ( n10848 , n10422 , n10426 );
and ( n10849 , n10426 , n10431 );
and ( n10850 , n10422 , n10431 );
or ( n10851 , n10848 , n10849 , n10850 );
xor ( n10852 , n10847 , n10851 );
and ( n10853 , n10432 , n10433 );
xor ( n10854 , n10852 , n10853 );
buf ( n10855 , n10854 );
buf ( n10856 , n10855 );
buf ( n10857 , n10856 );
and ( n10858 , n10857 , n4232 );
nor ( n10859 , n10797 , n10858 );
xnor ( n10860 , n10859 , n4230 );
xor ( n10861 , n10796 , n10860 );
and ( n10862 , n10481 , n10485 );
and ( n10863 , n10485 , n10490 );
and ( n10864 , n10481 , n10490 );
or ( n10865 , n10862 , n10863 , n10864 );
and ( n10866 , n7752 , n4788 );
and ( n10867 , n8179 , n4611 );
nor ( n10868 , n10866 , n10867 );
xnor ( n10869 , n10868 , n4784 );
xor ( n10870 , n10865 , n10869 );
and ( n10871 , n6907 , n5270 );
and ( n10872 , n7324 , n5021 );
nor ( n10873 , n10871 , n10872 );
xnor ( n10874 , n10873 , n5266 );
xor ( n10875 , n10870 , n10874 );
xor ( n10876 , n10861 , n10875 );
xor ( n10877 , n10792 , n10876 );
and ( n10878 , n10365 , n10369 );
and ( n10879 , n10369 , n10440 );
and ( n10880 , n10365 , n10440 );
or ( n10881 , n10878 , n10879 , n10880 );
and ( n10882 , n10472 , n10476 );
and ( n10883 , n10476 , n10491 );
and ( n10884 , n10472 , n10491 );
or ( n10885 , n10882 , n10883 , n10884 );
xor ( n10886 , n10881 , n10885 );
and ( n10887 , n9583 , n4319 );
and ( n10888 , n9989 , n4310 );
nor ( n10889 , n10887 , n10888 );
xnor ( n10890 , n10889 , n4315 );
and ( n10891 , n8640 , n4298 );
and ( n10892 , n9110 , n4287 );
nor ( n10893 , n10891 , n10892 );
xnor ( n10894 , n10893 , n4294 );
xor ( n10895 , n10890 , n10894 );
and ( n10896 , n10459 , n10463 );
and ( n10897 , n10463 , n10465 );
and ( n10898 , n10459 , n10465 );
or ( n10899 , n10896 , n10897 , n10898 );
and ( n10900 , n6168 , n5850 );
and ( n10901 , n6516 , n5566 );
nor ( n10902 , n10900 , n10901 );
xnor ( n10903 , n10902 , n5846 );
xor ( n10904 , n10899 , n10903 );
and ( n10905 , n5535 , n6554 );
and ( n10906 , n5818 , n6205 );
nor ( n10907 , n10905 , n10906 );
xnor ( n10908 , n10907 , n6550 );
and ( n10909 , n4999 , n7356 );
and ( n10910 , n5247 , n6953 );
nor ( n10911 , n10909 , n10910 );
xnor ( n10912 , n10911 , n7352 );
xor ( n10913 , n10908 , n10912 );
and ( n10914 , n4770 , n7349 );
xor ( n10915 , n10913 , n10914 );
xor ( n10916 , n10904 , n10915 );
xor ( n10917 , n10895 , n10916 );
xor ( n10918 , n10886 , n10917 );
xor ( n10919 , n10877 , n10918 );
and ( n10920 , n10361 , n10441 );
and ( n10921 , n10441 , n10493 );
and ( n10922 , n10361 , n10493 );
or ( n10923 , n10920 , n10921 , n10922 );
xor ( n10924 , n10919 , n10923 );
and ( n10925 , n10494 , n10498 );
and ( n10926 , n10499 , n10502 );
or ( n10927 , n10925 , n10926 );
xor ( n10928 , n10924 , n10927 );
buf ( n10929 , n10928 );
and ( n10930 , n10572 , n10576 );
and ( n10931 , n10576 , n10581 );
and ( n10932 , n10572 , n10581 );
or ( n10933 , n10930 , n10931 , n10932 );
and ( n10934 , n10542 , n10546 );
and ( n10935 , n10546 , n10560 );
and ( n10936 , n10542 , n10560 );
or ( n10937 , n10934 , n10935 , n10936 );
and ( n10938 , n10534 , n4418 );
buf ( n10939 , n3812 );
buf ( n10940 , n10939 );
and ( n10941 , n10940 , n4415 );
nor ( n10942 , n10938 , n10941 );
xnor ( n10943 , n10942 , n4413 );
xor ( n10944 , n10937 , n10943 );
and ( n10945 , n10515 , n10519 );
and ( n10946 , n10519 , n10524 );
and ( n10947 , n10515 , n10524 );
or ( n10948 , n10945 , n10946 , n10947 );
and ( n10949 , n10553 , n10554 );
and ( n10950 , n10554 , n10559 );
and ( n10951 , n10553 , n10559 );
or ( n10952 , n10949 , n10950 , n10951 );
xor ( n10953 , n10948 , n10952 );
and ( n10954 , n8728 , n4402 );
and ( n10955 , n9164 , n4391 );
nor ( n10956 , n10954 , n10955 );
xnor ( n10957 , n10956 , n4398 );
xor ( n10958 , n10953 , n10957 );
xor ( n10959 , n10944 , n10958 );
and ( n10960 , n10509 , n10513 );
and ( n10961 , n10513 , n10525 );
and ( n10962 , n10509 , n10525 );
or ( n10963 , n10960 , n10961 , n10962 );
and ( n10964 , n10531 , n10537 );
and ( n10965 , n10537 , n10561 );
and ( n10966 , n10531 , n10561 );
or ( n10967 , n10964 , n10965 , n10966 );
xor ( n10968 , n10963 , n10967 );
and ( n10969 , n9629 , n4433 );
and ( n10970 , n10072 , n4431 );
nor ( n10971 , n10969 , n10970 );
xnor ( n10972 , n10971 , n4441 );
and ( n10973 , n7857 , n4835 );
and ( n10974 , n8303 , n4648 );
nor ( n10975 , n10973 , n10974 );
xnor ( n10976 , n10975 , n4831 );
and ( n10977 , n6995 , n5323 );
and ( n10978 , n7417 , n5064 );
nor ( n10979 , n10977 , n10978 );
xnor ( n10980 , n10979 , n5319 );
xor ( n10981 , n10976 , n10980 );
and ( n10982 , n6235 , n5922 );
and ( n10983 , n6604 , n5616 );
nor ( n10984 , n10982 , n10983 );
xnor ( n10985 , n10984 , n5918 );
xor ( n10986 , n10981 , n10985 );
xor ( n10987 , n10972 , n10986 );
and ( n10988 , n5042 , n7444 );
and ( n10989 , n5300 , n7026 );
nor ( n10990 , n10988 , n10989 );
xnor ( n10991 , n10990 , n7440 );
and ( n10992 , n4817 , n7437 );
xor ( n10993 , n10991 , n10992 );
and ( n10994 , n10551 , n10552 );
xor ( n10995 , n10993 , n10994 );
and ( n10996 , n5588 , n6627 );
and ( n10997 , n5893 , n6272 );
nor ( n10998 , n10996 , n10997 );
xnor ( n10999 , n10998 , n6623 );
xor ( n11000 , n10995 , n10999 );
xor ( n11001 , n10987 , n11000 );
xor ( n11002 , n10968 , n11001 );
xor ( n11003 , n10959 , n11002 );
and ( n11004 , n10505 , n10526 );
and ( n11005 , n10526 , n10562 );
and ( n11006 , n10505 , n10562 );
or ( n11007 , n11004 , n11005 , n11006 );
xor ( n11008 , n11003 , n11007 );
xor ( n11009 , n10933 , n11008 );
and ( n11010 , n10563 , n10567 );
and ( n11011 , n10567 , n10582 );
and ( n11012 , n10563 , n10582 );
or ( n11013 , n11010 , n11011 , n11012 );
xor ( n11014 , n11009 , n11013 );
and ( n11015 , n10583 , n10587 );
and ( n11016 , n10588 , n10589 );
or ( n11017 , n11015 , n11016 );
xor ( n11018 , n11014 , n11017 );
buf ( n11019 , n11018 );
not ( n11020 , n454 );
and ( n11021 , n11020 , n10929 );
and ( n11022 , n11019 , n454 );
or ( n11023 , n11021 , n11022 );
buf ( n11024 , n11023 );
buf ( n11025 , n11024 );
and ( n11026 , n11025 , n4505 );
xor ( n11027 , n10788 , n11026 );
and ( n11028 , n9718 , n5089 );
and ( n11029 , n10156 , n4866 );
xor ( n11030 , n11028 , n11029 );
and ( n11031 , n10597 , n4557 );
xor ( n11032 , n11030 , n11031 );
xor ( n11033 , n11027 , n11032 );
and ( n11034 , n10352 , n10353 );
and ( n11035 , n10353 , n10599 );
and ( n11036 , n10352 , n10599 );
or ( n11037 , n11034 , n11035 , n11036 );
xor ( n11038 , n11033 , n11037 );
and ( n11039 , n10600 , n10604 );
and ( n11040 , n10604 , n10609 );
and ( n11041 , n10600 , n10609 );
or ( n11042 , n11039 , n11040 , n11041 );
xor ( n11043 , n11038 , n11042 );
or ( n11044 , n10610 , n10611 );
xnor ( n11045 , n11043 , n11044 );
and ( n11046 , n10612 , n10613 );
xor ( n11047 , n11045 , n11046 );
buf ( n11048 , n11047 );
not ( n11049 , n4509 );
and ( n11050 , n11049 , n10784 );
and ( n11051 , n11048 , n4509 );
or ( n11052 , n11050 , n11051 );
and ( n11053 , n10623 , n10725 );
and ( n11054 , n10725 , n10770 );
and ( n11055 , n10623 , n10770 );
or ( n11056 , n11053 , n11054 , n11055 );
and ( n11057 , n10627 , n10709 );
and ( n11058 , n10709 , n10724 );
and ( n11059 , n10627 , n10724 );
or ( n11060 , n11057 , n11058 , n11059 );
and ( n11061 , n10714 , n10718 );
and ( n11062 , n10718 , n10723 );
and ( n11063 , n10714 , n10723 );
or ( n11064 , n11061 , n11062 , n11063 );
and ( n11065 , n9885 , n4938 );
and ( n11066 , n10287 , n4711 );
nor ( n11067 , n11065 , n11066 );
xnor ( n11068 , n11067 , n4934 );
xor ( n11069 , n11064 , n11068 );
and ( n11070 , n10748 , n10752 );
and ( n11071 , n10752 , n10767 );
and ( n11072 , n10748 , n10767 );
or ( n11073 , n11070 , n11071 , n11072 );
and ( n11074 , n8057 , n6068 );
and ( n11075 , n8462 , n5730 );
nor ( n11076 , n11074 , n11075 );
xnor ( n11077 , n11076 , n6064 );
xor ( n11078 , n11073 , n11077 );
and ( n11079 , n7146 , n6711 );
and ( n11080 , n7587 , n6332 );
nor ( n11081 , n11079 , n11080 );
xnor ( n11082 , n11081 , n6707 );
xor ( n11083 , n11078 , n11082 );
xor ( n11084 , n11069 , n11083 );
xor ( n11085 , n11060 , n11084 );
and ( n11086 , n10730 , n10734 );
and ( n11087 , n10734 , n10769 );
and ( n11088 , n10730 , n10769 );
or ( n11089 , n11086 , n11087 , n11088 );
and ( n11090 , n10706 , n4524 );
and ( n11091 , n10675 , n10679 );
and ( n11092 , n10679 , n10694 );
and ( n11093 , n10675 , n10694 );
or ( n11094 , n11091 , n11092 , n11093 );
and ( n11095 , n10635 , n10639 );
and ( n11096 , n10639 , n10674 );
and ( n11097 , n10635 , n10674 );
or ( n11098 , n11095 , n11096 , n11097 );
and ( n11099 , n10684 , n10688 );
and ( n11100 , n10688 , n10693 );
and ( n11101 , n10684 , n10693 );
or ( n11102 , n11099 , n11100 , n11101 );
xor ( n11103 , n11098 , n11102 );
and ( n11104 , n10663 , n10667 );
and ( n11105 , n10667 , n10672 );
and ( n11106 , n10663 , n10672 );
or ( n11107 , n11104 , n11105 , n11106 );
and ( n11108 , n9848 , n4898 );
not ( n11109 , n11108 );
xnor ( n11110 , n11109 , n4904 );
not ( n11111 , n11110 );
xor ( n11112 , n11107 , n11111 );
and ( n11113 , n8001 , n6008 );
and ( n11114 , n8409 , n5689 );
nor ( n11115 , n11113 , n11114 );
xnor ( n11116 , n11115 , n6004 );
xor ( n11117 , n11112 , n11116 );
and ( n11118 , n10644 , n10658 );
and ( n11119 , n10658 , n10673 );
and ( n11120 , n10644 , n10673 );
or ( n11121 , n11118 , n11119 , n11120 );
xor ( n11122 , n11117 , n11121 );
and ( n11123 , n10648 , n10652 );
and ( n11124 , n10652 , n10657 );
and ( n11125 , n10648 , n10657 );
or ( n11126 , n11123 , n11124 , n11125 );
and ( n11127 , n8900 , n5405 );
and ( n11128 , n9297 , n5132 );
nor ( n11129 , n11127 , n11128 );
xnor ( n11130 , n11129 , n5401 );
and ( n11131 , n5672 , n8382 );
and ( n11132 , n5995 , n8042 );
nor ( n11133 , n11131 , n11132 );
xnor ( n11134 , n11133 , n8378 );
xor ( n11135 , n11130 , n11134 );
and ( n11136 , n5387 , n8375 );
xor ( n11137 , n11135 , n11136 );
xor ( n11138 , n11126 , n11137 );
or ( n11139 , n10633 , n10634 );
and ( n11140 , n7092 , n6761 );
and ( n11141 , n7531 , n6379 );
nor ( n11142 , n11140 , n11141 );
xnor ( n11143 , n11142 , n6757 );
xor ( n11144 , n11139 , n11143 );
and ( n11145 , n6353 , n7559 );
and ( n11146 , n6748 , n7107 );
nor ( n11147 , n11145 , n11146 );
xnor ( n11148 , n11147 , n7555 );
xor ( n11149 , n11144 , n11148 );
xor ( n11150 , n11138 , n11149 );
xor ( n11151 , n11122 , n11150 );
xor ( n11152 , n11103 , n11151 );
xor ( n11153 , n11094 , n11152 );
and ( n11154 , n10632 , n10695 );
and ( n11155 , n10695 , n10700 );
and ( n11156 , n10632 , n10700 );
or ( n11157 , n11154 , n11155 , n11156 );
xor ( n11158 , n11153 , n11157 );
and ( n11159 , n10701 , n10702 );
xor ( n11160 , n11158 , n11159 );
buf ( n11161 , n11160 );
buf ( n11162 , n11161 );
buf ( n11163 , n11162 );
and ( n11164 , n11163 , n4145 );
nor ( n11165 , n11090 , n11164 );
xnor ( n11166 , n11165 , n4521 );
xor ( n11167 , n11089 , n11166 );
and ( n11168 , n10739 , n10743 );
and ( n11169 , n10743 , n10768 );
and ( n11170 , n10739 , n10768 );
or ( n11171 , n11168 , n11169 , n11170 );
and ( n11172 , n8968 , n5441 );
and ( n11173 , n9367 , n5161 );
nor ( n11174 , n11172 , n11173 );
xnor ( n11175 , n11174 , n5437 );
xor ( n11176 , n11171 , n11175 );
and ( n11177 , n10757 , n10761 );
and ( n11178 , n10761 , n10766 );
and ( n11179 , n10757 , n10766 );
or ( n11180 , n11177 , n11178 , n11179 );
and ( n11181 , n6391 , n7630 );
and ( n11182 , n6796 , n7188 );
nor ( n11183 , n11181 , n11182 );
xnor ( n11184 , n11183 , n7626 );
xor ( n11185 , n11180 , n11184 );
and ( n11186 , n5700 , n8502 );
and ( n11187 , n6037 , n7970 );
nor ( n11188 , n11186 , n11187 );
xnor ( n11189 , n11188 , n8498 );
and ( n11190 , n5140 , n9407 );
and ( n11191 , n5419 , n8872 );
nor ( n11192 , n11190 , n11191 );
xnor ( n11193 , n11192 , n9403 );
xor ( n11194 , n11189 , n11193 );
and ( n11195 , n4696 , n10329 );
and ( n11196 , n4916 , n9791 );
nor ( n11197 , n11195 , n11196 );
not ( n11198 , n11197 );
xor ( n11199 , n11194 , n11198 );
xor ( n11200 , n11185 , n11199 );
xor ( n11201 , n11176 , n11200 );
xor ( n11202 , n11167 , n11201 );
xor ( n11203 , n11085 , n11202 );
xor ( n11204 , n11056 , n11203 );
and ( n11205 , n10771 , n10775 );
and ( n11206 , n10775 , n10780 );
and ( n11207 , n10771 , n10780 );
or ( n11208 , n11205 , n11206 , n11207 );
xor ( n11209 , n11204 , n11208 );
and ( n11210 , n10781 , n10782 );
xor ( n11211 , n11209 , n11210 );
buf ( n11212 , n11211 );
and ( n11213 , n10156 , n5089 );
and ( n11214 , n10597 , n4866 );
xor ( n11215 , n11213 , n11214 );
and ( n11216 , n11025 , n4557 );
xor ( n11217 , n11215 , n11216 );
and ( n11218 , n11028 , n11029 );
and ( n11219 , n11029 , n11031 );
and ( n11220 , n11028 , n11031 );
or ( n11221 , n11218 , n11219 , n11220 );
and ( n11222 , n10881 , n10885 );
and ( n11223 , n10885 , n10917 );
and ( n11224 , n10881 , n10917 );
or ( n11225 , n11222 , n11223 , n11224 );
and ( n11226 , n10796 , n10860 );
and ( n11227 , n10860 , n10875 );
and ( n11228 , n10796 , n10875 );
or ( n11229 , n11226 , n11227 , n11228 );
and ( n11230 , n10890 , n10894 );
and ( n11231 , n10894 , n10916 );
and ( n11232 , n10890 , n10916 );
or ( n11233 , n11230 , n11231 , n11232 );
xor ( n11234 , n11229 , n11233 );
and ( n11235 , n10899 , n10903 );
and ( n11236 , n10903 , n10915 );
and ( n11237 , n10899 , n10915 );
or ( n11238 , n11235 , n11236 , n11237 );
and ( n11239 , n10857 , n4235 );
and ( n11240 , n10826 , n10827 );
and ( n11241 , n10827 , n10839 );
and ( n11242 , n10826 , n10839 );
or ( n11243 , n11240 , n11241 , n11242 );
and ( n11244 , n10810 , n10821 );
and ( n11245 , n10821 , n10840 );
and ( n11246 , n10810 , n10840 );
or ( n11247 , n11244 , n11245 , n11246 );
xor ( n11248 , n11243 , n11247 );
and ( n11249 , n10811 , n10815 );
and ( n11250 , n10815 , n10820 );
and ( n11251 , n10811 , n10820 );
or ( n11252 , n11249 , n11250 , n11251 );
and ( n11253 , n7299 , n5208 );
not ( n11254 , n11253 );
xnor ( n11255 , n11254 , n5214 );
and ( n11256 , n5195 , n7277 );
and ( n11257 , n5487 , n6864 );
nor ( n11258 , n11256 , n11257 );
xnor ( n11259 , n11258 , n7283 );
xor ( n11260 , n11255 , n11259 );
and ( n11261 , n4965 , n7274 );
xor ( n11262 , n11260 , n11261 );
xor ( n11263 , n11252 , n11262 );
and ( n11264 , n10832 , n10836 );
and ( n11265 , n10836 , n10838 );
and ( n11266 , n10832 , n10838 );
or ( n11267 , n11264 , n11265 , n11266 );
and ( n11268 , n6444 , n5773 );
and ( n11269 , n6853 , n5519 );
nor ( n11270 , n11268 , n11269 );
xnor ( n11271 , n11270 , n5763 );
not ( n11272 , n11271 );
xor ( n11273 , n11267 , n11272 );
and ( n11274 , n5791 , n6496 );
and ( n11275 , n6120 , n6115 );
nor ( n11276 , n11274 , n11275 );
xnor ( n11277 , n11276 , n6453 );
xor ( n11278 , n11273 , n11277 );
xor ( n11279 , n11263 , n11278 );
xor ( n11280 , n11248 , n11279 );
and ( n11281 , n10801 , n10805 );
and ( n11282 , n10805 , n10841 );
and ( n11283 , n10801 , n10841 );
or ( n11284 , n11281 , n11282 , n11283 );
xor ( n11285 , n11280 , n11284 );
and ( n11286 , n10842 , n10846 );
and ( n11287 , n10846 , n10851 );
and ( n11288 , n10842 , n10851 );
or ( n11289 , n11286 , n11287 , n11288 );
xor ( n11290 , n11285 , n11289 );
and ( n11291 , n10852 , n10853 );
xor ( n11292 , n11290 , n11291 );
buf ( n11293 , n11292 );
buf ( n11294 , n11293 );
buf ( n11295 , n11294 );
and ( n11296 , n11295 , n4232 );
nor ( n11297 , n11239 , n11296 );
xnor ( n11298 , n11297 , n4230 );
xor ( n11299 , n11238 , n11298 );
and ( n11300 , n9989 , n4319 );
and ( n11301 , n10437 , n4310 );
nor ( n11302 , n11300 , n11301 );
xnor ( n11303 , n11302 , n4315 );
xor ( n11304 , n11299 , n11303 );
xor ( n11305 , n11234 , n11304 );
xor ( n11306 , n11225 , n11305 );
and ( n11307 , n10865 , n10869 );
and ( n11308 , n10869 , n10874 );
and ( n11309 , n10865 , n10874 );
or ( n11310 , n11307 , n11308 , n11309 );
and ( n11311 , n10908 , n10912 );
and ( n11312 , n10912 , n10914 );
and ( n11313 , n10908 , n10914 );
or ( n11314 , n11311 , n11312 , n11313 );
and ( n11315 , n7324 , n5270 );
and ( n11316 , n7752 , n5021 );
nor ( n11317 , n11315 , n11316 );
xnor ( n11318 , n11317 , n5266 );
xor ( n11319 , n11314 , n11318 );
and ( n11320 , n6516 , n5850 );
and ( n11321 , n6907 , n5566 );
nor ( n11322 , n11320 , n11321 );
xnor ( n11323 , n11322 , n5846 );
xor ( n11324 , n11319 , n11323 );
xor ( n11325 , n11310 , n11324 );
and ( n11326 , n5818 , n6554 );
and ( n11327 , n6168 , n6205 );
nor ( n11328 , n11326 , n11327 );
xnor ( n11329 , n11328 , n6550 );
and ( n11330 , n5247 , n7356 );
and ( n11331 , n5535 , n6953 );
nor ( n11332 , n11330 , n11331 );
xnor ( n11333 , n11332 , n7352 );
and ( n11334 , n4999 , n7349 );
xor ( n11335 , n11333 , n11334 );
xor ( n11336 , n11329 , n11335 );
and ( n11337 , n9110 , n4298 );
and ( n11338 , n9583 , n4287 );
nor ( n11339 , n11337 , n11338 );
xnor ( n11340 , n11339 , n4294 );
xor ( n11341 , n11336 , n11340 );
and ( n11342 , n8179 , n4788 );
and ( n11343 , n8640 , n4611 );
nor ( n11344 , n11342 , n11343 );
xnor ( n11345 , n11344 , n4784 );
xor ( n11346 , n11341 , n11345 );
xor ( n11347 , n11325 , n11346 );
xor ( n11348 , n11306 , n11347 );
and ( n11349 , n10792 , n10876 );
and ( n11350 , n10876 , n10918 );
and ( n11351 , n10792 , n10918 );
or ( n11352 , n11349 , n11350 , n11351 );
xor ( n11353 , n11348 , n11352 );
and ( n11354 , n10919 , n10923 );
and ( n11355 , n10924 , n10927 );
or ( n11356 , n11354 , n11355 );
xor ( n11357 , n11353 , n11356 );
buf ( n11358 , n11357 );
and ( n11359 , n10959 , n11002 );
and ( n11360 , n11002 , n11007 );
and ( n11361 , n10959 , n11007 );
or ( n11362 , n11359 , n11360 , n11361 );
and ( n11363 , n10963 , n10967 );
and ( n11364 , n10967 , n11001 );
and ( n11365 , n10963 , n11001 );
or ( n11366 , n11363 , n11364 , n11365 );
and ( n11367 , n10948 , n10952 );
and ( n11368 , n10952 , n10957 );
and ( n11369 , n10948 , n10957 );
or ( n11370 , n11367 , n11368 , n11369 );
and ( n11371 , n10972 , n10986 );
and ( n11372 , n10986 , n11000 );
and ( n11373 , n10972 , n11000 );
or ( n11374 , n11371 , n11372 , n11373 );
xor ( n11375 , n11370 , n11374 );
and ( n11376 , n10993 , n10994 );
and ( n11377 , n10994 , n10999 );
and ( n11378 , n10993 , n10999 );
or ( n11379 , n11376 , n11377 , n11378 );
and ( n11380 , n7417 , n5323 );
and ( n11381 , n7857 , n5064 );
nor ( n11382 , n11380 , n11381 );
xnor ( n11383 , n11382 , n5319 );
xor ( n11384 , n11379 , n11383 );
and ( n11385 , n5893 , n6627 );
and ( n11386 , n6235 , n6272 );
nor ( n11387 , n11385 , n11386 );
xnor ( n11388 , n11387 , n6623 );
xor ( n11389 , n11384 , n11388 );
xor ( n11390 , n11375 , n11389 );
xor ( n11391 , n11366 , n11390 );
and ( n11392 , n10937 , n10943 );
and ( n11393 , n10943 , n10958 );
and ( n11394 , n10937 , n10958 );
or ( n11395 , n11392 , n11393 , n11394 );
and ( n11396 , n10940 , n4418 );
buf ( n11397 , n3894 );
buf ( n11398 , n11397 );
and ( n11399 , n11398 , n4415 );
nor ( n11400 , n11396 , n11399 );
xnor ( n11401 , n11400 , n4413 );
and ( n11402 , n10072 , n4433 );
and ( n11403 , n10534 , n4431 );
nor ( n11404 , n11402 , n11403 );
xnor ( n11405 , n11404 , n4441 );
xor ( n11406 , n11401 , n11405 );
and ( n11407 , n9164 , n4402 );
and ( n11408 , n9629 , n4391 );
nor ( n11409 , n11407 , n11408 );
xnor ( n11410 , n11409 , n4398 );
xor ( n11411 , n11406 , n11410 );
xor ( n11412 , n11395 , n11411 );
and ( n11413 , n10976 , n10980 );
and ( n11414 , n10980 , n10985 );
and ( n11415 , n10976 , n10985 );
or ( n11416 , n11413 , n11414 , n11415 );
and ( n11417 , n8303 , n4835 );
and ( n11418 , n8728 , n4648 );
nor ( n11419 , n11417 , n11418 );
xnor ( n11420 , n11419 , n4831 );
xor ( n11421 , n11416 , n11420 );
and ( n11422 , n5300 , n7444 );
and ( n11423 , n5588 , n7026 );
nor ( n11424 , n11422 , n11423 );
xnor ( n11425 , n11424 , n7440 );
and ( n11426 , n5042 , n7437 );
xor ( n11427 , n11425 , n11426 );
and ( n11428 , n10991 , n10992 );
xor ( n11429 , n11427 , n11428 );
and ( n11430 , n6604 , n5922 );
and ( n11431 , n6995 , n5616 );
nor ( n11432 , n11430 , n11431 );
xnor ( n11433 , n11432 , n5918 );
xor ( n11434 , n11429 , n11433 );
xor ( n11435 , n11421 , n11434 );
xor ( n11436 , n11412 , n11435 );
xor ( n11437 , n11391 , n11436 );
xor ( n11438 , n11362 , n11437 );
and ( n11439 , n10933 , n11008 );
and ( n11440 , n11008 , n11013 );
and ( n11441 , n10933 , n11013 );
or ( n11442 , n11439 , n11440 , n11441 );
xor ( n11443 , n11438 , n11442 );
and ( n11444 , n11014 , n11017 );
xor ( n11445 , n11443 , n11444 );
buf ( n11446 , n11445 );
not ( n11447 , n454 );
and ( n11448 , n11447 , n11358 );
and ( n11449 , n11446 , n454 );
or ( n11450 , n11448 , n11449 );
buf ( n11451 , n11450 );
buf ( n11452 , n11451 );
and ( n11453 , n11452 , n4505 );
xor ( n11454 , n11221 , n11453 );
xor ( n11455 , n11217 , n11454 );
and ( n11456 , n10788 , n11026 );
and ( n11457 , n11026 , n11032 );
and ( n11458 , n10788 , n11032 );
or ( n11459 , n11456 , n11457 , n11458 );
xor ( n11460 , n11455 , n11459 );
and ( n11461 , n11033 , n11037 );
and ( n11462 , n11037 , n11042 );
and ( n11463 , n11033 , n11042 );
or ( n11464 , n11461 , n11462 , n11463 );
xor ( n11465 , n11460 , n11464 );
or ( n11466 , n11043 , n11044 );
xor ( n11467 , n11465 , n11466 );
not ( n11468 , n11467 );
and ( n11469 , n11045 , n11046 );
xor ( n11470 , n11468 , n11469 );
buf ( n11471 , n11470 );
not ( n11472 , n4509 );
and ( n11473 , n11472 , n11212 );
and ( n11474 , n11471 , n4509 );
or ( n11475 , n11473 , n11474 );
and ( n11476 , n11089 , n11166 );
and ( n11477 , n11166 , n11201 );
and ( n11478 , n11089 , n11201 );
or ( n11479 , n11476 , n11477 , n11478 );
and ( n11480 , n11073 , n11077 );
and ( n11481 , n11077 , n11082 );
and ( n11482 , n11073 , n11082 );
or ( n11483 , n11480 , n11481 , n11482 );
and ( n11484 , n11171 , n11175 );
and ( n11485 , n11175 , n11200 );
and ( n11486 , n11171 , n11200 );
or ( n11487 , n11484 , n11485 , n11486 );
xor ( n11488 , n11483 , n11487 );
and ( n11489 , n10287 , n4938 );
and ( n11490 , n10706 , n4711 );
nor ( n11491 , n11489 , n11490 );
xnor ( n11492 , n11491 , n4934 );
xor ( n11493 , n11488 , n11492 );
xor ( n11494 , n11479 , n11493 );
and ( n11495 , n11064 , n11068 );
and ( n11496 , n11068 , n11083 );
and ( n11497 , n11064 , n11083 );
or ( n11498 , n11495 , n11496 , n11497 );
and ( n11499 , n11163 , n4524 );
and ( n11500 , n11098 , n11102 );
and ( n11501 , n11102 , n11151 );
and ( n11502 , n11098 , n11151 );
or ( n11503 , n11500 , n11501 , n11502 );
and ( n11504 , n11126 , n11137 );
and ( n11505 , n11137 , n11149 );
and ( n11506 , n11126 , n11149 );
or ( n11507 , n11504 , n11505 , n11506 );
and ( n11508 , n11107 , n11111 );
and ( n11509 , n11111 , n11116 );
and ( n11510 , n11107 , n11116 );
or ( n11511 , n11508 , n11509 , n11510 );
and ( n11512 , n11130 , n11134 );
and ( n11513 , n11134 , n11136 );
and ( n11514 , n11130 , n11136 );
or ( n11515 , n11512 , n11513 , n11514 );
buf ( n11516 , n11110 );
xor ( n11517 , n11515 , n11516 );
and ( n11518 , n8409 , n6008 );
and ( n11519 , n8900 , n5689 );
nor ( n11520 , n11518 , n11519 );
xnor ( n11521 , n11520 , n6004 );
xor ( n11522 , n11517 , n11521 );
xor ( n11523 , n11511 , n11522 );
and ( n11524 , n11139 , n11143 );
and ( n11525 , n11143 , n11148 );
and ( n11526 , n11139 , n11148 );
or ( n11527 , n11524 , n11525 , n11526 );
not ( n11528 , n4904 );
and ( n11529 , n5995 , n8382 );
and ( n11530 , n6353 , n8042 );
nor ( n11531 , n11529 , n11530 );
xnor ( n11532 , n11531 , n8378 );
xor ( n11533 , n11528 , n11532 );
and ( n11534 , n5672 , n8375 );
xor ( n11535 , n11533 , n11534 );
xor ( n11536 , n11527 , n11535 );
and ( n11537 , n9297 , n5405 );
and ( n11538 , n9848 , n5132 );
nor ( n11539 , n11537 , n11538 );
xnor ( n11540 , n11539 , n5401 );
and ( n11541 , n7531 , n6761 );
and ( n11542 , n8001 , n6379 );
nor ( n11543 , n11541 , n11542 );
xnor ( n11544 , n11543 , n6757 );
xor ( n11545 , n11540 , n11544 );
and ( n11546 , n6748 , n7559 );
and ( n11547 , n7092 , n7107 );
nor ( n11548 , n11546 , n11547 );
xnor ( n11549 , n11548 , n7555 );
xor ( n11550 , n11545 , n11549 );
xor ( n11551 , n11536 , n11550 );
xor ( n11552 , n11523 , n11551 );
xor ( n11553 , n11507 , n11552 );
and ( n11554 , n11117 , n11121 );
and ( n11555 , n11121 , n11150 );
and ( n11556 , n11117 , n11150 );
or ( n11557 , n11554 , n11555 , n11556 );
xor ( n11558 , n11553 , n11557 );
xor ( n11559 , n11503 , n11558 );
and ( n11560 , n11094 , n11152 );
and ( n11561 , n11152 , n11157 );
and ( n11562 , n11094 , n11157 );
or ( n11563 , n11560 , n11561 , n11562 );
xor ( n11564 , n11559 , n11563 );
and ( n11565 , n11158 , n11159 );
xor ( n11566 , n11564 , n11565 );
buf ( n11567 , n11566 );
buf ( n11568 , n11567 );
buf ( n11569 , n11568 );
and ( n11570 , n11569 , n4145 );
nor ( n11571 , n11499 , n11570 );
xnor ( n11572 , n11571 , n4521 );
xor ( n11573 , n11498 , n11572 );
and ( n11574 , n9367 , n5441 );
and ( n11575 , n9885 , n5161 );
nor ( n11576 , n11574 , n11575 );
xnor ( n11577 , n11576 , n5437 );
and ( n11578 , n11180 , n11184 );
and ( n11579 , n11184 , n11199 );
and ( n11580 , n11180 , n11199 );
or ( n11581 , n11578 , n11579 , n11580 );
and ( n11582 , n8462 , n6068 );
and ( n11583 , n8968 , n5730 );
nor ( n11584 , n11582 , n11583 );
xnor ( n11585 , n11584 , n6064 );
xor ( n11586 , n11581 , n11585 );
and ( n11587 , n7587 , n6711 );
and ( n11588 , n8057 , n6332 );
nor ( n11589 , n11587 , n11588 );
xnor ( n11590 , n11589 , n6707 );
xor ( n11591 , n11586 , n11590 );
xor ( n11592 , n11577 , n11591 );
and ( n11593 , n11189 , n11193 );
and ( n11594 , n11193 , n11198 );
and ( n11595 , n11189 , n11198 );
or ( n11596 , n11593 , n11594 , n11595 );
and ( n11597 , n6796 , n7630 );
and ( n11598 , n7146 , n7188 );
nor ( n11599 , n11597 , n11598 );
xnor ( n11600 , n11599 , n7626 );
xor ( n11601 , n11596 , n11600 );
and ( n11602 , n6037 , n8502 );
and ( n11603 , n6391 , n7970 );
nor ( n11604 , n11602 , n11603 );
xnor ( n11605 , n11604 , n8498 );
and ( n11606 , n5419 , n9407 );
and ( n11607 , n5700 , n8872 );
nor ( n11608 , n11606 , n11607 );
xnor ( n11609 , n11608 , n9403 );
xor ( n11610 , n11605 , n11609 );
and ( n11611 , n4916 , n10329 );
and ( n11612 , n5140 , n9791 );
nor ( n11613 , n11611 , n11612 );
not ( n11614 , n11613 );
xor ( n11615 , n11610 , n11614 );
xor ( n11616 , n11601 , n11615 );
xor ( n11617 , n11592 , n11616 );
xor ( n11618 , n11573 , n11617 );
xor ( n11619 , n11494 , n11618 );
and ( n11620 , n11060 , n11084 );
and ( n11621 , n11084 , n11202 );
and ( n11622 , n11060 , n11202 );
or ( n11623 , n11620 , n11621 , n11622 );
xor ( n11624 , n11619 , n11623 );
and ( n11625 , n11056 , n11203 );
and ( n11626 , n11203 , n11208 );
and ( n11627 , n11056 , n11208 );
or ( n11628 , n11625 , n11626 , n11627 );
xor ( n11629 , n11624 , n11628 );
and ( n11630 , n11209 , n11210 );
xor ( n11631 , n11629 , n11630 );
buf ( n11632 , n11631 );
and ( n11633 , n11221 , n11453 );
and ( n11634 , n10597 , n5089 );
and ( n11635 , n11025 , n4866 );
xor ( n11636 , n11634 , n11635 );
and ( n11637 , n11452 , n4557 );
xor ( n11638 , n11636 , n11637 );
and ( n11639 , n11229 , n11233 );
and ( n11640 , n11233 , n11304 );
and ( n11641 , n11229 , n11304 );
or ( n11642 , n11639 , n11640 , n11641 );
and ( n11643 , n11238 , n11298 );
and ( n11644 , n11298 , n11303 );
and ( n11645 , n11238 , n11303 );
or ( n11646 , n11643 , n11644 , n11645 );
and ( n11647 , n11336 , n11340 );
and ( n11648 , n11340 , n11345 );
and ( n11649 , n11336 , n11345 );
or ( n11650 , n11647 , n11648 , n11649 );
xor ( n11651 , n11646 , n11650 );
and ( n11652 , n11295 , n4235 );
and ( n11653 , n11243 , n11247 );
and ( n11654 , n11247 , n11279 );
and ( n11655 , n11243 , n11279 );
or ( n11656 , n11653 , n11654 , n11655 );
and ( n11657 , n11267 , n11272 );
and ( n11658 , n11272 , n11277 );
and ( n11659 , n11267 , n11277 );
or ( n11660 , n11657 , n11658 , n11659 );
and ( n11661 , n11252 , n11262 );
and ( n11662 , n11262 , n11278 );
and ( n11663 , n11252 , n11278 );
or ( n11664 , n11661 , n11662 , n11663 );
xor ( n11665 , n11660 , n11664 );
and ( n11666 , n11255 , n11259 );
and ( n11667 , n11259 , n11261 );
and ( n11668 , n11255 , n11261 );
or ( n11669 , n11666 , n11667 , n11668 );
not ( n11670 , n5214 );
and ( n11671 , n6853 , n5773 );
and ( n11672 , n7299 , n5519 );
nor ( n11673 , n11671 , n11672 );
xnor ( n11674 , n11673 , n5763 );
xor ( n11675 , n11670 , n11674 );
and ( n11676 , n5487 , n7277 );
and ( n11677 , n5791 , n6864 );
nor ( n11678 , n11676 , n11677 );
xnor ( n11679 , n11678 , n7283 );
xor ( n11680 , n11675 , n11679 );
xor ( n11681 , n11669 , n11680 );
buf ( n11682 , n11271 );
and ( n11683 , n6120 , n6496 );
and ( n11684 , n6444 , n6115 );
nor ( n11685 , n11683 , n11684 );
xnor ( n11686 , n11685 , n6453 );
xor ( n11687 , n11682 , n11686 );
and ( n11688 , n5195 , n7274 );
xor ( n11689 , n11687 , n11688 );
xor ( n11690 , n11681 , n11689 );
xor ( n11691 , n11665 , n11690 );
xor ( n11692 , n11656 , n11691 );
and ( n11693 , n11280 , n11284 );
and ( n11694 , n11284 , n11289 );
and ( n11695 , n11280 , n11289 );
or ( n11696 , n11693 , n11694 , n11695 );
xor ( n11697 , n11692 , n11696 );
and ( n11698 , n11290 , n11291 );
xor ( n11699 , n11697 , n11698 );
buf ( n11700 , n11699 );
buf ( n11701 , n11700 );
buf ( n11702 , n11701 );
and ( n11703 , n11702 , n4232 );
nor ( n11704 , n11652 , n11703 );
xnor ( n11705 , n11704 , n4230 );
xor ( n11706 , n11651 , n11705 );
xor ( n11707 , n11642 , n11706 );
and ( n11708 , n11310 , n11324 );
and ( n11709 , n11324 , n11346 );
and ( n11710 , n11310 , n11346 );
or ( n11711 , n11708 , n11709 , n11710 );
and ( n11712 , n11314 , n11318 );
and ( n11713 , n11318 , n11323 );
and ( n11714 , n11314 , n11323 );
or ( n11715 , n11712 , n11713 , n11714 );
and ( n11716 , n8640 , n4788 );
and ( n11717 , n9110 , n4611 );
nor ( n11718 , n11716 , n11717 );
xnor ( n11719 , n11718 , n4784 );
xor ( n11720 , n11715 , n11719 );
and ( n11721 , n5535 , n7356 );
and ( n11722 , n5818 , n6953 );
nor ( n11723 , n11721 , n11722 );
xnor ( n11724 , n11723 , n7352 );
and ( n11725 , n5247 , n7349 );
xor ( n11726 , n11724 , n11725 );
and ( n11727 , n11333 , n11334 );
xor ( n11728 , n11726 , n11727 );
and ( n11729 , n6168 , n6554 );
and ( n11730 , n6516 , n6205 );
nor ( n11731 , n11729 , n11730 );
xnor ( n11732 , n11731 , n6550 );
xor ( n11733 , n11728 , n11732 );
xor ( n11734 , n11720 , n11733 );
xor ( n11735 , n11711 , n11734 );
and ( n11736 , n10437 , n4319 );
and ( n11737 , n10857 , n4310 );
nor ( n11738 , n11736 , n11737 );
xnor ( n11739 , n11738 , n4315 );
and ( n11740 , n9583 , n4298 );
and ( n11741 , n9989 , n4287 );
nor ( n11742 , n11740 , n11741 );
xnor ( n11743 , n11742 , n4294 );
xor ( n11744 , n11739 , n11743 );
and ( n11745 , n11329 , n11335 );
and ( n11746 , n7752 , n5270 );
and ( n11747 , n8179 , n5021 );
nor ( n11748 , n11746 , n11747 );
xnor ( n11749 , n11748 , n5266 );
xor ( n11750 , n11745 , n11749 );
and ( n11751 , n6907 , n5850 );
and ( n11752 , n7324 , n5566 );
nor ( n11753 , n11751 , n11752 );
xnor ( n11754 , n11753 , n5846 );
xor ( n11755 , n11750 , n11754 );
xor ( n11756 , n11744 , n11755 );
xor ( n11757 , n11735 , n11756 );
xor ( n11758 , n11707 , n11757 );
and ( n11759 , n11225 , n11305 );
and ( n11760 , n11305 , n11347 );
and ( n11761 , n11225 , n11347 );
or ( n11762 , n11759 , n11760 , n11761 );
xor ( n11763 , n11758 , n11762 );
and ( n11764 , n11348 , n11352 );
and ( n11765 , n11353 , n11356 );
or ( n11766 , n11764 , n11765 );
xor ( n11767 , n11763 , n11766 );
buf ( n11768 , n11767 );
and ( n11769 , n11395 , n11411 );
and ( n11770 , n11411 , n11435 );
and ( n11771 , n11395 , n11435 );
or ( n11772 , n11769 , n11770 , n11771 );
and ( n11773 , n11401 , n11405 );
and ( n11774 , n11405 , n11410 );
and ( n11775 , n11401 , n11410 );
or ( n11776 , n11773 , n11774 , n11775 );
and ( n11777 , n11370 , n11374 );
and ( n11778 , n11374 , n11389 );
and ( n11779 , n11370 , n11389 );
or ( n11780 , n11777 , n11778 , n11779 );
xor ( n11781 , n11776 , n11780 );
and ( n11782 , n11398 , n4418 );
buf ( n11783 , n3968 );
buf ( n11784 , n11783 );
and ( n11785 , n11784 , n4415 );
nor ( n11786 , n11782 , n11785 );
xnor ( n11787 , n11786 , n4413 );
and ( n11788 , n10534 , n4433 );
and ( n11789 , n10940 , n4431 );
nor ( n11790 , n11788 , n11789 );
xnor ( n11791 , n11790 , n4441 );
xor ( n11792 , n11787 , n11791 );
and ( n11793 , n9629 , n4402 );
and ( n11794 , n10072 , n4391 );
nor ( n11795 , n11793 , n11794 );
xnor ( n11796 , n11795 , n4398 );
xor ( n11797 , n11792 , n11796 );
xor ( n11798 , n11781 , n11797 );
xor ( n11799 , n11772 , n11798 );
and ( n11800 , n11416 , n11420 );
and ( n11801 , n11420 , n11434 );
and ( n11802 , n11416 , n11434 );
or ( n11803 , n11800 , n11801 , n11802 );
and ( n11804 , n8728 , n4835 );
and ( n11805 , n9164 , n4648 );
nor ( n11806 , n11804 , n11805 );
xnor ( n11807 , n11806 , n4831 );
and ( n11808 , n7857 , n5323 );
and ( n11809 , n8303 , n5064 );
nor ( n11810 , n11808 , n11809 );
xnor ( n11811 , n11810 , n5319 );
xor ( n11812 , n11807 , n11811 );
and ( n11813 , n6235 , n6627 );
and ( n11814 , n6604 , n6272 );
nor ( n11815 , n11813 , n11814 );
xnor ( n11816 , n11815 , n6623 );
xor ( n11817 , n11812 , n11816 );
xor ( n11818 , n11803 , n11817 );
and ( n11819 , n11379 , n11383 );
and ( n11820 , n11383 , n11388 );
and ( n11821 , n11379 , n11388 );
or ( n11822 , n11819 , n11820 , n11821 );
and ( n11823 , n11427 , n11428 );
and ( n11824 , n11428 , n11433 );
and ( n11825 , n11427 , n11433 );
or ( n11826 , n11823 , n11824 , n11825 );
xor ( n11827 , n11822 , n11826 );
and ( n11828 , n5588 , n7444 );
and ( n11829 , n5893 , n7026 );
nor ( n11830 , n11828 , n11829 );
xnor ( n11831 , n11830 , n7440 );
and ( n11832 , n5300 , n7437 );
xor ( n11833 , n11831 , n11832 );
and ( n11834 , n11425 , n11426 );
xor ( n11835 , n11833 , n11834 );
and ( n11836 , n6995 , n5922 );
and ( n11837 , n7417 , n5616 );
nor ( n11838 , n11836 , n11837 );
xnor ( n11839 , n11838 , n5918 );
xor ( n11840 , n11835 , n11839 );
xor ( n11841 , n11827 , n11840 );
xor ( n11842 , n11818 , n11841 );
xor ( n11843 , n11799 , n11842 );
and ( n11844 , n11366 , n11390 );
and ( n11845 , n11390 , n11436 );
and ( n11846 , n11366 , n11436 );
or ( n11847 , n11844 , n11845 , n11846 );
xor ( n11848 , n11843 , n11847 );
and ( n11849 , n11362 , n11437 );
and ( n11850 , n11437 , n11442 );
and ( n11851 , n11362 , n11442 );
or ( n11852 , n11849 , n11850 , n11851 );
xor ( n11853 , n11848 , n11852 );
and ( n11854 , n11443 , n11444 );
xor ( n11855 , n11853 , n11854 );
buf ( n11856 , n11855 );
not ( n11857 , n454 );
and ( n11858 , n11857 , n11768 );
and ( n11859 , n11856 , n454 );
or ( n11860 , n11858 , n11859 );
buf ( n11861 , n11860 );
buf ( n11862 , n11861 );
and ( n11863 , n11862 , n4505 );
not ( n11864 , n11863 );
xor ( n11865 , n11638 , n11864 );
and ( n11866 , n11213 , n11214 );
and ( n11867 , n11214 , n11216 );
and ( n11868 , n11213 , n11216 );
or ( n11869 , n11866 , n11867 , n11868 );
xor ( n11870 , n11865 , n11869 );
xor ( n11871 , n11633 , n11870 );
and ( n11872 , n11217 , n11454 );
and ( n11873 , n11454 , n11459 );
and ( n11874 , n11217 , n11459 );
or ( n11875 , n11872 , n11873 , n11874 );
xor ( n11876 , n11871 , n11875 );
and ( n11877 , n11460 , n11464 );
and ( n11878 , n11464 , n11466 );
and ( n11879 , n11460 , n11466 );
or ( n11880 , n11877 , n11878 , n11879 );
xor ( n11881 , n11876 , n11880 );
and ( n11882 , n11468 , n11469 );
or ( n11883 , n11467 , n11882 );
xor ( n11884 , n11881 , n11883 );
buf ( n11885 , n11884 );
not ( n11886 , n4509 );
and ( n11887 , n11886 , n11632 );
and ( n11888 , n11885 , n4509 );
or ( n11889 , n11887 , n11888 );
and ( n11890 , n11498 , n11572 );
and ( n11891 , n11572 , n11617 );
and ( n11892 , n11498 , n11617 );
or ( n11893 , n11890 , n11891 , n11892 );
and ( n11894 , n11577 , n11591 );
and ( n11895 , n11591 , n11616 );
and ( n11896 , n11577 , n11616 );
or ( n11897 , n11894 , n11895 , n11896 );
and ( n11898 , n10706 , n4938 );
and ( n11899 , n11163 , n4711 );
nor ( n11900 , n11898 , n11899 );
xnor ( n11901 , n11900 , n4934 );
xor ( n11902 , n11897 , n11901 );
and ( n11903 , n11596 , n11600 );
and ( n11904 , n11600 , n11615 );
and ( n11905 , n11596 , n11615 );
or ( n11906 , n11903 , n11904 , n11905 );
and ( n11907 , n8968 , n6068 );
and ( n11908 , n9367 , n5730 );
nor ( n11909 , n11907 , n11908 );
xnor ( n11910 , n11909 , n6064 );
xor ( n11911 , n11906 , n11910 );
and ( n11912 , n8057 , n6711 );
and ( n11913 , n8462 , n6332 );
nor ( n11914 , n11912 , n11913 );
xnor ( n11915 , n11914 , n6707 );
xor ( n11916 , n11911 , n11915 );
xor ( n11917 , n11902 , n11916 );
xor ( n11918 , n11893 , n11917 );
and ( n11919 , n11483 , n11487 );
and ( n11920 , n11487 , n11492 );
and ( n11921 , n11483 , n11492 );
or ( n11922 , n11919 , n11920 , n11921 );
and ( n11923 , n11569 , n4524 );
and ( n11924 , n11511 , n11522 );
and ( n11925 , n11522 , n11551 );
and ( n11926 , n11511 , n11551 );
or ( n11927 , n11924 , n11925 , n11926 );
and ( n11928 , n11528 , n11532 );
and ( n11929 , n11532 , n11534 );
and ( n11930 , n11528 , n11534 );
or ( n11931 , n11928 , n11929 , n11930 );
and ( n11932 , n11540 , n11544 );
and ( n11933 , n11544 , n11549 );
and ( n11934 , n11540 , n11549 );
or ( n11935 , n11932 , n11933 , n11934 );
xor ( n11936 , n11931 , n11935 );
and ( n11937 , n9848 , n5405 );
not ( n11938 , n11937 );
xnor ( n11939 , n11938 , n5401 );
not ( n11940 , n11939 );
and ( n11941 , n8001 , n6761 );
and ( n11942 , n8409 , n6379 );
nor ( n11943 , n11941 , n11942 );
xnor ( n11944 , n11943 , n6757 );
xor ( n11945 , n11940 , n11944 );
and ( n11946 , n6353 , n8382 );
and ( n11947 , n6748 , n8042 );
nor ( n11948 , n11946 , n11947 );
xnor ( n11949 , n11948 , n8378 );
xor ( n11950 , n11945 , n11949 );
xor ( n11951 , n11936 , n11950 );
xor ( n11952 , n11927 , n11951 );
and ( n11953 , n11515 , n11516 );
and ( n11954 , n11516 , n11521 );
and ( n11955 , n11515 , n11521 );
or ( n11956 , n11953 , n11954 , n11955 );
and ( n11957 , n11527 , n11535 );
and ( n11958 , n11535 , n11550 );
and ( n11959 , n11527 , n11550 );
or ( n11960 , n11957 , n11958 , n11959 );
xor ( n11961 , n11956 , n11960 );
and ( n11962 , n8900 , n6008 );
and ( n11963 , n9297 , n5689 );
nor ( n11964 , n11962 , n11963 );
xnor ( n11965 , n11964 , n6004 );
and ( n11966 , n7092 , n7559 );
and ( n11967 , n7531 , n7107 );
nor ( n11968 , n11966 , n11967 );
xnor ( n11969 , n11968 , n7555 );
xor ( n11970 , n11965 , n11969 );
and ( n11971 , n5995 , n8375 );
xor ( n11972 , n11970 , n11971 );
xor ( n11973 , n11961 , n11972 );
xor ( n11974 , n11952 , n11973 );
and ( n11975 , n11507 , n11552 );
and ( n11976 , n11552 , n11557 );
and ( n11977 , n11507 , n11557 );
or ( n11978 , n11975 , n11976 , n11977 );
xor ( n11979 , n11974 , n11978 );
and ( n11980 , n11503 , n11558 );
and ( n11981 , n11558 , n11563 );
and ( n11982 , n11503 , n11563 );
or ( n11983 , n11980 , n11981 , n11982 );
xor ( n11984 , n11979 , n11983 );
and ( n11985 , n11564 , n11565 );
xor ( n11986 , n11984 , n11985 );
buf ( n11987 , n11986 );
buf ( n11988 , n11987 );
buf ( n11989 , n11988 );
and ( n11990 , n11989 , n4145 );
nor ( n11991 , n11923 , n11990 );
xnor ( n11992 , n11991 , n4521 );
xor ( n11993 , n11922 , n11992 );
and ( n11994 , n11581 , n11585 );
and ( n11995 , n11585 , n11590 );
and ( n11996 , n11581 , n11590 );
or ( n11997 , n11994 , n11995 , n11996 );
and ( n11998 , n9885 , n5441 );
and ( n11999 , n10287 , n5161 );
nor ( n12000 , n11998 , n11999 );
xnor ( n12001 , n12000 , n5437 );
xor ( n12002 , n11997 , n12001 );
and ( n12003 , n11605 , n11609 );
and ( n12004 , n11609 , n11614 );
and ( n12005 , n11605 , n11614 );
or ( n12006 , n12003 , n12004 , n12005 );
and ( n12007 , n7146 , n7630 );
and ( n12008 , n7587 , n7188 );
nor ( n12009 , n12007 , n12008 );
xnor ( n12010 , n12009 , n7626 );
xor ( n12011 , n12006 , n12010 );
and ( n12012 , n6391 , n8502 );
and ( n12013 , n6796 , n7970 );
nor ( n12014 , n12012 , n12013 );
xnor ( n12015 , n12014 , n8498 );
and ( n12016 , n5700 , n9407 );
and ( n12017 , n6037 , n8872 );
nor ( n12018 , n12016 , n12017 );
xnor ( n12019 , n12018 , n9403 );
xor ( n12020 , n12015 , n12019 );
and ( n12021 , n5140 , n10329 );
and ( n12022 , n5419 , n9791 );
nor ( n12023 , n12021 , n12022 );
not ( n12024 , n12023 );
xor ( n12025 , n12020 , n12024 );
xor ( n12026 , n12011 , n12025 );
xor ( n12027 , n12002 , n12026 );
xor ( n12028 , n11993 , n12027 );
xor ( n12029 , n11918 , n12028 );
and ( n12030 , n11479 , n11493 );
and ( n12031 , n11493 , n11618 );
and ( n12032 , n11479 , n11618 );
or ( n12033 , n12030 , n12031 , n12032 );
xor ( n12034 , n12029 , n12033 );
and ( n12035 , n11619 , n11623 );
and ( n12036 , n11623 , n11628 );
and ( n12037 , n11619 , n11628 );
or ( n12038 , n12035 , n12036 , n12037 );
xor ( n12039 , n12034 , n12038 );
and ( n12040 , n11629 , n11630 );
xor ( n12041 , n12039 , n12040 );
buf ( n12042 , n12041 );
buf ( n12043 , n11863 );
and ( n12044 , n11634 , n11635 );
and ( n12045 , n11635 , n11637 );
and ( n12046 , n11634 , n11637 );
or ( n12047 , n12044 , n12045 , n12046 );
and ( n12048 , n11862 , n4557 );
xor ( n12049 , n12047 , n12048 );
and ( n12050 , n11025 , n5089 );
and ( n12051 , n11452 , n4866 );
xor ( n12052 , n12050 , n12051 );
and ( n12053 , n11642 , n11706 );
and ( n12054 , n11706 , n11757 );
and ( n12055 , n11642 , n11757 );
or ( n12056 , n12053 , n12054 , n12055 );
and ( n12057 , n11646 , n11650 );
and ( n12058 , n11650 , n11705 );
and ( n12059 , n11646 , n11705 );
or ( n12060 , n12057 , n12058 , n12059 );
and ( n12061 , n11711 , n11734 );
and ( n12062 , n11734 , n11756 );
and ( n12063 , n11711 , n11756 );
or ( n12064 , n12061 , n12062 , n12063 );
xor ( n12065 , n12060 , n12064 );
and ( n12066 , n11739 , n11743 );
and ( n12067 , n11743 , n11755 );
and ( n12068 , n11739 , n11755 );
or ( n12069 , n12066 , n12067 , n12068 );
and ( n12070 , n11702 , n4235 );
and ( n12071 , n11682 , n11686 );
and ( n12072 , n11686 , n11688 );
and ( n12073 , n11682 , n11688 );
or ( n12074 , n12071 , n12072 , n12073 );
and ( n12075 , n11669 , n11680 );
and ( n12076 , n11680 , n11689 );
and ( n12077 , n11669 , n11689 );
or ( n12078 , n12075 , n12076 , n12077 );
xor ( n12079 , n12074 , n12078 );
and ( n12080 , n11670 , n11674 );
and ( n12081 , n11674 , n11679 );
and ( n12082 , n11670 , n11679 );
or ( n12083 , n12080 , n12081 , n12082 );
and ( n12084 , n7299 , n5773 );
not ( n12085 , n12084 );
xnor ( n12086 , n12085 , n5763 );
not ( n12087 , n12086 );
xor ( n12088 , n12083 , n12087 );
and ( n12089 , n6444 , n6496 );
and ( n12090 , n6853 , n6115 );
nor ( n12091 , n12089 , n12090 );
xnor ( n12092 , n12091 , n6453 );
and ( n12093 , n5791 , n7277 );
and ( n12094 , n6120 , n6864 );
nor ( n12095 , n12093 , n12094 );
xnor ( n12096 , n12095 , n7283 );
xor ( n12097 , n12092 , n12096 );
and ( n12098 , n5487 , n7274 );
xor ( n12099 , n12097 , n12098 );
xor ( n12100 , n12088 , n12099 );
xor ( n12101 , n12079 , n12100 );
and ( n12102 , n11660 , n11664 );
and ( n12103 , n11664 , n11690 );
and ( n12104 , n11660 , n11690 );
or ( n12105 , n12102 , n12103 , n12104 );
xor ( n12106 , n12101 , n12105 );
and ( n12107 , n11656 , n11691 );
and ( n12108 , n11691 , n11696 );
and ( n12109 , n11656 , n11696 );
or ( n12110 , n12107 , n12108 , n12109 );
xor ( n12111 , n12106 , n12110 );
and ( n12112 , n11697 , n11698 );
xor ( n12113 , n12111 , n12112 );
buf ( n12114 , n12113 );
buf ( n12115 , n12114 );
buf ( n12116 , n12115 );
and ( n12117 , n12116 , n4232 );
nor ( n12118 , n12070 , n12117 );
xnor ( n12119 , n12118 , n4230 );
and ( n12120 , n10857 , n4319 );
and ( n12121 , n11295 , n4310 );
nor ( n12122 , n12120 , n12121 );
xnor ( n12123 , n12122 , n4315 );
xor ( n12124 , n12119 , n12123 );
and ( n12125 , n9989 , n4298 );
and ( n12126 , n10437 , n4287 );
nor ( n12127 , n12125 , n12126 );
xnor ( n12128 , n12127 , n4294 );
xor ( n12129 , n12124 , n12128 );
xor ( n12130 , n12069 , n12129 );
and ( n12131 , n11715 , n11719 );
and ( n12132 , n11719 , n11733 );
and ( n12133 , n11715 , n11733 );
or ( n12134 , n12131 , n12132 , n12133 );
and ( n12135 , n11726 , n11727 );
and ( n12136 , n11727 , n11732 );
and ( n12137 , n11726 , n11732 );
or ( n12138 , n12135 , n12136 , n12137 );
and ( n12139 , n8179 , n5270 );
and ( n12140 , n8640 , n5021 );
nor ( n12141 , n12139 , n12140 );
xnor ( n12142 , n12141 , n5266 );
xor ( n12143 , n12138 , n12142 );
and ( n12144 , n7324 , n5850 );
and ( n12145 , n7752 , n5566 );
nor ( n12146 , n12144 , n12145 );
xnor ( n12147 , n12146 , n5846 );
xor ( n12148 , n12143 , n12147 );
xor ( n12149 , n12134 , n12148 );
and ( n12150 , n11745 , n11749 );
and ( n12151 , n11749 , n11754 );
and ( n12152 , n11745 , n11754 );
or ( n12153 , n12150 , n12151 , n12152 );
and ( n12154 , n9110 , n4788 );
and ( n12155 , n9583 , n4611 );
nor ( n12156 , n12154 , n12155 );
xnor ( n12157 , n12156 , n4784 );
xor ( n12158 , n12153 , n12157 );
and ( n12159 , n5818 , n7356 );
and ( n12160 , n6168 , n6953 );
nor ( n12161 , n12159 , n12160 );
xnor ( n12162 , n12161 , n7352 );
and ( n12163 , n5535 , n7349 );
xor ( n12164 , n12162 , n12163 );
and ( n12165 , n11724 , n11725 );
xor ( n12166 , n12164 , n12165 );
and ( n12167 , n6516 , n6554 );
and ( n12168 , n6907 , n6205 );
nor ( n12169 , n12167 , n12168 );
xnor ( n12170 , n12169 , n6550 );
xor ( n12171 , n12166 , n12170 );
xor ( n12172 , n12158 , n12171 );
xor ( n12173 , n12149 , n12172 );
xor ( n12174 , n12130 , n12173 );
xor ( n12175 , n12065 , n12174 );
xor ( n12176 , n12056 , n12175 );
and ( n12177 , n11758 , n11762 );
and ( n12178 , n11763 , n11766 );
or ( n12179 , n12177 , n12178 );
xor ( n12180 , n12176 , n12179 );
buf ( n12181 , n12180 );
and ( n12182 , n11776 , n11780 );
and ( n12183 , n11780 , n11797 );
and ( n12184 , n11776 , n11797 );
or ( n12185 , n12182 , n12183 , n12184 );
and ( n12186 , n11787 , n11791 );
and ( n12187 , n11791 , n11796 );
and ( n12188 , n11787 , n11796 );
or ( n12189 , n12186 , n12187 , n12188 );
and ( n12190 , n11822 , n11826 );
and ( n12191 , n11826 , n11840 );
and ( n12192 , n11822 , n11840 );
or ( n12193 , n12190 , n12191 , n12192 );
xor ( n12194 , n12189 , n12193 );
and ( n12195 , n11833 , n11834 );
and ( n12196 , n11834 , n11839 );
and ( n12197 , n11833 , n11839 );
or ( n12198 , n12195 , n12196 , n12197 );
and ( n12199 , n8303 , n5323 );
and ( n12200 , n8728 , n5064 );
nor ( n12201 , n12199 , n12200 );
xnor ( n12202 , n12201 , n5319 );
xor ( n12203 , n12198 , n12202 );
and ( n12204 , n7417 , n5922 );
and ( n12205 , n7857 , n5616 );
nor ( n12206 , n12204 , n12205 );
xnor ( n12207 , n12206 , n5918 );
xor ( n12208 , n12203 , n12207 );
xor ( n12209 , n12194 , n12208 );
xor ( n12210 , n12185 , n12209 );
and ( n12211 , n11803 , n11817 );
and ( n12212 , n11817 , n11841 );
and ( n12213 , n11803 , n11841 );
or ( n12214 , n12211 , n12212 , n12213 );
and ( n12215 , n11784 , n4418 );
buf ( n12216 , n4030 );
buf ( n12217 , n12216 );
and ( n12218 , n12217 , n4415 );
nor ( n12219 , n12215 , n12218 );
xnor ( n12220 , n12219 , n4413 );
and ( n12221 , n10940 , n4433 );
and ( n12222 , n11398 , n4431 );
nor ( n12223 , n12221 , n12222 );
xnor ( n12224 , n12223 , n4441 );
xor ( n12225 , n12220 , n12224 );
and ( n12226 , n9164 , n4835 );
and ( n12227 , n9629 , n4648 );
nor ( n12228 , n12226 , n12227 );
xnor ( n12229 , n12228 , n4831 );
xor ( n12230 , n12225 , n12229 );
xor ( n12231 , n12214 , n12230 );
and ( n12232 , n11807 , n11811 );
and ( n12233 , n11811 , n11816 );
and ( n12234 , n11807 , n11816 );
or ( n12235 , n12232 , n12233 , n12234 );
and ( n12236 , n10072 , n4402 );
and ( n12237 , n10534 , n4391 );
nor ( n12238 , n12236 , n12237 );
xnor ( n12239 , n12238 , n4398 );
xor ( n12240 , n12235 , n12239 );
and ( n12241 , n6604 , n6627 );
and ( n12242 , n6995 , n6272 );
nor ( n12243 , n12241 , n12242 );
xnor ( n12244 , n12243 , n6623 );
and ( n12245 , n5588 , n7437 );
xor ( n12246 , n12244 , n12245 );
and ( n12247 , n11831 , n11832 );
xor ( n12248 , n12246 , n12247 );
and ( n12249 , n5893 , n7444 );
and ( n12250 , n6235 , n7026 );
nor ( n12251 , n12249 , n12250 );
xnor ( n12252 , n12251 , n7440 );
xor ( n12253 , n12248 , n12252 );
xor ( n12254 , n12240 , n12253 );
xor ( n12255 , n12231 , n12254 );
xor ( n12256 , n12210 , n12255 );
and ( n12257 , n11772 , n11798 );
and ( n12258 , n11798 , n11842 );
and ( n12259 , n11772 , n11842 );
or ( n12260 , n12257 , n12258 , n12259 );
xor ( n12261 , n12256 , n12260 );
and ( n12262 , n11843 , n11847 );
and ( n12263 , n11847 , n11852 );
and ( n12264 , n11843 , n11852 );
or ( n12265 , n12262 , n12263 , n12264 );
xor ( n12266 , n12261 , n12265 );
and ( n12267 , n11853 , n11854 );
xor ( n12268 , n12266 , n12267 );
buf ( n12269 , n12268 );
not ( n12270 , n454 );
and ( n12271 , n12270 , n12181 );
and ( n12272 , n12269 , n454 );
or ( n12273 , n12271 , n12272 );
buf ( n12274 , n12273 );
buf ( n12275 , n12274 );
and ( n12276 , n12275 , n4505 );
xor ( n12277 , n12052 , n12276 );
xor ( n12278 , n12049 , n12277 );
xor ( n12279 , n12043 , n12278 );
and ( n12280 , n11638 , n11864 );
and ( n12281 , n11864 , n11869 );
and ( n12282 , n11638 , n11869 );
or ( n12283 , n12280 , n12281 , n12282 );
xor ( n12284 , n12279 , n12283 );
and ( n12285 , n11633 , n11870 );
and ( n12286 , n11870 , n11875 );
and ( n12287 , n11633 , n11875 );
or ( n12288 , n12285 , n12286 , n12287 );
xnor ( n12289 , n12284 , n12288 );
and ( n12290 , n11876 , n11880 );
and ( n12291 , n11881 , n11883 );
or ( n12292 , n12290 , n12291 );
xor ( n12293 , n12289 , n12292 );
buf ( n12294 , n12293 );
not ( n12295 , n4509 );
and ( n12296 , n12295 , n12042 );
and ( n12297 , n12294 , n4509 );
or ( n12298 , n12296 , n12297 );
and ( n12299 , n11922 , n11992 );
and ( n12300 , n11992 , n12027 );
and ( n12301 , n11922 , n12027 );
or ( n12302 , n12299 , n12300 , n12301 );
and ( n12303 , n11906 , n11910 );
and ( n12304 , n11910 , n11915 );
and ( n12305 , n11906 , n11915 );
or ( n12306 , n12303 , n12304 , n12305 );
and ( n12307 , n11997 , n12001 );
and ( n12308 , n12001 , n12026 );
and ( n12309 , n11997 , n12026 );
or ( n12310 , n12307 , n12308 , n12309 );
xor ( n12311 , n12306 , n12310 );
and ( n12312 , n12006 , n12010 );
and ( n12313 , n12010 , n12025 );
and ( n12314 , n12006 , n12025 );
or ( n12315 , n12312 , n12313 , n12314 );
and ( n12316 , n9367 , n6068 );
and ( n12317 , n9885 , n5730 );
nor ( n12318 , n12316 , n12317 );
xnor ( n12319 , n12318 , n6064 );
xor ( n12320 , n12315 , n12319 );
and ( n12321 , n8462 , n6711 );
and ( n12322 , n8968 , n6332 );
nor ( n12323 , n12321 , n12322 );
xnor ( n12324 , n12323 , n6707 );
xor ( n12325 , n12320 , n12324 );
xor ( n12326 , n12311 , n12325 );
xor ( n12327 , n12302 , n12326 );
and ( n12328 , n11897 , n11901 );
and ( n12329 , n11901 , n11916 );
and ( n12330 , n11897 , n11916 );
or ( n12331 , n12328 , n12329 , n12330 );
and ( n12332 , n11989 , n4524 );
and ( n12333 , n11931 , n11935 );
and ( n12334 , n11935 , n11950 );
and ( n12335 , n11931 , n11950 );
or ( n12336 , n12333 , n12334 , n12335 );
and ( n12337 , n11956 , n11960 );
and ( n12338 , n11960 , n11972 );
and ( n12339 , n11956 , n11972 );
or ( n12340 , n12337 , n12338 , n12339 );
xor ( n12341 , n12336 , n12340 );
and ( n12342 , n11940 , n11944 );
and ( n12343 , n11944 , n11949 );
and ( n12344 , n11940 , n11949 );
or ( n12345 , n12342 , n12343 , n12344 );
and ( n12346 , n8409 , n6761 );
and ( n12347 , n8900 , n6379 );
nor ( n12348 , n12346 , n12347 );
xnor ( n12349 , n12348 , n6757 );
and ( n12350 , n7531 , n7559 );
and ( n12351 , n8001 , n7107 );
nor ( n12352 , n12350 , n12351 );
xnor ( n12353 , n12352 , n7555 );
xor ( n12354 , n12349 , n12353 );
and ( n12355 , n6748 , n8382 );
and ( n12356 , n7092 , n8042 );
nor ( n12357 , n12355 , n12356 );
xnor ( n12358 , n12357 , n8378 );
xor ( n12359 , n12354 , n12358 );
xor ( n12360 , n12345 , n12359 );
and ( n12361 , n11965 , n11969 );
and ( n12362 , n11969 , n11971 );
and ( n12363 , n11965 , n11971 );
or ( n12364 , n12361 , n12362 , n12363 );
buf ( n12365 , n11939 );
xor ( n12366 , n12364 , n12365 );
not ( n12367 , n5401 );
and ( n12368 , n9297 , n6008 );
and ( n12369 , n9848 , n5689 );
nor ( n12370 , n12368 , n12369 );
xnor ( n12371 , n12370 , n6004 );
xor ( n12372 , n12367 , n12371 );
and ( n12373 , n6353 , n8375 );
xor ( n12374 , n12372 , n12373 );
xor ( n12375 , n12366 , n12374 );
xor ( n12376 , n12360 , n12375 );
xor ( n12377 , n12341 , n12376 );
and ( n12378 , n11927 , n11951 );
and ( n12379 , n11951 , n11973 );
and ( n12380 , n11927 , n11973 );
or ( n12381 , n12378 , n12379 , n12380 );
xor ( n12382 , n12377 , n12381 );
and ( n12383 , n11974 , n11978 );
and ( n12384 , n11978 , n11983 );
and ( n12385 , n11974 , n11983 );
or ( n12386 , n12383 , n12384 , n12385 );
xor ( n12387 , n12382 , n12386 );
and ( n12388 , n11984 , n11985 );
xor ( n12389 , n12387 , n12388 );
buf ( n12390 , n12389 );
buf ( n12391 , n12390 );
buf ( n12392 , n12391 );
and ( n12393 , n12392 , n4145 );
nor ( n12394 , n12332 , n12393 );
xnor ( n12395 , n12394 , n4521 );
xor ( n12396 , n12331 , n12395 );
and ( n12397 , n11163 , n4938 );
and ( n12398 , n11569 , n4711 );
nor ( n12399 , n12397 , n12398 );
xnor ( n12400 , n12399 , n4934 );
and ( n12401 , n10287 , n5441 );
and ( n12402 , n10706 , n5161 );
nor ( n12403 , n12401 , n12402 );
xnor ( n12404 , n12403 , n5437 );
xor ( n12405 , n12400 , n12404 );
and ( n12406 , n12015 , n12019 );
and ( n12407 , n12019 , n12024 );
and ( n12408 , n12015 , n12024 );
or ( n12409 , n12406 , n12407 , n12408 );
and ( n12410 , n7587 , n7630 );
and ( n12411 , n8057 , n7188 );
nor ( n12412 , n12410 , n12411 );
xnor ( n12413 , n12412 , n7626 );
xor ( n12414 , n12409 , n12413 );
and ( n12415 , n6796 , n8502 );
and ( n12416 , n7146 , n7970 );
nor ( n12417 , n12415 , n12416 );
xnor ( n12418 , n12417 , n8498 );
and ( n12419 , n6037 , n9407 );
and ( n12420 , n6391 , n8872 );
nor ( n12421 , n12419 , n12420 );
xnor ( n12422 , n12421 , n9403 );
xor ( n12423 , n12418 , n12422 );
and ( n12424 , n5419 , n10329 );
and ( n12425 , n5700 , n9791 );
nor ( n12426 , n12424 , n12425 );
not ( n12427 , n12426 );
xor ( n12428 , n12423 , n12427 );
xor ( n12429 , n12414 , n12428 );
xor ( n12430 , n12405 , n12429 );
xor ( n12431 , n12396 , n12430 );
xor ( n12432 , n12327 , n12431 );
and ( n12433 , n11893 , n11917 );
and ( n12434 , n11917 , n12028 );
and ( n12435 , n11893 , n12028 );
or ( n12436 , n12433 , n12434 , n12435 );
xor ( n12437 , n12432 , n12436 );
and ( n12438 , n12029 , n12033 );
and ( n12439 , n12033 , n12038 );
and ( n12440 , n12029 , n12038 );
or ( n12441 , n12438 , n12439 , n12440 );
xor ( n12442 , n12437 , n12441 );
and ( n12443 , n12039 , n12040 );
xor ( n12444 , n12442 , n12443 );
buf ( n12445 , n12444 );
and ( n12446 , n12050 , n12051 );
and ( n12447 , n12051 , n12276 );
and ( n12448 , n12050 , n12276 );
or ( n12449 , n12446 , n12447 , n12448 );
and ( n12450 , n12069 , n12129 );
and ( n12451 , n12129 , n12173 );
and ( n12452 , n12069 , n12173 );
or ( n12453 , n12450 , n12451 , n12452 );
and ( n12454 , n12119 , n12123 );
and ( n12455 , n12123 , n12128 );
and ( n12456 , n12119 , n12128 );
or ( n12457 , n12454 , n12455 , n12456 );
and ( n12458 , n12153 , n12157 );
and ( n12459 , n12157 , n12171 );
and ( n12460 , n12153 , n12171 );
or ( n12461 , n12458 , n12459 , n12460 );
xor ( n12462 , n12457 , n12461 );
and ( n12463 , n12164 , n12165 );
and ( n12464 , n12165 , n12170 );
and ( n12465 , n12164 , n12170 );
or ( n12466 , n12463 , n12464 , n12465 );
and ( n12467 , n8640 , n5270 );
and ( n12468 , n9110 , n5021 );
nor ( n12469 , n12467 , n12468 );
xnor ( n12470 , n12469 , n5266 );
xor ( n12471 , n12466 , n12470 );
and ( n12472 , n7752 , n5850 );
and ( n12473 , n8179 , n5566 );
nor ( n12474 , n12472 , n12473 );
xnor ( n12475 , n12474 , n5846 );
xor ( n12476 , n12471 , n12475 );
xor ( n12477 , n12462 , n12476 );
xor ( n12478 , n12453 , n12477 );
and ( n12479 , n12134 , n12148 );
and ( n12480 , n12148 , n12172 );
and ( n12481 , n12134 , n12172 );
or ( n12482 , n12479 , n12480 , n12481 );
and ( n12483 , n12138 , n12142 );
and ( n12484 , n12142 , n12147 );
and ( n12485 , n12138 , n12147 );
or ( n12486 , n12483 , n12484 , n12485 );
and ( n12487 , n12116 , n4235 );
and ( n12488 , n12083 , n12087 );
and ( n12489 , n12087 , n12099 );
and ( n12490 , n12083 , n12099 );
or ( n12491 , n12488 , n12489 , n12490 );
not ( n12492 , n5763 );
and ( n12493 , n6853 , n6496 );
and ( n12494 , n7299 , n6115 );
nor ( n12495 , n12493 , n12494 );
xnor ( n12496 , n12495 , n6453 );
xor ( n12497 , n12492 , n12496 );
and ( n12498 , n5791 , n7274 );
xor ( n12499 , n12497 , n12498 );
xor ( n12500 , n12491 , n12499 );
and ( n12501 , n12092 , n12096 );
and ( n12502 , n12096 , n12098 );
and ( n12503 , n12092 , n12098 );
or ( n12504 , n12501 , n12502 , n12503 );
buf ( n12505 , n12086 );
xor ( n12506 , n12504 , n12505 );
and ( n12507 , n6120 , n7277 );
and ( n12508 , n6444 , n6864 );
nor ( n12509 , n12507 , n12508 );
xnor ( n12510 , n12509 , n7283 );
xor ( n12511 , n12506 , n12510 );
xor ( n12512 , n12500 , n12511 );
and ( n12513 , n12074 , n12078 );
and ( n12514 , n12078 , n12100 );
and ( n12515 , n12074 , n12100 );
or ( n12516 , n12513 , n12514 , n12515 );
xor ( n12517 , n12512 , n12516 );
and ( n12518 , n12101 , n12105 );
and ( n12519 , n12105 , n12110 );
and ( n12520 , n12101 , n12110 );
or ( n12521 , n12518 , n12519 , n12520 );
xor ( n12522 , n12517 , n12521 );
and ( n12523 , n12111 , n12112 );
xor ( n12524 , n12522 , n12523 );
buf ( n12525 , n12524 );
buf ( n12526 , n12525 );
buf ( n12527 , n12526 );
and ( n12528 , n12527 , n4232 );
nor ( n12529 , n12487 , n12528 );
xnor ( n12530 , n12529 , n4230 );
xor ( n12531 , n12486 , n12530 );
and ( n12532 , n11295 , n4319 );
and ( n12533 , n11702 , n4310 );
nor ( n12534 , n12532 , n12533 );
xnor ( n12535 , n12534 , n4315 );
xor ( n12536 , n12531 , n12535 );
xor ( n12537 , n12482 , n12536 );
and ( n12538 , n10437 , n4298 );
and ( n12539 , n10857 , n4287 );
nor ( n12540 , n12538 , n12539 );
xnor ( n12541 , n12540 , n4294 );
and ( n12542 , n9583 , n4788 );
and ( n12543 , n9989 , n4611 );
nor ( n12544 , n12542 , n12543 );
xnor ( n12545 , n12544 , n4784 );
xor ( n12546 , n12541 , n12545 );
and ( n12547 , n6168 , n7356 );
and ( n12548 , n6516 , n6953 );
nor ( n12549 , n12547 , n12548 );
xnor ( n12550 , n12549 , n7352 );
and ( n12551 , n5818 , n7349 );
xor ( n12552 , n12550 , n12551 );
and ( n12553 , n12162 , n12163 );
xor ( n12554 , n12552 , n12553 );
and ( n12555 , n6907 , n6554 );
and ( n12556 , n7324 , n6205 );
nor ( n12557 , n12555 , n12556 );
xnor ( n12558 , n12557 , n6550 );
xor ( n12559 , n12554 , n12558 );
xor ( n12560 , n12546 , n12559 );
xor ( n12561 , n12537 , n12560 );
xor ( n12562 , n12478 , n12561 );
and ( n12563 , n12060 , n12064 );
and ( n12564 , n12064 , n12174 );
and ( n12565 , n12060 , n12174 );
or ( n12566 , n12563 , n12564 , n12565 );
xor ( n12567 , n12562 , n12566 );
and ( n12568 , n12056 , n12175 );
and ( n12569 , n12176 , n12179 );
or ( n12570 , n12568 , n12569 );
xor ( n12571 , n12567 , n12570 );
buf ( n12572 , n12571 );
and ( n12573 , n12214 , n12230 );
and ( n12574 , n12230 , n12254 );
and ( n12575 , n12214 , n12254 );
or ( n12576 , n12573 , n12574 , n12575 );
and ( n12577 , n12220 , n12224 );
and ( n12578 , n12224 , n12229 );
and ( n12579 , n12220 , n12229 );
or ( n12580 , n12577 , n12578 , n12579 );
and ( n12581 , n12235 , n12239 );
and ( n12582 , n12239 , n12253 );
and ( n12583 , n12235 , n12253 );
or ( n12584 , n12581 , n12582 , n12583 );
xor ( n12585 , n12580 , n12584 );
and ( n12586 , n9629 , n4835 );
and ( n12587 , n10072 , n4648 );
nor ( n12588 , n12586 , n12587 );
xnor ( n12589 , n12588 , n4831 );
and ( n12590 , n8728 , n5323 );
and ( n12591 , n9164 , n5064 );
nor ( n12592 , n12590 , n12591 );
xnor ( n12593 , n12592 , n5319 );
xor ( n12594 , n12589 , n12593 );
and ( n12595 , n7857 , n5922 );
and ( n12596 , n8303 , n5616 );
nor ( n12597 , n12595 , n12596 );
xnor ( n12598 , n12597 , n5918 );
xor ( n12599 , n12594 , n12598 );
xor ( n12600 , n12585 , n12599 );
xor ( n12601 , n12576 , n12600 );
and ( n12602 , n12189 , n12193 );
and ( n12603 , n12193 , n12208 );
and ( n12604 , n12189 , n12208 );
or ( n12605 , n12602 , n12603 , n12604 );
and ( n12606 , n12246 , n12247 );
and ( n12607 , n12247 , n12252 );
and ( n12608 , n12246 , n12252 );
or ( n12609 , n12606 , n12607 , n12608 );
and ( n12610 , n12217 , n4418 );
buf ( n12611 , n4084 );
buf ( n12612 , n12611 );
and ( n12613 , n12612 , n4415 );
nor ( n12614 , n12610 , n12613 );
xnor ( n12615 , n12614 , n4413 );
xor ( n12616 , n12609 , n12615 );
and ( n12617 , n11398 , n4433 );
and ( n12618 , n11784 , n4431 );
nor ( n12619 , n12617 , n12618 );
xnor ( n12620 , n12619 , n4441 );
xor ( n12621 , n12616 , n12620 );
xor ( n12622 , n12605 , n12621 );
and ( n12623 , n12198 , n12202 );
and ( n12624 , n12202 , n12207 );
and ( n12625 , n12198 , n12207 );
or ( n12626 , n12623 , n12624 , n12625 );
and ( n12627 , n10534 , n4402 );
and ( n12628 , n10940 , n4391 );
nor ( n12629 , n12627 , n12628 );
xnor ( n12630 , n12629 , n4398 );
xor ( n12631 , n12626 , n12630 );
and ( n12632 , n6995 , n6627 );
and ( n12633 , n7417 , n6272 );
nor ( n12634 , n12632 , n12633 );
xnor ( n12635 , n12634 , n6623 );
and ( n12636 , n5893 , n7437 );
xor ( n12637 , n12635 , n12636 );
and ( n12638 , n12244 , n12245 );
xor ( n12639 , n12637 , n12638 );
and ( n12640 , n6235 , n7444 );
and ( n12641 , n6604 , n7026 );
nor ( n12642 , n12640 , n12641 );
xnor ( n12643 , n12642 , n7440 );
xor ( n12644 , n12639 , n12643 );
xor ( n12645 , n12631 , n12644 );
xor ( n12646 , n12622 , n12645 );
xor ( n12647 , n12601 , n12646 );
and ( n12648 , n12185 , n12209 );
and ( n12649 , n12209 , n12255 );
and ( n12650 , n12185 , n12255 );
or ( n12651 , n12648 , n12649 , n12650 );
xor ( n12652 , n12647 , n12651 );
and ( n12653 , n12256 , n12260 );
and ( n12654 , n12260 , n12265 );
and ( n12655 , n12256 , n12265 );
or ( n12656 , n12653 , n12654 , n12655 );
xor ( n12657 , n12652 , n12656 );
and ( n12658 , n12266 , n12267 );
xor ( n12659 , n12657 , n12658 );
buf ( n12660 , n12659 );
not ( n12661 , n454 );
and ( n12662 , n12661 , n12572 );
and ( n12663 , n12660 , n454 );
or ( n12664 , n12662 , n12663 );
buf ( n12665 , n12664 );
buf ( n12666 , n12665 );
and ( n12667 , n12666 , n4505 );
xor ( n12668 , n12449 , n12667 );
and ( n12669 , n11452 , n5089 );
and ( n12670 , n11862 , n4866 );
xor ( n12671 , n12669 , n12670 );
and ( n12672 , n12275 , n4557 );
xor ( n12673 , n12671 , n12672 );
xor ( n12674 , n12668 , n12673 );
and ( n12675 , n12047 , n12048 );
and ( n12676 , n12048 , n12277 );
and ( n12677 , n12047 , n12277 );
or ( n12678 , n12675 , n12676 , n12677 );
xor ( n12679 , n12674 , n12678 );
and ( n12680 , n12043 , n12278 );
and ( n12681 , n12278 , n12283 );
and ( n12682 , n12043 , n12283 );
or ( n12683 , n12680 , n12681 , n12682 );
xor ( n12684 , n12679 , n12683 );
or ( n12685 , n12284 , n12288 );
xnor ( n12686 , n12684 , n12685 );
and ( n12687 , n12289 , n12292 );
xor ( n12688 , n12686 , n12687 );
buf ( n12689 , n12688 );
not ( n12690 , n4509 );
and ( n12691 , n12690 , n12445 );
and ( n12692 , n12689 , n4509 );
or ( n12693 , n12691 , n12692 );
and ( n12694 , n12331 , n12395 );
and ( n12695 , n12395 , n12430 );
and ( n12696 , n12331 , n12430 );
or ( n12697 , n12694 , n12695 , n12696 );
and ( n12698 , n12392 , n4524 );
and ( n12699 , n12345 , n12359 );
and ( n12700 , n12359 , n12375 );
and ( n12701 , n12345 , n12375 );
or ( n12702 , n12699 , n12700 , n12701 );
and ( n12703 , n12349 , n12353 );
and ( n12704 , n12353 , n12358 );
and ( n12705 , n12349 , n12358 );
or ( n12706 , n12703 , n12704 , n12705 );
and ( n12707 , n9848 , n6008 );
not ( n12708 , n12707 );
xnor ( n12709 , n12708 , n6004 );
not ( n12710 , n12709 );
xor ( n12711 , n12706 , n12710 );
and ( n12712 , n8001 , n7559 );
and ( n12713 , n8409 , n7107 );
nor ( n12714 , n12712 , n12713 );
xnor ( n12715 , n12714 , n7555 );
xor ( n12716 , n12711 , n12715 );
xor ( n12717 , n12702 , n12716 );
and ( n12718 , n12367 , n12371 );
and ( n12719 , n12371 , n12373 );
and ( n12720 , n12367 , n12373 );
or ( n12721 , n12718 , n12719 , n12720 );
and ( n12722 , n12364 , n12365 );
and ( n12723 , n12365 , n12374 );
and ( n12724 , n12364 , n12374 );
or ( n12725 , n12722 , n12723 , n12724 );
xor ( n12726 , n12721 , n12725 );
and ( n12727 , n8900 , n6761 );
and ( n12728 , n9297 , n6379 );
nor ( n12729 , n12727 , n12728 );
xnor ( n12730 , n12729 , n6757 );
and ( n12731 , n7092 , n8382 );
and ( n12732 , n7531 , n8042 );
nor ( n12733 , n12731 , n12732 );
xnor ( n12734 , n12733 , n8378 );
xor ( n12735 , n12730 , n12734 );
and ( n12736 , n6748 , n8375 );
xor ( n12737 , n12735 , n12736 );
xor ( n12738 , n12726 , n12737 );
xor ( n12739 , n12717 , n12738 );
and ( n12740 , n12336 , n12340 );
and ( n12741 , n12340 , n12376 );
and ( n12742 , n12336 , n12376 );
or ( n12743 , n12740 , n12741 , n12742 );
xor ( n12744 , n12739 , n12743 );
and ( n12745 , n12377 , n12381 );
and ( n12746 , n12381 , n12386 );
and ( n12747 , n12377 , n12386 );
or ( n12748 , n12745 , n12746 , n12747 );
xor ( n12749 , n12744 , n12748 );
and ( n12750 , n12387 , n12388 );
xor ( n12751 , n12749 , n12750 );
buf ( n12752 , n12751 );
buf ( n12753 , n12752 );
buf ( n12754 , n12753 );
and ( n12755 , n12754 , n4145 );
nor ( n12756 , n12698 , n12755 );
xnor ( n12757 , n12756 , n4521 );
and ( n12758 , n11569 , n4938 );
and ( n12759 , n11989 , n4711 );
nor ( n12760 , n12758 , n12759 );
xnor ( n12761 , n12760 , n4934 );
xor ( n12762 , n12757 , n12761 );
and ( n12763 , n12409 , n12413 );
and ( n12764 , n12413 , n12428 );
and ( n12765 , n12409 , n12428 );
or ( n12766 , n12763 , n12764 , n12765 );
and ( n12767 , n9885 , n6068 );
and ( n12768 , n10287 , n5730 );
nor ( n12769 , n12767 , n12768 );
xnor ( n12770 , n12769 , n6064 );
xor ( n12771 , n12766 , n12770 );
and ( n12772 , n8968 , n6711 );
and ( n12773 , n9367 , n6332 );
nor ( n12774 , n12772 , n12773 );
xnor ( n12775 , n12774 , n6707 );
xor ( n12776 , n12771 , n12775 );
xor ( n12777 , n12762 , n12776 );
xor ( n12778 , n12697 , n12777 );
and ( n12779 , n12306 , n12310 );
and ( n12780 , n12310 , n12325 );
and ( n12781 , n12306 , n12325 );
or ( n12782 , n12779 , n12780 , n12781 );
and ( n12783 , n12400 , n12404 );
and ( n12784 , n12404 , n12429 );
and ( n12785 , n12400 , n12429 );
or ( n12786 , n12783 , n12784 , n12785 );
xor ( n12787 , n12782 , n12786 );
and ( n12788 , n12315 , n12319 );
and ( n12789 , n12319 , n12324 );
and ( n12790 , n12315 , n12324 );
or ( n12791 , n12788 , n12789 , n12790 );
and ( n12792 , n10706 , n5441 );
and ( n12793 , n11163 , n5161 );
nor ( n12794 , n12792 , n12793 );
xnor ( n12795 , n12794 , n5437 );
xor ( n12796 , n12791 , n12795 );
and ( n12797 , n12418 , n12422 );
and ( n12798 , n12422 , n12427 );
and ( n12799 , n12418 , n12427 );
or ( n12800 , n12797 , n12798 , n12799 );
and ( n12801 , n8057 , n7630 );
and ( n12802 , n8462 , n7188 );
nor ( n12803 , n12801 , n12802 );
xnor ( n12804 , n12803 , n7626 );
xor ( n12805 , n12800 , n12804 );
and ( n12806 , n7146 , n8502 );
and ( n12807 , n7587 , n7970 );
nor ( n12808 , n12806 , n12807 );
xnor ( n12809 , n12808 , n8498 );
and ( n12810 , n6391 , n9407 );
and ( n12811 , n6796 , n8872 );
nor ( n12812 , n12810 , n12811 );
xnor ( n12813 , n12812 , n9403 );
xor ( n12814 , n12809 , n12813 );
and ( n12815 , n5700 , n10329 );
and ( n12816 , n6037 , n9791 );
nor ( n12817 , n12815 , n12816 );
not ( n12818 , n12817 );
xor ( n12819 , n12814 , n12818 );
xor ( n12820 , n12805 , n12819 );
xor ( n12821 , n12796 , n12820 );
xor ( n12822 , n12787 , n12821 );
xor ( n12823 , n12778 , n12822 );
and ( n12824 , n12302 , n12326 );
and ( n12825 , n12326 , n12431 );
and ( n12826 , n12302 , n12431 );
or ( n12827 , n12824 , n12825 , n12826 );
xor ( n12828 , n12823 , n12827 );
and ( n12829 , n12432 , n12436 );
and ( n12830 , n12436 , n12441 );
and ( n12831 , n12432 , n12441 );
or ( n12832 , n12829 , n12830 , n12831 );
xor ( n12833 , n12828 , n12832 );
and ( n12834 , n12442 , n12443 );
xor ( n12835 , n12833 , n12834 );
buf ( n12836 , n12835 );
and ( n12837 , n12669 , n12670 );
and ( n12838 , n12670 , n12672 );
and ( n12839 , n12669 , n12672 );
or ( n12840 , n12837 , n12838 , n12839 );
and ( n12841 , n12666 , n4557 );
xor ( n12842 , n12840 , n12841 );
and ( n12843 , n11862 , n5089 );
and ( n12844 , n12275 , n4866 );
xor ( n12845 , n12843 , n12844 );
and ( n12846 , n12457 , n12461 );
and ( n12847 , n12461 , n12476 );
and ( n12848 , n12457 , n12476 );
or ( n12849 , n12846 , n12847 , n12848 );
and ( n12850 , n12482 , n12536 );
and ( n12851 , n12536 , n12560 );
and ( n12852 , n12482 , n12560 );
or ( n12853 , n12850 , n12851 , n12852 );
xor ( n12854 , n12849 , n12853 );
and ( n12855 , n12466 , n12470 );
and ( n12856 , n12470 , n12475 );
and ( n12857 , n12466 , n12475 );
or ( n12858 , n12855 , n12856 , n12857 );
and ( n12859 , n12527 , n4235 );
and ( n12860 , n12492 , n12496 );
and ( n12861 , n12496 , n12498 );
and ( n12862 , n12492 , n12498 );
or ( n12863 , n12860 , n12861 , n12862 );
and ( n12864 , n12504 , n12505 );
and ( n12865 , n12505 , n12510 );
and ( n12866 , n12504 , n12510 );
or ( n12867 , n12864 , n12865 , n12866 );
xor ( n12868 , n12863 , n12867 );
and ( n12869 , n7299 , n6496 );
not ( n12870 , n12869 );
xnor ( n12871 , n12870 , n6453 );
not ( n12872 , n12871 );
and ( n12873 , n6444 , n7277 );
and ( n12874 , n6853 , n6864 );
nor ( n12875 , n12873 , n12874 );
xnor ( n12876 , n12875 , n7283 );
xor ( n12877 , n12872 , n12876 );
and ( n12878 , n6120 , n7274 );
xor ( n12879 , n12877 , n12878 );
xor ( n12880 , n12868 , n12879 );
and ( n12881 , n12491 , n12499 );
and ( n12882 , n12499 , n12511 );
and ( n12883 , n12491 , n12511 );
or ( n12884 , n12881 , n12882 , n12883 );
xor ( n12885 , n12880 , n12884 );
and ( n12886 , n12512 , n12516 );
and ( n12887 , n12516 , n12521 );
and ( n12888 , n12512 , n12521 );
or ( n12889 , n12886 , n12887 , n12888 );
xor ( n12890 , n12885 , n12889 );
and ( n12891 , n12522 , n12523 );
xor ( n12892 , n12890 , n12891 );
buf ( n12893 , n12892 );
buf ( n12894 , n12893 );
buf ( n12895 , n12894 );
and ( n12896 , n12895 , n4232 );
nor ( n12897 , n12859 , n12896 );
xnor ( n12898 , n12897 , n4230 );
xor ( n12899 , n12858 , n12898 );
and ( n12900 , n11702 , n4319 );
and ( n12901 , n12116 , n4310 );
nor ( n12902 , n12900 , n12901 );
xnor ( n12903 , n12902 , n4315 );
xor ( n12904 , n12899 , n12903 );
and ( n12905 , n10857 , n4298 );
and ( n12906 , n11295 , n4287 );
nor ( n12907 , n12905 , n12906 );
xnor ( n12908 , n12907 , n4294 );
and ( n12909 , n9989 , n4788 );
and ( n12910 , n10437 , n4611 );
nor ( n12911 , n12909 , n12910 );
xnor ( n12912 , n12911 , n4784 );
xor ( n12913 , n12908 , n12912 );
and ( n12914 , n6516 , n7356 );
and ( n12915 , n6907 , n6953 );
nor ( n12916 , n12914 , n12915 );
xnor ( n12917 , n12916 , n7352 );
and ( n12918 , n6168 , n7349 );
xor ( n12919 , n12917 , n12918 );
and ( n12920 , n12550 , n12551 );
xor ( n12921 , n12919 , n12920 );
and ( n12922 , n7324 , n6554 );
and ( n12923 , n7752 , n6205 );
nor ( n12924 , n12922 , n12923 );
xnor ( n12925 , n12924 , n6550 );
xor ( n12926 , n12921 , n12925 );
xor ( n12927 , n12913 , n12926 );
xor ( n12928 , n12904 , n12927 );
and ( n12929 , n12486 , n12530 );
and ( n12930 , n12530 , n12535 );
and ( n12931 , n12486 , n12535 );
or ( n12932 , n12929 , n12930 , n12931 );
and ( n12933 , n12541 , n12545 );
and ( n12934 , n12545 , n12559 );
and ( n12935 , n12541 , n12559 );
or ( n12936 , n12933 , n12934 , n12935 );
xor ( n12937 , n12932 , n12936 );
and ( n12938 , n12552 , n12553 );
and ( n12939 , n12553 , n12558 );
and ( n12940 , n12552 , n12558 );
or ( n12941 , n12938 , n12939 , n12940 );
and ( n12942 , n9110 , n5270 );
and ( n12943 , n9583 , n5021 );
nor ( n12944 , n12942 , n12943 );
xnor ( n12945 , n12944 , n5266 );
xor ( n12946 , n12941 , n12945 );
and ( n12947 , n8179 , n5850 );
and ( n12948 , n8640 , n5566 );
nor ( n12949 , n12947 , n12948 );
xnor ( n12950 , n12949 , n5846 );
xor ( n12951 , n12946 , n12950 );
xor ( n12952 , n12937 , n12951 );
xor ( n12953 , n12928 , n12952 );
xor ( n12954 , n12854 , n12953 );
and ( n12955 , n12453 , n12477 );
and ( n12956 , n12477 , n12561 );
and ( n12957 , n12453 , n12561 );
or ( n12958 , n12955 , n12956 , n12957 );
xor ( n12959 , n12954 , n12958 );
and ( n12960 , n12562 , n12566 );
and ( n12961 , n12567 , n12570 );
or ( n12962 , n12960 , n12961 );
xor ( n12963 , n12959 , n12962 );
buf ( n12964 , n12963 );
and ( n12965 , n12580 , n12584 );
and ( n12966 , n12584 , n12599 );
and ( n12967 , n12580 , n12599 );
or ( n12968 , n12965 , n12966 , n12967 );
and ( n12969 , n12626 , n12630 );
and ( n12970 , n12630 , n12644 );
and ( n12971 , n12626 , n12644 );
or ( n12972 , n12969 , n12970 , n12971 );
xor ( n12973 , n12968 , n12972 );
and ( n12974 , n12612 , n4418 );
buf ( n12975 , n4126 );
buf ( n12976 , n12975 );
and ( n12977 , n12976 , n4415 );
nor ( n12978 , n12974 , n12977 );
xnor ( n12979 , n12978 , n4413 );
and ( n12980 , n6604 , n7444 );
and ( n12981 , n6995 , n7026 );
nor ( n12982 , n12980 , n12981 );
xnor ( n12983 , n12982 , n7440 );
xor ( n12984 , n12979 , n12983 );
and ( n12985 , n6235 , n7437 );
xor ( n12986 , n12984 , n12985 );
and ( n12987 , n12635 , n12636 );
and ( n12988 , n7417 , n6627 );
and ( n12989 , n7857 , n6272 );
nor ( n12990 , n12988 , n12989 );
xnor ( n12991 , n12990 , n6623 );
xor ( n12992 , n12987 , n12991 );
xor ( n12993 , n12986 , n12992 );
and ( n12994 , n12609 , n12615 );
and ( n12995 , n12615 , n12620 );
and ( n12996 , n12609 , n12620 );
or ( n12997 , n12994 , n12995 , n12996 );
xor ( n12998 , n12993 , n12997 );
xor ( n12999 , n12973 , n12998 );
and ( n13000 , n12605 , n12621 );
and ( n13001 , n12621 , n12645 );
and ( n13002 , n12605 , n12645 );
or ( n13003 , n13000 , n13001 , n13002 );
and ( n13004 , n12589 , n12593 );
and ( n13005 , n12593 , n12598 );
and ( n13006 , n12589 , n12598 );
or ( n13007 , n13004 , n13005 , n13006 );
and ( n13008 , n11784 , n4433 );
and ( n13009 , n12217 , n4431 );
nor ( n13010 , n13008 , n13009 );
xnor ( n13011 , n13010 , n4441 );
and ( n13012 , n10072 , n4835 );
and ( n13013 , n10534 , n4648 );
nor ( n13014 , n13012 , n13013 );
xnor ( n13015 , n13014 , n4831 );
xor ( n13016 , n13011 , n13015 );
and ( n13017 , n8303 , n5922 );
and ( n13018 , n8728 , n5616 );
nor ( n13019 , n13017 , n13018 );
xnor ( n13020 , n13019 , n5918 );
xor ( n13021 , n13016 , n13020 );
xor ( n13022 , n13007 , n13021 );
and ( n13023 , n12637 , n12638 );
and ( n13024 , n12638 , n12643 );
and ( n13025 , n12637 , n12643 );
or ( n13026 , n13023 , n13024 , n13025 );
and ( n13027 , n10940 , n4402 );
and ( n13028 , n11398 , n4391 );
nor ( n13029 , n13027 , n13028 );
xnor ( n13030 , n13029 , n4398 );
xor ( n13031 , n13026 , n13030 );
and ( n13032 , n9164 , n5323 );
and ( n13033 , n9629 , n5064 );
nor ( n13034 , n13032 , n13033 );
xnor ( n13035 , n13034 , n5319 );
xor ( n13036 , n13031 , n13035 );
xor ( n13037 , n13022 , n13036 );
xor ( n13038 , n13003 , n13037 );
xor ( n13039 , n12999 , n13038 );
and ( n13040 , n12576 , n12600 );
and ( n13041 , n12600 , n12646 );
and ( n13042 , n12576 , n12646 );
or ( n13043 , n13040 , n13041 , n13042 );
xor ( n13044 , n13039 , n13043 );
and ( n13045 , n12647 , n12651 );
and ( n13046 , n12651 , n12656 );
and ( n13047 , n12647 , n12656 );
or ( n13048 , n13045 , n13046 , n13047 );
xor ( n13049 , n13044 , n13048 );
and ( n13050 , n12657 , n12658 );
xor ( n13051 , n13049 , n13050 );
buf ( n13052 , n13051 );
not ( n13053 , n454 );
and ( n13054 , n13053 , n12964 );
and ( n13055 , n13052 , n454 );
or ( n13056 , n13054 , n13055 );
buf ( n13057 , n13056 );
buf ( n13058 , n13057 );
and ( n13059 , n13058 , n4505 );
xor ( n13060 , n12845 , n13059 );
xor ( n13061 , n12842 , n13060 );
and ( n13062 , n12449 , n12667 );
and ( n13063 , n12667 , n12673 );
and ( n13064 , n12449 , n12673 );
or ( n13065 , n13062 , n13063 , n13064 );
xor ( n13066 , n13061 , n13065 );
and ( n13067 , n12674 , n12678 );
and ( n13068 , n12678 , n12683 );
and ( n13069 , n12674 , n12683 );
or ( n13070 , n13067 , n13068 , n13069 );
xor ( n13071 , n13066 , n13070 );
or ( n13072 , n12684 , n12685 );
xnor ( n13073 , n13071 , n13072 );
and ( n13074 , n12686 , n12687 );
xor ( n13075 , n13073 , n13074 );
buf ( n13076 , n13075 );
not ( n13077 , n4509 );
and ( n13078 , n13077 , n12836 );
and ( n13079 , n13076 , n4509 );
or ( n13080 , n13078 , n13079 );
and ( n13081 , n12782 , n12786 );
and ( n13082 , n12786 , n12821 );
and ( n13083 , n12782 , n12821 );
or ( n13084 , n13081 , n13082 , n13083 );
and ( n13085 , n12766 , n12770 );
and ( n13086 , n12770 , n12775 );
and ( n13087 , n12766 , n12775 );
or ( n13088 , n13085 , n13086 , n13087 );
and ( n13089 , n12791 , n12795 );
and ( n13090 , n12795 , n12820 );
and ( n13091 , n12791 , n12820 );
or ( n13092 , n13089 , n13090 , n13091 );
xor ( n13093 , n13088 , n13092 );
and ( n13094 , n12754 , n4524 );
and ( n13095 , n12702 , n12716 );
and ( n13096 , n12716 , n12738 );
and ( n13097 , n12702 , n12738 );
or ( n13098 , n13095 , n13096 , n13097 );
and ( n13099 , n12706 , n12710 );
and ( n13100 , n12710 , n12715 );
and ( n13101 , n12706 , n12715 );
or ( n13102 , n13099 , n13100 , n13101 );
and ( n13103 , n12721 , n12725 );
and ( n13104 , n12725 , n12737 );
and ( n13105 , n12721 , n12737 );
or ( n13106 , n13103 , n13104 , n13105 );
xor ( n13107 , n13102 , n13106 );
and ( n13108 , n12730 , n12734 );
and ( n13109 , n12734 , n12736 );
and ( n13110 , n12730 , n12736 );
or ( n13111 , n13108 , n13109 , n13110 );
not ( n13112 , n6004 );
and ( n13113 , n9297 , n6761 );
and ( n13114 , n9848 , n6379 );
nor ( n13115 , n13113 , n13114 );
xnor ( n13116 , n13115 , n6757 );
xor ( n13117 , n13112 , n13116 );
and ( n13118 , n7531 , n8382 );
and ( n13119 , n8001 , n8042 );
nor ( n13120 , n13118 , n13119 );
xnor ( n13121 , n13120 , n8378 );
xor ( n13122 , n13117 , n13121 );
xor ( n13123 , n13111 , n13122 );
buf ( n13124 , n12709 );
and ( n13125 , n8409 , n7559 );
and ( n13126 , n8900 , n7107 );
nor ( n13127 , n13125 , n13126 );
xnor ( n13128 , n13127 , n7555 );
xor ( n13129 , n13124 , n13128 );
and ( n13130 , n7092 , n8375 );
xor ( n13131 , n13129 , n13130 );
xor ( n13132 , n13123 , n13131 );
xor ( n13133 , n13107 , n13132 );
xor ( n13134 , n13098 , n13133 );
and ( n13135 , n12739 , n12743 );
and ( n13136 , n12743 , n12748 );
and ( n13137 , n12739 , n12748 );
or ( n13138 , n13135 , n13136 , n13137 );
xor ( n13139 , n13134 , n13138 );
and ( n13140 , n12749 , n12750 );
xor ( n13141 , n13139 , n13140 );
buf ( n13142 , n13141 );
buf ( n13143 , n13142 );
buf ( n13144 , n13143 );
and ( n13145 , n13144 , n4145 );
nor ( n13146 , n13094 , n13145 );
xnor ( n13147 , n13146 , n4521 );
xor ( n13148 , n13093 , n13147 );
xor ( n13149 , n13084 , n13148 );
and ( n13150 , n12757 , n12761 );
and ( n13151 , n12761 , n12776 );
and ( n13152 , n12757 , n12776 );
or ( n13153 , n13150 , n13151 , n13152 );
and ( n13154 , n11989 , n4938 );
and ( n13155 , n12392 , n4711 );
nor ( n13156 , n13154 , n13155 );
xnor ( n13157 , n13156 , n4934 );
and ( n13158 , n11163 , n5441 );
and ( n13159 , n11569 , n5161 );
nor ( n13160 , n13158 , n13159 );
xnor ( n13161 , n13160 , n5437 );
xor ( n13162 , n13157 , n13161 );
and ( n13163 , n12809 , n12813 );
and ( n13164 , n12813 , n12818 );
and ( n13165 , n12809 , n12818 );
or ( n13166 , n13163 , n13164 , n13165 );
and ( n13167 , n9367 , n6711 );
and ( n13168 , n9885 , n6332 );
nor ( n13169 , n13167 , n13168 );
xnor ( n13170 , n13169 , n6707 );
xor ( n13171 , n13166 , n13170 );
and ( n13172 , n8462 , n7630 );
and ( n13173 , n8968 , n7188 );
nor ( n13174 , n13172 , n13173 );
xnor ( n13175 , n13174 , n7626 );
xor ( n13176 , n13171 , n13175 );
xor ( n13177 , n13162 , n13176 );
xor ( n13178 , n13153 , n13177 );
and ( n13179 , n7587 , n8502 );
and ( n13180 , n8057 , n7970 );
nor ( n13181 , n13179 , n13180 );
xnor ( n13182 , n13181 , n8498 );
and ( n13183 , n6796 , n9407 );
and ( n13184 , n7146 , n8872 );
nor ( n13185 , n13183 , n13184 );
xnor ( n13186 , n13185 , n9403 );
and ( n13187 , n6037 , n10329 );
and ( n13188 , n6391 , n9791 );
nor ( n13189 , n13187 , n13188 );
not ( n13190 , n13189 );
xor ( n13191 , n13186 , n13190 );
xor ( n13192 , n13182 , n13191 );
and ( n13193 , n12800 , n12804 );
and ( n13194 , n12804 , n12819 );
and ( n13195 , n12800 , n12819 );
or ( n13196 , n13193 , n13194 , n13195 );
xor ( n13197 , n13192 , n13196 );
and ( n13198 , n10287 , n6068 );
and ( n13199 , n10706 , n5730 );
nor ( n13200 , n13198 , n13199 );
xnor ( n13201 , n13200 , n6064 );
xor ( n13202 , n13197 , n13201 );
xor ( n13203 , n13178 , n13202 );
xor ( n13204 , n13149 , n13203 );
and ( n13205 , n12697 , n12777 );
and ( n13206 , n12777 , n12822 );
and ( n13207 , n12697 , n12822 );
or ( n13208 , n13205 , n13206 , n13207 );
xor ( n13209 , n13204 , n13208 );
and ( n13210 , n12823 , n12827 );
and ( n13211 , n12827 , n12832 );
and ( n13212 , n12823 , n12832 );
or ( n13213 , n13210 , n13211 , n13212 );
xor ( n13214 , n13209 , n13213 );
and ( n13215 , n12833 , n12834 );
xor ( n13216 , n13214 , n13215 );
buf ( n13217 , n13216 );
and ( n13218 , n12843 , n12844 );
and ( n13219 , n12844 , n13059 );
and ( n13220 , n12843 , n13059 );
or ( n13221 , n13218 , n13219 , n13220 );
and ( n13222 , n12904 , n12927 );
and ( n13223 , n12927 , n12952 );
and ( n13224 , n12904 , n12952 );
or ( n13225 , n13222 , n13223 , n13224 );
and ( n13226 , n12849 , n12853 );
and ( n13227 , n12853 , n12953 );
and ( n13228 , n12849 , n12953 );
or ( n13229 , n13226 , n13227 , n13228 );
xor ( n13230 , n13225 , n13229 );
and ( n13231 , n12908 , n12912 );
and ( n13232 , n12912 , n12926 );
and ( n13233 , n12908 , n12926 );
or ( n13234 , n13231 , n13232 , n13233 );
and ( n13235 , n12919 , n12920 );
and ( n13236 , n12920 , n12925 );
and ( n13237 , n12919 , n12925 );
or ( n13238 , n13235 , n13236 , n13237 );
and ( n13239 , n9583 , n5270 );
and ( n13240 , n9989 , n5021 );
nor ( n13241 , n13239 , n13240 );
xnor ( n13242 , n13241 , n5266 );
xor ( n13243 , n13238 , n13242 );
and ( n13244 , n8640 , n5850 );
and ( n13245 , n9110 , n5566 );
nor ( n13246 , n13244 , n13245 );
xnor ( n13247 , n13246 , n5846 );
xor ( n13248 , n13243 , n13247 );
xor ( n13249 , n13234 , n13248 );
and ( n13250 , n12917 , n12918 );
and ( n13251 , n11295 , n4298 );
and ( n13252 , n11702 , n4287 );
nor ( n13253 , n13251 , n13252 );
xnor ( n13254 , n13253 , n4294 );
and ( n13255 , n7752 , n6554 );
and ( n13256 , n8179 , n6205 );
nor ( n13257 , n13255 , n13256 );
xnor ( n13258 , n13257 , n6550 );
xor ( n13259 , n13254 , n13258 );
and ( n13260 , n6907 , n7356 );
and ( n13261 , n7324 , n6953 );
nor ( n13262 , n13260 , n13261 );
xnor ( n13263 , n13262 , n7352 );
and ( n13264 , n6516 , n7349 );
xor ( n13265 , n13263 , n13264 );
xor ( n13266 , n13259 , n13265 );
xor ( n13267 , n13250 , n13266 );
and ( n13268 , n12941 , n12945 );
and ( n13269 , n12945 , n12950 );
and ( n13270 , n12941 , n12950 );
or ( n13271 , n13268 , n13269 , n13270 );
xor ( n13272 , n13267 , n13271 );
xor ( n13273 , n13249 , n13272 );
and ( n13274 , n12858 , n12898 );
and ( n13275 , n12898 , n12903 );
and ( n13276 , n12858 , n12903 );
or ( n13277 , n13274 , n13275 , n13276 );
and ( n13278 , n12932 , n12936 );
and ( n13279 , n12936 , n12951 );
and ( n13280 , n12932 , n12951 );
or ( n13281 , n13278 , n13279 , n13280 );
xor ( n13282 , n13277 , n13281 );
and ( n13283 , n12895 , n4235 );
and ( n13284 , n12872 , n12876 );
and ( n13285 , n12876 , n12878 );
and ( n13286 , n12872 , n12878 );
or ( n13287 , n13284 , n13285 , n13286 );
buf ( n13288 , n12871 );
xor ( n13289 , n13287 , n13288 );
not ( n13290 , n6453 );
and ( n13291 , n6853 , n7277 );
and ( n13292 , n7299 , n6864 );
nor ( n13293 , n13291 , n13292 );
xnor ( n13294 , n13293 , n7283 );
xor ( n13295 , n13290 , n13294 );
and ( n13296 , n6444 , n7274 );
xor ( n13297 , n13295 , n13296 );
xor ( n13298 , n13289 , n13297 );
and ( n13299 , n12863 , n12867 );
and ( n13300 , n12867 , n12879 );
and ( n13301 , n12863 , n12879 );
or ( n13302 , n13299 , n13300 , n13301 );
xor ( n13303 , n13298 , n13302 );
and ( n13304 , n12880 , n12884 );
and ( n13305 , n12884 , n12889 );
and ( n13306 , n12880 , n12889 );
or ( n13307 , n13304 , n13305 , n13306 );
xor ( n13308 , n13303 , n13307 );
and ( n13309 , n12890 , n12891 );
xor ( n13310 , n13308 , n13309 );
buf ( n13311 , n13310 );
buf ( n13312 , n13311 );
buf ( n13313 , n13312 );
and ( n13314 , n13313 , n4232 );
nor ( n13315 , n13283 , n13314 );
xnor ( n13316 , n13315 , n4230 );
and ( n13317 , n12116 , n4319 );
and ( n13318 , n12527 , n4310 );
nor ( n13319 , n13317 , n13318 );
xnor ( n13320 , n13319 , n4315 );
xor ( n13321 , n13316 , n13320 );
and ( n13322 , n10437 , n4788 );
and ( n13323 , n10857 , n4611 );
nor ( n13324 , n13322 , n13323 );
xnor ( n13325 , n13324 , n4784 );
xor ( n13326 , n13321 , n13325 );
xor ( n13327 , n13282 , n13326 );
xor ( n13328 , n13273 , n13327 );
xor ( n13329 , n13230 , n13328 );
and ( n13330 , n12954 , n12958 );
and ( n13331 , n12959 , n12962 );
or ( n13332 , n13330 , n13331 );
xor ( n13333 , n13329 , n13332 );
buf ( n13334 , n13333 );
and ( n13335 , n12999 , n13038 );
and ( n13336 , n13038 , n13043 );
and ( n13337 , n12999 , n13043 );
or ( n13338 , n13335 , n13336 , n13337 );
and ( n13339 , n12968 , n12972 );
and ( n13340 , n12972 , n12998 );
and ( n13341 , n12968 , n12998 );
or ( n13342 , n13339 , n13340 , n13341 );
and ( n13343 , n13007 , n13021 );
and ( n13344 , n13021 , n13036 );
and ( n13345 , n13007 , n13036 );
or ( n13346 , n13343 , n13344 , n13345 );
and ( n13347 , n12986 , n12992 );
and ( n13348 , n12992 , n12997 );
and ( n13349 , n12986 , n12997 );
or ( n13350 , n13347 , n13348 , n13349 );
xor ( n13351 , n13346 , n13350 );
and ( n13352 , n7857 , n6627 );
and ( n13353 , n8303 , n6272 );
nor ( n13354 , n13352 , n13353 );
xnor ( n13355 , n13354 , n6623 );
and ( n13356 , n6995 , n7444 );
and ( n13357 , n7417 , n7026 );
nor ( n13358 , n13356 , n13357 );
xnor ( n13359 , n13358 , n7440 );
and ( n13360 , n6604 , n7437 );
xor ( n13361 , n13359 , n13360 );
xor ( n13362 , n13355 , n13361 );
and ( n13363 , n12979 , n12983 );
and ( n13364 , n12983 , n12985 );
and ( n13365 , n12979 , n12985 );
or ( n13366 , n13363 , n13364 , n13365 );
xor ( n13367 , n13362 , n13366 );
and ( n13368 , n13026 , n13030 );
and ( n13369 , n13030 , n13035 );
and ( n13370 , n13026 , n13035 );
or ( n13371 , n13368 , n13369 , n13370 );
xor ( n13372 , n13367 , n13371 );
and ( n13373 , n12976 , n4418 );
not ( n13374 , n13373 );
xnor ( n13375 , n13374 , n4413 );
and ( n13376 , n11398 , n4402 );
and ( n13377 , n11784 , n4391 );
nor ( n13378 , n13376 , n13377 );
xnor ( n13379 , n13378 , n4398 );
xor ( n13380 , n13375 , n13379 );
and ( n13381 , n9629 , n5323 );
and ( n13382 , n10072 , n5064 );
nor ( n13383 , n13381 , n13382 );
xnor ( n13384 , n13383 , n5319 );
xor ( n13385 , n13380 , n13384 );
and ( n13386 , n13011 , n13015 );
and ( n13387 , n13015 , n13020 );
and ( n13388 , n13011 , n13020 );
or ( n13389 , n13386 , n13387 , n13388 );
and ( n13390 , n12217 , n4433 );
and ( n13391 , n12612 , n4431 );
nor ( n13392 , n13390 , n13391 );
xnor ( n13393 , n13392 , n4441 );
and ( n13394 , n10534 , n4835 );
and ( n13395 , n10940 , n4648 );
nor ( n13396 , n13394 , n13395 );
xnor ( n13397 , n13396 , n4831 );
xor ( n13398 , n13393 , n13397 );
and ( n13399 , n8728 , n5922 );
and ( n13400 , n9164 , n5616 );
nor ( n13401 , n13399 , n13400 );
xnor ( n13402 , n13401 , n5918 );
xor ( n13403 , n13398 , n13402 );
xor ( n13404 , n13389 , n13403 );
xor ( n13405 , n13385 , n13404 );
and ( n13406 , n12987 , n12991 );
xor ( n13407 , n13405 , n13406 );
xor ( n13408 , n13372 , n13407 );
xor ( n13409 , n13351 , n13408 );
xor ( n13410 , n13342 , n13409 );
and ( n13411 , n13003 , n13037 );
xor ( n13412 , n13410 , n13411 );
xor ( n13413 , n13338 , n13412 );
and ( n13414 , n13044 , n13048 );
and ( n13415 , n13049 , n13050 );
or ( n13416 , n13414 , n13415 );
xor ( n13417 , n13413 , n13416 );
buf ( n13418 , n13417 );
not ( n13419 , n454 );
and ( n13420 , n13419 , n13334 );
and ( n13421 , n13418 , n454 );
or ( n13422 , n13420 , n13421 );
buf ( n13423 , n13422 );
buf ( n13424 , n13423 );
and ( n13425 , n13424 , n4505 );
xor ( n13426 , n13221 , n13425 );
and ( n13427 , n12275 , n5089 );
and ( n13428 , n12666 , n4866 );
xor ( n13429 , n13427 , n13428 );
and ( n13430 , n13058 , n4557 );
xor ( n13431 , n13429 , n13430 );
xor ( n13432 , n13426 , n13431 );
and ( n13433 , n12840 , n12841 );
and ( n13434 , n12841 , n13060 );
and ( n13435 , n12840 , n13060 );
or ( n13436 , n13433 , n13434 , n13435 );
xor ( n13437 , n13432 , n13436 );
and ( n13438 , n13061 , n13065 );
and ( n13439 , n13065 , n13070 );
and ( n13440 , n13061 , n13070 );
or ( n13441 , n13438 , n13439 , n13440 );
xor ( n13442 , n13437 , n13441 );
or ( n13443 , n13071 , n13072 );
xnor ( n13444 , n13442 , n13443 );
and ( n13445 , n13073 , n13074 );
xor ( n13446 , n13444 , n13445 );
buf ( n13447 , n13446 );
not ( n13448 , n4509 );
and ( n13449 , n13448 , n13217 );
and ( n13450 , n13447 , n4509 );
or ( n13451 , n13449 , n13450 );
and ( n13452 , n13153 , n13177 );
and ( n13453 , n13177 , n13202 );
and ( n13454 , n13153 , n13202 );
or ( n13455 , n13452 , n13453 , n13454 );
and ( n13456 , n13192 , n13196 );
and ( n13457 , n13196 , n13201 );
and ( n13458 , n13192 , n13201 );
or ( n13459 , n13456 , n13457 , n13458 );
and ( n13460 , n13144 , n4524 );
and ( n13461 , n13111 , n13122 );
and ( n13462 , n13122 , n13131 );
and ( n13463 , n13111 , n13131 );
or ( n13464 , n13461 , n13462 , n13463 );
and ( n13465 , n8900 , n7559 );
and ( n13466 , n9297 , n7107 );
nor ( n13467 , n13465 , n13466 );
xnor ( n13468 , n13467 , n7555 );
and ( n13469 , n8001 , n8382 );
and ( n13470 , n8409 , n8042 );
nor ( n13471 , n13469 , n13470 );
xnor ( n13472 , n13471 , n8378 );
xor ( n13473 , n13468 , n13472 );
and ( n13474 , n7531 , n8375 );
xor ( n13475 , n13473 , n13474 );
xor ( n13476 , n13464 , n13475 );
and ( n13477 , n13112 , n13116 );
and ( n13478 , n13116 , n13121 );
and ( n13479 , n13112 , n13121 );
or ( n13480 , n13477 , n13478 , n13479 );
and ( n13481 , n13124 , n13128 );
and ( n13482 , n13128 , n13130 );
and ( n13483 , n13124 , n13130 );
or ( n13484 , n13481 , n13482 , n13483 );
xor ( n13485 , n13480 , n13484 );
and ( n13486 , n9848 , n6761 );
not ( n13487 , n13486 );
xnor ( n13488 , n13487 , n6757 );
not ( n13489 , n13488 );
xor ( n13490 , n13485 , n13489 );
xor ( n13491 , n13476 , n13490 );
and ( n13492 , n13102 , n13106 );
and ( n13493 , n13106 , n13132 );
and ( n13494 , n13102 , n13132 );
or ( n13495 , n13492 , n13493 , n13494 );
xor ( n13496 , n13491 , n13495 );
and ( n13497 , n13098 , n13133 );
and ( n13498 , n13133 , n13138 );
and ( n13499 , n13098 , n13138 );
or ( n13500 , n13497 , n13498 , n13499 );
xor ( n13501 , n13496 , n13500 );
and ( n13502 , n13139 , n13140 );
xor ( n13503 , n13501 , n13502 );
buf ( n13504 , n13503 );
buf ( n13505 , n13504 );
buf ( n13506 , n13505 );
and ( n13507 , n13506 , n4145 );
nor ( n13508 , n13460 , n13507 );
xnor ( n13509 , n13508 , n4521 );
xor ( n13510 , n13459 , n13509 );
and ( n13511 , n13166 , n13170 );
and ( n13512 , n13170 , n13175 );
and ( n13513 , n13166 , n13175 );
or ( n13514 , n13511 , n13512 , n13513 );
and ( n13515 , n10706 , n6068 );
and ( n13516 , n11163 , n5730 );
nor ( n13517 , n13515 , n13516 );
xnor ( n13518 , n13517 , n6064 );
xor ( n13519 , n13514 , n13518 );
and ( n13520 , n9885 , n6711 );
and ( n13521 , n10287 , n6332 );
nor ( n13522 , n13520 , n13521 );
xnor ( n13523 , n13522 , n6707 );
xor ( n13524 , n13519 , n13523 );
xor ( n13525 , n13510 , n13524 );
xor ( n13526 , n13455 , n13525 );
and ( n13527 , n13088 , n13092 );
and ( n13528 , n13092 , n13147 );
and ( n13529 , n13088 , n13147 );
or ( n13530 , n13527 , n13528 , n13529 );
and ( n13531 , n13157 , n13161 );
and ( n13532 , n13161 , n13176 );
and ( n13533 , n13157 , n13176 );
or ( n13534 , n13531 , n13532 , n13533 );
xor ( n13535 , n13530 , n13534 );
and ( n13536 , n12392 , n4938 );
and ( n13537 , n12754 , n4711 );
nor ( n13538 , n13536 , n13537 );
xnor ( n13539 , n13538 , n4934 );
and ( n13540 , n11569 , n5441 );
and ( n13541 , n11989 , n5161 );
nor ( n13542 , n13540 , n13541 );
xnor ( n13543 , n13542 , n5437 );
xor ( n13544 , n13539 , n13543 );
and ( n13545 , n13182 , n13191 );
and ( n13546 , n8968 , n7630 );
and ( n13547 , n9367 , n7188 );
nor ( n13548 , n13546 , n13547 );
xnor ( n13549 , n13548 , n7626 );
xor ( n13550 , n13545 , n13549 );
and ( n13551 , n7146 , n9407 );
and ( n13552 , n7587 , n8872 );
nor ( n13553 , n13551 , n13552 );
xnor ( n13554 , n13553 , n9403 );
and ( n13555 , n6391 , n10329 );
and ( n13556 , n6796 , n9791 );
nor ( n13557 , n13555 , n13556 );
not ( n13558 , n13557 );
xor ( n13559 , n13554 , n13558 );
and ( n13560 , n13186 , n13190 );
xor ( n13561 , n13559 , n13560 );
and ( n13562 , n8057 , n8502 );
and ( n13563 , n8462 , n7970 );
nor ( n13564 , n13562 , n13563 );
xnor ( n13565 , n13564 , n8498 );
xor ( n13566 , n13561 , n13565 );
xor ( n13567 , n13550 , n13566 );
xor ( n13568 , n13544 , n13567 );
xor ( n13569 , n13535 , n13568 );
xor ( n13570 , n13526 , n13569 );
and ( n13571 , n13084 , n13148 );
and ( n13572 , n13148 , n13203 );
and ( n13573 , n13084 , n13203 );
or ( n13574 , n13571 , n13572 , n13573 );
xor ( n13575 , n13570 , n13574 );
and ( n13576 , n13204 , n13208 );
and ( n13577 , n13208 , n13213 );
and ( n13578 , n13204 , n13213 );
or ( n13579 , n13576 , n13577 , n13578 );
xor ( n13580 , n13575 , n13579 );
and ( n13581 , n13214 , n13215 );
xor ( n13582 , n13580 , n13581 );
buf ( n13583 , n13582 );
and ( n13584 , n13427 , n13428 );
and ( n13585 , n13428 , n13430 );
and ( n13586 , n13427 , n13430 );
or ( n13587 , n13584 , n13585 , n13586 );
and ( n13588 , n13424 , n4557 );
xor ( n13589 , n13587 , n13588 );
and ( n13590 , n12666 , n5089 );
and ( n13591 , n13058 , n4866 );
xor ( n13592 , n13590 , n13591 );
and ( n13593 , n13225 , n13229 );
and ( n13594 , n13229 , n13328 );
and ( n13595 , n13225 , n13328 );
or ( n13596 , n13593 , n13594 , n13595 );
and ( n13597 , n13234 , n13248 );
and ( n13598 , n13250 , n13266 );
and ( n13599 , n13266 , n13271 );
and ( n13600 , n13250 , n13271 );
or ( n13601 , n13598 , n13599 , n13600 );
xor ( n13602 , n13597 , n13601 );
and ( n13603 , n8179 , n6554 );
and ( n13604 , n8640 , n6205 );
nor ( n13605 , n13603 , n13604 );
xnor ( n13606 , n13605 , n6550 );
and ( n13607 , n7324 , n7356 );
and ( n13608 , n7752 , n6953 );
nor ( n13609 , n13607 , n13608 );
xnor ( n13610 , n13609 , n7352 );
and ( n13611 , n6907 , n7349 );
xor ( n13612 , n13610 , n13611 );
xor ( n13613 , n13606 , n13612 );
and ( n13614 , n13263 , n13264 );
xor ( n13615 , n13613 , n13614 );
and ( n13616 , n13238 , n13242 );
and ( n13617 , n13242 , n13247 );
and ( n13618 , n13238 , n13247 );
or ( n13619 , n13616 , n13617 , n13618 );
xor ( n13620 , n13615 , n13619 );
and ( n13621 , n13313 , n4235 );
and ( n13622 , n13290 , n13294 );
and ( n13623 , n13294 , n13296 );
and ( n13624 , n13290 , n13296 );
or ( n13625 , n13622 , n13623 , n13624 );
and ( n13626 , n7299 , n7277 );
not ( n13627 , n13626 );
xnor ( n13628 , n13627 , n7283 );
xor ( n13629 , n13625 , n13628 );
and ( n13630 , n6853 , n7274 );
not ( n13631 , n13630 );
xor ( n13632 , n13629 , n13631 );
and ( n13633 , n13287 , n13288 );
and ( n13634 , n13288 , n13297 );
and ( n13635 , n13287 , n13297 );
or ( n13636 , n13633 , n13634 , n13635 );
xor ( n13637 , n13632 , n13636 );
and ( n13638 , n13298 , n13302 );
and ( n13639 , n13302 , n13307 );
and ( n13640 , n13298 , n13307 );
or ( n13641 , n13638 , n13639 , n13640 );
xor ( n13642 , n13637 , n13641 );
and ( n13643 , n13308 , n13309 );
xor ( n13644 , n13642 , n13643 );
buf ( n13645 , n13644 );
buf ( n13646 , n13645 );
buf ( n13647 , n13646 );
and ( n13648 , n13647 , n4232 );
nor ( n13649 , n13621 , n13648 );
xnor ( n13650 , n13649 , n4230 );
and ( n13651 , n12527 , n4319 );
and ( n13652 , n12895 , n4310 );
nor ( n13653 , n13651 , n13652 );
xnor ( n13654 , n13653 , n4315 );
xor ( n13655 , n13650 , n13654 );
and ( n13656 , n11702 , n4298 );
and ( n13657 , n12116 , n4287 );
nor ( n13658 , n13656 , n13657 );
xnor ( n13659 , n13658 , n4294 );
xor ( n13660 , n13655 , n13659 );
and ( n13661 , n13316 , n13320 );
and ( n13662 , n13320 , n13325 );
and ( n13663 , n13316 , n13325 );
or ( n13664 , n13661 , n13662 , n13663 );
and ( n13665 , n10857 , n4788 );
and ( n13666 , n11295 , n4611 );
nor ( n13667 , n13665 , n13666 );
xnor ( n13668 , n13667 , n4784 );
and ( n13669 , n9989 , n5270 );
and ( n13670 , n10437 , n5021 );
nor ( n13671 , n13669 , n13670 );
xnor ( n13672 , n13671 , n5266 );
xor ( n13673 , n13668 , n13672 );
and ( n13674 , n9110 , n5850 );
and ( n13675 , n9583 , n5566 );
nor ( n13676 , n13674 , n13675 );
xnor ( n13677 , n13676 , n5846 );
xor ( n13678 , n13673 , n13677 );
xor ( n13679 , n13664 , n13678 );
xor ( n13680 , n13660 , n13679 );
and ( n13681 , n13254 , n13258 );
and ( n13682 , n13258 , n13265 );
and ( n13683 , n13254 , n13265 );
or ( n13684 , n13681 , n13682 , n13683 );
xor ( n13685 , n13680 , n13684 );
xor ( n13686 , n13620 , n13685 );
xor ( n13687 , n13602 , n13686 );
and ( n13688 , n13277 , n13281 );
and ( n13689 , n13281 , n13326 );
and ( n13690 , n13277 , n13326 );
or ( n13691 , n13688 , n13689 , n13690 );
xor ( n13692 , n13687 , n13691 );
and ( n13693 , n13249 , n13272 );
and ( n13694 , n13272 , n13327 );
and ( n13695 , n13249 , n13327 );
or ( n13696 , n13693 , n13694 , n13695 );
xor ( n13697 , n13692 , n13696 );
xor ( n13698 , n13596 , n13697 );
and ( n13699 , n13329 , n13332 );
xor ( n13700 , n13698 , n13699 );
buf ( n13701 , n13700 );
and ( n13702 , n13346 , n13350 );
and ( n13703 , n13350 , n13408 );
and ( n13704 , n13346 , n13408 );
or ( n13705 , n13702 , n13703 , n13704 );
and ( n13706 , n13375 , n13379 );
and ( n13707 , n13379 , n13384 );
and ( n13708 , n13375 , n13384 );
or ( n13709 , n13706 , n13707 , n13708 );
and ( n13710 , n13389 , n13403 );
xor ( n13711 , n13709 , n13710 );
and ( n13712 , n13355 , n13361 );
and ( n13713 , n13361 , n13366 );
and ( n13714 , n13355 , n13366 );
or ( n13715 , n13712 , n13713 , n13714 );
xor ( n13716 , n13711 , n13715 );
and ( n13717 , n13367 , n13371 );
and ( n13718 , n13371 , n13407 );
and ( n13719 , n13367 , n13407 );
or ( n13720 , n13717 , n13718 , n13719 );
xor ( n13721 , n13716 , n13720 );
and ( n13722 , n12612 , n4433 );
and ( n13723 , n12976 , n4431 );
nor ( n13724 , n13722 , n13723 );
xnor ( n13725 , n13724 , n4441 );
and ( n13726 , n10940 , n4835 );
and ( n13727 , n11398 , n4648 );
nor ( n13728 , n13726 , n13727 );
xnor ( n13729 , n13728 , n4831 );
xor ( n13730 , n13725 , n13729 );
and ( n13731 , n8303 , n6627 );
and ( n13732 , n8728 , n6272 );
nor ( n13733 , n13731 , n13732 );
xnor ( n13734 , n13733 , n6623 );
xor ( n13735 , n13730 , n13734 );
and ( n13736 , n10072 , n5323 );
and ( n13737 , n10534 , n5064 );
nor ( n13738 , n13736 , n13737 );
xnor ( n13739 , n13738 , n5319 );
and ( n13740 , n9164 , n5922 );
and ( n13741 , n9629 , n5616 );
nor ( n13742 , n13740 , n13741 );
xnor ( n13743 , n13742 , n5918 );
xor ( n13744 , n13739 , n13743 );
xor ( n13745 , n13735 , n13744 );
and ( n13746 , n13393 , n13397 );
and ( n13747 , n13397 , n13402 );
and ( n13748 , n13393 , n13402 );
or ( n13749 , n13746 , n13747 , n13748 );
xor ( n13750 , n13745 , n13749 );
and ( n13751 , n11784 , n4402 );
and ( n13752 , n12217 , n4391 );
nor ( n13753 , n13751 , n13752 );
xnor ( n13754 , n13753 , n4398 );
not ( n13755 , n4413 );
and ( n13756 , n6995 , n7437 );
xnor ( n13757 , n13755 , n13756 );
and ( n13758 , n13359 , n13360 );
xor ( n13759 , n13757 , n13758 );
and ( n13760 , n7417 , n7444 );
and ( n13761 , n7857 , n7026 );
nor ( n13762 , n13760 , n13761 );
xnor ( n13763 , n13762 , n7440 );
xor ( n13764 , n13759 , n13763 );
xor ( n13765 , n13754 , n13764 );
xor ( n13766 , n13750 , n13765 );
and ( n13767 , n13385 , n13404 );
and ( n13768 , n13404 , n13406 );
and ( n13769 , n13385 , n13406 );
or ( n13770 , n13767 , n13768 , n13769 );
xor ( n13771 , n13766 , n13770 );
xor ( n13772 , n13721 , n13771 );
xor ( n13773 , n13705 , n13772 );
and ( n13774 , n13342 , n13409 );
and ( n13775 , n13409 , n13411 );
and ( n13776 , n13342 , n13411 );
or ( n13777 , n13774 , n13775 , n13776 );
xor ( n13778 , n13773 , n13777 );
and ( n13779 , n13338 , n13412 );
and ( n13780 , n13413 , n13416 );
or ( n13781 , n13779 , n13780 );
xor ( n13782 , n13778 , n13781 );
buf ( n13783 , n13782 );
not ( n13784 , n454 );
and ( n13785 , n13784 , n13701 );
and ( n13786 , n13783 , n454 );
or ( n13787 , n13785 , n13786 );
buf ( n13788 , n13787 );
buf ( n13789 , n13788 );
and ( n13790 , n13789 , n4505 );
xor ( n13791 , n13592 , n13790 );
xor ( n13792 , n13589 , n13791 );
and ( n13793 , n13221 , n13425 );
and ( n13794 , n13425 , n13431 );
and ( n13795 , n13221 , n13431 );
or ( n13796 , n13793 , n13794 , n13795 );
xor ( n13797 , n13792 , n13796 );
and ( n13798 , n13432 , n13436 );
and ( n13799 , n13436 , n13441 );
and ( n13800 , n13432 , n13441 );
or ( n13801 , n13798 , n13799 , n13800 );
xor ( n13802 , n13797 , n13801 );
or ( n13803 , n13442 , n13443 );
xnor ( n13804 , n13802 , n13803 );
and ( n13805 , n13444 , n13445 );
xor ( n13806 , n13804 , n13805 );
buf ( n13807 , n13806 );
not ( n13808 , n4509 );
and ( n13809 , n13808 , n13583 );
and ( n13810 , n13807 , n4509 );
or ( n13811 , n13809 , n13810 );
and ( n13812 , n13530 , n13534 );
and ( n13813 , n13534 , n13568 );
and ( n13814 , n13530 , n13568 );
or ( n13815 , n13812 , n13813 , n13814 );
and ( n13816 , n13514 , n13518 );
and ( n13817 , n13518 , n13523 );
and ( n13818 , n13514 , n13523 );
or ( n13819 , n13816 , n13817 , n13818 );
and ( n13820 , n13539 , n13543 );
and ( n13821 , n13543 , n13567 );
and ( n13822 , n13539 , n13567 );
or ( n13823 , n13820 , n13821 , n13822 );
xor ( n13824 , n13819 , n13823 );
and ( n13825 , n13506 , n4524 );
and ( n13826 , n13464 , n13475 );
and ( n13827 , n13475 , n13490 );
and ( n13828 , n13464 , n13490 );
or ( n13829 , n13826 , n13827 , n13828 );
and ( n13830 , n13480 , n13484 );
and ( n13831 , n13484 , n13489 );
and ( n13832 , n13480 , n13489 );
or ( n13833 , n13830 , n13831 , n13832 );
not ( n13834 , n6757 );
and ( n13835 , n9297 , n7559 );
and ( n13836 , n9848 , n7107 );
nor ( n13837 , n13835 , n13836 );
xnor ( n13838 , n13837 , n7555 );
xor ( n13839 , n13834 , n13838 );
and ( n13840 , n8001 , n8375 );
xor ( n13841 , n13839 , n13840 );
xor ( n13842 , n13833 , n13841 );
and ( n13843 , n13468 , n13472 );
and ( n13844 , n13472 , n13474 );
and ( n13845 , n13468 , n13474 );
or ( n13846 , n13843 , n13844 , n13845 );
buf ( n13847 , n13488 );
xor ( n13848 , n13846 , n13847 );
and ( n13849 , n8409 , n8382 );
and ( n13850 , n8900 , n8042 );
nor ( n13851 , n13849 , n13850 );
xnor ( n13852 , n13851 , n8378 );
xor ( n13853 , n13848 , n13852 );
xor ( n13854 , n13842 , n13853 );
xor ( n13855 , n13829 , n13854 );
and ( n13856 , n13491 , n13495 );
and ( n13857 , n13495 , n13500 );
and ( n13858 , n13491 , n13500 );
or ( n13859 , n13856 , n13857 , n13858 );
xor ( n13860 , n13855 , n13859 );
and ( n13861 , n13501 , n13502 );
xor ( n13862 , n13860 , n13861 );
buf ( n13863 , n13862 );
buf ( n13864 , n13863 );
buf ( n13865 , n13864 );
and ( n13866 , n13865 , n4145 );
nor ( n13867 , n13825 , n13866 );
xnor ( n13868 , n13867 , n4521 );
xor ( n13869 , n13824 , n13868 );
xor ( n13870 , n13815 , n13869 );
and ( n13871 , n13459 , n13509 );
and ( n13872 , n13509 , n13524 );
and ( n13873 , n13459 , n13524 );
or ( n13874 , n13871 , n13872 , n13873 );
and ( n13875 , n13545 , n13549 );
and ( n13876 , n13549 , n13566 );
and ( n13877 , n13545 , n13566 );
or ( n13878 , n13875 , n13876 , n13877 );
and ( n13879 , n12754 , n4938 );
and ( n13880 , n13144 , n4711 );
nor ( n13881 , n13879 , n13880 );
xnor ( n13882 , n13881 , n4934 );
xor ( n13883 , n13878 , n13882 );
and ( n13884 , n11989 , n5441 );
and ( n13885 , n12392 , n5161 );
nor ( n13886 , n13884 , n13885 );
xnor ( n13887 , n13886 , n5437 );
xor ( n13888 , n13883 , n13887 );
xor ( n13889 , n13874 , n13888 );
and ( n13890 , n11163 , n6068 );
and ( n13891 , n11569 , n5730 );
nor ( n13892 , n13890 , n13891 );
xnor ( n13893 , n13892 , n6064 );
and ( n13894 , n13559 , n13560 );
and ( n13895 , n13560 , n13565 );
and ( n13896 , n13559 , n13565 );
or ( n13897 , n13894 , n13895 , n13896 );
and ( n13898 , n10287 , n6711 );
and ( n13899 , n10706 , n6332 );
nor ( n13900 , n13898 , n13899 );
xnor ( n13901 , n13900 , n6707 );
xor ( n13902 , n13897 , n13901 );
and ( n13903 , n9367 , n7630 );
and ( n13904 , n9885 , n7188 );
nor ( n13905 , n13903 , n13904 );
xnor ( n13906 , n13905 , n7626 );
xor ( n13907 , n13902 , n13906 );
xor ( n13908 , n13893 , n13907 );
and ( n13909 , n7587 , n9407 );
and ( n13910 , n8057 , n8872 );
nor ( n13911 , n13909 , n13910 );
xnor ( n13912 , n13911 , n9403 );
and ( n13913 , n6796 , n10329 );
and ( n13914 , n7146 , n9791 );
nor ( n13915 , n13913 , n13914 );
not ( n13916 , n13915 );
xor ( n13917 , n13912 , n13916 );
and ( n13918 , n13554 , n13558 );
xor ( n13919 , n13917 , n13918 );
and ( n13920 , n8462 , n8502 );
and ( n13921 , n8968 , n7970 );
nor ( n13922 , n13920 , n13921 );
xnor ( n13923 , n13922 , n8498 );
xor ( n13924 , n13919 , n13923 );
xor ( n13925 , n13908 , n13924 );
xor ( n13926 , n13889 , n13925 );
xor ( n13927 , n13870 , n13926 );
and ( n13928 , n13455 , n13525 );
and ( n13929 , n13525 , n13569 );
and ( n13930 , n13455 , n13569 );
or ( n13931 , n13928 , n13929 , n13930 );
xor ( n13932 , n13927 , n13931 );
and ( n13933 , n13570 , n13574 );
and ( n13934 , n13574 , n13579 );
and ( n13935 , n13570 , n13579 );
or ( n13936 , n13933 , n13934 , n13935 );
xor ( n13937 , n13932 , n13936 );
and ( n13938 , n13580 , n13581 );
xor ( n13939 , n13937 , n13938 );
buf ( n13940 , n13939 );
and ( n13941 , n13590 , n13591 );
and ( n13942 , n13591 , n13790 );
and ( n13943 , n13590 , n13790 );
or ( n13944 , n13941 , n13942 , n13943 );
and ( n13945 , n13597 , n13601 );
and ( n13946 , n13601 , n13686 );
and ( n13947 , n13597 , n13686 );
or ( n13948 , n13945 , n13946 , n13947 );
and ( n13949 , n13650 , n13654 );
and ( n13950 , n13654 , n13659 );
and ( n13951 , n13650 , n13659 );
or ( n13952 , n13949 , n13950 , n13951 );
and ( n13953 , n13664 , n13678 );
xor ( n13954 , n13952 , n13953 );
and ( n13955 , n13606 , n13612 );
and ( n13956 , n13612 , n13614 );
and ( n13957 , n13606 , n13614 );
or ( n13958 , n13955 , n13956 , n13957 );
xor ( n13959 , n13954 , n13958 );
and ( n13960 , n13615 , n13619 );
and ( n13961 , n13619 , n13685 );
and ( n13962 , n13615 , n13685 );
or ( n13963 , n13960 , n13961 , n13962 );
xor ( n13964 , n13959 , n13963 );
and ( n13965 , n12116 , n4298 );
and ( n13966 , n12527 , n4287 );
nor ( n13967 , n13965 , n13966 );
xnor ( n13968 , n13967 , n4294 );
and ( n13969 , n11295 , n4788 );
and ( n13970 , n11702 , n4611 );
nor ( n13971 , n13969 , n13970 );
xnor ( n13972 , n13971 , n4784 );
xor ( n13973 , n13968 , n13972 );
and ( n13974 , n12895 , n4319 );
and ( n13975 , n13313 , n4310 );
nor ( n13976 , n13974 , n13975 );
xnor ( n13977 , n13976 , n4315 );
and ( n13978 , n10437 , n5270 );
and ( n13979 , n10857 , n5021 );
nor ( n13980 , n13978 , n13979 );
xnor ( n13981 , n13980 , n5266 );
xor ( n13982 , n13977 , n13981 );
and ( n13983 , n9583 , n5850 );
and ( n13984 , n9989 , n5566 );
nor ( n13985 , n13983 , n13984 );
xnor ( n13986 , n13985 , n5846 );
xor ( n13987 , n13982 , n13986 );
xor ( n13988 , n13973 , n13987 );
and ( n13989 , n13668 , n13672 );
and ( n13990 , n13672 , n13677 );
and ( n13991 , n13668 , n13677 );
or ( n13992 , n13989 , n13990 , n13991 );
and ( n13993 , n13647 , n4235 );
and ( n13994 , n13625 , n13628 );
and ( n13995 , n13628 , n13631 );
and ( n13996 , n13625 , n13631 );
or ( n13997 , n13994 , n13995 , n13996 );
buf ( n13998 , n13630 );
not ( n13999 , n7283 );
xor ( n14000 , n13998 , n13999 );
and ( n14001 , n7299 , n7274 );
xor ( n14002 , n14000 , n14001 );
xor ( n14003 , n13997 , n14002 );
and ( n14004 , n13632 , n13636 );
and ( n14005 , n13636 , n13641 );
and ( n14006 , n13632 , n13641 );
or ( n14007 , n14004 , n14005 , n14006 );
xor ( n14008 , n14003 , n14007 );
and ( n14009 , n13642 , n13643 );
xor ( n14010 , n14008 , n14009 );
buf ( n14011 , n14010 );
buf ( n14012 , n14011 );
buf ( n14013 , n14012 );
and ( n14014 , n14013 , n4232 );
nor ( n14015 , n13993 , n14014 );
xnor ( n14016 , n14015 , n4230 );
xor ( n14017 , n13992 , n14016 );
and ( n14018 , n7752 , n7356 );
and ( n14019 , n8179 , n6953 );
nor ( n14020 , n14018 , n14019 );
xnor ( n14021 , n14020 , n7352 );
and ( n14022 , n7324 , n7349 );
xor ( n14023 , n14021 , n14022 );
and ( n14024 , n13610 , n13611 );
xor ( n14025 , n14023 , n14024 );
and ( n14026 , n8640 , n6554 );
and ( n14027 , n9110 , n6205 );
nor ( n14028 , n14026 , n14027 );
xnor ( n14029 , n14028 , n6550 );
xor ( n14030 , n14025 , n14029 );
xor ( n14031 , n14017 , n14030 );
xor ( n14032 , n13988 , n14031 );
and ( n14033 , n13660 , n13679 );
and ( n14034 , n13679 , n13684 );
and ( n14035 , n13660 , n13684 );
or ( n14036 , n14033 , n14034 , n14035 );
xor ( n14037 , n14032 , n14036 );
xor ( n14038 , n13964 , n14037 );
xor ( n14039 , n13948 , n14038 );
and ( n14040 , n13687 , n13691 );
and ( n14041 , n13691 , n13696 );
and ( n14042 , n13687 , n13696 );
or ( n14043 , n14040 , n14041 , n14042 );
xor ( n14044 , n14039 , n14043 );
and ( n14045 , n13596 , n13697 );
and ( n14046 , n13698 , n13699 );
or ( n14047 , n14045 , n14046 );
xor ( n14048 , n14044 , n14047 );
buf ( n14049 , n14048 );
and ( n14050 , n13716 , n13720 );
and ( n14051 , n13720 , n13771 );
and ( n14052 , n13716 , n13771 );
or ( n14053 , n14050 , n14051 , n14052 );
and ( n14054 , n13739 , n13743 );
and ( n14055 , n13725 , n13729 );
and ( n14056 , n13729 , n13734 );
and ( n14057 , n13725 , n13734 );
or ( n14058 , n14055 , n14056 , n14057 );
and ( n14059 , n12976 , n4433 );
not ( n14060 , n14059 );
xnor ( n14061 , n14060 , n4441 );
and ( n14062 , n11398 , n4835 );
and ( n14063 , n11784 , n4648 );
nor ( n14064 , n14062 , n14063 );
xnor ( n14065 , n14064 , n4831 );
xor ( n14066 , n14061 , n14065 );
and ( n14067 , n9629 , n5922 );
and ( n14068 , n10072 , n5616 );
nor ( n14069 , n14067 , n14068 );
xnor ( n14070 , n14069 , n5918 );
xor ( n14071 , n14066 , n14070 );
xor ( n14072 , n14058 , n14071 );
and ( n14073 , n12217 , n4402 );
and ( n14074 , n12612 , n4391 );
nor ( n14075 , n14073 , n14074 );
xnor ( n14076 , n14075 , n4398 );
and ( n14077 , n10534 , n5323 );
and ( n14078 , n10940 , n5064 );
nor ( n14079 , n14077 , n14078 );
xnor ( n14080 , n14079 , n5319 );
xor ( n14081 , n14076 , n14080 );
and ( n14082 , n8728 , n6627 );
and ( n14083 , n9164 , n6272 );
nor ( n14084 , n14082 , n14083 );
xnor ( n14085 , n14084 , n6623 );
xor ( n14086 , n14081 , n14085 );
xor ( n14087 , n14072 , n14086 );
xor ( n14088 , n14054 , n14087 );
and ( n14089 , n13735 , n13744 );
and ( n14090 , n13744 , n13749 );
and ( n14091 , n13735 , n13749 );
or ( n14092 , n14089 , n14090 , n14091 );
xor ( n14093 , n14088 , n14092 );
and ( n14094 , n13750 , n13765 );
and ( n14095 , n13765 , n13770 );
and ( n14096 , n13750 , n13770 );
or ( n14097 , n14094 , n14095 , n14096 );
xor ( n14098 , n14093 , n14097 );
and ( n14099 , n13757 , n13758 );
and ( n14100 , n13758 , n13763 );
and ( n14101 , n13757 , n13763 );
or ( n14102 , n14099 , n14100 , n14101 );
or ( n14103 , n13755 , n13756 );
and ( n14104 , n7857 , n7444 );
and ( n14105 , n8303 , n7026 );
nor ( n14106 , n14104 , n14105 );
xnor ( n14107 , n14106 , n7440 );
xor ( n14108 , n14103 , n14107 );
and ( n14109 , n7417 , n7437 );
not ( n14110 , n14109 );
xor ( n14111 , n14108 , n14110 );
xor ( n14112 , n14102 , n14111 );
and ( n14113 , n13754 , n13764 );
xor ( n14114 , n14112 , n14113 );
and ( n14115 , n13709 , n13710 );
and ( n14116 , n13710 , n13715 );
and ( n14117 , n13709 , n13715 );
or ( n14118 , n14115 , n14116 , n14117 );
xor ( n14119 , n14114 , n14118 );
xor ( n14120 , n14098 , n14119 );
xor ( n14121 , n14053 , n14120 );
and ( n14122 , n13705 , n13772 );
and ( n14123 , n13772 , n13777 );
and ( n14124 , n13705 , n13777 );
or ( n14125 , n14122 , n14123 , n14124 );
xor ( n14126 , n14121 , n14125 );
and ( n14127 , n13778 , n13781 );
xor ( n14128 , n14126 , n14127 );
buf ( n14129 , n14128 );
not ( n14130 , n454 );
and ( n14131 , n14130 , n14049 );
and ( n14132 , n14129 , n454 );
or ( n14133 , n14131 , n14132 );
buf ( n14134 , n14133 );
buf ( n14135 , n14134 );
and ( n14136 , n14135 , n4505 );
xor ( n14137 , n13944 , n14136 );
and ( n14138 , n13058 , n5089 );
and ( n14139 , n13424 , n4866 );
xor ( n14140 , n14138 , n14139 );
and ( n14141 , n13789 , n4557 );
xor ( n14142 , n14140 , n14141 );
xor ( n14143 , n14137 , n14142 );
and ( n14144 , n13587 , n13588 );
and ( n14145 , n13588 , n13791 );
and ( n14146 , n13587 , n13791 );
or ( n14147 , n14144 , n14145 , n14146 );
xor ( n14148 , n14143 , n14147 );
and ( n14149 , n13792 , n13796 );
and ( n14150 , n13796 , n13801 );
and ( n14151 , n13792 , n13801 );
or ( n14152 , n14149 , n14150 , n14151 );
xor ( n14153 , n14148 , n14152 );
or ( n14154 , n13802 , n13803 );
xnor ( n14155 , n14153 , n14154 );
and ( n14156 , n13804 , n13805 );
xor ( n14157 , n14155 , n14156 );
buf ( n14158 , n14157 );
not ( n14159 , n4509 );
and ( n14160 , n14159 , n13940 );
and ( n14161 , n14158 , n4509 );
or ( n14162 , n14160 , n14161 );
and ( n14163 , n13874 , n13888 );
and ( n14164 , n13888 , n13925 );
and ( n14165 , n13874 , n13925 );
or ( n14166 , n14163 , n14164 , n14165 );
and ( n14167 , n13878 , n13882 );
and ( n14168 , n13882 , n13887 );
and ( n14169 , n13878 , n13887 );
or ( n14170 , n14167 , n14168 , n14169 );
and ( n14171 , n13893 , n13907 );
and ( n14172 , n13907 , n13924 );
and ( n14173 , n13893 , n13924 );
or ( n14174 , n14171 , n14172 , n14173 );
xor ( n14175 , n14170 , n14174 );
and ( n14176 , n13865 , n4524 );
and ( n14177 , n13834 , n13838 );
and ( n14178 , n13838 , n13840 );
and ( n14179 , n13834 , n13840 );
or ( n14180 , n14177 , n14178 , n14179 );
and ( n14181 , n13846 , n13847 );
and ( n14182 , n13847 , n13852 );
and ( n14183 , n13846 , n13852 );
or ( n14184 , n14181 , n14182 , n14183 );
xor ( n14185 , n14180 , n14184 );
and ( n14186 , n9848 , n7559 );
not ( n14187 , n14186 );
xnor ( n14188 , n14187 , n7555 );
not ( n14189 , n14188 );
and ( n14190 , n8900 , n8382 );
and ( n14191 , n9297 , n8042 );
nor ( n14192 , n14190 , n14191 );
xnor ( n14193 , n14192 , n8378 );
xor ( n14194 , n14189 , n14193 );
and ( n14195 , n8409 , n8375 );
xor ( n14196 , n14194 , n14195 );
xor ( n14197 , n14185 , n14196 );
and ( n14198 , n13833 , n13841 );
and ( n14199 , n13841 , n13853 );
and ( n14200 , n13833 , n13853 );
or ( n14201 , n14198 , n14199 , n14200 );
xor ( n14202 , n14197 , n14201 );
and ( n14203 , n13829 , n13854 );
and ( n14204 , n13854 , n13859 );
and ( n14205 , n13829 , n13859 );
or ( n14206 , n14203 , n14204 , n14205 );
xor ( n14207 , n14202 , n14206 );
and ( n14208 , n13860 , n13861 );
xor ( n14209 , n14207 , n14208 );
buf ( n14210 , n14209 );
buf ( n14211 , n14210 );
buf ( n14212 , n14211 );
and ( n14213 , n14212 , n4145 );
nor ( n14214 , n14176 , n14213 );
xnor ( n14215 , n14214 , n4521 );
xor ( n14216 , n14175 , n14215 );
xor ( n14217 , n14166 , n14216 );
and ( n14218 , n13819 , n13823 );
and ( n14219 , n13823 , n13868 );
and ( n14220 , n13819 , n13868 );
or ( n14221 , n14218 , n14219 , n14220 );
and ( n14222 , n12392 , n5441 );
and ( n14223 , n12754 , n5161 );
nor ( n14224 , n14222 , n14223 );
xnor ( n14225 , n14224 , n5437 );
and ( n14226 , n11569 , n6068 );
and ( n14227 , n11989 , n5730 );
nor ( n14228 , n14226 , n14227 );
xnor ( n14229 , n14228 , n6064 );
xor ( n14230 , n14225 , n14229 );
and ( n14231 , n8057 , n9407 );
and ( n14232 , n8462 , n8872 );
nor ( n14233 , n14231 , n14232 );
xnor ( n14234 , n14233 , n9403 );
and ( n14235 , n7146 , n10329 );
and ( n14236 , n7587 , n9791 );
nor ( n14237 , n14235 , n14236 );
not ( n14238 , n14237 );
xor ( n14239 , n14234 , n14238 );
and ( n14240 , n13912 , n13916 );
xor ( n14241 , n14239 , n14240 );
and ( n14242 , n8968 , n8502 );
and ( n14243 , n9367 , n7970 );
nor ( n14244 , n14242 , n14243 );
xnor ( n14245 , n14244 , n8498 );
xor ( n14246 , n14241 , n14245 );
xor ( n14247 , n14230 , n14246 );
xor ( n14248 , n14221 , n14247 );
and ( n14249 , n13897 , n13901 );
and ( n14250 , n13901 , n13906 );
and ( n14251 , n13897 , n13906 );
or ( n14252 , n14249 , n14250 , n14251 );
and ( n14253 , n13144 , n4938 );
and ( n14254 , n13506 , n4711 );
nor ( n14255 , n14253 , n14254 );
xnor ( n14256 , n14255 , n4934 );
xor ( n14257 , n14252 , n14256 );
and ( n14258 , n13917 , n13918 );
and ( n14259 , n13918 , n13923 );
and ( n14260 , n13917 , n13923 );
or ( n14261 , n14258 , n14259 , n14260 );
and ( n14262 , n10706 , n6711 );
and ( n14263 , n11163 , n6332 );
nor ( n14264 , n14262 , n14263 );
xnor ( n14265 , n14264 , n6707 );
xor ( n14266 , n14261 , n14265 );
and ( n14267 , n9885 , n7630 );
and ( n14268 , n10287 , n7188 );
nor ( n14269 , n14267 , n14268 );
xnor ( n14270 , n14269 , n7626 );
xor ( n14271 , n14266 , n14270 );
xor ( n14272 , n14257 , n14271 );
xor ( n14273 , n14248 , n14272 );
xor ( n14274 , n14217 , n14273 );
and ( n14275 , n13815 , n13869 );
and ( n14276 , n13869 , n13926 );
and ( n14277 , n13815 , n13926 );
or ( n14278 , n14275 , n14276 , n14277 );
xor ( n14279 , n14274 , n14278 );
and ( n14280 , n13927 , n13931 );
and ( n14281 , n13931 , n13936 );
and ( n14282 , n13927 , n13936 );
or ( n14283 , n14280 , n14281 , n14282 );
xor ( n14284 , n14279 , n14283 );
and ( n14285 , n13937 , n13938 );
xor ( n14286 , n14284 , n14285 );
buf ( n14287 , n14286 );
and ( n14288 , n13424 , n5089 );
and ( n14289 , n13789 , n4866 );
xor ( n14290 , n14288 , n14289 );
and ( n14291 , n13968 , n13972 );
and ( n14292 , n13972 , n13987 );
and ( n14293 , n13968 , n13987 );
or ( n14294 , n14291 , n14292 , n14293 );
and ( n14295 , n14023 , n14024 );
and ( n14296 , n14024 , n14029 );
and ( n14297 , n14023 , n14029 );
or ( n14298 , n14295 , n14296 , n14297 );
and ( n14299 , n13313 , n4319 );
and ( n14300 , n13647 , n4310 );
nor ( n14301 , n14299 , n14300 );
xnor ( n14302 , n14301 , n4315 );
xor ( n14303 , n14298 , n14302 );
and ( n14304 , n11702 , n4788 );
and ( n14305 , n12116 , n4611 );
nor ( n14306 , n14304 , n14305 );
xnor ( n14307 , n14306 , n4784 );
xor ( n14308 , n14303 , n14307 );
xor ( n14309 , n14294 , n14308 );
and ( n14310 , n14013 , n4235 );
not ( n14311 , n14310 );
xnor ( n14312 , n14311 , n4230 );
and ( n14313 , n8179 , n7356 );
and ( n14314 , n8640 , n6953 );
nor ( n14315 , n14313 , n14314 );
xnor ( n14316 , n14315 , n7352 );
and ( n14317 , n7752 , n7349 );
xor ( n14318 , n14316 , n14317 );
and ( n14319 , n14021 , n14022 );
xor ( n14320 , n14318 , n14319 );
and ( n14321 , n9110 , n6554 );
and ( n14322 , n9583 , n6205 );
nor ( n14323 , n14321 , n14322 );
xnor ( n14324 , n14323 , n6550 );
xor ( n14325 , n14320 , n14324 );
xor ( n14326 , n14312 , n14325 );
xor ( n14327 , n14309 , n14326 );
and ( n14328 , n13959 , n13963 );
and ( n14329 , n13963 , n14037 );
and ( n14330 , n13959 , n14037 );
or ( n14331 , n14328 , n14329 , n14330 );
xor ( n14332 , n14327 , n14331 );
and ( n14333 , n13952 , n13953 );
and ( n14334 , n13953 , n13958 );
and ( n14335 , n13952 , n13958 );
or ( n14336 , n14333 , n14334 , n14335 );
and ( n14337 , n13977 , n13981 );
and ( n14338 , n13981 , n13986 );
and ( n14339 , n13977 , n13986 );
or ( n14340 , n14337 , n14338 , n14339 );
and ( n14341 , n13992 , n14016 );
and ( n14342 , n14016 , n14030 );
and ( n14343 , n13992 , n14030 );
or ( n14344 , n14341 , n14342 , n14343 );
xor ( n14345 , n14340 , n14344 );
and ( n14346 , n12527 , n4298 );
and ( n14347 , n12895 , n4287 );
nor ( n14348 , n14346 , n14347 );
xnor ( n14349 , n14348 , n4294 );
and ( n14350 , n10857 , n5270 );
and ( n14351 , n11295 , n5021 );
nor ( n14352 , n14350 , n14351 );
xnor ( n14353 , n14352 , n5266 );
xor ( n14354 , n14349 , n14353 );
and ( n14355 , n9989 , n5850 );
and ( n14356 , n10437 , n5566 );
nor ( n14357 , n14355 , n14356 );
xnor ( n14358 , n14357 , n5846 );
xor ( n14359 , n14354 , n14358 );
xor ( n14360 , n14345 , n14359 );
xor ( n14361 , n14336 , n14360 );
and ( n14362 , n13988 , n14031 );
and ( n14363 , n14031 , n14036 );
and ( n14364 , n13988 , n14036 );
or ( n14365 , n14362 , n14363 , n14364 );
xor ( n14366 , n14361 , n14365 );
xor ( n14367 , n14332 , n14366 );
and ( n14368 , n13948 , n14038 );
and ( n14369 , n14038 , n14043 );
and ( n14370 , n13948 , n14043 );
or ( n14371 , n14368 , n14369 , n14370 );
xor ( n14372 , n14367 , n14371 );
and ( n14373 , n14044 , n14047 );
xor ( n14374 , n14372 , n14373 );
buf ( n14375 , n14374 );
and ( n14376 , n14061 , n14065 );
and ( n14377 , n14065 , n14070 );
and ( n14378 , n14061 , n14070 );
or ( n14379 , n14376 , n14377 , n14378 );
and ( n14380 , n11784 , n4835 );
and ( n14381 , n12217 , n4648 );
nor ( n14382 , n14380 , n14381 );
xnor ( n14383 , n14382 , n4831 );
and ( n14384 , n10072 , n5922 );
and ( n14385 , n10534 , n5616 );
nor ( n14386 , n14384 , n14385 );
xnor ( n14387 , n14386 , n5918 );
xor ( n14388 , n14383 , n14387 );
and ( n14389 , n9164 , n6627 );
and ( n14390 , n9629 , n6272 );
nor ( n14391 , n14389 , n14390 );
xnor ( n14392 , n14391 , n6623 );
xor ( n14393 , n14388 , n14392 );
xor ( n14394 , n14379 , n14393 );
and ( n14395 , n12612 , n4402 );
and ( n14396 , n12976 , n4391 );
nor ( n14397 , n14395 , n14396 );
xnor ( n14398 , n14397 , n4398 );
and ( n14399 , n10940 , n5323 );
and ( n14400 , n11398 , n5064 );
nor ( n14401 , n14399 , n14400 );
xnor ( n14402 , n14401 , n5319 );
xor ( n14403 , n14398 , n14402 );
and ( n14404 , n8303 , n7444 );
and ( n14405 , n8728 , n7026 );
nor ( n14406 , n14404 , n14405 );
xnor ( n14407 , n14406 , n7440 );
xor ( n14408 , n14403 , n14407 );
xor ( n14409 , n14394 , n14408 );
and ( n14410 , n14058 , n14071 );
and ( n14411 , n14071 , n14086 );
and ( n14412 , n14058 , n14086 );
or ( n14413 , n14410 , n14411 , n14412 );
xor ( n14414 , n14409 , n14413 );
and ( n14415 , n14102 , n14111 );
xor ( n14416 , n14414 , n14415 );
and ( n14417 , n14093 , n14097 );
and ( n14418 , n14097 , n14119 );
and ( n14419 , n14093 , n14119 );
or ( n14420 , n14417 , n14418 , n14419 );
xor ( n14421 , n14416 , n14420 );
and ( n14422 , n14054 , n14087 );
and ( n14423 , n14087 , n14092 );
and ( n14424 , n14054 , n14092 );
or ( n14425 , n14422 , n14423 , n14424 );
and ( n14426 , n14076 , n14080 );
and ( n14427 , n14080 , n14085 );
and ( n14428 , n14076 , n14085 );
or ( n14429 , n14426 , n14427 , n14428 );
and ( n14430 , n14103 , n14107 );
and ( n14431 , n14107 , n14110 );
and ( n14432 , n14103 , n14110 );
or ( n14433 , n14430 , n14431 , n14432 );
xor ( n14434 , n14429 , n14433 );
buf ( n14435 , n14109 );
not ( n14436 , n4441 );
xor ( n14437 , n14435 , n14436 );
and ( n14438 , n7857 , n7437 );
xor ( n14439 , n14437 , n14438 );
xor ( n14440 , n14434 , n14439 );
xor ( n14441 , n14425 , n14440 );
and ( n14442 , n14112 , n14113 );
and ( n14443 , n14113 , n14118 );
and ( n14444 , n14112 , n14118 );
or ( n14445 , n14442 , n14443 , n14444 );
xor ( n14446 , n14441 , n14445 );
xor ( n14447 , n14421 , n14446 );
and ( n14448 , n14053 , n14120 );
and ( n14449 , n14120 , n14125 );
and ( n14450 , n14053 , n14125 );
or ( n14451 , n14448 , n14449 , n14450 );
xor ( n14452 , n14447 , n14451 );
and ( n14453 , n14126 , n14127 );
xor ( n14454 , n14452 , n14453 );
buf ( n14455 , n14454 );
not ( n14456 , n454 );
and ( n14457 , n14456 , n14375 );
and ( n14458 , n14455 , n454 );
or ( n14459 , n14457 , n14458 );
buf ( n14460 , n14459 );
buf ( n14461 , n14460 );
and ( n14462 , n14461 , n4505 );
xor ( n14463 , n14290 , n14462 );
and ( n14464 , n14138 , n14139 );
and ( n14465 , n14139 , n14141 );
and ( n14466 , n14138 , n14141 );
or ( n14467 , n14464 , n14465 , n14466 );
and ( n14468 , n14135 , n4557 );
xor ( n14469 , n14467 , n14468 );
xor ( n14470 , n14463 , n14469 );
and ( n14471 , n13944 , n14136 );
and ( n14472 , n14136 , n14142 );
and ( n14473 , n13944 , n14142 );
or ( n14474 , n14471 , n14472 , n14473 );
xor ( n14475 , n14470 , n14474 );
and ( n14476 , n14143 , n14147 );
and ( n14477 , n14147 , n14152 );
and ( n14478 , n14143 , n14152 );
or ( n14479 , n14476 , n14477 , n14478 );
xor ( n14480 , n14475 , n14479 );
or ( n14481 , n14153 , n14154 );
xor ( n14482 , n14480 , n14481 );
not ( n14483 , n14482 );
and ( n14484 , n14155 , n14156 );
xor ( n14485 , n14483 , n14484 );
buf ( n14486 , n14485 );
not ( n14487 , n4509 );
and ( n14488 , n14487 , n14287 );
and ( n14489 , n14486 , n4509 );
or ( n14490 , n14488 , n14489 );
and ( n14491 , n14221 , n14247 );
and ( n14492 , n14247 , n14272 );
and ( n14493 , n14221 , n14272 );
or ( n14494 , n14491 , n14492 , n14493 );
and ( n14495 , n14225 , n14229 );
and ( n14496 , n14229 , n14246 );
and ( n14497 , n14225 , n14246 );
or ( n14498 , n14495 , n14496 , n14497 );
and ( n14499 , n14252 , n14256 );
and ( n14500 , n14256 , n14271 );
and ( n14501 , n14252 , n14271 );
or ( n14502 , n14499 , n14500 , n14501 );
xor ( n14503 , n14498 , n14502 );
and ( n14504 , n14239 , n14240 );
and ( n14505 , n14240 , n14245 );
and ( n14506 , n14239 , n14245 );
or ( n14507 , n14504 , n14505 , n14506 );
and ( n14508 , n11163 , n6711 );
and ( n14509 , n11569 , n6332 );
nor ( n14510 , n14508 , n14509 );
xnor ( n14511 , n14510 , n6707 );
xor ( n14512 , n14507 , n14511 );
and ( n14513 , n10287 , n7630 );
and ( n14514 , n10706 , n7188 );
nor ( n14515 , n14513 , n14514 );
xnor ( n14516 , n14515 , n7626 );
xor ( n14517 , n14512 , n14516 );
xor ( n14518 , n14503 , n14517 );
xor ( n14519 , n14494 , n14518 );
and ( n14520 , n14170 , n14174 );
and ( n14521 , n14174 , n14215 );
and ( n14522 , n14170 , n14215 );
or ( n14523 , n14520 , n14521 , n14522 );
and ( n14524 , n14261 , n14265 );
and ( n14525 , n14265 , n14270 );
and ( n14526 , n14261 , n14270 );
or ( n14527 , n14524 , n14525 , n14526 );
and ( n14528 , n14212 , n4524 );
and ( n14529 , n14189 , n14193 );
and ( n14530 , n14193 , n14195 );
and ( n14531 , n14189 , n14195 );
or ( n14532 , n14529 , n14530 , n14531 );
buf ( n14533 , n14188 );
xor ( n14534 , n14532 , n14533 );
not ( n14535 , n7555 );
and ( n14536 , n9297 , n8382 );
and ( n14537 , n9848 , n8042 );
nor ( n14538 , n14536 , n14537 );
xnor ( n14539 , n14538 , n8378 );
xor ( n14540 , n14535 , n14539 );
and ( n14541 , n8900 , n8375 );
xor ( n14542 , n14540 , n14541 );
xor ( n14543 , n14534 , n14542 );
and ( n14544 , n14180 , n14184 );
and ( n14545 , n14184 , n14196 );
and ( n14546 , n14180 , n14196 );
or ( n14547 , n14544 , n14545 , n14546 );
xor ( n14548 , n14543 , n14547 );
and ( n14549 , n14197 , n14201 );
and ( n14550 , n14201 , n14206 );
and ( n14551 , n14197 , n14206 );
or ( n14552 , n14549 , n14550 , n14551 );
xor ( n14553 , n14548 , n14552 );
and ( n14554 , n14207 , n14208 );
xor ( n14555 , n14553 , n14554 );
buf ( n14556 , n14555 );
buf ( n14557 , n14556 );
buf ( n14558 , n14557 );
and ( n14559 , n14558 , n4145 );
nor ( n14560 , n14528 , n14559 );
xnor ( n14561 , n14560 , n4521 );
xor ( n14562 , n14527 , n14561 );
and ( n14563 , n13506 , n4938 );
and ( n14564 , n13865 , n4711 );
nor ( n14565 , n14563 , n14564 );
xnor ( n14566 , n14565 , n4934 );
xor ( n14567 , n14562 , n14566 );
xor ( n14568 , n14523 , n14567 );
and ( n14569 , n12754 , n5441 );
and ( n14570 , n13144 , n5161 );
nor ( n14571 , n14569 , n14570 );
xnor ( n14572 , n14571 , n5437 );
and ( n14573 , n11989 , n6068 );
and ( n14574 , n12392 , n5730 );
nor ( n14575 , n14573 , n14574 );
xnor ( n14576 , n14575 , n6064 );
xor ( n14577 , n14572 , n14576 );
and ( n14578 , n8462 , n9407 );
and ( n14579 , n8968 , n8872 );
nor ( n14580 , n14578 , n14579 );
xnor ( n14581 , n14580 , n9403 );
and ( n14582 , n7587 , n10329 );
and ( n14583 , n8057 , n9791 );
nor ( n14584 , n14582 , n14583 );
not ( n14585 , n14584 );
xor ( n14586 , n14581 , n14585 );
and ( n14587 , n14234 , n14238 );
xor ( n14588 , n14586 , n14587 );
and ( n14589 , n9367 , n8502 );
and ( n14590 , n9885 , n7970 );
nor ( n14591 , n14589 , n14590 );
xnor ( n14592 , n14591 , n8498 );
xor ( n14593 , n14588 , n14592 );
xor ( n14594 , n14577 , n14593 );
xor ( n14595 , n14568 , n14594 );
xor ( n14596 , n14519 , n14595 );
and ( n14597 , n14166 , n14216 );
and ( n14598 , n14216 , n14273 );
and ( n14599 , n14166 , n14273 );
or ( n14600 , n14597 , n14598 , n14599 );
xor ( n14601 , n14596 , n14600 );
and ( n14602 , n14274 , n14278 );
and ( n14603 , n14278 , n14283 );
and ( n14604 , n14274 , n14283 );
or ( n14605 , n14602 , n14603 , n14604 );
xor ( n14606 , n14601 , n14605 );
and ( n14607 , n14284 , n14285 );
xor ( n14608 , n14606 , n14607 );
buf ( n14609 , n14608 );
and ( n14610 , n14467 , n14468 );
and ( n14611 , n14349 , n14353 );
and ( n14612 , n14353 , n14358 );
and ( n14613 , n14349 , n14358 );
or ( n14614 , n14611 , n14612 , n14613 );
and ( n14615 , n14318 , n14319 );
and ( n14616 , n14319 , n14324 );
and ( n14617 , n14318 , n14324 );
or ( n14618 , n14615 , n14616 , n14617 );
xor ( n14619 , n14614 , n14618 );
not ( n14620 , n4230 );
and ( n14621 , n8179 , n7349 );
xnor ( n14622 , n14620 , n14621 );
and ( n14623 , n14316 , n14317 );
xor ( n14624 , n14622 , n14623 );
and ( n14625 , n8640 , n7356 );
and ( n14626 , n9110 , n6953 );
nor ( n14627 , n14625 , n14626 );
xnor ( n14628 , n14627 , n7352 );
xor ( n14629 , n14624 , n14628 );
xor ( n14630 , n14619 , n14629 );
and ( n14631 , n14312 , n14325 );
xor ( n14632 , n14630 , n14631 );
and ( n14633 , n14298 , n14302 );
and ( n14634 , n14302 , n14307 );
and ( n14635 , n14298 , n14307 );
or ( n14636 , n14633 , n14634 , n14635 );
and ( n14637 , n12116 , n4788 );
and ( n14638 , n12527 , n4611 );
nor ( n14639 , n14637 , n14638 );
xnor ( n14640 , n14639 , n4784 );
and ( n14641 , n10437 , n5850 );
and ( n14642 , n10857 , n5566 );
nor ( n14643 , n14641 , n14642 );
xnor ( n14644 , n14643 , n5846 );
xor ( n14645 , n14640 , n14644 );
and ( n14646 , n9583 , n6554 );
and ( n14647 , n9989 , n6205 );
nor ( n14648 , n14646 , n14647 );
xnor ( n14649 , n14648 , n6550 );
xor ( n14650 , n14645 , n14649 );
xor ( n14651 , n14636 , n14650 );
and ( n14652 , n13647 , n4319 );
and ( n14653 , n14013 , n4310 );
nor ( n14654 , n14652 , n14653 );
xnor ( n14655 , n14654 , n4315 );
and ( n14656 , n12895 , n4298 );
and ( n14657 , n13313 , n4287 );
nor ( n14658 , n14656 , n14657 );
xnor ( n14659 , n14658 , n4294 );
xor ( n14660 , n14655 , n14659 );
and ( n14661 , n11295 , n5270 );
and ( n14662 , n11702 , n5021 );
nor ( n14663 , n14661 , n14662 );
xnor ( n14664 , n14663 , n5266 );
xor ( n14665 , n14660 , n14664 );
xor ( n14666 , n14651 , n14665 );
xor ( n14667 , n14632 , n14666 );
and ( n14668 , n14327 , n14331 );
and ( n14669 , n14331 , n14366 );
and ( n14670 , n14327 , n14366 );
or ( n14671 , n14668 , n14669 , n14670 );
xor ( n14672 , n14667 , n14671 );
and ( n14673 , n14340 , n14344 );
and ( n14674 , n14344 , n14359 );
and ( n14675 , n14340 , n14359 );
or ( n14676 , n14673 , n14674 , n14675 );
and ( n14677 , n14294 , n14308 );
and ( n14678 , n14308 , n14326 );
and ( n14679 , n14294 , n14326 );
or ( n14680 , n14677 , n14678 , n14679 );
xor ( n14681 , n14676 , n14680 );
and ( n14682 , n14336 , n14360 );
and ( n14683 , n14360 , n14365 );
and ( n14684 , n14336 , n14365 );
or ( n14685 , n14682 , n14683 , n14684 );
xor ( n14686 , n14681 , n14685 );
xor ( n14687 , n14672 , n14686 );
and ( n14688 , n14367 , n14371 );
and ( n14689 , n14372 , n14373 );
or ( n14690 , n14688 , n14689 );
xor ( n14691 , n14687 , n14690 );
buf ( n14692 , n14691 );
and ( n14693 , n14425 , n14440 );
and ( n14694 , n14440 , n14445 );
and ( n14695 , n14425 , n14445 );
or ( n14696 , n14693 , n14694 , n14695 );
and ( n14697 , n14416 , n14420 );
and ( n14698 , n14420 , n14446 );
and ( n14699 , n14416 , n14446 );
or ( n14700 , n14697 , n14698 , n14699 );
xor ( n14701 , n14696 , n14700 );
and ( n14702 , n14409 , n14413 );
and ( n14703 , n14413 , n14415 );
and ( n14704 , n14409 , n14415 );
or ( n14705 , n14702 , n14703 , n14704 );
and ( n14706 , n14398 , n14402 );
and ( n14707 , n14402 , n14407 );
and ( n14708 , n14398 , n14407 );
or ( n14709 , n14706 , n14707 , n14708 );
and ( n14710 , n14435 , n14436 );
and ( n14711 , n14436 , n14438 );
and ( n14712 , n14435 , n14438 );
or ( n14713 , n14710 , n14711 , n14712 );
and ( n14714 , n10534 , n5922 );
and ( n14715 , n10940 , n5616 );
nor ( n14716 , n14714 , n14715 );
xnor ( n14717 , n14716 , n5918 );
xor ( n14718 , n14713 , n14717 );
and ( n14719 , n9629 , n6627 );
and ( n14720 , n10072 , n6272 );
nor ( n14721 , n14719 , n14720 );
xnor ( n14722 , n14721 , n6623 );
xor ( n14723 , n14718 , n14722 );
xor ( n14724 , n14709 , n14723 );
and ( n14725 , n12217 , n4835 );
and ( n14726 , n12612 , n4648 );
nor ( n14727 , n14725 , n14726 );
xnor ( n14728 , n14727 , n4831 );
and ( n14729 , n8728 , n7444 );
and ( n14730 , n9164 , n7026 );
nor ( n14731 , n14729 , n14730 );
xnor ( n14732 , n14731 , n7440 );
xor ( n14733 , n14728 , n14732 );
and ( n14734 , n8303 , n7437 );
not ( n14735 , n14734 );
xor ( n14736 , n14733 , n14735 );
xor ( n14737 , n14724 , n14736 );
xor ( n14738 , n14705 , n14737 );
and ( n14739 , n14379 , n14393 );
and ( n14740 , n14393 , n14408 );
and ( n14741 , n14379 , n14408 );
or ( n14742 , n14739 , n14740 , n14741 );
and ( n14743 , n14429 , n14433 );
and ( n14744 , n14433 , n14439 );
and ( n14745 , n14429 , n14439 );
or ( n14746 , n14743 , n14744 , n14745 );
xor ( n14747 , n14742 , n14746 );
and ( n14748 , n14383 , n14387 );
and ( n14749 , n14387 , n14392 );
and ( n14750 , n14383 , n14392 );
or ( n14751 , n14748 , n14749 , n14750 );
and ( n14752 , n12976 , n4402 );
not ( n14753 , n14752 );
xnor ( n14754 , n14753 , n4398 );
xor ( n14755 , n14751 , n14754 );
and ( n14756 , n11398 , n5323 );
and ( n14757 , n11784 , n5064 );
nor ( n14758 , n14756 , n14757 );
xnor ( n14759 , n14758 , n5319 );
xor ( n14760 , n14755 , n14759 );
xor ( n14761 , n14747 , n14760 );
xor ( n14762 , n14738 , n14761 );
xor ( n14763 , n14701 , n14762 );
and ( n14764 , n14447 , n14451 );
and ( n14765 , n14452 , n14453 );
or ( n14766 , n14764 , n14765 );
xor ( n14767 , n14763 , n14766 );
buf ( n14768 , n14767 );
not ( n14769 , n454 );
and ( n14770 , n14769 , n14692 );
and ( n14771 , n14768 , n454 );
or ( n14772 , n14770 , n14771 );
buf ( n14773 , n14772 );
buf ( n14774 , n14773 );
and ( n14775 , n14774 , n4505 );
and ( n14776 , n14288 , n14289 );
and ( n14777 , n14289 , n14462 );
and ( n14778 , n14288 , n14462 );
or ( n14779 , n14776 , n14777 , n14778 );
xor ( n14780 , n14775 , n14779 );
and ( n14781 , n13789 , n5089 );
and ( n14782 , n14135 , n4866 );
xor ( n14783 , n14781 , n14782 );
and ( n14784 , n14461 , n4557 );
xor ( n14785 , n14783 , n14784 );
xor ( n14786 , n14780 , n14785 );
xor ( n14787 , n14610 , n14786 );
and ( n14788 , n14463 , n14469 );
and ( n14789 , n14469 , n14474 );
and ( n14790 , n14463 , n14474 );
or ( n14791 , n14788 , n14789 , n14790 );
xor ( n14792 , n14787 , n14791 );
and ( n14793 , n14475 , n14479 );
and ( n14794 , n14479 , n14481 );
and ( n14795 , n14475 , n14481 );
or ( n14796 , n14793 , n14794 , n14795 );
xnor ( n14797 , n14792 , n14796 );
and ( n14798 , n14483 , n14484 );
or ( n14799 , n14482 , n14798 );
xor ( n14800 , n14797 , n14799 );
buf ( n14801 , n14800 );
not ( n14802 , n4509 );
and ( n14803 , n14802 , n14609 );
and ( n14804 , n14801 , n4509 );
or ( n14805 , n14803 , n14804 );
and ( n14806 , n14523 , n14567 );
and ( n14807 , n14567 , n14594 );
and ( n14808 , n14523 , n14594 );
or ( n14809 , n14806 , n14807 , n14808 );
and ( n14810 , n14527 , n14561 );
and ( n14811 , n14561 , n14566 );
and ( n14812 , n14527 , n14566 );
or ( n14813 , n14810 , n14811 , n14812 );
and ( n14814 , n14572 , n14576 );
and ( n14815 , n14576 , n14593 );
and ( n14816 , n14572 , n14593 );
or ( n14817 , n14814 , n14815 , n14816 );
xor ( n14818 , n14813 , n14817 );
and ( n14819 , n14586 , n14587 );
and ( n14820 , n14587 , n14592 );
and ( n14821 , n14586 , n14592 );
or ( n14822 , n14819 , n14820 , n14821 );
and ( n14823 , n11569 , n6711 );
and ( n14824 , n11989 , n6332 );
nor ( n14825 , n14823 , n14824 );
xnor ( n14826 , n14825 , n6707 );
xor ( n14827 , n14822 , n14826 );
and ( n14828 , n10706 , n7630 );
and ( n14829 , n11163 , n7188 );
nor ( n14830 , n14828 , n14829 );
xnor ( n14831 , n14830 , n7626 );
xor ( n14832 , n14827 , n14831 );
xor ( n14833 , n14818 , n14832 );
xor ( n14834 , n14809 , n14833 );
and ( n14835 , n14498 , n14502 );
and ( n14836 , n14502 , n14517 );
and ( n14837 , n14498 , n14517 );
or ( n14838 , n14835 , n14836 , n14837 );
and ( n14839 , n14558 , n4524 );
and ( n14840 , n14535 , n14539 );
and ( n14841 , n14539 , n14541 );
and ( n14842 , n14535 , n14541 );
or ( n14843 , n14840 , n14841 , n14842 );
and ( n14844 , n9848 , n8382 );
not ( n14845 , n14844 );
xnor ( n14846 , n14845 , n8378 );
not ( n14847 , n14846 );
xor ( n14848 , n14843 , n14847 );
and ( n14849 , n9297 , n8375 );
xor ( n14850 , n14848 , n14849 );
and ( n14851 , n14532 , n14533 );
and ( n14852 , n14533 , n14542 );
and ( n14853 , n14532 , n14542 );
or ( n14854 , n14851 , n14852 , n14853 );
xor ( n14855 , n14850 , n14854 );
and ( n14856 , n14543 , n14547 );
and ( n14857 , n14547 , n14552 );
and ( n14858 , n14543 , n14552 );
or ( n14859 , n14856 , n14857 , n14858 );
xor ( n14860 , n14855 , n14859 );
and ( n14861 , n14553 , n14554 );
xor ( n14862 , n14860 , n14861 );
buf ( n14863 , n14862 );
buf ( n14864 , n14863 );
buf ( n14865 , n14864 );
and ( n14866 , n14865 , n4145 );
nor ( n14867 , n14839 , n14866 );
xnor ( n14868 , n14867 , n4521 );
and ( n14869 , n13865 , n4938 );
and ( n14870 , n14212 , n4711 );
nor ( n14871 , n14869 , n14870 );
xnor ( n14872 , n14871 , n4934 );
xor ( n14873 , n14868 , n14872 );
and ( n14874 , n12392 , n6068 );
and ( n14875 , n12754 , n5730 );
nor ( n14876 , n14874 , n14875 );
xnor ( n14877 , n14876 , n6064 );
xor ( n14878 , n14873 , n14877 );
xor ( n14879 , n14838 , n14878 );
and ( n14880 , n14507 , n14511 );
and ( n14881 , n14511 , n14516 );
and ( n14882 , n14507 , n14516 );
or ( n14883 , n14880 , n14881 , n14882 );
and ( n14884 , n13144 , n5441 );
and ( n14885 , n13506 , n5161 );
nor ( n14886 , n14884 , n14885 );
xnor ( n14887 , n14886 , n5437 );
xor ( n14888 , n14883 , n14887 );
and ( n14889 , n8968 , n9407 );
and ( n14890 , n9367 , n8872 );
nor ( n14891 , n14889 , n14890 );
xnor ( n14892 , n14891 , n9403 );
and ( n14893 , n8057 , n10329 );
and ( n14894 , n8462 , n9791 );
nor ( n14895 , n14893 , n14894 );
not ( n14896 , n14895 );
xor ( n14897 , n14892 , n14896 );
and ( n14898 , n14581 , n14585 );
xor ( n14899 , n14897 , n14898 );
and ( n14900 , n9885 , n8502 );
and ( n14901 , n10287 , n7970 );
nor ( n14902 , n14900 , n14901 );
xnor ( n14903 , n14902 , n8498 );
xor ( n14904 , n14899 , n14903 );
xor ( n14905 , n14888 , n14904 );
xor ( n14906 , n14879 , n14905 );
xor ( n14907 , n14834 , n14906 );
and ( n14908 , n14494 , n14518 );
and ( n14909 , n14518 , n14595 );
and ( n14910 , n14494 , n14595 );
or ( n14911 , n14908 , n14909 , n14910 );
xor ( n14912 , n14907 , n14911 );
and ( n14913 , n14596 , n14600 );
and ( n14914 , n14600 , n14605 );
and ( n14915 , n14596 , n14605 );
or ( n14916 , n14913 , n14914 , n14915 );
xor ( n14917 , n14912 , n14916 );
and ( n14918 , n14606 , n14607 );
xor ( n14919 , n14917 , n14918 );
buf ( n14920 , n14919 );
and ( n14921 , n14775 , n14779 );
and ( n14922 , n14779 , n14785 );
and ( n14923 , n14775 , n14785 );
or ( n14924 , n14921 , n14922 , n14923 );
and ( n14925 , n14135 , n5089 );
and ( n14926 , n14461 , n4866 );
xor ( n14927 , n14925 , n14926 );
and ( n14928 , n14676 , n14680 );
and ( n14929 , n14680 , n14685 );
and ( n14930 , n14676 , n14685 );
or ( n14931 , n14928 , n14929 , n14930 );
and ( n14932 , n14640 , n14644 );
and ( n14933 , n14644 , n14649 );
and ( n14934 , n14640 , n14649 );
or ( n14935 , n14932 , n14933 , n14934 );
and ( n14936 , n14655 , n14659 );
and ( n14937 , n14659 , n14664 );
and ( n14938 , n14655 , n14664 );
or ( n14939 , n14936 , n14937 , n14938 );
xor ( n14940 , n14935 , n14939 );
and ( n14941 , n14013 , n4319 );
not ( n14942 , n14941 );
xnor ( n14943 , n14942 , n4315 );
and ( n14944 , n13313 , n4298 );
and ( n14945 , n13647 , n4287 );
nor ( n14946 , n14944 , n14945 );
xnor ( n14947 , n14946 , n4294 );
xor ( n14948 , n14943 , n14947 );
and ( n14949 , n11702 , n5270 );
and ( n14950 , n12116 , n5021 );
nor ( n14951 , n14949 , n14950 );
xnor ( n14952 , n14951 , n5266 );
xor ( n14953 , n14948 , n14952 );
xor ( n14954 , n14940 , n14953 );
and ( n14955 , n14614 , n14618 );
and ( n14956 , n14618 , n14629 );
and ( n14957 , n14614 , n14629 );
or ( n14958 , n14955 , n14956 , n14957 );
and ( n14959 , n14636 , n14650 );
and ( n14960 , n14650 , n14665 );
and ( n14961 , n14636 , n14665 );
or ( n14962 , n14959 , n14960 , n14961 );
xor ( n14963 , n14958 , n14962 );
and ( n14964 , n14622 , n14623 );
and ( n14965 , n14623 , n14628 );
and ( n14966 , n14622 , n14628 );
or ( n14967 , n14964 , n14965 , n14966 );
and ( n14968 , n12527 , n4788 );
and ( n14969 , n12895 , n4611 );
nor ( n14970 , n14968 , n14969 );
xnor ( n14971 , n14970 , n4784 );
and ( n14972 , n10857 , n5850 );
and ( n14973 , n11295 , n5566 );
nor ( n14974 , n14972 , n14973 );
xnor ( n14975 , n14974 , n5846 );
xor ( n14976 , n14971 , n14975 );
and ( n14977 , n9989 , n6554 );
and ( n14978 , n10437 , n6205 );
nor ( n14979 , n14977 , n14978 );
xnor ( n14980 , n14979 , n6550 );
xor ( n14981 , n14976 , n14980 );
xor ( n14982 , n14967 , n14981 );
or ( n14983 , n14620 , n14621 );
and ( n14984 , n9110 , n7356 );
and ( n14985 , n9583 , n6953 );
nor ( n14986 , n14984 , n14985 );
xnor ( n14987 , n14986 , n7352 );
xor ( n14988 , n14983 , n14987 );
and ( n14989 , n8640 , n7349 );
not ( n14990 , n14989 );
xor ( n14991 , n14988 , n14990 );
xor ( n14992 , n14982 , n14991 );
xor ( n14993 , n14963 , n14992 );
xor ( n14994 , n14954 , n14993 );
and ( n14995 , n14630 , n14631 );
and ( n14996 , n14631 , n14666 );
and ( n14997 , n14630 , n14666 );
or ( n14998 , n14995 , n14996 , n14997 );
xor ( n14999 , n14994 , n14998 );
xor ( n15000 , n14931 , n14999 );
and ( n15001 , n14667 , n14671 );
and ( n15002 , n14671 , n14686 );
and ( n15003 , n14667 , n14686 );
or ( n15004 , n15001 , n15002 , n15003 );
xor ( n15005 , n15000 , n15004 );
and ( n15006 , n14687 , n14690 );
xor ( n15007 , n15005 , n15006 );
buf ( n15008 , n15007 );
and ( n15009 , n14705 , n14737 );
and ( n15010 , n14737 , n14761 );
and ( n15011 , n14705 , n14761 );
or ( n15012 , n15009 , n15010 , n15011 );
and ( n15013 , n14709 , n14723 );
and ( n15014 , n14723 , n14736 );
and ( n15015 , n14709 , n14736 );
or ( n15016 , n15013 , n15014 , n15015 );
and ( n15017 , n14742 , n14746 );
and ( n15018 , n14746 , n14760 );
and ( n15019 , n14742 , n14760 );
or ( n15020 , n15017 , n15018 , n15019 );
xor ( n15021 , n15016 , n15020 );
and ( n15022 , n14751 , n14754 );
and ( n15023 , n14754 , n14759 );
and ( n15024 , n14751 , n14759 );
or ( n15025 , n15022 , n15023 , n15024 );
and ( n15026 , n11784 , n5323 );
and ( n15027 , n12217 , n5064 );
nor ( n15028 , n15026 , n15027 );
xnor ( n15029 , n15028 , n5319 );
and ( n15030 , n9164 , n7444 );
and ( n15031 , n9629 , n7026 );
nor ( n15032 , n15030 , n15031 );
xnor ( n15033 , n15032 , n7440 );
xor ( n15034 , n15029 , n15033 );
buf ( n15035 , n14734 );
not ( n15036 , n4398 );
xor ( n15037 , n15035 , n15036 );
and ( n15038 , n8728 , n7437 );
xor ( n15039 , n15037 , n15038 );
xor ( n15040 , n15034 , n15039 );
xor ( n15041 , n15025 , n15040 );
and ( n15042 , n14713 , n14717 );
and ( n15043 , n14717 , n14722 );
and ( n15044 , n14713 , n14722 );
or ( n15045 , n15042 , n15043 , n15044 );
and ( n15046 , n14728 , n14732 );
and ( n15047 , n14732 , n14735 );
and ( n15048 , n14728 , n14735 );
or ( n15049 , n15046 , n15047 , n15048 );
xor ( n15050 , n15045 , n15049 );
and ( n15051 , n12612 , n4835 );
and ( n15052 , n12976 , n4648 );
nor ( n15053 , n15051 , n15052 );
xnor ( n15054 , n15053 , n4831 );
and ( n15055 , n10940 , n5922 );
and ( n15056 , n11398 , n5616 );
nor ( n15057 , n15055 , n15056 );
xnor ( n15058 , n15057 , n5918 );
xor ( n15059 , n15054 , n15058 );
and ( n15060 , n10072 , n6627 );
and ( n15061 , n10534 , n6272 );
nor ( n15062 , n15060 , n15061 );
xnor ( n15063 , n15062 , n6623 );
xor ( n15064 , n15059 , n15063 );
xor ( n15065 , n15050 , n15064 );
xor ( n15066 , n15041 , n15065 );
xor ( n15067 , n15021 , n15066 );
xor ( n15068 , n15012 , n15067 );
and ( n15069 , n14696 , n14700 );
and ( n15070 , n14700 , n14762 );
and ( n15071 , n14696 , n14762 );
or ( n15072 , n15069 , n15070 , n15071 );
xor ( n15073 , n15068 , n15072 );
and ( n15074 , n14763 , n14766 );
xor ( n15075 , n15073 , n15074 );
buf ( n15076 , n15075 );
not ( n15077 , n454 );
and ( n15078 , n15077 , n15008 );
and ( n15079 , n15076 , n454 );
or ( n15080 , n15078 , n15079 );
buf ( n15081 , n15080 );
buf ( n15082 , n15081 );
and ( n15083 , n15082 , n4505 );
xor ( n15084 , n14927 , n15083 );
and ( n15085 , n14774 , n4557 );
not ( n15086 , n15085 );
xor ( n15087 , n15084 , n15086 );
and ( n15088 , n14781 , n14782 );
and ( n15089 , n14782 , n14784 );
and ( n15090 , n14781 , n14784 );
or ( n15091 , n15088 , n15089 , n15090 );
xor ( n15092 , n15087 , n15091 );
xor ( n15093 , n14924 , n15092 );
and ( n15094 , n14610 , n14786 );
and ( n15095 , n14786 , n14791 );
and ( n15096 , n14610 , n14791 );
or ( n15097 , n15094 , n15095 , n15096 );
xor ( n15098 , n15093 , n15097 );
or ( n15099 , n14792 , n14796 );
xor ( n15100 , n15098 , n15099 );
and ( n15101 , n14797 , n14799 );
xor ( n15102 , n15100 , n15101 );
buf ( n15103 , n15102 );
not ( n15104 , n4509 );
and ( n15105 , n15104 , n14920 );
and ( n15106 , n15103 , n4509 );
or ( n15107 , n15105 , n15106 );
and ( n15108 , n14838 , n14878 );
and ( n15109 , n14878 , n14905 );
and ( n15110 , n14838 , n14905 );
or ( n15111 , n15108 , n15109 , n15110 );
and ( n15112 , n14868 , n14872 );
and ( n15113 , n14872 , n14877 );
and ( n15114 , n14868 , n14877 );
or ( n15115 , n15112 , n15113 , n15114 );
and ( n15116 , n14883 , n14887 );
and ( n15117 , n14887 , n14904 );
and ( n15118 , n14883 , n14904 );
or ( n15119 , n15116 , n15117 , n15118 );
xor ( n15120 , n15115 , n15119 );
and ( n15121 , n14897 , n14898 );
and ( n15122 , n14898 , n14903 );
and ( n15123 , n14897 , n14903 );
or ( n15124 , n15121 , n15122 , n15123 );
and ( n15125 , n11989 , n6711 );
and ( n15126 , n12392 , n6332 );
nor ( n15127 , n15125 , n15126 );
xnor ( n15128 , n15127 , n6707 );
xor ( n15129 , n15124 , n15128 );
and ( n15130 , n11163 , n7630 );
and ( n15131 , n11569 , n7188 );
nor ( n15132 , n15130 , n15131 );
xnor ( n15133 , n15132 , n7626 );
xor ( n15134 , n15129 , n15133 );
xor ( n15135 , n15120 , n15134 );
xor ( n15136 , n15111 , n15135 );
and ( n15137 , n14813 , n14817 );
and ( n15138 , n14817 , n14832 );
and ( n15139 , n14813 , n14832 );
or ( n15140 , n15137 , n15138 , n15139 );
and ( n15141 , n14865 , n4524 );
and ( n15142 , n14843 , n14847 );
and ( n15143 , n14847 , n14849 );
and ( n15144 , n14843 , n14849 );
or ( n15145 , n15142 , n15143 , n15144 );
buf ( n15146 , n14846 );
not ( n15147 , n8378 );
xor ( n15148 , n15146 , n15147 );
and ( n15149 , n9848 , n8375 );
xor ( n15150 , n15148 , n15149 );
xor ( n15151 , n15145 , n15150 );
and ( n15152 , n14850 , n14854 );
and ( n15153 , n14854 , n14859 );
and ( n15154 , n14850 , n14859 );
or ( n15155 , n15152 , n15153 , n15154 );
xor ( n15156 , n15151 , n15155 );
and ( n15157 , n14860 , n14861 );
xor ( n15158 , n15156 , n15157 );
buf ( n15159 , n15158 );
buf ( n15160 , n15159 );
buf ( n15161 , n15160 );
and ( n15162 , n15161 , n4145 );
nor ( n15163 , n15141 , n15162 );
xnor ( n15164 , n15163 , n4521 );
and ( n15165 , n14212 , n4938 );
and ( n15166 , n14558 , n4711 );
nor ( n15167 , n15165 , n15166 );
xnor ( n15168 , n15167 , n4934 );
xor ( n15169 , n15164 , n15168 );
and ( n15170 , n12754 , n6068 );
and ( n15171 , n13144 , n5730 );
nor ( n15172 , n15170 , n15171 );
xnor ( n15173 , n15172 , n6064 );
xor ( n15174 , n15169 , n15173 );
xor ( n15175 , n15140 , n15174 );
and ( n15176 , n14822 , n14826 );
and ( n15177 , n14826 , n14831 );
and ( n15178 , n14822 , n14831 );
or ( n15179 , n15176 , n15177 , n15178 );
and ( n15180 , n13506 , n5441 );
and ( n15181 , n13865 , n5161 );
nor ( n15182 , n15180 , n15181 );
xnor ( n15183 , n15182 , n5437 );
xor ( n15184 , n15179 , n15183 );
and ( n15185 , n9367 , n9407 );
and ( n15186 , n9885 , n8872 );
nor ( n15187 , n15185 , n15186 );
xnor ( n15188 , n15187 , n9403 );
and ( n15189 , n8462 , n10329 );
and ( n15190 , n8968 , n9791 );
nor ( n15191 , n15189 , n15190 );
not ( n15192 , n15191 );
xor ( n15193 , n15188 , n15192 );
and ( n15194 , n14892 , n14896 );
xor ( n15195 , n15193 , n15194 );
and ( n15196 , n10287 , n8502 );
and ( n15197 , n10706 , n7970 );
nor ( n15198 , n15196 , n15197 );
xnor ( n15199 , n15198 , n8498 );
xor ( n15200 , n15195 , n15199 );
xor ( n15201 , n15184 , n15200 );
xor ( n15202 , n15175 , n15201 );
xor ( n15203 , n15136 , n15202 );
and ( n15204 , n14809 , n14833 );
and ( n15205 , n14833 , n14906 );
and ( n15206 , n14809 , n14906 );
or ( n15207 , n15204 , n15205 , n15206 );
xor ( n15208 , n15203 , n15207 );
and ( n15209 , n14907 , n14911 );
and ( n15210 , n14911 , n14916 );
and ( n15211 , n14907 , n14916 );
or ( n15212 , n15209 , n15210 , n15211 );
xor ( n15213 , n15208 , n15212 );
and ( n15214 , n14917 , n14918 );
xor ( n15215 , n15213 , n15214 );
buf ( n15216 , n15215 );
buf ( n15217 , n15085 );
and ( n15218 , n14925 , n14926 );
and ( n15219 , n14926 , n15083 );
and ( n15220 , n14925 , n15083 );
or ( n15221 , n15218 , n15219 , n15220 );
and ( n15222 , n14958 , n14962 );
and ( n15223 , n14962 , n14992 );
and ( n15224 , n14958 , n14992 );
or ( n15225 , n15222 , n15223 , n15224 );
and ( n15226 , n14943 , n14947 );
and ( n15227 , n14947 , n14952 );
and ( n15228 , n14943 , n14952 );
or ( n15229 , n15226 , n15227 , n15228 );
and ( n15230 , n12116 , n5270 );
and ( n15231 , n12527 , n5021 );
nor ( n15232 , n15230 , n15231 );
xnor ( n15233 , n15232 , n5266 );
and ( n15234 , n10437 , n6554 );
and ( n15235 , n10857 , n6205 );
nor ( n15236 , n15234 , n15235 );
xnor ( n15237 , n15236 , n6550 );
xor ( n15238 , n15233 , n15237 );
and ( n15239 , n9583 , n7356 );
and ( n15240 , n9989 , n6953 );
nor ( n15241 , n15239 , n15240 );
xnor ( n15242 , n15241 , n7352 );
xor ( n15243 , n15238 , n15242 );
xor ( n15244 , n15229 , n15243 );
and ( n15245 , n13647 , n4298 );
and ( n15246 , n14013 , n4287 );
nor ( n15247 , n15245 , n15246 );
xnor ( n15248 , n15247 , n4294 );
and ( n15249 , n12895 , n4788 );
and ( n15250 , n13313 , n4611 );
nor ( n15251 , n15249 , n15250 );
xnor ( n15252 , n15251 , n4784 );
xor ( n15253 , n15248 , n15252 );
and ( n15254 , n11295 , n5850 );
and ( n15255 , n11702 , n5566 );
nor ( n15256 , n15254 , n15255 );
xnor ( n15257 , n15256 , n5846 );
xor ( n15258 , n15253 , n15257 );
xor ( n15259 , n15244 , n15258 );
xor ( n15260 , n15225 , n15259 );
and ( n15261 , n14935 , n14939 );
and ( n15262 , n14939 , n14953 );
and ( n15263 , n14935 , n14953 );
or ( n15264 , n15261 , n15262 , n15263 );
and ( n15265 , n14967 , n14981 );
and ( n15266 , n14981 , n14991 );
and ( n15267 , n14967 , n14991 );
or ( n15268 , n15265 , n15266 , n15267 );
xor ( n15269 , n15264 , n15268 );
and ( n15270 , n14971 , n14975 );
and ( n15271 , n14975 , n14980 );
and ( n15272 , n14971 , n14980 );
or ( n15273 , n15270 , n15271 , n15272 );
and ( n15274 , n14983 , n14987 );
and ( n15275 , n14987 , n14990 );
and ( n15276 , n14983 , n14990 );
or ( n15277 , n15274 , n15275 , n15276 );
xor ( n15278 , n15273 , n15277 );
buf ( n15279 , n14989 );
not ( n15280 , n4315 );
xor ( n15281 , n15279 , n15280 );
and ( n15282 , n9110 , n7349 );
xor ( n15283 , n15281 , n15282 );
xor ( n15284 , n15278 , n15283 );
xor ( n15285 , n15269 , n15284 );
xor ( n15286 , n15260 , n15285 );
and ( n15287 , n14954 , n14993 );
and ( n15288 , n14993 , n14998 );
and ( n15289 , n14954 , n14998 );
or ( n15290 , n15287 , n15288 , n15289 );
xor ( n15291 , n15286 , n15290 );
and ( n15292 , n14931 , n14999 );
and ( n15293 , n14999 , n15004 );
and ( n15294 , n14931 , n15004 );
or ( n15295 , n15292 , n15293 , n15294 );
xor ( n15296 , n15291 , n15295 );
and ( n15297 , n15005 , n15006 );
xor ( n15298 , n15296 , n15297 );
buf ( n15299 , n15298 );
and ( n15300 , n15025 , n15040 );
and ( n15301 , n15040 , n15065 );
and ( n15302 , n15025 , n15065 );
or ( n15303 , n15300 , n15301 , n15302 );
and ( n15304 , n15054 , n15058 );
and ( n15305 , n15058 , n15063 );
and ( n15306 , n15054 , n15063 );
or ( n15307 , n15304 , n15305 , n15306 );
and ( n15308 , n15035 , n15036 );
and ( n15309 , n15036 , n15038 );
and ( n15310 , n15035 , n15038 );
or ( n15311 , n15308 , n15309 , n15310 );
xor ( n15312 , n15307 , n15311 );
and ( n15313 , n12976 , n4835 );
not ( n15314 , n15313 );
xnor ( n15315 , n15314 , n4831 );
and ( n15316 , n11398 , n5922 );
and ( n15317 , n11784 , n5616 );
nor ( n15318 , n15316 , n15317 );
xnor ( n15319 , n15318 , n5918 );
xor ( n15320 , n15315 , n15319 );
and ( n15321 , n9164 , n7437 );
not ( n15322 , n15321 );
xor ( n15323 , n15320 , n15322 );
xor ( n15324 , n15312 , n15323 );
xor ( n15325 , n15303 , n15324 );
and ( n15326 , n15029 , n15033 );
and ( n15327 , n15033 , n15039 );
and ( n15328 , n15029 , n15039 );
or ( n15329 , n15326 , n15327 , n15328 );
and ( n15330 , n15045 , n15049 );
and ( n15331 , n15049 , n15064 );
and ( n15332 , n15045 , n15064 );
or ( n15333 , n15330 , n15331 , n15332 );
xor ( n15334 , n15329 , n15333 );
and ( n15335 , n12217 , n5323 );
and ( n15336 , n12612 , n5064 );
nor ( n15337 , n15335 , n15336 );
xnor ( n15338 , n15337 , n5319 );
and ( n15339 , n10534 , n6627 );
and ( n15340 , n10940 , n6272 );
nor ( n15341 , n15339 , n15340 );
xnor ( n15342 , n15341 , n6623 );
xor ( n15343 , n15338 , n15342 );
and ( n15344 , n9629 , n7444 );
and ( n15345 , n10072 , n7026 );
nor ( n15346 , n15344 , n15345 );
xnor ( n15347 , n15346 , n7440 );
xor ( n15348 , n15343 , n15347 );
xor ( n15349 , n15334 , n15348 );
xor ( n15350 , n15325 , n15349 );
and ( n15351 , n15016 , n15020 );
and ( n15352 , n15020 , n15066 );
and ( n15353 , n15016 , n15066 );
or ( n15354 , n15351 , n15352 , n15353 );
xor ( n15355 , n15350 , n15354 );
and ( n15356 , n15012 , n15067 );
and ( n15357 , n15067 , n15072 );
and ( n15358 , n15012 , n15072 );
or ( n15359 , n15356 , n15357 , n15358 );
xor ( n15360 , n15355 , n15359 );
and ( n15361 , n15073 , n15074 );
xor ( n15362 , n15360 , n15361 );
buf ( n15363 , n15362 );
not ( n15364 , n454 );
and ( n15365 , n15364 , n15299 );
and ( n15366 , n15363 , n454 );
or ( n15367 , n15365 , n15366 );
buf ( n15368 , n15367 );
buf ( n15369 , n15368 );
and ( n15370 , n15369 , n4505 );
xor ( n15371 , n15221 , n15370 );
and ( n15372 , n14461 , n5089 );
and ( n15373 , n14774 , n4866 );
xor ( n15374 , n15372 , n15373 );
and ( n15375 , n15082 , n4557 );
xor ( n15376 , n15374 , n15375 );
xor ( n15377 , n15371 , n15376 );
xor ( n15378 , n15217 , n15377 );
and ( n15379 , n15084 , n15086 );
and ( n15380 , n15086 , n15091 );
and ( n15381 , n15084 , n15091 );
or ( n15382 , n15379 , n15380 , n15381 );
xor ( n15383 , n15378 , n15382 );
and ( n15384 , n14924 , n15092 );
and ( n15385 , n15092 , n15097 );
and ( n15386 , n14924 , n15097 );
or ( n15387 , n15384 , n15385 , n15386 );
xnor ( n15388 , n15383 , n15387 );
and ( n15389 , n15098 , n15099 );
and ( n15390 , n15100 , n15101 );
or ( n15391 , n15389 , n15390 );
xor ( n15392 , n15388 , n15391 );
buf ( n15393 , n15392 );
not ( n15394 , n4509 );
and ( n15395 , n15394 , n15216 );
and ( n15396 , n15393 , n4509 );
or ( n15397 , n15395 , n15396 );
and ( n15398 , n15140 , n15174 );
and ( n15399 , n15174 , n15201 );
and ( n15400 , n15140 , n15201 );
or ( n15401 , n15398 , n15399 , n15400 );
and ( n15402 , n15164 , n15168 );
and ( n15403 , n15168 , n15173 );
and ( n15404 , n15164 , n15173 );
or ( n15405 , n15402 , n15403 , n15404 );
and ( n15406 , n15161 , n4524 );
not ( n15407 , n15406 );
xnor ( n15408 , n15407 , n4521 );
and ( n15409 , n14558 , n4938 );
and ( n15410 , n14865 , n4711 );
nor ( n15411 , n15409 , n15410 );
xnor ( n15412 , n15411 , n4934 );
xor ( n15413 , n15408 , n15412 );
and ( n15414 , n13144 , n6068 );
and ( n15415 , n13506 , n5730 );
nor ( n15416 , n15414 , n15415 );
xnor ( n15417 , n15416 , n6064 );
xor ( n15418 , n15413 , n15417 );
xor ( n15419 , n15405 , n15418 );
and ( n15420 , n15193 , n15194 );
and ( n15421 , n15194 , n15199 );
and ( n15422 , n15193 , n15199 );
or ( n15423 , n15420 , n15421 , n15422 );
and ( n15424 , n12392 , n6711 );
and ( n15425 , n12754 , n6332 );
nor ( n15426 , n15424 , n15425 );
xnor ( n15427 , n15426 , n6707 );
xor ( n15428 , n15423 , n15427 );
and ( n15429 , n11569 , n7630 );
and ( n15430 , n11989 , n7188 );
nor ( n15431 , n15429 , n15430 );
xnor ( n15432 , n15431 , n7626 );
xor ( n15433 , n15428 , n15432 );
xor ( n15434 , n15419 , n15433 );
xor ( n15435 , n15401 , n15434 );
and ( n15436 , n15179 , n15183 );
and ( n15437 , n15183 , n15200 );
and ( n15438 , n15179 , n15200 );
or ( n15439 , n15436 , n15437 , n15438 );
and ( n15440 , n15115 , n15119 );
and ( n15441 , n15119 , n15134 );
and ( n15442 , n15115 , n15134 );
or ( n15443 , n15440 , n15441 , n15442 );
xor ( n15444 , n15439 , n15443 );
and ( n15445 , n15124 , n15128 );
and ( n15446 , n15128 , n15133 );
and ( n15447 , n15124 , n15133 );
or ( n15448 , n15445 , n15446 , n15447 );
and ( n15449 , n13865 , n5441 );
and ( n15450 , n14212 , n5161 );
nor ( n15451 , n15449 , n15450 );
xnor ( n15452 , n15451 , n5437 );
xor ( n15453 , n15448 , n15452 );
and ( n15454 , n9885 , n9407 );
and ( n15455 , n10287 , n8872 );
nor ( n15456 , n15454 , n15455 );
xnor ( n15457 , n15456 , n9403 );
and ( n15458 , n8968 , n10329 );
and ( n15459 , n9367 , n9791 );
nor ( n15460 , n15458 , n15459 );
not ( n15461 , n15460 );
xor ( n15462 , n15457 , n15461 );
and ( n15463 , n15188 , n15192 );
xor ( n15464 , n15462 , n15463 );
and ( n15465 , n10706 , n8502 );
and ( n15466 , n11163 , n7970 );
nor ( n15467 , n15465 , n15466 );
xnor ( n15468 , n15467 , n8498 );
xor ( n15469 , n15464 , n15468 );
xor ( n15470 , n15453 , n15469 );
xor ( n15471 , n15444 , n15470 );
xor ( n15472 , n15435 , n15471 );
and ( n15473 , n15111 , n15135 );
and ( n15474 , n15135 , n15202 );
and ( n15475 , n15111 , n15202 );
or ( n15476 , n15473 , n15474 , n15475 );
xor ( n15477 , n15472 , n15476 );
and ( n15478 , n15203 , n15207 );
and ( n15479 , n15207 , n15212 );
and ( n15480 , n15203 , n15212 );
or ( n15481 , n15478 , n15479 , n15480 );
xor ( n15482 , n15477 , n15481 );
and ( n15483 , n15213 , n15214 );
xor ( n15484 , n15482 , n15483 );
buf ( n15485 , n15484 );
and ( n15486 , n15372 , n15373 );
and ( n15487 , n15373 , n15375 );
and ( n15488 , n15372 , n15375 );
or ( n15489 , n15486 , n15487 , n15488 );
and ( n15490 , n15369 , n4557 );
xor ( n15491 , n15489 , n15490 );
and ( n15492 , n14774 , n5089 );
and ( n15493 , n15082 , n4866 );
xor ( n15494 , n15492 , n15493 );
and ( n15495 , n15264 , n15268 );
and ( n15496 , n15268 , n15284 );
and ( n15497 , n15264 , n15284 );
or ( n15498 , n15495 , n15496 , n15497 );
and ( n15499 , n15248 , n15252 );
and ( n15500 , n15252 , n15257 );
and ( n15501 , n15248 , n15257 );
or ( n15502 , n15499 , n15500 , n15501 );
and ( n15503 , n12527 , n5270 );
and ( n15504 , n12895 , n5021 );
nor ( n15505 , n15503 , n15504 );
xnor ( n15506 , n15505 , n5266 );
and ( n15507 , n10857 , n6554 );
and ( n15508 , n11295 , n6205 );
nor ( n15509 , n15507 , n15508 );
xnor ( n15510 , n15509 , n6550 );
xor ( n15511 , n15506 , n15510 );
and ( n15512 , n9989 , n7356 );
and ( n15513 , n10437 , n6953 );
nor ( n15514 , n15512 , n15513 );
xnor ( n15515 , n15514 , n7352 );
xor ( n15516 , n15511 , n15515 );
xor ( n15517 , n15502 , n15516 );
and ( n15518 , n13313 , n4788 );
and ( n15519 , n13647 , n4611 );
nor ( n15520 , n15518 , n15519 );
xnor ( n15521 , n15520 , n4784 );
and ( n15522 , n11702 , n5850 );
and ( n15523 , n12116 , n5566 );
nor ( n15524 , n15522 , n15523 );
xnor ( n15525 , n15524 , n5846 );
xor ( n15526 , n15521 , n15525 );
and ( n15527 , n9583 , n7349 );
not ( n15528 , n15527 );
xor ( n15529 , n15526 , n15528 );
xor ( n15530 , n15517 , n15529 );
xor ( n15531 , n15498 , n15530 );
and ( n15532 , n15229 , n15243 );
and ( n15533 , n15243 , n15258 );
and ( n15534 , n15229 , n15258 );
or ( n15535 , n15532 , n15533 , n15534 );
and ( n15536 , n15273 , n15277 );
and ( n15537 , n15277 , n15283 );
and ( n15538 , n15273 , n15283 );
or ( n15539 , n15536 , n15537 , n15538 );
xor ( n15540 , n15535 , n15539 );
and ( n15541 , n15233 , n15237 );
and ( n15542 , n15237 , n15242 );
and ( n15543 , n15233 , n15242 );
or ( n15544 , n15541 , n15542 , n15543 );
and ( n15545 , n15279 , n15280 );
and ( n15546 , n15280 , n15282 );
and ( n15547 , n15279 , n15282 );
or ( n15548 , n15545 , n15546 , n15547 );
xor ( n15549 , n15544 , n15548 );
and ( n15550 , n14013 , n4298 );
not ( n15551 , n15550 );
xnor ( n15552 , n15551 , n4294 );
xor ( n15553 , n15549 , n15552 );
xor ( n15554 , n15540 , n15553 );
xor ( n15555 , n15531 , n15554 );
and ( n15556 , n15225 , n15259 );
and ( n15557 , n15259 , n15285 );
and ( n15558 , n15225 , n15285 );
or ( n15559 , n15556 , n15557 , n15558 );
xor ( n15560 , n15555 , n15559 );
and ( n15561 , n15286 , n15290 );
and ( n15562 , n15290 , n15295 );
and ( n15563 , n15286 , n15295 );
or ( n15564 , n15561 , n15562 , n15563 );
xor ( n15565 , n15560 , n15564 );
and ( n15566 , n15296 , n15297 );
xor ( n15567 , n15565 , n15566 );
buf ( n15568 , n15567 );
and ( n15569 , n15307 , n15311 );
and ( n15570 , n15311 , n15323 );
and ( n15571 , n15307 , n15323 );
or ( n15572 , n15569 , n15570 , n15571 );
and ( n15573 , n15329 , n15333 );
and ( n15574 , n15333 , n15348 );
and ( n15575 , n15329 , n15348 );
or ( n15576 , n15573 , n15574 , n15575 );
xor ( n15577 , n15572 , n15576 );
and ( n15578 , n11784 , n5922 );
and ( n15579 , n12217 , n5616 );
nor ( n15580 , n15578 , n15579 );
xnor ( n15581 , n15580 , n5918 );
and ( n15582 , n10072 , n7444 );
and ( n15583 , n10534 , n7026 );
nor ( n15584 , n15582 , n15583 );
xnor ( n15585 , n15584 , n7440 );
xor ( n15586 , n15581 , n15585 );
and ( n15587 , n9629 , n7437 );
xor ( n15588 , n15586 , n15587 );
not ( n15589 , n4831 );
and ( n15590 , n12612 , n5323 );
and ( n15591 , n12976 , n5064 );
nor ( n15592 , n15590 , n15591 );
xnor ( n15593 , n15592 , n5319 );
xor ( n15594 , n15589 , n15593 );
and ( n15595 , n10940 , n6627 );
and ( n15596 , n11398 , n6272 );
nor ( n15597 , n15595 , n15596 );
xnor ( n15598 , n15597 , n6623 );
xor ( n15599 , n15594 , n15598 );
xor ( n15600 , n15588 , n15599 );
and ( n15601 , n15338 , n15342 );
and ( n15602 , n15342 , n15347 );
and ( n15603 , n15338 , n15347 );
or ( n15604 , n15601 , n15602 , n15603 );
and ( n15605 , n15315 , n15319 );
and ( n15606 , n15319 , n15322 );
and ( n15607 , n15315 , n15322 );
or ( n15608 , n15605 , n15606 , n15607 );
xor ( n15609 , n15604 , n15608 );
buf ( n15610 , n15321 );
xor ( n15611 , n15609 , n15610 );
xor ( n15612 , n15600 , n15611 );
xor ( n15613 , n15577 , n15612 );
and ( n15614 , n15303 , n15324 );
and ( n15615 , n15324 , n15349 );
and ( n15616 , n15303 , n15349 );
or ( n15617 , n15614 , n15615 , n15616 );
xor ( n15618 , n15613 , n15617 );
and ( n15619 , n15350 , n15354 );
and ( n15620 , n15354 , n15359 );
and ( n15621 , n15350 , n15359 );
or ( n15622 , n15619 , n15620 , n15621 );
xor ( n15623 , n15618 , n15622 );
and ( n15624 , n15360 , n15361 );
xor ( n15625 , n15623 , n15624 );
buf ( n15626 , n15625 );
not ( n15627 , n454 );
and ( n15628 , n15627 , n15568 );
and ( n15629 , n15626 , n454 );
or ( n15630 , n15628 , n15629 );
buf ( n15631 , n15630 );
buf ( n15632 , n15631 );
and ( n15633 , n15632 , n4505 );
xor ( n15634 , n15494 , n15633 );
xor ( n15635 , n15491 , n15634 );
and ( n15636 , n15221 , n15370 );
and ( n15637 , n15370 , n15376 );
and ( n15638 , n15221 , n15376 );
or ( n15639 , n15636 , n15637 , n15638 );
xor ( n15640 , n15635 , n15639 );
and ( n15641 , n15217 , n15377 );
and ( n15642 , n15377 , n15382 );
and ( n15643 , n15217 , n15382 );
or ( n15644 , n15641 , n15642 , n15643 );
xor ( n15645 , n15640 , n15644 );
or ( n15646 , n15383 , n15387 );
xnor ( n15647 , n15645 , n15646 );
and ( n15648 , n15388 , n15391 );
xor ( n15649 , n15647 , n15648 );
buf ( n15650 , n15649 );
not ( n15651 , n4509 );
and ( n15652 , n15651 , n15485 );
and ( n15653 , n15650 , n4509 );
or ( n15654 , n15652 , n15653 );
and ( n15655 , n15423 , n15427 );
and ( n15656 , n15427 , n15432 );
and ( n15657 , n15423 , n15432 );
or ( n15658 , n15655 , n15656 , n15657 );
and ( n15659 , n15448 , n15452 );
and ( n15660 , n15452 , n15469 );
and ( n15661 , n15448 , n15469 );
or ( n15662 , n15659 , n15660 , n15661 );
xor ( n15663 , n15658 , n15662 );
and ( n15664 , n15462 , n15463 );
and ( n15665 , n15463 , n15468 );
and ( n15666 , n15462 , n15468 );
or ( n15667 , n15664 , n15665 , n15666 );
and ( n15668 , n11163 , n8502 );
and ( n15669 , n11569 , n7970 );
nor ( n15670 , n15668 , n15669 );
xnor ( n15671 , n15670 , n8498 );
and ( n15672 , n10287 , n9407 );
and ( n15673 , n10706 , n8872 );
nor ( n15674 , n15672 , n15673 );
xnor ( n15675 , n15674 , n9403 );
xor ( n15676 , n15671 , n15675 );
not ( n15677 , n4521 );
and ( n15678 , n9367 , n10329 );
and ( n15679 , n9885 , n9791 );
nor ( n15680 , n15678 , n15679 );
not ( n15681 , n15680 );
xnor ( n15682 , n15677 , n15681 );
xor ( n15683 , n15676 , n15682 );
xor ( n15684 , n15667 , n15683 );
and ( n15685 , n15408 , n15412 );
and ( n15686 , n15412 , n15417 );
and ( n15687 , n15408 , n15417 );
or ( n15688 , n15685 , n15686 , n15687 );
and ( n15689 , n14865 , n4938 );
and ( n15690 , n15161 , n4711 );
nor ( n15691 , n15689 , n15690 );
xnor ( n15692 , n15691 , n4934 );
and ( n15693 , n14212 , n5441 );
and ( n15694 , n14558 , n5161 );
nor ( n15695 , n15693 , n15694 );
xnor ( n15696 , n15695 , n5437 );
xor ( n15697 , n15692 , n15696 );
and ( n15698 , n13506 , n6068 );
and ( n15699 , n13865 , n5730 );
nor ( n15700 , n15698 , n15699 );
xnor ( n15701 , n15700 , n6064 );
xor ( n15702 , n15697 , n15701 );
xor ( n15703 , n15688 , n15702 );
and ( n15704 , n15457 , n15461 );
and ( n15705 , n12754 , n6711 );
and ( n15706 , n13144 , n6332 );
nor ( n15707 , n15705 , n15706 );
xnor ( n15708 , n15707 , n6707 );
xor ( n15709 , n15704 , n15708 );
and ( n15710 , n11989 , n7630 );
and ( n15711 , n12392 , n7188 );
nor ( n15712 , n15710 , n15711 );
xnor ( n15713 , n15712 , n7626 );
xor ( n15714 , n15709 , n15713 );
xor ( n15715 , n15703 , n15714 );
xor ( n15716 , n15684 , n15715 );
xor ( n15717 , n15663 , n15716 );
and ( n15718 , n15405 , n15418 );
and ( n15719 , n15418 , n15433 );
and ( n15720 , n15405 , n15433 );
or ( n15721 , n15718 , n15719 , n15720 );
and ( n15722 , n15439 , n15443 );
and ( n15723 , n15443 , n15470 );
and ( n15724 , n15439 , n15470 );
or ( n15725 , n15722 , n15723 , n15724 );
xor ( n15726 , n15721 , n15725 );
xor ( n15727 , n15717 , n15726 );
and ( n15728 , n15401 , n15434 );
and ( n15729 , n15434 , n15471 );
and ( n15730 , n15401 , n15471 );
or ( n15731 , n15728 , n15729 , n15730 );
xor ( n15732 , n15727 , n15731 );
and ( n15733 , n15472 , n15476 );
and ( n15734 , n15476 , n15481 );
and ( n15735 , n15472 , n15481 );
or ( n15736 , n15733 , n15734 , n15735 );
xor ( n15737 , n15732 , n15736 );
and ( n15738 , n15482 , n15483 );
xor ( n15739 , n15737 , n15738 );
buf ( n15740 , n15739 );
and ( n15741 , n15492 , n15493 );
and ( n15742 , n15493 , n15633 );
and ( n15743 , n15492 , n15633 );
or ( n15744 , n15741 , n15742 , n15743 );
and ( n15745 , n15535 , n15539 );
and ( n15746 , n15539 , n15553 );
and ( n15747 , n15535 , n15553 );
or ( n15748 , n15745 , n15746 , n15747 );
and ( n15749 , n15521 , n15525 );
and ( n15750 , n15525 , n15528 );
and ( n15751 , n15521 , n15528 );
or ( n15752 , n15749 , n15750 , n15751 );
not ( n15753 , n4294 );
and ( n15754 , n10437 , n7356 );
and ( n15755 , n10857 , n6953 );
nor ( n15756 , n15754 , n15755 );
xnor ( n15757 , n15756 , n7352 );
xor ( n15758 , n15753 , n15757 );
and ( n15759 , n9989 , n7349 );
xor ( n15760 , n15758 , n15759 );
xor ( n15761 , n15752 , n15760 );
buf ( n15762 , n15527 );
and ( n15763 , n12116 , n5850 );
and ( n15764 , n12527 , n5566 );
nor ( n15765 , n15763 , n15764 );
xnor ( n15766 , n15765 , n5846 );
xor ( n15767 , n15762 , n15766 );
and ( n15768 , n11295 , n6554 );
and ( n15769 , n11702 , n6205 );
nor ( n15770 , n15768 , n15769 );
xnor ( n15771 , n15770 , n6550 );
xor ( n15772 , n15767 , n15771 );
xor ( n15773 , n15761 , n15772 );
xor ( n15774 , n15748 , n15773 );
and ( n15775 , n15544 , n15548 );
and ( n15776 , n15548 , n15552 );
and ( n15777 , n15544 , n15552 );
or ( n15778 , n15775 , n15776 , n15777 );
and ( n15779 , n15502 , n15516 );
and ( n15780 , n15516 , n15529 );
and ( n15781 , n15502 , n15529 );
or ( n15782 , n15779 , n15780 , n15781 );
xor ( n15783 , n15778 , n15782 );
and ( n15784 , n15506 , n15510 );
and ( n15785 , n15510 , n15515 );
and ( n15786 , n15506 , n15515 );
or ( n15787 , n15784 , n15785 , n15786 );
and ( n15788 , n13647 , n4788 );
and ( n15789 , n14013 , n4611 );
nor ( n15790 , n15788 , n15789 );
xnor ( n15791 , n15790 , n4784 );
xor ( n15792 , n15787 , n15791 );
and ( n15793 , n12895 , n5270 );
and ( n15794 , n13313 , n5021 );
nor ( n15795 , n15793 , n15794 );
xnor ( n15796 , n15795 , n5266 );
xor ( n15797 , n15792 , n15796 );
xor ( n15798 , n15783 , n15797 );
xor ( n15799 , n15774 , n15798 );
and ( n15800 , n15498 , n15530 );
and ( n15801 , n15530 , n15554 );
and ( n15802 , n15498 , n15554 );
or ( n15803 , n15800 , n15801 , n15802 );
xor ( n15804 , n15799 , n15803 );
and ( n15805 , n15555 , n15559 );
and ( n15806 , n15559 , n15564 );
and ( n15807 , n15555 , n15564 );
or ( n15808 , n15805 , n15806 , n15807 );
xor ( n15809 , n15804 , n15808 );
and ( n15810 , n15565 , n15566 );
xor ( n15811 , n15809 , n15810 );
buf ( n15812 , n15811 );
and ( n15813 , n15604 , n15608 );
and ( n15814 , n15608 , n15610 );
and ( n15815 , n15604 , n15610 );
or ( n15816 , n15813 , n15814 , n15815 );
and ( n15817 , n15588 , n15599 );
and ( n15818 , n15599 , n15611 );
and ( n15819 , n15588 , n15611 );
or ( n15820 , n15817 , n15818 , n15819 );
xor ( n15821 , n15816 , n15820 );
and ( n15822 , n15589 , n15593 );
and ( n15823 , n15593 , n15598 );
and ( n15824 , n15589 , n15598 );
or ( n15825 , n15822 , n15823 , n15824 );
and ( n15826 , n12976 , n5323 );
not ( n15827 , n15826 );
xnor ( n15828 , n15827 , n5319 );
and ( n15829 , n10534 , n7444 );
and ( n15830 , n10940 , n7026 );
nor ( n15831 , n15829 , n15830 );
xnor ( n15832 , n15831 , n7440 );
xor ( n15833 , n15828 , n15832 );
and ( n15834 , n10072 , n7437 );
xor ( n15835 , n15833 , n15834 );
xor ( n15836 , n15825 , n15835 );
and ( n15837 , n15581 , n15585 );
and ( n15838 , n15585 , n15587 );
and ( n15839 , n15581 , n15587 );
or ( n15840 , n15837 , n15838 , n15839 );
and ( n15841 , n12217 , n5922 );
and ( n15842 , n12612 , n5616 );
nor ( n15843 , n15841 , n15842 );
xnor ( n15844 , n15843 , n5918 );
not ( n15845 , n15844 );
xor ( n15846 , n15840 , n15845 );
and ( n15847 , n11398 , n6627 );
and ( n15848 , n11784 , n6272 );
nor ( n15849 , n15847 , n15848 );
xnor ( n15850 , n15849 , n6623 );
xor ( n15851 , n15846 , n15850 );
xor ( n15852 , n15836 , n15851 );
xor ( n15853 , n15821 , n15852 );
and ( n15854 , n15572 , n15576 );
and ( n15855 , n15576 , n15612 );
and ( n15856 , n15572 , n15612 );
or ( n15857 , n15854 , n15855 , n15856 );
xor ( n15858 , n15853 , n15857 );
and ( n15859 , n15613 , n15617 );
and ( n15860 , n15617 , n15622 );
and ( n15861 , n15613 , n15622 );
or ( n15862 , n15859 , n15860 , n15861 );
xor ( n15863 , n15858 , n15862 );
and ( n15864 , n15623 , n15624 );
xor ( n15865 , n15863 , n15864 );
buf ( n15866 , n15865 );
not ( n15867 , n454 );
and ( n15868 , n15867 , n15812 );
and ( n15869 , n15866 , n454 );
or ( n15870 , n15868 , n15869 );
buf ( n15871 , n15870 );
buf ( n15872 , n15871 );
and ( n15873 , n15872 , n4505 );
xor ( n15874 , n15744 , n15873 );
and ( n15875 , n15082 , n5089 );
and ( n15876 , n15369 , n4866 );
xor ( n15877 , n15875 , n15876 );
and ( n15878 , n15632 , n4557 );
xor ( n15879 , n15877 , n15878 );
xor ( n15880 , n15874 , n15879 );
and ( n15881 , n15489 , n15490 );
and ( n15882 , n15490 , n15634 );
and ( n15883 , n15489 , n15634 );
or ( n15884 , n15881 , n15882 , n15883 );
xor ( n15885 , n15880 , n15884 );
and ( n15886 , n15635 , n15639 );
and ( n15887 , n15639 , n15644 );
and ( n15888 , n15635 , n15644 );
or ( n15889 , n15886 , n15887 , n15888 );
xor ( n15890 , n15885 , n15889 );
or ( n15891 , n15645 , n15646 );
xnor ( n15892 , n15890 , n15891 );
and ( n15893 , n15647 , n15648 );
xor ( n15894 , n15892 , n15893 );
buf ( n15895 , n15894 );
not ( n15896 , n4509 );
and ( n15897 , n15896 , n15740 );
and ( n15898 , n15895 , n4509 );
or ( n15899 , n15897 , n15898 );
and ( n15900 , n15667 , n15683 );
and ( n15901 , n15683 , n15715 );
and ( n15902 , n15667 , n15715 );
or ( n15903 , n15900 , n15901 , n15902 );
and ( n15904 , n15688 , n15702 );
and ( n15905 , n15702 , n15714 );
and ( n15906 , n15688 , n15714 );
or ( n15907 , n15904 , n15905 , n15906 );
and ( n15908 , n10706 , n9407 );
and ( n15909 , n11163 , n8872 );
nor ( n15910 , n15908 , n15909 );
xnor ( n15911 , n15910 , n9403 );
and ( n15912 , n15161 , n4938 );
not ( n15913 , n15912 );
xnor ( n15914 , n15913 , n4934 );
and ( n15915 , n14558 , n5441 );
and ( n15916 , n14865 , n5161 );
nor ( n15917 , n15915 , n15916 );
xnor ( n15918 , n15917 , n5437 );
xor ( n15919 , n15914 , n15918 );
and ( n15920 , n13865 , n6068 );
and ( n15921 , n14212 , n5730 );
nor ( n15922 , n15920 , n15921 );
xnor ( n15923 , n15922 , n6064 );
xor ( n15924 , n15919 , n15923 );
xor ( n15925 , n15911 , n15924 );
and ( n15926 , n15692 , n15696 );
and ( n15927 , n15696 , n15701 );
and ( n15928 , n15692 , n15701 );
or ( n15929 , n15926 , n15927 , n15928 );
and ( n15930 , n13144 , n6711 );
and ( n15931 , n13506 , n6332 );
nor ( n15932 , n15930 , n15931 );
xnor ( n15933 , n15932 , n6707 );
and ( n15934 , n12392 , n7630 );
and ( n15935 , n12754 , n7188 );
nor ( n15936 , n15934 , n15935 );
xnor ( n15937 , n15936 , n7626 );
xor ( n15938 , n15933 , n15937 );
and ( n15939 , n11569 , n8502 );
and ( n15940 , n11989 , n7970 );
nor ( n15941 , n15939 , n15940 );
xnor ( n15942 , n15941 , n8498 );
xor ( n15943 , n15938 , n15942 );
xor ( n15944 , n15929 , n15943 );
xor ( n15945 , n15925 , n15944 );
xor ( n15946 , n15907 , n15945 );
or ( n15947 , n15677 , n15681 );
and ( n15948 , n9885 , n10329 );
and ( n15949 , n10287 , n9791 );
nor ( n15950 , n15948 , n15949 );
xor ( n15951 , n15947 , n15950 );
and ( n15952 , n15704 , n15708 );
and ( n15953 , n15708 , n15713 );
and ( n15954 , n15704 , n15713 );
or ( n15955 , n15952 , n15953 , n15954 );
xor ( n15956 , n15951 , n15955 );
and ( n15957 , n15671 , n15675 );
and ( n15958 , n15675 , n15682 );
and ( n15959 , n15671 , n15682 );
or ( n15960 , n15957 , n15958 , n15959 );
xor ( n15961 , n15956 , n15960 );
xor ( n15962 , n15946 , n15961 );
xor ( n15963 , n15903 , n15962 );
and ( n15964 , n15658 , n15662 );
and ( n15965 , n15662 , n15716 );
and ( n15966 , n15658 , n15716 );
or ( n15967 , n15964 , n15965 , n15966 );
xor ( n15968 , n15963 , n15967 );
and ( n15969 , n15721 , n15725 );
xor ( n15970 , n15968 , n15969 );
and ( n15971 , n15717 , n15726 );
and ( n15972 , n15726 , n15731 );
and ( n15973 , n15717 , n15731 );
or ( n15974 , n15971 , n15972 , n15973 );
xor ( n15975 , n15970 , n15974 );
and ( n15976 , n15732 , n15736 );
and ( n15977 , n15737 , n15738 );
or ( n15978 , n15976 , n15977 );
xor ( n15979 , n15975 , n15978 );
buf ( n15980 , n15979 );
and ( n15981 , n15369 , n5089 );
and ( n15982 , n15632 , n4866 );
xor ( n15983 , n15981 , n15982 );
and ( n15984 , n15778 , n15782 );
and ( n15985 , n15782 , n15797 );
and ( n15986 , n15778 , n15797 );
or ( n15987 , n15984 , n15985 , n15986 );
and ( n15988 , n15753 , n15757 );
and ( n15989 , n15757 , n15759 );
and ( n15990 , n15753 , n15759 );
or ( n15991 , n15988 , n15989 , n15990 );
and ( n15992 , n15762 , n15766 );
and ( n15993 , n15766 , n15771 );
and ( n15994 , n15762 , n15771 );
or ( n15995 , n15992 , n15993 , n15994 );
xor ( n15996 , n15991 , n15995 );
and ( n15997 , n12527 , n5850 );
and ( n15998 , n12895 , n5566 );
nor ( n15999 , n15997 , n15998 );
xnor ( n16000 , n15999 , n5846 );
and ( n16001 , n11702 , n6554 );
and ( n16002 , n12116 , n6205 );
nor ( n16003 , n16001 , n16002 );
xnor ( n16004 , n16003 , n6550 );
xor ( n16005 , n16000 , n16004 );
and ( n16006 , n10437 , n7349 );
xor ( n16007 , n16005 , n16006 );
xor ( n16008 , n15996 , n16007 );
xor ( n16009 , n15987 , n16008 );
and ( n16010 , n15787 , n15791 );
and ( n16011 , n15791 , n15796 );
and ( n16012 , n15787 , n15796 );
or ( n16013 , n16010 , n16011 , n16012 );
and ( n16014 , n15752 , n15760 );
and ( n16015 , n15760 , n15772 );
and ( n16016 , n15752 , n15772 );
or ( n16017 , n16014 , n16015 , n16016 );
xor ( n16018 , n16013 , n16017 );
and ( n16019 , n14013 , n4788 );
not ( n16020 , n16019 );
xnor ( n16021 , n16020 , n4784 );
and ( n16022 , n13313 , n5270 );
and ( n16023 , n13647 , n5021 );
nor ( n16024 , n16022 , n16023 );
xnor ( n16025 , n16024 , n5266 );
xor ( n16026 , n16021 , n16025 );
and ( n16027 , n10857 , n7356 );
and ( n16028 , n11295 , n6953 );
nor ( n16029 , n16027 , n16028 );
xnor ( n16030 , n16029 , n7352 );
not ( n16031 , n16030 );
xor ( n16032 , n16026 , n16031 );
xor ( n16033 , n16018 , n16032 );
xor ( n16034 , n16009 , n16033 );
and ( n16035 , n15748 , n15773 );
and ( n16036 , n15773 , n15798 );
and ( n16037 , n15748 , n15798 );
or ( n16038 , n16035 , n16036 , n16037 );
xor ( n16039 , n16034 , n16038 );
and ( n16040 , n15799 , n15803 );
and ( n16041 , n15803 , n15808 );
and ( n16042 , n15799 , n15808 );
or ( n16043 , n16040 , n16041 , n16042 );
xor ( n16044 , n16039 , n16043 );
and ( n16045 , n15809 , n15810 );
xor ( n16046 , n16044 , n16045 );
buf ( n16047 , n16046 );
and ( n16048 , n15816 , n15820 );
and ( n16049 , n15820 , n15852 );
and ( n16050 , n15816 , n15852 );
or ( n16051 , n16048 , n16049 , n16050 );
and ( n16052 , n15840 , n15845 );
and ( n16053 , n15845 , n15850 );
and ( n16054 , n15840 , n15850 );
or ( n16055 , n16052 , n16053 , n16054 );
and ( n16056 , n15825 , n15835 );
and ( n16057 , n15835 , n15851 );
and ( n16058 , n15825 , n15851 );
or ( n16059 , n16056 , n16057 , n16058 );
xor ( n16060 , n16055 , n16059 );
and ( n16061 , n15828 , n15832 );
and ( n16062 , n15832 , n15834 );
and ( n16063 , n15828 , n15834 );
or ( n16064 , n16061 , n16062 , n16063 );
not ( n16065 , n5319 );
and ( n16066 , n12612 , n5922 );
and ( n16067 , n12976 , n5616 );
nor ( n16068 , n16066 , n16067 );
xnor ( n16069 , n16068 , n5918 );
xor ( n16070 , n16065 , n16069 );
and ( n16071 , n10940 , n7444 );
and ( n16072 , n11398 , n7026 );
nor ( n16073 , n16071 , n16072 );
xnor ( n16074 , n16073 , n7440 );
xor ( n16075 , n16070 , n16074 );
xor ( n16076 , n16064 , n16075 );
buf ( n16077 , n15844 );
and ( n16078 , n11784 , n6627 );
and ( n16079 , n12217 , n6272 );
nor ( n16080 , n16078 , n16079 );
xnor ( n16081 , n16080 , n6623 );
xor ( n16082 , n16077 , n16081 );
and ( n16083 , n10534 , n7437 );
xor ( n16084 , n16082 , n16083 );
xor ( n16085 , n16076 , n16084 );
xor ( n16086 , n16060 , n16085 );
xor ( n16087 , n16051 , n16086 );
and ( n16088 , n15853 , n15857 );
and ( n16089 , n15857 , n15862 );
and ( n16090 , n15853 , n15862 );
or ( n16091 , n16088 , n16089 , n16090 );
xor ( n16092 , n16087 , n16091 );
and ( n16093 , n15863 , n15864 );
xor ( n16094 , n16092 , n16093 );
buf ( n16095 , n16094 );
not ( n16096 , n454 );
and ( n16097 , n16096 , n16047 );
and ( n16098 , n16095 , n454 );
or ( n16099 , n16097 , n16098 );
buf ( n16100 , n16099 );
buf ( n16101 , n16100 );
and ( n16102 , n16101 , n4505 );
xor ( n16103 , n15983 , n16102 );
and ( n16104 , n15875 , n15876 );
and ( n16105 , n15876 , n15878 );
and ( n16106 , n15875 , n15878 );
or ( n16107 , n16104 , n16105 , n16106 );
and ( n16108 , n15872 , n4557 );
xor ( n16109 , n16107 , n16108 );
xor ( n16110 , n16103 , n16109 );
and ( n16111 , n15744 , n15873 );
and ( n16112 , n15873 , n15879 );
and ( n16113 , n15744 , n15879 );
or ( n16114 , n16111 , n16112 , n16113 );
xor ( n16115 , n16110 , n16114 );
and ( n16116 , n15880 , n15884 );
and ( n16117 , n15884 , n15889 );
and ( n16118 , n15880 , n15889 );
or ( n16119 , n16116 , n16117 , n16118 );
xor ( n16120 , n16115 , n16119 );
or ( n16121 , n15890 , n15891 );
xor ( n16122 , n16120 , n16121 );
not ( n16123 , n16122 );
and ( n16124 , n15892 , n15893 );
xor ( n16125 , n16123 , n16124 );
buf ( n16126 , n16125 );
not ( n16127 , n4509 );
and ( n16128 , n16127 , n15980 );
and ( n16129 , n16126 , n4509 );
or ( n16130 , n16128 , n16129 );
not ( n16131 , n4934 );
and ( n16132 , n11163 , n9407 );
and ( n16133 , n11569 , n8872 );
nor ( n16134 , n16132 , n16133 );
xnor ( n16135 , n16134 , n9403 );
xor ( n16136 , n16131 , n16135 );
and ( n16137 , n10287 , n10329 );
and ( n16138 , n10706 , n9791 );
nor ( n16139 , n16137 , n16138 );
not ( n16140 , n16139 );
xor ( n16141 , n16136 , n16140 );
and ( n16142 , n14865 , n5441 );
and ( n16143 , n15161 , n5161 );
nor ( n16144 , n16142 , n16143 );
xnor ( n16145 , n16144 , n5437 );
and ( n16146 , n14212 , n6068 );
and ( n16147 , n14558 , n5730 );
nor ( n16148 , n16146 , n16147 );
xnor ( n16149 , n16148 , n6064 );
xor ( n16150 , n16145 , n16149 );
and ( n16151 , n13506 , n6711 );
and ( n16152 , n13865 , n6332 );
nor ( n16153 , n16151 , n16152 );
xnor ( n16154 , n16153 , n6707 );
xor ( n16155 , n16150 , n16154 );
xor ( n16156 , n16141 , n16155 );
and ( n16157 , n15933 , n15937 );
and ( n16158 , n15937 , n15942 );
and ( n16159 , n15933 , n15942 );
or ( n16160 , n16157 , n16158 , n16159 );
xor ( n16161 , n16156 , n16160 );
not ( n16162 , n15950 );
buf ( n16163 , n16162 );
and ( n16164 , n12754 , n7630 );
and ( n16165 , n13144 , n7188 );
nor ( n16166 , n16164 , n16165 );
xnor ( n16167 , n16166 , n7626 );
xor ( n16168 , n16163 , n16167 );
and ( n16169 , n11989 , n8502 );
and ( n16170 , n12392 , n7970 );
nor ( n16171 , n16169 , n16170 );
xnor ( n16172 , n16171 , n8498 );
xor ( n16173 , n16168 , n16172 );
xor ( n16174 , n16161 , n16173 );
and ( n16175 , n15911 , n15924 );
and ( n16176 , n15924 , n15944 );
and ( n16177 , n15911 , n15944 );
or ( n16178 , n16175 , n16176 , n16177 );
xor ( n16179 , n16174 , n16178 );
and ( n16180 , n15951 , n15955 );
and ( n16181 , n15955 , n15960 );
and ( n16182 , n15951 , n15960 );
or ( n16183 , n16180 , n16181 , n16182 );
and ( n16184 , n15914 , n15918 );
and ( n16185 , n15918 , n15923 );
and ( n16186 , n15914 , n15923 );
or ( n16187 , n16184 , n16185 , n16186 );
and ( n16188 , n15929 , n15943 );
xor ( n16189 , n16187 , n16188 );
and ( n16190 , n15947 , n15950 );
xor ( n16191 , n16189 , n16190 );
xor ( n16192 , n16183 , n16191 );
and ( n16193 , n15907 , n15945 );
and ( n16194 , n15945 , n15961 );
and ( n16195 , n15907 , n15961 );
or ( n16196 , n16193 , n16194 , n16195 );
xor ( n16197 , n16192 , n16196 );
xor ( n16198 , n16179 , n16197 );
and ( n16199 , n15903 , n15962 );
and ( n16200 , n15962 , n15967 );
and ( n16201 , n15903 , n15967 );
or ( n16202 , n16199 , n16200 , n16201 );
xor ( n16203 , n16198 , n16202 );
and ( n16204 , n15968 , n15969 );
and ( n16205 , n15969 , n15974 );
and ( n16206 , n15968 , n15974 );
or ( n16207 , n16204 , n16205 , n16206 );
xor ( n16208 , n16203 , n16207 );
and ( n16209 , n15975 , n15978 );
xor ( n16210 , n16208 , n16209 );
buf ( n16211 , n16210 );
and ( n16212 , n16107 , n16108 );
and ( n16213 , n15991 , n15995 );
and ( n16214 , n15995 , n16007 );
and ( n16215 , n15991 , n16007 );
or ( n16216 , n16213 , n16214 , n16215 );
and ( n16217 , n16013 , n16017 );
and ( n16218 , n16017 , n16032 );
and ( n16219 , n16013 , n16032 );
or ( n16220 , n16217 , n16218 , n16219 );
xor ( n16221 , n16216 , n16220 );
and ( n16222 , n16021 , n16025 );
and ( n16223 , n16025 , n16031 );
and ( n16224 , n16021 , n16031 );
or ( n16225 , n16222 , n16223 , n16224 );
and ( n16226 , n13647 , n5270 );
and ( n16227 , n14013 , n5021 );
nor ( n16228 , n16226 , n16227 );
xnor ( n16229 , n16228 , n5266 );
and ( n16230 , n12895 , n5850 );
and ( n16231 , n13313 , n5566 );
nor ( n16232 , n16230 , n16231 );
xnor ( n16233 , n16232 , n5846 );
xor ( n16234 , n16229 , n16233 );
and ( n16235 , n11295 , n7356 );
and ( n16236 , n11702 , n6953 );
nor ( n16237 , n16235 , n16236 );
xnor ( n16238 , n16237 , n7352 );
xor ( n16239 , n16234 , n16238 );
xor ( n16240 , n16225 , n16239 );
and ( n16241 , n16000 , n16004 );
and ( n16242 , n16004 , n16006 );
and ( n16243 , n16000 , n16006 );
or ( n16244 , n16241 , n16242 , n16243 );
buf ( n16245 , n16030 );
xor ( n16246 , n16244 , n16245 );
not ( n16247 , n4784 );
and ( n16248 , n12116 , n6554 );
and ( n16249 , n12527 , n6205 );
nor ( n16250 , n16248 , n16249 );
xnor ( n16251 , n16250 , n6550 );
xor ( n16252 , n16247 , n16251 );
and ( n16253 , n10857 , n7349 );
xor ( n16254 , n16252 , n16253 );
xor ( n16255 , n16246 , n16254 );
xor ( n16256 , n16240 , n16255 );
xor ( n16257 , n16221 , n16256 );
and ( n16258 , n15987 , n16008 );
and ( n16259 , n16008 , n16033 );
and ( n16260 , n15987 , n16033 );
or ( n16261 , n16258 , n16259 , n16260 );
xor ( n16262 , n16257 , n16261 );
and ( n16263 , n16034 , n16038 );
and ( n16264 , n16038 , n16043 );
and ( n16265 , n16034 , n16043 );
or ( n16266 , n16263 , n16264 , n16265 );
xor ( n16267 , n16262 , n16266 );
and ( n16268 , n16044 , n16045 );
xor ( n16269 , n16267 , n16268 );
buf ( n16270 , n16269 );
and ( n16271 , n16077 , n16081 );
and ( n16272 , n16081 , n16083 );
and ( n16273 , n16077 , n16083 );
or ( n16274 , n16271 , n16272 , n16273 );
and ( n16275 , n16064 , n16075 );
and ( n16276 , n16075 , n16084 );
and ( n16277 , n16064 , n16084 );
or ( n16278 , n16275 , n16276 , n16277 );
xor ( n16279 , n16274 , n16278 );
and ( n16280 , n16065 , n16069 );
and ( n16281 , n16069 , n16074 );
and ( n16282 , n16065 , n16074 );
or ( n16283 , n16280 , n16281 , n16282 );
and ( n16284 , n12976 , n5922 );
not ( n16285 , n16284 );
xnor ( n16286 , n16285 , n5918 );
not ( n16287 , n16286 );
xor ( n16288 , n16283 , n16287 );
and ( n16289 , n12217 , n6627 );
and ( n16290 , n12612 , n6272 );
nor ( n16291 , n16289 , n16290 );
xnor ( n16292 , n16291 , n6623 );
and ( n16293 , n11398 , n7444 );
and ( n16294 , n11784 , n7026 );
nor ( n16295 , n16293 , n16294 );
xnor ( n16296 , n16295 , n7440 );
xor ( n16297 , n16292 , n16296 );
and ( n16298 , n10940 , n7437 );
xor ( n16299 , n16297 , n16298 );
xor ( n16300 , n16288 , n16299 );
xor ( n16301 , n16279 , n16300 );
and ( n16302 , n16055 , n16059 );
and ( n16303 , n16059 , n16085 );
and ( n16304 , n16055 , n16085 );
or ( n16305 , n16302 , n16303 , n16304 );
xor ( n16306 , n16301 , n16305 );
and ( n16307 , n16051 , n16086 );
and ( n16308 , n16086 , n16091 );
and ( n16309 , n16051 , n16091 );
or ( n16310 , n16307 , n16308 , n16309 );
xor ( n16311 , n16306 , n16310 );
and ( n16312 , n16092 , n16093 );
xor ( n16313 , n16311 , n16312 );
buf ( n16314 , n16313 );
not ( n16315 , n454 );
and ( n16316 , n16315 , n16270 );
and ( n16317 , n16314 , n454 );
or ( n16318 , n16316 , n16317 );
buf ( n16319 , n16318 );
buf ( n16320 , n16319 );
and ( n16321 , n16320 , n4505 );
and ( n16322 , n15632 , n5089 );
and ( n16323 , n15872 , n4866 );
xor ( n16324 , n16322 , n16323 );
and ( n16325 , n16101 , n4557 );
xor ( n16326 , n16324 , n16325 );
xor ( n16327 , n16321 , n16326 );
and ( n16328 , n15981 , n15982 );
and ( n16329 , n15982 , n16102 );
and ( n16330 , n15981 , n16102 );
or ( n16331 , n16328 , n16329 , n16330 );
xor ( n16332 , n16327 , n16331 );
xor ( n16333 , n16212 , n16332 );
and ( n16334 , n16103 , n16109 );
and ( n16335 , n16109 , n16114 );
and ( n16336 , n16103 , n16114 );
or ( n16337 , n16334 , n16335 , n16336 );
xor ( n16338 , n16333 , n16337 );
and ( n16339 , n16115 , n16119 );
and ( n16340 , n16119 , n16121 );
and ( n16341 , n16115 , n16121 );
or ( n16342 , n16339 , n16340 , n16341 );
xnor ( n16343 , n16338 , n16342 );
and ( n16344 , n16123 , n16124 );
or ( n16345 , n16122 , n16344 );
xor ( n16346 , n16343 , n16345 );
buf ( n16347 , n16346 );
not ( n16348 , n4509 );
and ( n16349 , n16348 , n16211 );
and ( n16350 , n16347 , n4509 );
or ( n16351 , n16349 , n16350 );
and ( n16352 , n16183 , n16191 );
and ( n16353 , n16191 , n16196 );
and ( n16354 , n16183 , n16196 );
or ( n16355 , n16352 , n16353 , n16354 );
and ( n16356 , n16163 , n16167 );
and ( n16357 , n16167 , n16172 );
and ( n16358 , n16163 , n16172 );
or ( n16359 , n16356 , n16357 , n16358 );
and ( n16360 , n14558 , n6068 );
and ( n16361 , n14865 , n5730 );
nor ( n16362 , n16360 , n16361 );
xnor ( n16363 , n16362 , n6064 );
xor ( n16364 , n16359 , n16363 );
and ( n16365 , n13865 , n6711 );
and ( n16366 , n14212 , n6332 );
nor ( n16367 , n16365 , n16366 );
xnor ( n16368 , n16367 , n6707 );
xor ( n16369 , n16364 , n16368 );
and ( n16370 , n16161 , n16173 );
and ( n16371 , n16173 , n16178 );
and ( n16372 , n16161 , n16178 );
or ( n16373 , n16370 , n16371 , n16372 );
xor ( n16374 , n16369 , n16373 );
and ( n16375 , n16141 , n16155 );
and ( n16376 , n16155 , n16160 );
and ( n16377 , n16141 , n16160 );
or ( n16378 , n16375 , n16376 , n16377 );
and ( n16379 , n16145 , n16149 );
and ( n16380 , n16149 , n16154 );
and ( n16381 , n16145 , n16154 );
or ( n16382 , n16379 , n16380 , n16381 );
and ( n16383 , n16131 , n16135 );
and ( n16384 , n16135 , n16140 );
and ( n16385 , n16131 , n16140 );
or ( n16386 , n16383 , n16384 , n16385 );
and ( n16387 , n15161 , n5441 );
not ( n16388 , n16387 );
xnor ( n16389 , n16388 , n5437 );
xor ( n16390 , n16386 , n16389 );
and ( n16391 , n13144 , n7630 );
and ( n16392 , n13506 , n7188 );
nor ( n16393 , n16391 , n16392 );
xnor ( n16394 , n16393 , n7626 );
xor ( n16395 , n16390 , n16394 );
xor ( n16396 , n16382 , n16395 );
and ( n16397 , n12392 , n8502 );
and ( n16398 , n12754 , n7970 );
nor ( n16399 , n16397 , n16398 );
xnor ( n16400 , n16399 , n8498 );
and ( n16401 , n11569 , n9407 );
and ( n16402 , n11989 , n8872 );
nor ( n16403 , n16401 , n16402 );
xnor ( n16404 , n16403 , n9403 );
xor ( n16405 , n16400 , n16404 );
and ( n16406 , n10706 , n10329 );
and ( n16407 , n11163 , n9791 );
nor ( n16408 , n16406 , n16407 );
xor ( n16409 , n16405 , n16408 );
xor ( n16410 , n16396 , n16409 );
xor ( n16411 , n16378 , n16410 );
and ( n16412 , n16187 , n16188 );
and ( n16413 , n16188 , n16190 );
and ( n16414 , n16187 , n16190 );
or ( n16415 , n16412 , n16413 , n16414 );
xor ( n16416 , n16411 , n16415 );
xor ( n16417 , n16374 , n16416 );
xor ( n16418 , n16355 , n16417 );
and ( n16419 , n16179 , n16197 );
and ( n16420 , n16197 , n16202 );
and ( n16421 , n16179 , n16202 );
or ( n16422 , n16419 , n16420 , n16421 );
xor ( n16423 , n16418 , n16422 );
and ( n16424 , n16203 , n16207 );
and ( n16425 , n16208 , n16209 );
or ( n16426 , n16424 , n16425 );
xor ( n16427 , n16423 , n16426 );
buf ( n16428 , n16427 );
and ( n16429 , n15872 , n5089 );
and ( n16430 , n16101 , n4866 );
xor ( n16431 , n16429 , n16430 );
and ( n16432 , n16225 , n16239 );
and ( n16433 , n16239 , n16255 );
and ( n16434 , n16225 , n16255 );
or ( n16435 , n16432 , n16433 , n16434 );
and ( n16436 , n16247 , n16251 );
and ( n16437 , n16251 , n16253 );
and ( n16438 , n16247 , n16253 );
or ( n16439 , n16436 , n16437 , n16438 );
and ( n16440 , n14013 , n5270 );
not ( n16441 , n16440 );
xnor ( n16442 , n16441 , n5266 );
xor ( n16443 , n16439 , n16442 );
and ( n16444 , n11295 , n7349 );
not ( n16445 , n16444 );
xor ( n16446 , n16443 , n16445 );
xor ( n16447 , n16435 , n16446 );
and ( n16448 , n16229 , n16233 );
and ( n16449 , n16233 , n16238 );
and ( n16450 , n16229 , n16238 );
or ( n16451 , n16448 , n16449 , n16450 );
and ( n16452 , n16244 , n16245 );
and ( n16453 , n16245 , n16254 );
and ( n16454 , n16244 , n16254 );
or ( n16455 , n16452 , n16453 , n16454 );
xor ( n16456 , n16451 , n16455 );
and ( n16457 , n13313 , n5850 );
and ( n16458 , n13647 , n5566 );
nor ( n16459 , n16457 , n16458 );
xnor ( n16460 , n16459 , n5846 );
and ( n16461 , n12527 , n6554 );
and ( n16462 , n12895 , n6205 );
nor ( n16463 , n16461 , n16462 );
xnor ( n16464 , n16463 , n6550 );
xor ( n16465 , n16460 , n16464 );
and ( n16466 , n11702 , n7356 );
and ( n16467 , n12116 , n6953 );
nor ( n16468 , n16466 , n16467 );
xnor ( n16469 , n16468 , n7352 );
xor ( n16470 , n16465 , n16469 );
xor ( n16471 , n16456 , n16470 );
xor ( n16472 , n16447 , n16471 );
and ( n16473 , n16216 , n16220 );
and ( n16474 , n16220 , n16256 );
and ( n16475 , n16216 , n16256 );
or ( n16476 , n16473 , n16474 , n16475 );
xor ( n16477 , n16472 , n16476 );
and ( n16478 , n16257 , n16261 );
and ( n16479 , n16261 , n16266 );
and ( n16480 , n16257 , n16266 );
or ( n16481 , n16478 , n16479 , n16480 );
xor ( n16482 , n16477 , n16481 );
and ( n16483 , n16267 , n16268 );
xor ( n16484 , n16482 , n16483 );
buf ( n16485 , n16484 );
and ( n16486 , n16283 , n16287 );
and ( n16487 , n16287 , n16299 );
and ( n16488 , n16283 , n16299 );
or ( n16489 , n16486 , n16487 , n16488 );
not ( n16490 , n5918 );
and ( n16491 , n12612 , n6627 );
and ( n16492 , n12976 , n6272 );
nor ( n16493 , n16491 , n16492 );
xnor ( n16494 , n16493 , n6623 );
xor ( n16495 , n16490 , n16494 );
and ( n16496 , n11398 , n7437 );
xor ( n16497 , n16495 , n16496 );
xor ( n16498 , n16489 , n16497 );
and ( n16499 , n16292 , n16296 );
and ( n16500 , n16296 , n16298 );
and ( n16501 , n16292 , n16298 );
or ( n16502 , n16499 , n16500 , n16501 );
buf ( n16503 , n16286 );
xor ( n16504 , n16502 , n16503 );
and ( n16505 , n11784 , n7444 );
and ( n16506 , n12217 , n7026 );
nor ( n16507 , n16505 , n16506 );
xnor ( n16508 , n16507 , n7440 );
xor ( n16509 , n16504 , n16508 );
xor ( n16510 , n16498 , n16509 );
and ( n16511 , n16274 , n16278 );
and ( n16512 , n16278 , n16300 );
and ( n16513 , n16274 , n16300 );
or ( n16514 , n16511 , n16512 , n16513 );
xor ( n16515 , n16510 , n16514 );
and ( n16516 , n16301 , n16305 );
and ( n16517 , n16305 , n16310 );
and ( n16518 , n16301 , n16310 );
or ( n16519 , n16516 , n16517 , n16518 );
xor ( n16520 , n16515 , n16519 );
and ( n16521 , n16311 , n16312 );
xor ( n16522 , n16520 , n16521 );
buf ( n16523 , n16522 );
not ( n16524 , n454 );
and ( n16525 , n16524 , n16485 );
and ( n16526 , n16523 , n454 );
or ( n16527 , n16525 , n16526 );
buf ( n16528 , n16527 );
buf ( n16529 , n16528 );
and ( n16530 , n16529 , n4505 );
xor ( n16531 , n16431 , n16530 );
and ( n16532 , n16322 , n16323 );
and ( n16533 , n16323 , n16325 );
and ( n16534 , n16322 , n16325 );
or ( n16535 , n16532 , n16533 , n16534 );
and ( n16536 , n16320 , n4557 );
xor ( n16537 , n16535 , n16536 );
xor ( n16538 , n16531 , n16537 );
and ( n16539 , n16321 , n16326 );
and ( n16540 , n16326 , n16331 );
and ( n16541 , n16321 , n16331 );
or ( n16542 , n16539 , n16540 , n16541 );
xor ( n16543 , n16538 , n16542 );
and ( n16544 , n16212 , n16332 );
and ( n16545 , n16332 , n16337 );
and ( n16546 , n16212 , n16337 );
or ( n16547 , n16544 , n16545 , n16546 );
xor ( n16548 , n16543 , n16547 );
or ( n16549 , n16338 , n16342 );
xor ( n16550 , n16548 , n16549 );
not ( n16551 , n16550 );
and ( n16552 , n16343 , n16345 );
xor ( n16553 , n16551 , n16552 );
buf ( n16554 , n16553 );
not ( n16555 , n4509 );
and ( n16556 , n16555 , n16428 );
and ( n16557 , n16554 , n4509 );
or ( n16558 , n16556 , n16557 );
and ( n16559 , n16369 , n16373 );
and ( n16560 , n16373 , n16416 );
and ( n16561 , n16369 , n16416 );
or ( n16562 , n16559 , n16560 , n16561 );
and ( n16563 , n16386 , n16389 );
and ( n16564 , n16389 , n16394 );
and ( n16565 , n16386 , n16394 );
or ( n16566 , n16563 , n16564 , n16565 );
not ( n16567 , n5437 );
and ( n16568 , n12754 , n8502 );
and ( n16569 , n13144 , n7970 );
nor ( n16570 , n16568 , n16569 );
xnor ( n16571 , n16570 , n8498 );
xor ( n16572 , n16567 , n16571 );
and ( n16573 , n11163 , n10329 );
and ( n16574 , n11569 , n9791 );
nor ( n16575 , n16573 , n16574 );
not ( n16576 , n16575 );
xor ( n16577 , n16572 , n16576 );
xor ( n16578 , n16566 , n16577 );
not ( n16579 , n16408 );
buf ( n16580 , n16579 );
and ( n16581 , n13506 , n7630 );
and ( n16582 , n13865 , n7188 );
nor ( n16583 , n16581 , n16582 );
xnor ( n16584 , n16583 , n7626 );
xor ( n16585 , n16580 , n16584 );
and ( n16586 , n11989 , n9407 );
and ( n16587 , n12392 , n8872 );
nor ( n16588 , n16586 , n16587 );
xnor ( n16589 , n16588 , n9403 );
xor ( n16590 , n16585 , n16589 );
xor ( n16591 , n16578 , n16590 );
and ( n16592 , n16378 , n16410 );
and ( n16593 , n16410 , n16415 );
and ( n16594 , n16378 , n16415 );
or ( n16595 , n16592 , n16593 , n16594 );
xor ( n16596 , n16591 , n16595 );
and ( n16597 , n16359 , n16363 );
and ( n16598 , n16363 , n16368 );
and ( n16599 , n16359 , n16368 );
or ( n16600 , n16597 , n16598 , n16599 );
and ( n16601 , n16382 , n16395 );
and ( n16602 , n16395 , n16409 );
and ( n16603 , n16382 , n16409 );
or ( n16604 , n16601 , n16602 , n16603 );
xor ( n16605 , n16600 , n16604 );
and ( n16606 , n16400 , n16404 );
and ( n16607 , n16404 , n16408 );
and ( n16608 , n16400 , n16408 );
or ( n16609 , n16606 , n16607 , n16608 );
and ( n16610 , n14865 , n6068 );
and ( n16611 , n15161 , n5730 );
nor ( n16612 , n16610 , n16611 );
xnor ( n16613 , n16612 , n6064 );
xor ( n16614 , n16609 , n16613 );
and ( n16615 , n14212 , n6711 );
and ( n16616 , n14558 , n6332 );
nor ( n16617 , n16615 , n16616 );
xnor ( n16618 , n16617 , n6707 );
xor ( n16619 , n16614 , n16618 );
xor ( n16620 , n16605 , n16619 );
xor ( n16621 , n16596 , n16620 );
xor ( n16622 , n16562 , n16621 );
and ( n16623 , n16355 , n16417 );
and ( n16624 , n16417 , n16422 );
and ( n16625 , n16355 , n16422 );
or ( n16626 , n16623 , n16624 , n16625 );
xor ( n16627 , n16622 , n16626 );
and ( n16628 , n16423 , n16426 );
xor ( n16629 , n16627 , n16628 );
buf ( n16630 , n16629 );
and ( n16631 , n16535 , n16536 );
and ( n16632 , n16101 , n5089 );
and ( n16633 , n16320 , n4866 );
xor ( n16634 , n16632 , n16633 );
and ( n16635 , n16529 , n4557 );
xor ( n16636 , n16634 , n16635 );
and ( n16637 , n16435 , n16446 );
and ( n16638 , n16446 , n16471 );
and ( n16639 , n16435 , n16471 );
or ( n16640 , n16637 , n16638 , n16639 );
and ( n16641 , n16439 , n16442 );
and ( n16642 , n16442 , n16445 );
and ( n16643 , n16439 , n16445 );
or ( n16644 , n16641 , n16642 , n16643 );
and ( n16645 , n16451 , n16455 );
and ( n16646 , n16455 , n16470 );
and ( n16647 , n16451 , n16470 );
or ( n16648 , n16645 , n16646 , n16647 );
xor ( n16649 , n16644 , n16648 );
and ( n16650 , n16460 , n16464 );
and ( n16651 , n16464 , n16469 );
and ( n16652 , n16460 , n16469 );
or ( n16653 , n16650 , n16651 , n16652 );
not ( n16654 , n5266 );
and ( n16655 , n12116 , n7356 );
and ( n16656 , n12527 , n6953 );
nor ( n16657 , n16655 , n16656 );
xnor ( n16658 , n16657 , n7352 );
xor ( n16659 , n16654 , n16658 );
and ( n16660 , n11702 , n7349 );
xor ( n16661 , n16659 , n16660 );
xor ( n16662 , n16653 , n16661 );
buf ( n16663 , n16444 );
and ( n16664 , n13647 , n5850 );
and ( n16665 , n14013 , n5566 );
nor ( n16666 , n16664 , n16665 );
xnor ( n16667 , n16666 , n5846 );
xor ( n16668 , n16663 , n16667 );
and ( n16669 , n12895 , n6554 );
and ( n16670 , n13313 , n6205 );
nor ( n16671 , n16669 , n16670 );
xnor ( n16672 , n16671 , n6550 );
xor ( n16673 , n16668 , n16672 );
xor ( n16674 , n16662 , n16673 );
xor ( n16675 , n16649 , n16674 );
xor ( n16676 , n16640 , n16675 );
and ( n16677 , n16472 , n16476 );
and ( n16678 , n16476 , n16481 );
and ( n16679 , n16472 , n16481 );
or ( n16680 , n16677 , n16678 , n16679 );
xor ( n16681 , n16676 , n16680 );
and ( n16682 , n16482 , n16483 );
xor ( n16683 , n16681 , n16682 );
buf ( n16684 , n16683 );
and ( n16685 , n16490 , n16494 );
and ( n16686 , n16494 , n16496 );
and ( n16687 , n16490 , n16496 );
or ( n16688 , n16685 , n16686 , n16687 );
and ( n16689 , n16502 , n16503 );
and ( n16690 , n16503 , n16508 );
and ( n16691 , n16502 , n16508 );
or ( n16692 , n16689 , n16690 , n16691 );
xor ( n16693 , n16688 , n16692 );
and ( n16694 , n12976 , n6627 );
not ( n16695 , n16694 );
xnor ( n16696 , n16695 , n6623 );
not ( n16697 , n16696 );
and ( n16698 , n12217 , n7444 );
and ( n16699 , n12612 , n7026 );
nor ( n16700 , n16698 , n16699 );
xnor ( n16701 , n16700 , n7440 );
xor ( n16702 , n16697 , n16701 );
and ( n16703 , n11784 , n7437 );
xor ( n16704 , n16702 , n16703 );
xor ( n16705 , n16693 , n16704 );
and ( n16706 , n16489 , n16497 );
and ( n16707 , n16497 , n16509 );
and ( n16708 , n16489 , n16509 );
or ( n16709 , n16706 , n16707 , n16708 );
xor ( n16710 , n16705 , n16709 );
and ( n16711 , n16510 , n16514 );
and ( n16712 , n16514 , n16519 );
and ( n16713 , n16510 , n16519 );
or ( n16714 , n16711 , n16712 , n16713 );
xor ( n16715 , n16710 , n16714 );
and ( n16716 , n16520 , n16521 );
xor ( n16717 , n16715 , n16716 );
buf ( n16718 , n16717 );
not ( n16719 , n454 );
and ( n16720 , n16719 , n16684 );
and ( n16721 , n16718 , n454 );
or ( n16722 , n16720 , n16721 );
buf ( n16723 , n16722 );
buf ( n16724 , n16723 );
and ( n16725 , n16724 , n4505 );
not ( n16726 , n16725 );
xor ( n16727 , n16636 , n16726 );
and ( n16728 , n16429 , n16430 );
and ( n16729 , n16430 , n16530 );
and ( n16730 , n16429 , n16530 );
or ( n16731 , n16728 , n16729 , n16730 );
xor ( n16732 , n16727 , n16731 );
xor ( n16733 , n16631 , n16732 );
and ( n16734 , n16531 , n16537 );
and ( n16735 , n16537 , n16542 );
and ( n16736 , n16531 , n16542 );
or ( n16737 , n16734 , n16735 , n16736 );
xor ( n16738 , n16733 , n16737 );
and ( n16739 , n16543 , n16547 );
and ( n16740 , n16547 , n16549 );
and ( n16741 , n16543 , n16549 );
or ( n16742 , n16739 , n16740 , n16741 );
xor ( n16743 , n16738 , n16742 );
and ( n16744 , n16551 , n16552 );
or ( n16745 , n16550 , n16744 );
xor ( n16746 , n16743 , n16745 );
buf ( n16747 , n16746 );
not ( n16748 , n4509 );
and ( n16749 , n16748 , n16630 );
and ( n16750 , n16747 , n4509 );
or ( n16751 , n16749 , n16750 );
and ( n16752 , n16600 , n16604 );
and ( n16753 , n16604 , n16619 );
and ( n16754 , n16600 , n16619 );
or ( n16755 , n16752 , n16753 , n16754 );
and ( n16756 , n16567 , n16571 );
and ( n16757 , n16571 , n16576 );
and ( n16758 , n16567 , n16576 );
or ( n16759 , n16756 , n16757 , n16758 );
and ( n16760 , n16580 , n16584 );
and ( n16761 , n16584 , n16589 );
and ( n16762 , n16580 , n16589 );
or ( n16763 , n16760 , n16761 , n16762 );
xor ( n16764 , n16759 , n16763 );
and ( n16765 , n14558 , n6711 );
and ( n16766 , n14865 , n6332 );
nor ( n16767 , n16765 , n16766 );
xnor ( n16768 , n16767 , n6707 );
and ( n16769 , n13865 , n7630 );
and ( n16770 , n14212 , n7188 );
nor ( n16771 , n16769 , n16770 );
xnor ( n16772 , n16771 , n7626 );
xor ( n16773 , n16768 , n16772 );
and ( n16774 , n12392 , n9407 );
and ( n16775 , n12754 , n8872 );
nor ( n16776 , n16774 , n16775 );
xnor ( n16777 , n16776 , n9403 );
not ( n16778 , n16777 );
xor ( n16779 , n16773 , n16778 );
xor ( n16780 , n16764 , n16779 );
xor ( n16781 , n16755 , n16780 );
and ( n16782 , n16609 , n16613 );
and ( n16783 , n16613 , n16618 );
and ( n16784 , n16609 , n16618 );
or ( n16785 , n16782 , n16783 , n16784 );
and ( n16786 , n16566 , n16577 );
and ( n16787 , n16577 , n16590 );
and ( n16788 , n16566 , n16590 );
or ( n16789 , n16786 , n16787 , n16788 );
xor ( n16790 , n16785 , n16789 );
and ( n16791 , n15161 , n6068 );
not ( n16792 , n16791 );
xnor ( n16793 , n16792 , n6064 );
and ( n16794 , n13144 , n8502 );
and ( n16795 , n13506 , n7970 );
nor ( n16796 , n16794 , n16795 );
xnor ( n16797 , n16796 , n8498 );
xor ( n16798 , n16793 , n16797 );
and ( n16799 , n11569 , n10329 );
and ( n16800 , n11989 , n9791 );
nor ( n16801 , n16799 , n16800 );
not ( n16802 , n16801 );
xor ( n16803 , n16798 , n16802 );
xor ( n16804 , n16790 , n16803 );
xor ( n16805 , n16781 , n16804 );
and ( n16806 , n16591 , n16595 );
and ( n16807 , n16595 , n16620 );
and ( n16808 , n16591 , n16620 );
or ( n16809 , n16806 , n16807 , n16808 );
xor ( n16810 , n16805 , n16809 );
and ( n16811 , n16562 , n16621 );
and ( n16812 , n16621 , n16626 );
and ( n16813 , n16562 , n16626 );
or ( n16814 , n16811 , n16812 , n16813 );
xor ( n16815 , n16810 , n16814 );
and ( n16816 , n16627 , n16628 );
xor ( n16817 , n16815 , n16816 );
buf ( n16818 , n16817 );
buf ( n16819 , n16725 );
and ( n16820 , n16632 , n16633 );
and ( n16821 , n16633 , n16635 );
and ( n16822 , n16632 , n16635 );
or ( n16823 , n16820 , n16821 , n16822 );
and ( n16824 , n16724 , n4557 );
xor ( n16825 , n16823 , n16824 );
and ( n16826 , n16320 , n5089 );
and ( n16827 , n16529 , n4866 );
xor ( n16828 , n16826 , n16827 );
and ( n16829 , n16653 , n16661 );
and ( n16830 , n16661 , n16673 );
and ( n16831 , n16653 , n16673 );
or ( n16832 , n16829 , n16830 , n16831 );
and ( n16833 , n14013 , n5850 );
not ( n16834 , n16833 );
xnor ( n16835 , n16834 , n5846 );
and ( n16836 , n13313 , n6554 );
and ( n16837 , n13647 , n6205 );
nor ( n16838 , n16836 , n16837 );
xnor ( n16839 , n16838 , n6550 );
xor ( n16840 , n16835 , n16839 );
and ( n16841 , n12116 , n7349 );
xor ( n16842 , n16840 , n16841 );
xor ( n16843 , n16832 , n16842 );
and ( n16844 , n16654 , n16658 );
and ( n16845 , n16658 , n16660 );
and ( n16846 , n16654 , n16660 );
or ( n16847 , n16844 , n16845 , n16846 );
and ( n16848 , n16663 , n16667 );
and ( n16849 , n16667 , n16672 );
and ( n16850 , n16663 , n16672 );
or ( n16851 , n16848 , n16849 , n16850 );
xor ( n16852 , n16847 , n16851 );
and ( n16853 , n12527 , n7356 );
and ( n16854 , n12895 , n6953 );
nor ( n16855 , n16853 , n16854 );
xnor ( n16856 , n16855 , n7352 );
not ( n16857 , n16856 );
xor ( n16858 , n16852 , n16857 );
xor ( n16859 , n16843 , n16858 );
and ( n16860 , n16644 , n16648 );
and ( n16861 , n16648 , n16674 );
and ( n16862 , n16644 , n16674 );
or ( n16863 , n16860 , n16861 , n16862 );
xor ( n16864 , n16859 , n16863 );
and ( n16865 , n16640 , n16675 );
and ( n16866 , n16675 , n16680 );
and ( n16867 , n16640 , n16680 );
or ( n16868 , n16865 , n16866 , n16867 );
xor ( n16869 , n16864 , n16868 );
and ( n16870 , n16681 , n16682 );
xor ( n16871 , n16869 , n16870 );
buf ( n16872 , n16871 );
and ( n16873 , n16697 , n16701 );
and ( n16874 , n16701 , n16703 );
and ( n16875 , n16697 , n16703 );
or ( n16876 , n16873 , n16874 , n16875 );
buf ( n16877 , n16696 );
xor ( n16878 , n16876 , n16877 );
not ( n16879 , n6623 );
and ( n16880 , n12612 , n7444 );
and ( n16881 , n12976 , n7026 );
nor ( n16882 , n16880 , n16881 );
xnor ( n16883 , n16882 , n7440 );
xor ( n16884 , n16879 , n16883 );
and ( n16885 , n12217 , n7437 );
xor ( n16886 , n16884 , n16885 );
xor ( n16887 , n16878 , n16886 );
and ( n16888 , n16688 , n16692 );
and ( n16889 , n16692 , n16704 );
and ( n16890 , n16688 , n16704 );
or ( n16891 , n16888 , n16889 , n16890 );
xor ( n16892 , n16887 , n16891 );
and ( n16893 , n16705 , n16709 );
and ( n16894 , n16709 , n16714 );
and ( n16895 , n16705 , n16714 );
or ( n16896 , n16893 , n16894 , n16895 );
xor ( n16897 , n16892 , n16896 );
and ( n16898 , n16715 , n16716 );
xor ( n16899 , n16897 , n16898 );
buf ( n16900 , n16899 );
not ( n16901 , n454 );
and ( n16902 , n16901 , n16872 );
and ( n16903 , n16900 , n454 );
or ( n16904 , n16902 , n16903 );
buf ( n16905 , n16904 );
buf ( n16906 , n16905 );
and ( n16907 , n16906 , n4505 );
xor ( n16908 , n16828 , n16907 );
xor ( n16909 , n16825 , n16908 );
xor ( n16910 , n16819 , n16909 );
and ( n16911 , n16636 , n16726 );
and ( n16912 , n16726 , n16731 );
and ( n16913 , n16636 , n16731 );
or ( n16914 , n16911 , n16912 , n16913 );
xor ( n16915 , n16910 , n16914 );
and ( n16916 , n16631 , n16732 );
and ( n16917 , n16732 , n16737 );
and ( n16918 , n16631 , n16737 );
or ( n16919 , n16916 , n16917 , n16918 );
xnor ( n16920 , n16915 , n16919 );
and ( n16921 , n16738 , n16742 );
and ( n16922 , n16743 , n16745 );
or ( n16923 , n16921 , n16922 );
xor ( n16924 , n16920 , n16923 );
buf ( n16925 , n16924 );
not ( n16926 , n4509 );
and ( n16927 , n16926 , n16818 );
and ( n16928 , n16925 , n4509 );
or ( n16929 , n16927 , n16928 );
and ( n16930 , n16759 , n16763 );
and ( n16931 , n16763 , n16779 );
and ( n16932 , n16759 , n16779 );
or ( n16933 , n16930 , n16931 , n16932 );
and ( n16934 , n16785 , n16789 );
and ( n16935 , n16789 , n16803 );
and ( n16936 , n16785 , n16803 );
or ( n16937 , n16934 , n16935 , n16936 );
xor ( n16938 , n16933 , n16937 );
and ( n16939 , n16768 , n16772 );
and ( n16940 , n16772 , n16778 );
and ( n16941 , n16768 , n16778 );
or ( n16942 , n16939 , n16940 , n16941 );
and ( n16943 , n14865 , n6711 );
and ( n16944 , n15161 , n6332 );
nor ( n16945 , n16943 , n16944 );
xnor ( n16946 , n16945 , n6707 );
and ( n16947 , n14212 , n7630 );
and ( n16948 , n14558 , n7188 );
nor ( n16949 , n16947 , n16948 );
xnor ( n16950 , n16949 , n7626 );
xor ( n16951 , n16946 , n16950 );
and ( n16952 , n13506 , n8502 );
and ( n16953 , n13865 , n7970 );
nor ( n16954 , n16952 , n16953 );
xnor ( n16955 , n16954 , n8498 );
xor ( n16956 , n16951 , n16955 );
xor ( n16957 , n16942 , n16956 );
and ( n16958 , n16793 , n16797 );
and ( n16959 , n16797 , n16802 );
and ( n16960 , n16793 , n16802 );
or ( n16961 , n16958 , n16959 , n16960 );
buf ( n16962 , n16777 );
xor ( n16963 , n16961 , n16962 );
not ( n16964 , n6064 );
and ( n16965 , n12754 , n9407 );
and ( n16966 , n13144 , n8872 );
nor ( n16967 , n16965 , n16966 );
xnor ( n16968 , n16967 , n9403 );
xor ( n16969 , n16964 , n16968 );
and ( n16970 , n11989 , n10329 );
and ( n16971 , n12392 , n9791 );
nor ( n16972 , n16970 , n16971 );
not ( n16973 , n16972 );
xor ( n16974 , n16969 , n16973 );
xor ( n16975 , n16963 , n16974 );
xor ( n16976 , n16957 , n16975 );
xor ( n16977 , n16938 , n16976 );
and ( n16978 , n16755 , n16780 );
and ( n16979 , n16780 , n16804 );
and ( n16980 , n16755 , n16804 );
or ( n16981 , n16978 , n16979 , n16980 );
xor ( n16982 , n16977 , n16981 );
and ( n16983 , n16805 , n16809 );
and ( n16984 , n16809 , n16814 );
and ( n16985 , n16805 , n16814 );
or ( n16986 , n16983 , n16984 , n16985 );
xor ( n16987 , n16982 , n16986 );
and ( n16988 , n16815 , n16816 );
xor ( n16989 , n16987 , n16988 );
buf ( n16990 , n16989 );
and ( n16991 , n16826 , n16827 );
and ( n16992 , n16827 , n16907 );
and ( n16993 , n16826 , n16907 );
or ( n16994 , n16991 , n16992 , n16993 );
and ( n16995 , n16832 , n16842 );
and ( n16996 , n16842 , n16858 );
and ( n16997 , n16832 , n16858 );
or ( n16998 , n16995 , n16996 , n16997 );
and ( n16999 , n16835 , n16839 );
and ( n17000 , n16839 , n16841 );
and ( n17001 , n16835 , n16841 );
or ( n17002 , n16999 , n17000 , n17001 );
and ( n17003 , n16847 , n16851 );
and ( n17004 , n16851 , n16857 );
and ( n17005 , n16847 , n16857 );
or ( n17006 , n17003 , n17004 , n17005 );
xor ( n17007 , n17002 , n17006 );
buf ( n17008 , n16856 );
and ( n17009 , n13647 , n6554 );
and ( n17010 , n14013 , n6205 );
nor ( n17011 , n17009 , n17010 );
xnor ( n17012 , n17011 , n6550 );
xor ( n17013 , n17008 , n17012 );
not ( n17014 , n5846 );
and ( n17015 , n12895 , n7356 );
and ( n17016 , n13313 , n6953 );
nor ( n17017 , n17015 , n17016 );
xnor ( n17018 , n17017 , n7352 );
xor ( n17019 , n17014 , n17018 );
and ( n17020 , n12527 , n7349 );
xor ( n17021 , n17019 , n17020 );
xor ( n17022 , n17013 , n17021 );
xor ( n17023 , n17007 , n17022 );
xor ( n17024 , n16998 , n17023 );
and ( n17025 , n16859 , n16863 );
and ( n17026 , n16863 , n16868 );
and ( n17027 , n16859 , n16868 );
or ( n17028 , n17025 , n17026 , n17027 );
xor ( n17029 , n17024 , n17028 );
and ( n17030 , n16869 , n16870 );
xor ( n17031 , n17029 , n17030 );
buf ( n17032 , n17031 );
and ( n17033 , n16879 , n16883 );
and ( n17034 , n16883 , n16885 );
and ( n17035 , n16879 , n16885 );
or ( n17036 , n17033 , n17034 , n17035 );
and ( n17037 , n12976 , n7444 );
not ( n17038 , n17037 );
xnor ( n17039 , n17038 , n7440 );
xor ( n17040 , n17036 , n17039 );
and ( n17041 , n12612 , n7437 );
not ( n17042 , n17041 );
xor ( n17043 , n17040 , n17042 );
and ( n17044 , n16876 , n16877 );
and ( n17045 , n16877 , n16886 );
and ( n17046 , n16876 , n16886 );
or ( n17047 , n17044 , n17045 , n17046 );
xor ( n17048 , n17043 , n17047 );
and ( n17049 , n16887 , n16891 );
and ( n17050 , n16891 , n16896 );
and ( n17051 , n16887 , n16896 );
or ( n17052 , n17049 , n17050 , n17051 );
xor ( n17053 , n17048 , n17052 );
and ( n17054 , n16897 , n16898 );
xor ( n17055 , n17053 , n17054 );
buf ( n17056 , n17055 );
not ( n17057 , n454 );
and ( n17058 , n17057 , n17032 );
and ( n17059 , n17056 , n454 );
or ( n17060 , n17058 , n17059 );
buf ( n17061 , n17060 );
buf ( n17062 , n17061 );
and ( n17063 , n17062 , n4505 );
xor ( n17064 , n16994 , n17063 );
and ( n17065 , n16529 , n5089 );
and ( n17066 , n16724 , n4866 );
xor ( n17067 , n17065 , n17066 );
and ( n17068 , n16906 , n4557 );
xor ( n17069 , n17067 , n17068 );
xor ( n17070 , n17064 , n17069 );
and ( n17071 , n16823 , n16824 );
and ( n17072 , n16824 , n16908 );
and ( n17073 , n16823 , n16908 );
or ( n17074 , n17071 , n17072 , n17073 );
xor ( n17075 , n17070 , n17074 );
and ( n17076 , n16819 , n16909 );
and ( n17077 , n16909 , n16914 );
and ( n17078 , n16819 , n16914 );
or ( n17079 , n17076 , n17077 , n17078 );
xor ( n17080 , n17075 , n17079 );
or ( n17081 , n16915 , n16919 );
xnor ( n17082 , n17080 , n17081 );
and ( n17083 , n16920 , n16923 );
xor ( n17084 , n17082 , n17083 );
buf ( n17085 , n17084 );
not ( n17086 , n4509 );
and ( n17087 , n17086 , n16990 );
and ( n17088 , n17085 , n4509 );
or ( n17089 , n17087 , n17088 );
and ( n17090 , n16961 , n16962 );
and ( n17091 , n16962 , n16974 );
and ( n17092 , n16961 , n16974 );
or ( n17093 , n17090 , n17091 , n17092 );
and ( n17094 , n16942 , n16956 );
and ( n17095 , n16956 , n16975 );
and ( n17096 , n16942 , n16975 );
or ( n17097 , n17094 , n17095 , n17096 );
xor ( n17098 , n17093 , n17097 );
and ( n17099 , n16946 , n16950 );
and ( n17100 , n16950 , n16955 );
and ( n17101 , n16946 , n16955 );
or ( n17102 , n17099 , n17100 , n17101 );
and ( n17103 , n15161 , n6711 );
not ( n17104 , n17103 );
xnor ( n17105 , n17104 , n6707 );
and ( n17106 , n14558 , n7630 );
and ( n17107 , n14865 , n7188 );
nor ( n17108 , n17106 , n17107 );
xnor ( n17109 , n17108 , n7626 );
xor ( n17110 , n17105 , n17109 );
and ( n17111 , n13144 , n9407 );
and ( n17112 , n13506 , n8872 );
nor ( n17113 , n17111 , n17112 );
xnor ( n17114 , n17113 , n9403 );
xor ( n17115 , n17110 , n17114 );
xor ( n17116 , n17102 , n17115 );
and ( n17117 , n16964 , n16968 );
and ( n17118 , n16968 , n16973 );
and ( n17119 , n16964 , n16973 );
or ( n17120 , n17117 , n17118 , n17119 );
and ( n17121 , n13865 , n8502 );
and ( n17122 , n14212 , n7970 );
nor ( n17123 , n17121 , n17122 );
xnor ( n17124 , n17123 , n8498 );
xor ( n17125 , n17120 , n17124 );
and ( n17126 , n12392 , n10329 );
and ( n17127 , n12754 , n9791 );
nor ( n17128 , n17126 , n17127 );
xor ( n17129 , n17125 , n17128 );
xor ( n17130 , n17116 , n17129 );
xor ( n17131 , n17098 , n17130 );
and ( n17132 , n16933 , n16937 );
and ( n17133 , n16937 , n16976 );
and ( n17134 , n16933 , n16976 );
or ( n17135 , n17132 , n17133 , n17134 );
xor ( n17136 , n17131 , n17135 );
and ( n17137 , n16977 , n16981 );
and ( n17138 , n16981 , n16986 );
and ( n17139 , n16977 , n16986 );
or ( n17140 , n17137 , n17138 , n17139 );
xor ( n17141 , n17136 , n17140 );
and ( n17142 , n16987 , n16988 );
xor ( n17143 , n17141 , n17142 );
buf ( n17144 , n17143 );
and ( n17145 , n17065 , n17066 );
and ( n17146 , n17066 , n17068 );
and ( n17147 , n17065 , n17068 );
or ( n17148 , n17145 , n17146 , n17147 );
and ( n17149 , n17062 , n4557 );
xor ( n17150 , n17148 , n17149 );
and ( n17151 , n16724 , n5089 );
and ( n17152 , n16906 , n4866 );
xor ( n17153 , n17151 , n17152 );
and ( n17154 , n17014 , n17018 );
and ( n17155 , n17018 , n17020 );
and ( n17156 , n17014 , n17020 );
or ( n17157 , n17154 , n17155 , n17156 );
and ( n17158 , n17008 , n17012 );
and ( n17159 , n17012 , n17021 );
and ( n17160 , n17008 , n17021 );
or ( n17161 , n17158 , n17159 , n17160 );
xor ( n17162 , n17157 , n17161 );
and ( n17163 , n14013 , n6554 );
not ( n17164 , n17163 );
xnor ( n17165 , n17164 , n6550 );
and ( n17166 , n13313 , n7356 );
and ( n17167 , n13647 , n6953 );
nor ( n17168 , n17166 , n17167 );
xnor ( n17169 , n17168 , n7352 );
xor ( n17170 , n17165 , n17169 );
and ( n17171 , n12895 , n7349 );
not ( n17172 , n17171 );
xor ( n17173 , n17170 , n17172 );
xor ( n17174 , n17162 , n17173 );
and ( n17175 , n17002 , n17006 );
and ( n17176 , n17006 , n17022 );
and ( n17177 , n17002 , n17022 );
or ( n17178 , n17175 , n17176 , n17177 );
xor ( n17179 , n17174 , n17178 );
and ( n17180 , n16998 , n17023 );
and ( n17181 , n17023 , n17028 );
and ( n17182 , n16998 , n17028 );
or ( n17183 , n17180 , n17181 , n17182 );
xor ( n17184 , n17179 , n17183 );
and ( n17185 , n17029 , n17030 );
xor ( n17186 , n17184 , n17185 );
buf ( n17187 , n17186 );
and ( n17188 , n17036 , n17039 );
and ( n17189 , n17039 , n17042 );
and ( n17190 , n17036 , n17042 );
or ( n17191 , n17188 , n17189 , n17190 );
buf ( n17192 , n17041 );
not ( n17193 , n7440 );
xor ( n17194 , n17192 , n17193 );
and ( n17195 , n12976 , n7437 );
xor ( n17196 , n17194 , n17195 );
xor ( n17197 , n17191 , n17196 );
and ( n17198 , n17043 , n17047 );
and ( n17199 , n17047 , n17052 );
and ( n17200 , n17043 , n17052 );
or ( n17201 , n17198 , n17199 , n17200 );
xor ( n17202 , n17197 , n17201 );
and ( n17203 , n17053 , n17054 );
xor ( n17204 , n17202 , n17203 );
buf ( n17205 , n17204 );
not ( n17206 , n454 );
and ( n17207 , n17206 , n17187 );
and ( n17208 , n17205 , n454 );
or ( n17209 , n17207 , n17208 );
buf ( n17210 , n17209 );
buf ( n17211 , n17210 );
and ( n17212 , n17211 , n4505 );
xor ( n17213 , n17153 , n17212 );
xor ( n17214 , n17150 , n17213 );
and ( n17215 , n16994 , n17063 );
and ( n17216 , n17063 , n17069 );
and ( n17217 , n16994 , n17069 );
or ( n17218 , n17215 , n17216 , n17217 );
xor ( n17219 , n17214 , n17218 );
and ( n17220 , n17070 , n17074 );
and ( n17221 , n17074 , n17079 );
and ( n17222 , n17070 , n17079 );
or ( n17223 , n17220 , n17221 , n17222 );
xor ( n17224 , n17219 , n17223 );
or ( n17225 , n17080 , n17081 );
xnor ( n17226 , n17224 , n17225 );
and ( n17227 , n17082 , n17083 );
xor ( n17228 , n17226 , n17227 );
buf ( n17229 , n17228 );
not ( n17230 , n4509 );
and ( n17231 , n17230 , n17144 );
and ( n17232 , n17229 , n4509 );
or ( n17233 , n17231 , n17232 );
and ( n17234 , n17093 , n17097 );
and ( n17235 , n17097 , n17130 );
and ( n17236 , n17093 , n17130 );
or ( n17237 , n17234 , n17235 , n17236 );
and ( n17238 , n17120 , n17124 );
and ( n17239 , n17124 , n17128 );
and ( n17240 , n17120 , n17128 );
or ( n17241 , n17238 , n17239 , n17240 );
and ( n17242 , n17102 , n17115 );
and ( n17243 , n17115 , n17129 );
and ( n17244 , n17102 , n17129 );
or ( n17245 , n17242 , n17243 , n17244 );
xor ( n17246 , n17241 , n17245 );
and ( n17247 , n17105 , n17109 );
and ( n17248 , n17109 , n17114 );
and ( n17249 , n17105 , n17114 );
or ( n17250 , n17247 , n17248 , n17249 );
not ( n17251 , n6707 );
and ( n17252 , n13506 , n9407 );
and ( n17253 , n13865 , n8872 );
nor ( n17254 , n17252 , n17253 );
xnor ( n17255 , n17254 , n9403 );
xor ( n17256 , n17251 , n17255 );
and ( n17257 , n12754 , n10329 );
and ( n17258 , n13144 , n9791 );
nor ( n17259 , n17257 , n17258 );
not ( n17260 , n17259 );
xor ( n17261 , n17256 , n17260 );
xor ( n17262 , n17250 , n17261 );
not ( n17263 , n17128 );
buf ( n17264 , n17263 );
and ( n17265 , n14865 , n7630 );
and ( n17266 , n15161 , n7188 );
nor ( n17267 , n17265 , n17266 );
xnor ( n17268 , n17267 , n7626 );
xor ( n17269 , n17264 , n17268 );
and ( n17270 , n14212 , n8502 );
and ( n17271 , n14558 , n7970 );
nor ( n17272 , n17270 , n17271 );
xnor ( n17273 , n17272 , n8498 );
xor ( n17274 , n17269 , n17273 );
xor ( n17275 , n17262 , n17274 );
xor ( n17276 , n17246 , n17275 );
xor ( n17277 , n17237 , n17276 );
and ( n17278 , n17131 , n17135 );
and ( n17279 , n17135 , n17140 );
and ( n17280 , n17131 , n17140 );
or ( n17281 , n17278 , n17279 , n17280 );
xor ( n17282 , n17277 , n17281 );
and ( n17283 , n17141 , n17142 );
xor ( n17284 , n17282 , n17283 );
buf ( n17285 , n17284 );
and ( n17286 , n16906 , n5089 );
and ( n17287 , n17062 , n4866 );
xor ( n17288 , n17286 , n17287 );
and ( n17289 , n17165 , n17169 );
and ( n17290 , n17169 , n17172 );
and ( n17291 , n17165 , n17172 );
or ( n17292 , n17289 , n17290 , n17291 );
buf ( n17293 , n17171 );
xor ( n17294 , n17292 , n17293 );
not ( n17295 , n6550 );
and ( n17296 , n13647 , n7356 );
and ( n17297 , n14013 , n6953 );
nor ( n17298 , n17296 , n17297 );
xnor ( n17299 , n17298 , n7352 );
xor ( n17300 , n17295 , n17299 );
and ( n17301 , n13313 , n7349 );
xor ( n17302 , n17300 , n17301 );
xor ( n17303 , n17294 , n17302 );
and ( n17304 , n17157 , n17161 );
and ( n17305 , n17161 , n17173 );
and ( n17306 , n17157 , n17173 );
or ( n17307 , n17304 , n17305 , n17306 );
xor ( n17308 , n17303 , n17307 );
and ( n17309 , n17174 , n17178 );
and ( n17310 , n17178 , n17183 );
and ( n17311 , n17174 , n17183 );
or ( n17312 , n17309 , n17310 , n17311 );
xor ( n17313 , n17308 , n17312 );
and ( n17314 , n17184 , n17185 );
xor ( n17315 , n17313 , n17314 );
buf ( n17316 , n17315 );
not ( n17317 , n454 );
and ( n17318 , n17317 , n17316 );
and ( n17319 , C0 , n454 );
or ( n17320 , n17318 , n17319 );
buf ( n17321 , n17320 );
buf ( n17322 , n17321 );
and ( n17323 , n17322 , n4505 );
xor ( n17324 , n17288 , n17323 );
and ( n17325 , n17151 , n17152 );
and ( n17326 , n17152 , n17212 );
and ( n17327 , n17151 , n17212 );
or ( n17328 , n17325 , n17326 , n17327 );
and ( n17329 , n17211 , n4557 );
xor ( n17330 , n17328 , n17329 );
xor ( n17331 , n17324 , n17330 );
and ( n17332 , n17148 , n17149 );
and ( n17333 , n17149 , n17213 );
and ( n17334 , n17148 , n17213 );
or ( n17335 , n17332 , n17333 , n17334 );
xor ( n17336 , n17331 , n17335 );
and ( n17337 , n17214 , n17218 );
and ( n17338 , n17218 , n17223 );
and ( n17339 , n17214 , n17223 );
or ( n17340 , n17337 , n17338 , n17339 );
xor ( n17341 , n17336 , n17340 );
or ( n17342 , n17224 , n17225 );
xor ( n17343 , n17341 , n17342 );
not ( n17344 , n17343 );
and ( n17345 , n17226 , n17227 );
xor ( n17346 , n17344 , n17345 );
buf ( n17347 , n17346 );
not ( n17348 , n4509 );
and ( n17349 , n17348 , n17285 );
and ( n17350 , n17347 , n4509 );
or ( n17351 , n17349 , n17350 );
and ( n17352 , n17250 , n17261 );
and ( n17353 , n17261 , n17274 );
and ( n17354 , n17250 , n17274 );
or ( n17355 , n17352 , n17353 , n17354 );
and ( n17356 , n14558 , n8502 );
and ( n17357 , n14865 , n7970 );
nor ( n17358 , n17356 , n17357 );
xnor ( n17359 , n17358 , n8498 );
and ( n17360 , n13865 , n9407 );
and ( n17361 , n14212 , n8872 );
nor ( n17362 , n17360 , n17361 );
xnor ( n17363 , n17362 , n9403 );
xor ( n17364 , n17359 , n17363 );
and ( n17365 , n13144 , n10329 );
and ( n17366 , n13506 , n9791 );
nor ( n17367 , n17365 , n17366 );
not ( n17368 , n17367 );
xor ( n17369 , n17364 , n17368 );
xor ( n17370 , n17355 , n17369 );
and ( n17371 , n17251 , n17255 );
and ( n17372 , n17255 , n17260 );
and ( n17373 , n17251 , n17260 );
or ( n17374 , n17371 , n17372 , n17373 );
and ( n17375 , n17264 , n17268 );
and ( n17376 , n17268 , n17273 );
and ( n17377 , n17264 , n17273 );
or ( n17378 , n17375 , n17376 , n17377 );
xor ( n17379 , n17374 , n17378 );
and ( n17380 , n15161 , n7630 );
not ( n17381 , n17380 );
xnor ( n17382 , n17381 , n7626 );
not ( n17383 , n17382 );
xor ( n17384 , n17379 , n17383 );
xor ( n17385 , n17370 , n17384 );
and ( n17386 , n17241 , n17245 );
and ( n17387 , n17245 , n17275 );
and ( n17388 , n17241 , n17275 );
or ( n17389 , n17386 , n17387 , n17388 );
xor ( n17390 , n17385 , n17389 );
and ( n17391 , n17237 , n17276 );
and ( n17392 , n17276 , n17281 );
and ( n17393 , n17237 , n17281 );
or ( n17394 , n17391 , n17392 , n17393 );
xor ( n17395 , n17390 , n17394 );
and ( n17396 , n17282 , n17283 );
xor ( n17397 , n17395 , n17396 );
buf ( n17398 , n17397 );
and ( n17399 , n17328 , n17329 );
and ( n17400 , n17211 , n4866 );
not ( n17401 , n17400 );
and ( n17402 , n17286 , n17287 );
and ( n17403 , n17287 , n17323 );
and ( n17404 , n17286 , n17323 );
or ( n17405 , n17402 , n17403 , n17404 );
xor ( n17406 , n17401 , n17405 );
and ( n17407 , n17062 , n5089 );
and ( n17408 , n17322 , n4557 );
xor ( n17409 , n17407 , n17408 );
and ( n17410 , n17295 , n17299 );
and ( n17411 , n17299 , n17301 );
and ( n17412 , n17295 , n17301 );
or ( n17413 , n17410 , n17411 , n17412 );
and ( n17414 , n14013 , n7356 );
not ( n17415 , n17414 );
xnor ( n17416 , n17415 , n7352 );
xor ( n17417 , n17413 , n17416 );
and ( n17418 , n13647 , n7349 );
not ( n17419 , n17418 );
xor ( n17420 , n17417 , n17419 );
and ( n17421 , n17292 , n17293 );
and ( n17422 , n17293 , n17302 );
and ( n17423 , n17292 , n17302 );
or ( n17424 , n17421 , n17422 , n17423 );
xor ( n17425 , n17420 , n17424 );
and ( n17426 , n17303 , n17307 );
and ( n17427 , n17307 , n17312 );
and ( n17428 , n17303 , n17312 );
or ( n17429 , n17426 , n17427 , n17428 );
xor ( n17430 , n17425 , n17429 );
and ( n17431 , n17313 , n17314 );
xor ( n17432 , n17430 , n17431 );
buf ( n17433 , n17432 );
not ( n17434 , n454 );
and ( n17435 , n17434 , n17433 );
and ( n17436 , C0 , n454 );
or ( n17437 , n17435 , n17436 );
buf ( n17438 , n17437 );
buf ( n17439 , n17438 );
and ( n17440 , n17439 , n4505 );
xor ( n17441 , n17409 , n17440 );
xor ( n17442 , n17406 , n17441 );
xor ( n17443 , n17399 , n17442 );
and ( n17444 , n17324 , n17330 );
and ( n17445 , n17330 , n17335 );
and ( n17446 , n17324 , n17335 );
or ( n17447 , n17444 , n17445 , n17446 );
xor ( n17448 , n17443 , n17447 );
and ( n17449 , n17336 , n17340 );
and ( n17450 , n17340 , n17342 );
and ( n17451 , n17336 , n17342 );
or ( n17452 , n17449 , n17450 , n17451 );
xor ( n17453 , n17448 , n17452 );
and ( n17454 , n17344 , n17345 );
or ( n17455 , n17343 , n17454 );
xor ( n17456 , n17453 , n17455 );
buf ( n17457 , n17456 );
not ( n17458 , n4509 );
and ( n17459 , n17458 , n17398 );
and ( n17460 , n17457 , n4509 );
or ( n17461 , n17459 , n17460 );
and ( n17462 , n17355 , n17369 );
and ( n17463 , n17369 , n17384 );
and ( n17464 , n17355 , n17384 );
or ( n17465 , n17462 , n17463 , n17464 );
and ( n17466 , n17374 , n17378 );
and ( n17467 , n17378 , n17383 );
and ( n17468 , n17374 , n17383 );
or ( n17469 , n17466 , n17467 , n17468 );
not ( n17470 , n7626 );
and ( n17471 , n14865 , n8502 );
and ( n17472 , n15161 , n7970 );
nor ( n17473 , n17471 , n17472 );
xnor ( n17474 , n17473 , n8498 );
xor ( n17475 , n17470 , n17474 );
and ( n17476 , n13506 , n10329 );
and ( n17477 , n13865 , n9791 );
nor ( n17478 , n17476 , n17477 );
not ( n17479 , n17478 );
xor ( n17480 , n17475 , n17479 );
xor ( n17481 , n17469 , n17480 );
and ( n17482 , n17359 , n17363 );
and ( n17483 , n17363 , n17368 );
and ( n17484 , n17359 , n17368 );
or ( n17485 , n17482 , n17483 , n17484 );
buf ( n17486 , n17382 );
xor ( n17487 , n17485 , n17486 );
and ( n17488 , n14212 , n9407 );
and ( n17489 , n14558 , n8872 );
nor ( n17490 , n17488 , n17489 );
xnor ( n17491 , n17490 , n9403 );
xor ( n17492 , n17487 , n17491 );
xor ( n17493 , n17481 , n17492 );
xor ( n17494 , n17465 , n17493 );
and ( n17495 , n17385 , n17389 );
and ( n17496 , n17389 , n17394 );
and ( n17497 , n17385 , n17394 );
or ( n17498 , n17495 , n17496 , n17497 );
xor ( n17499 , n17494 , n17498 );
and ( n17500 , n17395 , n17396 );
xor ( n17501 , n17499 , n17500 );
buf ( n17502 , n17501 );
and ( n17503 , n17401 , n17405 );
and ( n17504 , n17405 , n17441 );
and ( n17505 , n17401 , n17441 );
or ( n17506 , n17503 , n17504 , n17505 );
buf ( n17507 , n17400 );
and ( n17508 , n17407 , n17408 );
and ( n17509 , n17408 , n17440 );
and ( n17510 , n17407 , n17440 );
or ( n17511 , n17508 , n17509 , n17510 );
xor ( n17512 , n17507 , n17511 );
and ( n17513 , n17211 , n5089 );
and ( n17514 , n17322 , n4866 );
and ( n17515 , n17439 , n4557 );
xor ( n17516 , n17514 , n17515 );
and ( n17517 , n17413 , n17416 );
and ( n17518 , n17416 , n17419 );
and ( n17519 , n17413 , n17419 );
or ( n17520 , n17517 , n17518 , n17519 );
buf ( n17521 , n17418 );
not ( n17522 , n7352 );
xor ( n17523 , n17521 , n17522 );
and ( n17524 , n14013 , n7349 );
xor ( n17525 , n17523 , n17524 );
xor ( n17526 , n17520 , n17525 );
and ( n17527 , n17420 , n17424 );
and ( n17528 , n17424 , n17429 );
and ( n17529 , n17420 , n17429 );
or ( n17530 , n17527 , n17528 , n17529 );
xor ( n17531 , n17526 , n17530 );
and ( n17532 , n17430 , n17431 );
xor ( n17533 , n17531 , n17532 );
buf ( n17534 , n17533 );
not ( n17535 , n454 );
and ( n17536 , n17535 , n17534 );
and ( n17537 , C0 , n454 );
or ( n17538 , n17536 , n17537 );
buf ( n17539 , n17538 );
buf ( n17540 , n17539 );
and ( n17541 , n17540 , n4505 );
xor ( n17542 , n17516 , n17541 );
xor ( n17543 , n17513 , n17542 );
xor ( n17544 , n17512 , n17543 );
xor ( n17545 , n17506 , n17544 );
and ( n17546 , n17399 , n17442 );
and ( n17547 , n17442 , n17447 );
and ( n17548 , n17399 , n17447 );
or ( n17549 , n17546 , n17547 , n17548 );
xor ( n17550 , n17545 , n17549 );
not ( n17551 , n17550 );
and ( n17552 , n17448 , n17452 );
and ( n17553 , n17453 , n17455 );
or ( n17554 , n17552 , n17553 );
xor ( n17555 , n17551 , n17554 );
buf ( n17556 , n17555 );
not ( n17557 , n4509 );
and ( n17558 , n17557 , n17502 );
and ( n17559 , n17556 , n4509 );
or ( n17560 , n17558 , n17559 );
and ( n17561 , n17470 , n17474 );
and ( n17562 , n17474 , n17479 );
and ( n17563 , n17470 , n17479 );
or ( n17564 , n17561 , n17562 , n17563 );
and ( n17565 , n17485 , n17486 );
and ( n17566 , n17486 , n17491 );
and ( n17567 , n17485 , n17491 );
or ( n17568 , n17565 , n17566 , n17567 );
xor ( n17569 , n17564 , n17568 );
and ( n17570 , n15161 , n8502 );
not ( n17571 , n17570 );
xnor ( n17572 , n17571 , n8498 );
not ( n17573 , n17572 );
and ( n17574 , n14558 , n9407 );
and ( n17575 , n14865 , n8872 );
nor ( n17576 , n17574 , n17575 );
xnor ( n17577 , n17576 , n9403 );
xor ( n17578 , n17573 , n17577 );
and ( n17579 , n13865 , n10329 );
and ( n17580 , n14212 , n9791 );
nor ( n17581 , n17579 , n17580 );
not ( n17582 , n17581 );
xor ( n17583 , n17578 , n17582 );
xor ( n17584 , n17569 , n17583 );
and ( n17585 , n17469 , n17480 );
and ( n17586 , n17480 , n17492 );
and ( n17587 , n17469 , n17492 );
or ( n17588 , n17585 , n17586 , n17587 );
xor ( n17589 , n17584 , n17588 );
and ( n17590 , n17465 , n17493 );
and ( n17591 , n17493 , n17498 );
and ( n17592 , n17465 , n17498 );
or ( n17593 , n17590 , n17591 , n17592 );
xor ( n17594 , n17589 , n17593 );
and ( n17595 , n17499 , n17500 );
xor ( n17596 , n17594 , n17595 );
buf ( n17597 , n17596 );
and ( n17598 , n17322 , n5089 );
and ( n17599 , n17540 , n4557 );
xor ( n17600 , n17598 , n17599 );
and ( n17601 , n17514 , n17515 );
and ( n17602 , n17515 , n17541 );
and ( n17603 , n17514 , n17541 );
or ( n17604 , n17601 , n17602 , n17603 );
xor ( n17605 , n17600 , n17604 );
and ( n17606 , n17439 , n4866 );
xor ( n17607 , n17605 , n17606 );
and ( n17608 , n17513 , n17542 );
xor ( n17609 , n17607 , n17608 );
and ( n17610 , n17507 , n17511 );
and ( n17611 , n17511 , n17543 );
and ( n17612 , n17507 , n17543 );
or ( n17613 , n17610 , n17611 , n17612 );
xor ( n17614 , n17609 , n17613 );
and ( n17615 , n17506 , n17544 );
and ( n17616 , n17544 , n17549 );
and ( n17617 , n17506 , n17549 );
or ( n17618 , n17615 , n17616 , n17617 );
xnor ( n17619 , n17614 , n17618 );
and ( n17620 , n17551 , n17554 );
or ( n17621 , n17550 , n17620 );
xor ( n17622 , n17619 , n17621 );
buf ( n17623 , n17622 );
not ( n17624 , n4509 );
and ( n17625 , n17624 , n17597 );
and ( n17626 , n17623 , n4509 );
or ( n17627 , n17625 , n17626 );
and ( n17628 , n17573 , n17577 );
and ( n17629 , n17577 , n17582 );
and ( n17630 , n17573 , n17582 );
or ( n17631 , n17628 , n17629 , n17630 );
buf ( n17632 , n17572 );
xor ( n17633 , n17631 , n17632 );
not ( n17634 , n8498 );
and ( n17635 , n14865 , n9407 );
and ( n17636 , n15161 , n8872 );
nor ( n17637 , n17635 , n17636 );
xnor ( n17638 , n17637 , n9403 );
xor ( n17639 , n17634 , n17638 );
and ( n17640 , n14212 , n10329 );
and ( n17641 , n14558 , n9791 );
nor ( n17642 , n17640 , n17641 );
not ( n17643 , n17642 );
xor ( n17644 , n17639 , n17643 );
xor ( n17645 , n17633 , n17644 );
and ( n17646 , n17564 , n17568 );
and ( n17647 , n17568 , n17583 );
and ( n17648 , n17564 , n17583 );
or ( n17649 , n17646 , n17647 , n17648 );
xor ( n17650 , n17645 , n17649 );
and ( n17651 , n17584 , n17588 );
and ( n17652 , n17588 , n17593 );
and ( n17653 , n17584 , n17593 );
or ( n17654 , n17651 , n17652 , n17653 );
xor ( n17655 , n17650 , n17654 );
and ( n17656 , n17594 , n17595 );
xor ( n17657 , n17655 , n17656 );
buf ( n17658 , n17657 );
and ( n17659 , n17598 , n17599 );
and ( n17660 , n17439 , n5089 );
xor ( n17661 , n17659 , n17660 );
and ( n17662 , n17540 , n4866 );
xor ( n17663 , n17661 , n17662 );
and ( n17664 , n17600 , n17604 );
and ( n17665 , n17604 , n17606 );
and ( n17666 , n17600 , n17606 );
or ( n17667 , n17664 , n17665 , n17666 );
xor ( n17668 , n17663 , n17667 );
and ( n17669 , n17607 , n17608 );
and ( n17670 , n17608 , n17613 );
and ( n17671 , n17607 , n17613 );
or ( n17672 , n17669 , n17670 , n17671 );
xor ( n17673 , n17668 , n17672 );
or ( n17674 , n17614 , n17618 );
xnor ( n17675 , n17673 , n17674 );
and ( n17676 , n17619 , n17621 );
xor ( n17677 , n17675 , n17676 );
buf ( n17678 , n17677 );
not ( n17679 , n4509 );
and ( n17680 , n17679 , n17658 );
and ( n17681 , n17678 , n4509 );
or ( n17682 , n17680 , n17681 );
and ( n17683 , n17634 , n17638 );
and ( n17684 , n17638 , n17643 );
and ( n17685 , n17634 , n17643 );
or ( n17686 , n17683 , n17684 , n17685 );
and ( n17687 , n15161 , n9407 );
not ( n17688 , n17687 );
xnor ( n17689 , n17688 , n9403 );
xor ( n17690 , n17686 , n17689 );
and ( n17691 , n14558 , n10329 );
and ( n17692 , n14865 , n9791 );
nor ( n17693 , n17691 , n17692 );
xor ( n17694 , n17690 , n17693 );
and ( n17695 , n17631 , n17632 );
and ( n17696 , n17632 , n17644 );
and ( n17697 , n17631 , n17644 );
or ( n17698 , n17695 , n17696 , n17697 );
xor ( n17699 , n17694 , n17698 );
and ( n17700 , n17645 , n17649 );
and ( n17701 , n17649 , n17654 );
and ( n17702 , n17645 , n17654 );
or ( n17703 , n17700 , n17701 , n17702 );
xor ( n17704 , n17699 , n17703 );
and ( n17705 , n17655 , n17656 );
xor ( n17706 , n17704 , n17705 );
buf ( n17707 , n17706 );
and ( n17708 , n17540 , n5089 );
and ( n17709 , n17659 , n17660 );
and ( n17710 , n17660 , n17662 );
and ( n17711 , n17659 , n17662 );
or ( n17712 , n17709 , n17710 , n17711 );
xor ( n17713 , n17708 , n17712 );
and ( n17714 , n17663 , n17667 );
and ( n17715 , n17667 , n17672 );
and ( n17716 , n17663 , n17672 );
or ( n17717 , n17714 , n17715 , n17716 );
xor ( n17718 , n17713 , n17717 );
or ( n17719 , n17673 , n17674 );
xnor ( n17720 , n17718 , n17719 );
and ( n17721 , n17675 , n17676 );
xor ( n17722 , n17720 , n17721 );
buf ( n17723 , n17722 );
not ( n17724 , n4509 );
and ( n17725 , n17724 , n17707 );
and ( n17726 , n17723 , n4509 );
or ( n17727 , n17725 , n17726 );
and ( n17728 , n17686 , n17689 );
and ( n17729 , n17689 , n17693 );
and ( n17730 , n17686 , n17693 );
or ( n17731 , n17728 , n17729 , n17730 );
not ( n17732 , n17693 );
buf ( n17733 , n17732 );
not ( n17734 , n9403 );
xor ( n17735 , n17733 , n17734 );
and ( n17736 , n14865 , n10329 );
and ( n17737 , n15161 , n9791 );
nor ( n17738 , n17736 , n17737 );
not ( n17739 , n17738 );
xor ( n17740 , n17735 , n17739 );
xor ( n17741 , n17731 , n17740 );
and ( n17742 , n17694 , n17698 );
and ( n17743 , n17698 , n17703 );
and ( n17744 , n17694 , n17703 );
or ( n17745 , n17742 , n17743 , n17744 );
xor ( n17746 , n17741 , n17745 );
and ( n17747 , n17704 , n17705 );
xor ( n17748 , n17746 , n17747 );
buf ( n17749 , n17748 );
and ( n17750 , n17708 , n17712 );
and ( n17751 , n17712 , n17717 );
and ( n17752 , n17708 , n17717 );
or ( n17753 , n17750 , n17751 , n17752 );
or ( n17754 , n17718 , n17719 );
xnor ( n17755 , n17753 , n17754 );
and ( n17756 , n17720 , n17721 );
xor ( n17757 , n17755 , n17756 );
buf ( n17758 , n17757 );
not ( n17759 , n4509 );
and ( n17760 , n17759 , n17749 );
and ( n17761 , n17758 , n4509 );
or ( n17762 , n17760 , n17761 );
and ( n17763 , n15161 , n10329 );
and ( n17764 , n17733 , n17734 );
and ( n17765 , n17734 , n17739 );
and ( n17766 , n17733 , n17739 );
or ( n17767 , n17764 , n17765 , n17766 );
xor ( n17768 , n17763 , n17767 );
and ( n17769 , n17731 , n17740 );
and ( n17770 , n17740 , n17745 );
and ( n17771 , n17731 , n17745 );
or ( n17772 , n17769 , n17770 , n17771 );
xor ( n17773 , n17768 , n17772 );
not ( n17774 , n17773 );
and ( n17775 , n17746 , n17747 );
xor ( n17776 , n17774 , n17775 );
buf ( n17777 , n17776 );
not ( n17778 , n4509 );
and ( n17779 , n17778 , n17777 );
and ( n17780 , C0 , n4509 );
or ( n17781 , n17779 , n17780 );
buf ( n17782 , n4373 );
buf ( n17783 , n17782 );
buf ( n17784 , n4486 );
buf ( n17785 , n17784 );
not ( n17786 , n454 );
and ( n17787 , n17786 , n17783 );
and ( n17788 , n17785 , n454 );
or ( n17789 , n17787 , n17788 );
xor ( n17790 , n4372 , n4375 );
buf ( n17791 , n17790 );
xor ( n17792 , n4485 , n4488 );
buf ( n17793 , n17792 );
not ( n17794 , n454 );
and ( n17795 , n17794 , n17791 );
and ( n17796 , n17793 , n454 );
or ( n17797 , n17795 , n17796 );
xor ( n17798 , n4368 , n4376 );
buf ( n17799 , n17798 );
xor ( n17800 , n4481 , n4489 );
buf ( n17801 , n17800 );
not ( n17802 , n454 );
and ( n17803 , n17802 , n17799 );
and ( n17804 , n17801 , n454 );
or ( n17805 , n17803 , n17804 );
xor ( n17806 , n4362 , n4378 );
buf ( n17807 , n17806 );
xor ( n17808 , n4475 , n4491 );
buf ( n17809 , n17808 );
not ( n17810 , n454 );
and ( n17811 , n17810 , n17807 );
and ( n17812 , n17809 , n454 );
or ( n17813 , n17811 , n17812 );
xor ( n17814 , n4355 , n4380 );
buf ( n17815 , n17814 );
xor ( n17816 , n4468 , n4493 );
buf ( n17817 , n17816 );
not ( n17818 , n454 );
and ( n17819 , n17818 , n17815 );
and ( n17820 , n17817 , n454 );
or ( n17821 , n17819 , n17820 );
not ( C0n , n4509 );
and ( C0 , C0n , n4509 );
endmodule
