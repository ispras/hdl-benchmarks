//NOTE: no-implementation module stub

module lx1 (
    input wire SYSCLK,
    input wire SYSCLKF,
    input wire SL_SLEEPSYS_C2_R,
    input wire SL_SLEEPSYS_C3_R,
    input wire BUSCLK,
    input wire BUSCLKF,
    input wire SL_SLEEPBUS_C2_BR,
    input wire SL_SLEEPBUS_C3_BR,
    input wire ResetN,
    input wire RESET_PWRON_N,
    input wire RESET_D1_R_N,
    input wire CFG_MEMSEQUENTIAL,
    input wire CFG_MEMZEROFIRST,
    input wire CFG_MEMFULLWORD,
    input wire CFG_LBCSYNCMODE,
    input wire CFG_LBCWBDISABLE,
    input wire CFG_EJTNMINUS1,
    input wire CFG_EJTMLOG2,
    input wire CFG_EJTBIT0M16,
    input wire JTAG_TDO_NR,
    input wire JTAG_TDI,
    input wire JTAG_TMS,
    input wire JTAG_CLOCK,
    input wire JTAG_TRST_N,
    input wire JTAG_RST_N,
    input wire JPT_PCST_DR,
    input wire JPT_TPC_DR,
    input wire EJT_DCLK,
    input wire CFG_EJDIS,
    input wire CFG_DWDISW,
    input wire Cond_in1,
    input wire [31:0] C1rd_data,
    input wire [31:0] C1rd_addr,
    input wire C1rhold,
    input wire C1rd_gen,
    input wire C1rd_con,
    input wire [31:0] C1wr_addr,
    input wire C1wr_gen,
    input wire C1wr_con,
    input wire [31:0] C1wr_data,
    input wire Cond_in2,
    input wire [31:0] C2rd_data,
    input wire [31:0] C2rd_addr,
    input wire C2rhold,
    input wire C2rd_gen,
    input wire C2rd_con,
    input wire [31:0] C2wr_addr,
    input wire C2wr_gen,
    input wire C2wr_con,
    input wire [31:0] C2wr_data,
    input wire Cond_in3,
    input wire [31:0] C3rd_data,
    input wire [31:0] C3rd_addr,
    input wire C3rhold,
    input wire C3rd_gen,
    input wire C3rd_con,
    input wire [31:0] C3wr_addr,
    input wire C3wr_gen,
    input wire C3wr_con,
    input wire [31:0] C3wr_data,
    input wire [31:0] C3cnt_inst,
    input wire [31:0] C3cnt_imiss,
    input wire [31:0] C3cnt_istall,
    input wire [31:0] C3cnt_dmiss,
    input wire [31:0] C3cnt_dstall,
    input wire [31:0] C3cnt_dload,
    input wire [31:0] C3cnt_dstore,
    input wire CEI_INSTM32_S_R_N,
    input wire CE1_RES_E,
    input wire CEI_CE1HOLD,
    input wire CEI_XCPN_M_C1,
    input wire CE1_SEL_E_R,
    input wire CE1_HALT_E_R,
    input wire CEI_CE1OP_S_R,
    input wire CEI_CE1AOP_E_R,
    input wire CEI_CE1BOP_E_R,
    input wire [31:0] LDataI,
    input wire LIrdyI,
    input wire LFrameI,
    input wire LSel,
    input wire LAbort,
    input wire LTrdy,
    input wire [31:0] LId,
    input wire [31:0] LUc,
    input wire LReq,
    input wire LGnt,
    input wire [31:0] LAddrO,
    input wire [31:0] LDataO,
    input wire LIrdy,
    input wire LFrame,
    input wire [31:0] LCmd,
    input wire [31:0] LCoe,
    input wire [31:0] LToe,
    input wire [31:0] LXoe,
    input wire [31:0] LDoe,
    input wire EXT_ICREQRAM_R,
    input wire IC_GNTRAM_R,
    input wire [31:0] IC_TAGINDEX,
    input wire [31:0] ICR_TAGRD0,
    input wire [31:0] IC_TAGWR0,
    input wire IC_TAG0WE,
    input wire IC_TAG0WEN,
    input wire IC_TAG0RE,
    input wire IC_TAG0REN,
    input wire IC_TAG0CS,
    input wire IC_TAG0CSN,
    input wire [31:0] IC_INSTINDEX,
    input wire IC_INSTWR,
    input wire IC_INST0WE,
    input wire IC_INST0WEN,
    input wire IC_INST0RE,
    input wire IC_INST0REN,
    input wire IC_INST0CS,
    input wire IC_INST0CSN,
    input wire CFG_ICOFF,
    input wire ICR_TAGMASK,
    input wire ICR_INST0RD,
    input wire IW_VALIDINDEX,
    input wire IWR_VALIDRD,
    input wire IW_VALIDWR,
    input wire IW_VALIDWE,
    input wire IW_VALIDWEN,
    input wire IW_VALIDRE,
    input wire IW_VALIDREN,
    input wire IW_VALIDCS,
    input wire IW_VALIDCSN,
    input wire IW_INSTINDEX,
    input wire IWR_INSTRD,
    input wire IW_INSTWR,
    input wire IW_INSTWE,
    input wire IW_INSTWEN,
    input wire IW_INSTRE,
    input wire IW_INSTREN,
    input wire IW_INSTCS,
    input wire IW_INSTCSN,
    input wire EXT_IWREQRAM_R,
    input wire IW_GNTRAM_R,
    input wire CFG_IWBASE,
    input wire CFG_IWTOP,
    input wire EXT_DCREQRAM_R,
    input wire DC_GNTRAM_R,
    input wire [31:0] DC_TAGINDEX,
    input wire [31:0] DC_TAGWR,
    input wire DC_TAGWE,
    input wire DC_TAGWEN,
    input wire DC_TAGRE,
    input wire DC_TAGREN,
    input wire DC_TAGCS,
    input wire DC_TAGCSN,
    input wire DCC_TAGMASK,
    input wire [31:0] DC_DATAINDEX,
    input wire [31:0] DC_DATAWR,
    input wire DC_DATAWE,
    input wire DC_DATAWEN,
    input wire DC_DATARE,
    input wire DC_DATAREN,
    input wire DC_DATACS,
    input wire DC_DATACSN,
    input wire CFG_DCOFF,
    input wire [31:0] DCR_TAGRD,
    input wire DCR_DATARD,
    input wire [31:0] DW_DATAINDEX,
    input wire DWR_DATARD,
    input wire DW_DATAWR,
    input wire DW_DATAWE,
    input wire DW_DATAWEN,
    input wire DW_DATARE,
    input wire DW_DATAREN,
    input wire DW_DATACS,
    input wire DW_DATACSN,
    input wire EXT_DWREQRAM_R,
    input wire DW_GNTRAM_R,
    input wire CFG_DWBASE,
    input wire CFG_DWTOP,
    input wire EXT_SLEEPREQ_R,
    input wire CFG_SLEEPENABLE,
    input wire IntreqN
);

endmodule
