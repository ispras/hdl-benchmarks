//NOTE: no-implementation module stub

module SW10201A (
    input  wire [4:0] A0,
    input  wire [4:0] A1,
    input  wire [4:0] A2,
    input  wire [4:0] A3,
    input  wire [4:0] A4,
    input  wire [4:0] B0,
    input  wire [4:0] B1,
    input  wire [4:0] B2,
    input  wire [4:0] B3,
    input  wire [4:0] B4,
    input  wire CKA,
    input  wire CKB,
    input  wire CSA,
    input  wire CSB,
    input  wire [11:0] DI0,
    input  wire [11:0] DI1,
    input  wire [11:0] DI2,
    input  wire [11:0] DI3,
    input  wire [11:0] DI4,
    input  wire [11:0] DI5,
    input  wire [11:0] DI6,
    input  wire [11:0] DI7,
    input  wire [11:0] DI8,
    input  wire [11:0] DI9,
    input  wire [11:0] DI10,
    input  wire [11:0] DI11,
    input  wire [11:0] DI12,
    input  wire [11:0] DI13,
    input  wire [11:0] DI14,
    input  wire [11:0] DI15,
    input  wire [11:0] DI16,
    input  wire [11:0] DI17,
    input  wire [11:0] DI18,
    input  wire [11:0] DI19,
    input  wire [11:0] DI20,
    input  wire [11:0] DI21,
    input  wire [11:0] DI22,
    input  wire [11:0] DI23,
    input  wire [11:0] DI24,
    input  wire [11:0] DI25,
    output reg [11:0] DO0,
    output reg [11:0] DO1,
    output reg [11:0] DO2,
    output reg [11:0] DO3,
    output reg [11:0] DO4,
    output reg [11:0] DO5,
    output reg [11:0] DO6,
    output reg [11:0] DO7,
    output reg [11:0] DO8,
    output reg [11:0] DO9,
    output reg [11:0] DO10,
    output reg [11:0] DO11,
    output reg [11:0] DO12,
    output reg [11:0] DO13,
    output reg [11:0] DO14,
    output reg [11:0] DO15,
    output reg [11:0] DO16,
    output reg [11:0] DO17,
    output reg [11:0] DO18,
    output reg [11:0] DO19,
    output reg [11:0] DO20,
    output reg [11:0] DO21,
    output reg [11:0] DO22,
    output reg [11:0] DO23,
    output reg [11:0] DO24,
    output reg [11:0] DO25,
    input  wire WEB,
    input  wire OE
);

endmodule
