module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 ;
output n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , 
 n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , 
 n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , 
 n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , 
 n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , 
 n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , 
 n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , 
 n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , 
 n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , 
 n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , 
 n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , 
 n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , 
 n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , 
 n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , 
 n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , 
 n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , 
 n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , 
 n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , 
 n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , 
 n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , 
 n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , 
 n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , 
 n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , 
 n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , 
 n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , 
 n379 , n380 , n381 , n382 , n383 ;
wire n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , 
 n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , 
 n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , 
 n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , 
 n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , 
 n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
 n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , 
 n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , 
 n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , 
 n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , 
 n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , 
 n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , 
 n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , 
 n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , 
 n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , 
 n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , 
 n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , 
 n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , 
 n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , 
 n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , 
 n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , 
 n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
 n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
 n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
 n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
 n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , 
 n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , 
 n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , 
 n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , 
 n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , 
 n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , 
 n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , 
 n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , 
 n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , 
 n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , 
 n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
 n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , 
 n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , 
 n1149 , n1150 , n1151 , n291647 , n291648 , n1221 , n291650 , n291651 , n291652 , n291653 , 
 n291654 , n291655 , n291656 , n291657 , n291658 , n291659 , n291660 , n291661 , n291662 , n291663 , 
 n291664 , n291665 , n1238 , n291667 , n291668 , n1241 , n291670 , n1243 , n291672 , n291673 , 
 n291674 , n291675 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , 
 n291684 , n291685 , n291686 , n291687 , n291688 , n291689 , n291690 , n1263 , n1264 , n1265 , 
 n1266 , n1267 , n1268 , n291697 , n1270 , n1271 , n291700 , n291701 , n1274 , n291703 , 
 n291704 , n291705 , n291706 , n291707 , n291708 , n291709 , n291710 , n291711 , n291712 , n291713 , 
 n291714 , n291715 , n291716 , n1289 , n291718 , n291719 , n1292 , n291721 , n291722 , n291723 , 
 n291724 , n1297 , n291726 , n1299 , n291728 , n1301 , n291730 , n291731 , n291732 , n291733 , 
 n291734 , n291735 , n291736 , n291737 , n291738 , n291739 , n1312 , n1313 , n1314 , n291743 , 
 n1316 , n1317 , n291746 , n1319 , n291748 , n291749 , n1322 , n1323 , n1324 , n1325 , 
 n1326 , n291755 , n1328 , n291757 , n1330 , n291759 , n1332 , n291761 , n291762 , n291763 , 
 n1336 , n291765 , n1338 , n1339 , n291768 , n291769 , n1342 , n1343 , n1344 , n291773 , 
 n1346 , n291775 , n291776 , n1349 , n1350 , n1351 , n291780 , n291781 , n1354 , n1355 , 
 n1356 , n1357 , n291786 , n291787 , n291788 , n291789 , n291790 , n291791 , n291792 , n291793 , 
 n291794 , n291795 , n291796 , n291797 , n291798 , n291799 , n291800 , n1373 , n291802 , n1375 , 
 n1376 , n291805 , n291806 , n291807 , n291808 , n291809 , n291810 , n1383 , n291812 , n291813 , 
 n1386 , n1387 , n1388 , n1389 , n291818 , n1391 , n291820 , n291821 , n291822 , n291823 , 
 n291824 , n1397 , n291826 , n291827 , n291828 , n291829 , n1402 , n291831 , n291832 , n1405 , 
 n1406 , n291835 , n291836 , n291837 , n291838 , n291839 , n291840 , n1413 , n291842 , n291843 , 
 n291844 , n291845 , n291846 , n1419 , n1420 , n291849 , n1422 , n291851 , n291852 , n1425 , 
 n291854 , n291855 , n291856 , n291857 , n291858 , n291859 , n291860 , n291861 , n1434 , n291863 , 
 n291864 , n291865 , n291866 , n291867 , n291868 , n291869 , n1442 , n291871 , n291872 , n1445 , 
 n291874 , n291875 , n1448 , n291877 , n291878 , n291879 , n291880 , n1453 , n291882 , n291883 , 
 n1456 , n291885 , n291886 , n291887 , n291888 , n291889 , n1462 , n291891 , n291892 , n1465 , 
 n291894 , n291895 , n1468 , n1469 , n291898 , n291899 , n1472 , n291901 , n1474 , n291903 , 
 n291904 , n1477 , n291906 , n291907 , n291908 , n291909 , n291910 , n291911 , n291912 , n291913 , 
 n291914 , n291915 , n291916 , n1489 , n291918 , n291919 , n291920 , n291921 , n291922 , n291923 , 
 n291924 , n291925 , n1498 , n291927 , n291928 , n291929 , n291930 , n291931 , n291932 , n291933 , 
 n1506 , n1507 , n1508 , n291937 , n291938 , n291939 , n291940 , n291941 , n291942 , n291943 , 
 n291944 , n291945 , n291946 , n291947 , n291948 , n1521 , n291950 , n291951 , n1524 , n1525 , 
 n291954 , n1527 , n291956 , n291957 , n291958 , n1531 , n291960 , n291961 , n291962 , n291963 , 
 n291964 , n291965 , n291966 , n1539 , n291968 , n291969 , n291970 , n1543 , n291972 , n291973 , 
 n291974 , n291975 , n1548 , n291977 , n1550 , n291979 , n291980 , n1553 , n291982 , n291983 , 
 n291984 , n291985 , n291986 , n1559 , n291988 , n291989 , n1562 , n291991 , n291992 , n291993 , 
 n291994 , n291995 , n291996 , n291997 , n1570 , n291999 , n1572 , n1573 , n292002 , n292003 , 
 n1576 , n292005 , n292006 , n1579 , n1580 , n292009 , n1582 , n292011 , n292012 , n292013 , 
 n292014 , n1587 , n292016 , n1589 , n292018 , n292019 , n292020 , n292021 , n292022 , n292023 , 
 n292024 , n1597 , n292026 , n1599 , n1600 , n1601 , n292030 , n1603 , n1604 , n1605 , 
 n292034 , n292035 , n292036 , n292037 , n292038 , n1611 , n292040 , n1613 , n292042 , n1615 , 
 n292044 , n1617 , n292046 , n1619 , n292048 , n292049 , n292050 , n292051 , n292052 , n292053 , 
 n292054 , n292055 , n292056 , n292057 , n1630 , n292059 , n292060 , n1633 , n292062 , n1635 , 
 n1636 , n1637 , n292066 , n1639 , n292068 , n292069 , n292070 , n292071 , n292072 , n292073 , 
 n1646 , n1647 , n292076 , n292077 , n292078 , n292079 , n292080 , n1653 , n1654 , n292083 , 
 n292084 , n292085 , n1658 , n1659 , n292088 , n292089 , n1662 , n292091 , n292092 , n292093 , 
 n1666 , n1667 , n292096 , n1669 , n292098 , n292099 , n1672 , n292101 , n292102 , n1675 , 
 n292104 , n292105 , n1678 , n292107 , n292108 , n292109 , n292110 , n1683 , n292112 , n292113 , 
 n1686 , n292115 , n292116 , n292117 , n292118 , n292119 , n1692 , n1693 , n1694 , n1695 , 
 n292124 , n292125 , n1698 , n292127 , n292128 , n292129 , n292130 , n292131 , n292132 , n1705 , 
 n1706 , n1707 , n292136 , n292137 , n1710 , n1711 , n1712 , n292141 , n292142 , n292143 , 
 n292144 , n292145 , n292146 , n1719 , n292148 , n1721 , n292150 , n292151 , n292152 , n292153 , 
 n292154 , n292155 , n292156 , n1729 , n292158 , n292159 , n1732 , n292161 , n292162 , n1735 , 
 n292164 , n1737 , n292166 , n1739 , n292168 , n292169 , n292170 , n1743 , n292172 , n292173 , 
 n292174 , n292175 , n292176 , n1749 , n1750 , n1751 , n292180 , n1753 , n292182 , n292183 , 
 n1756 , n292185 , n1758 , n292187 , n1760 , n292189 , n292190 , n292191 , n292192 , n292193 , 
 n292194 , n292195 , n292196 , n292197 , n1770 , n292199 , n1772 , n1773 , n292202 , n1775 , 
 n292204 , n292205 , n1778 , n1779 , n1780 , n292209 , n1782 , n292211 , n292212 , n292213 , 
 n292214 , n292215 , n1788 , n1789 , n1790 , n292219 , n292220 , n292221 , n1794 , n292223 , 
 n292224 , n1797 , n292226 , n1799 , n292228 , n1801 , n292230 , n292231 , n292232 , n292233 , 
 n292234 , n292235 , n292236 , n292237 , n292238 , n292239 , n292240 , n292241 , n292242 , n292243 , 
 n292244 , n1817 , n292246 , n1819 , n292248 , n292249 , n292250 , n292251 , n292252 , n292253 , 
 n1826 , n292255 , n292256 , n1829 , n292258 , n292259 , n1832 , n292261 , n292262 , n1835 , 
 n292264 , n292265 , n1838 , n292267 , n1840 , n292269 , n1842 , n292271 , n292272 , n292273 , 
 n292274 , n1847 , n292276 , n292277 , n1850 , n292279 , n1852 , n292281 , n292282 , n292283 , 
 n292284 , n292285 , n292286 , n292287 , n292288 , n1861 , n292290 , n292291 , n1864 , n292293 , 
 n1866 , n1867 , n1868 , n292297 , n292298 , n292299 , n292300 , n292301 , n292302 , n292303 , 
 n292304 , n1877 , n292306 , n292307 , n1880 , n292309 , n292310 , n292311 , n292312 , n292313 , 
 n292314 , n1887 , n292316 , n292317 , n292318 , n292319 , n292320 , n292321 , n292322 , n292323 , 
 n1896 , n292325 , n292326 , n292327 , n1900 , n1901 , n292330 , n1903 , n292332 , n292333 , 
 n292334 , n292335 , n292336 , n292337 , n1910 , n292339 , n1912 , n1913 , n1914 , n292343 , 
 n1916 , n292345 , n292346 , n292347 , n292348 , n292349 , n292350 , n292351 , n292352 , n1925 , 
 n292354 , n292355 , n292356 , n292357 , n292358 , n292359 , n292360 , n1933 , n1934 , n292363 , 
 n1936 , n292365 , n292366 , n292367 , n292368 , n292369 , n292370 , n292371 , n292372 , n292373 , 
 n292374 , n292375 , n292376 , n292377 , n1950 , n1951 , n292380 , n292381 , n292382 , n292383 , 
 n292384 , n292385 , n1958 , n1959 , n1960 , n1961 , n1962 , n292391 , n1964 , n292393 , 
 n1966 , n1967 , n1968 , n1969 , n292398 , n292399 , n292400 , n292401 , n292402 , n292403 , 
 n292404 , n292405 , n1978 , n292407 , n292408 , n292409 , n292410 , n292411 , n292412 , n292413 , 
 n292414 , n292415 , n292416 , n292417 , n292418 , n292419 , n1992 , n292421 , n292422 , n1995 , 
 n292424 , n1997 , n1998 , n1999 , n292428 , n292429 , n292430 , n292431 , n292432 , n292433 , 
 n292434 , n292435 , n292436 , n292437 , n292438 , n292439 , n292440 , n292441 , n2014 , n292443 , 
 n292444 , n2017 , n292446 , n292447 , n2020 , n292449 , n292450 , n2023 , n292452 , n292453 , 
 n2026 , n292455 , n292456 , n2029 , n292458 , n292459 , n2032 , n292461 , n2034 , n292463 , 
 n292464 , n2037 , n2038 , n292467 , n292468 , n2041 , n292470 , n292471 , n2044 , n292473 , 
 n2046 , n2047 , n2048 , n292477 , n292478 , n292479 , n292480 , n292481 , n292482 , n292483 , 
 n292484 , n292485 , n2058 , n292487 , n292488 , n2061 , n2062 , n2063 , n2064 , n2065 , 
 n2066 , n292495 , n2068 , n292497 , n292498 , n292499 , n292500 , n292501 , n292502 , n2075 , 
 n292504 , n292505 , n2078 , n2079 , n292508 , n292509 , n292510 , n292511 , n2084 , n2085 , 
 n2086 , n2087 , n2088 , n2089 , n292518 , n292519 , n292520 , n292521 , n292522 , n292523 , 
 n292524 , n2097 , n292526 , n292527 , n2100 , n292529 , n292530 , n2103 , n2104 , n292533 , 
 n2106 , n292535 , n292536 , n2109 , n292538 , n292539 , n2112 , n292541 , n292542 , n292543 , 
 n292544 , n2117 , n2118 , n292547 , n2120 , n292549 , n292550 , n292551 , n292552 , n292553 , 
 n292554 , n2127 , n292556 , n292557 , n292558 , n292559 , n292560 , n292561 , n2134 , n292563 , 
 n292564 , n292565 , n292566 , n292567 , n2140 , n2141 , n2142 , n2143 , n292572 , n2145 , 
 n2146 , n2147 , n292576 , n292577 , n2150 , n292579 , n2152 , n292581 , n2154 , n2155 , 
 n292584 , n2157 , n292586 , n2159 , n2160 , n292589 , n2162 , n292591 , n292592 , n292593 , 
 n292594 , n292595 , n292596 , n292597 , n2170 , n292599 , n292600 , n292601 , n292602 , n292603 , 
 n292604 , n2177 , n292606 , n292607 , n292608 , n292609 , n2182 , n292611 , n292612 , n2185 , 
 n292614 , n2187 , n292616 , n292617 , n2190 , n292619 , n292620 , n292621 , n292622 , n292623 , 
 n292624 , n2197 , n292626 , n292627 , n2200 , n292629 , n2202 , n292631 , n292632 , n292633 , 
 n2206 , n292635 , n292636 , n292637 , n292638 , n292639 , n292640 , n2213 , n292642 , n292643 , 
 n292644 , n292645 , n292646 , n2219 , n2220 , n292649 , n2222 , n292651 , n292652 , n292653 , 
 n292654 , n292655 , n292656 , n292657 , n292658 , n2231 , n292660 , n292661 , n2234 , n292663 , 
 n292664 , n2237 , n2238 , n292667 , n292668 , n292669 , n292670 , n292671 , n292672 , n292673 , 
 n292674 , n292675 , n2248 , n292677 , n2250 , n292679 , n292680 , n292681 , n292682 , n292683 , 
 n292684 , n292685 , n292686 , n292687 , n2260 , n2261 , n2262 , n2263 , n2264 , n292693 , 
 n2266 , n292695 , n292696 , n2269 , n292698 , n292699 , n292700 , n292701 , n2274 , n292703 , 
 n292704 , n2277 , n2278 , n292707 , n2280 , n292709 , n292710 , n2283 , n2284 , n292713 , 
 n292714 , n292715 , n292716 , n2289 , n292718 , n292719 , n292720 , n292721 , n292722 , n2295 , 
 n292724 , n292725 , n292726 , n292727 , n292728 , n292729 , n292730 , n292731 , n292732 , n292733 , 
 n292734 , n292735 , n292736 , n2309 , n292738 , n292739 , n2312 , n292741 , n292742 , n2315 , 
 n292744 , n292745 , n2318 , n292747 , n292748 , n292749 , n292750 , n292751 , n2324 , n292753 , 
 n292754 , n292755 , n2328 , n292757 , n2330 , n292759 , n2332 , n2333 , n2334 , n2335 , 
 n292764 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n292771 , n292772 , n2345 , 
 n292774 , n2347 , n292776 , n292777 , n292778 , n292779 , n2352 , n2353 , n292782 , n2355 , 
 n292784 , n292785 , n2358 , n292787 , n2360 , n2361 , n2362 , n292791 , n292792 , n292793 , 
 n2366 , n2367 , n2368 , n292797 , n2370 , n292799 , n2372 , n2373 , n292802 , n2375 , 
 n2376 , n292805 , n2378 , n292807 , n292808 , n2381 , n292810 , n2383 , n292812 , n292813 , 
 n292814 , n292815 , n2388 , n292817 , n292818 , n292819 , n292820 , n2393 , n292822 , n292823 , 
 n2396 , n292825 , n292826 , n292827 , n2400 , n2401 , n292830 , n292831 , n2404 , n2405 , 
 n292834 , n292835 , n292836 , n292837 , n2410 , n292839 , n2412 , n292841 , n2414 , n292843 , 
 n292844 , n292845 , n292846 , n292847 , n2420 , n292849 , n2422 , n292851 , n292852 , n292853 , 
 n292854 , n292855 , n292856 , n292857 , n292858 , n292859 , n292860 , n292861 , n292862 , n292863 , 
 n292864 , n292865 , n2438 , n292867 , n292868 , n2441 , n292870 , n292871 , n292872 , n292873 , 
 n2446 , n292875 , n292876 , n292877 , n292878 , n292879 , n292880 , n292881 , n292882 , n292883 , 
 n2456 , n292885 , n292886 , n2459 , n292888 , n292889 , n2462 , n292891 , n292892 , n292893 , 
 n292894 , n2467 , n292896 , n292897 , n292898 , n292899 , n292900 , n292901 , n2474 , n292903 , 
 n292904 , n292905 , n292906 , n292907 , n2480 , n292909 , n2482 , n292911 , n292912 , n292913 , 
 n292914 , n292915 , n292916 , n292917 , n292918 , n292919 , n292920 , n292921 , n292922 , n292923 , 
 n2496 , n292925 , n292926 , n2499 , n292928 , n292929 , n2502 , n292931 , n2504 , n292933 , 
 n2506 , n292935 , n292936 , n2509 , n292938 , n292939 , n2512 , n2513 , n292942 , n2515 , 
 n2516 , n292945 , n2518 , n292947 , n2520 , n292949 , n2522 , n292951 , n292952 , n292953 , 
 n292954 , n292955 , n292956 , n2529 , n292958 , n2531 , n2532 , n292961 , n2534 , n2535 , 
 n292964 , n292965 , n292966 , n2539 , n292968 , n292969 , n292970 , n292971 , n292972 , n292973 , 
 n292974 , n292975 , n292976 , n292977 , n292978 , n292979 , n292980 , n292981 , n292982 , n2555 , 
 n292984 , n292985 , n292986 , n292987 , n292988 , n292989 , n292990 , n292991 , n292992 , n292993 , 
 n292994 , n2567 , n292996 , n292997 , n292998 , n292999 , n293000 , n293001 , n293002 , n2575 , 
 n2576 , n293005 , n293006 , n2579 , n2580 , n293009 , n293010 , n2583 , n2584 , n293013 , 
 n293014 , n2587 , n293016 , n293017 , n293018 , n293019 , n293020 , n293021 , n2594 , n293023 , 
 n293024 , n2597 , n293026 , n293027 , n293028 , n2601 , n293030 , n293031 , n293032 , n293033 , 
 n293034 , n293035 , n293036 , n2609 , n293038 , n2611 , n293040 , n293041 , n293042 , n2615 , 
 n293044 , n293045 , n293046 , n293047 , n2620 , n293049 , n293050 , n293051 , n293052 , n293053 , 
 n293054 , n293055 , n293056 , n293057 , n293058 , n2631 , n293060 , n293061 , n2634 , n293063 , 
 n293064 , n293065 , n2638 , n293067 , n293068 , n293069 , n2642 , n2643 , n2644 , n2645 , 
 n2646 , n293075 , n293076 , n293077 , n293078 , n2651 , n2652 , n293081 , n293082 , n293083 , 
 n293084 , n293085 , n2658 , n293087 , n2660 , n2661 , n293090 , n293091 , n293092 , n293093 , 
 n293094 , n2667 , n2668 , n293097 , n2670 , n2671 , n293100 , n2673 , n293102 , n2675 , 
 n293104 , n293105 , n293106 , n293107 , n2680 , n2681 , n293110 , n2683 , n2684 , n293113 , 
 n2686 , n293115 , n2688 , n293117 , n293118 , n2691 , n293120 , n293121 , n293122 , n293123 , 
 n2696 , n293125 , n293126 , n2699 , n293128 , n293129 , n293130 , n293131 , n293132 , n293133 , 
 n2706 , n293135 , n293136 , n293137 , n293138 , n2711 , n293140 , n2713 , n293142 , n293143 , 
 n293144 , n293145 , n293146 , n293147 , n293148 , n293149 , n2722 , n293151 , n293152 , n2725 , 
 n2726 , n2727 , n2728 , n2729 , n293158 , n293159 , n293160 , n293161 , n293162 , n293163 , 
 n293164 , n293165 , n293166 , n293167 , n2740 , n293169 , n2742 , n2743 , n293172 , n293173 , 
 n293174 , n293175 , n293176 , n293177 , n2750 , n293179 , n293180 , n2753 , n293182 , n293183 , 
 n2756 , n293185 , n293186 , n2759 , n293188 , n293189 , n2762 , n293191 , n2764 , n293193 , 
 n293194 , n293195 , n293196 , n293197 , n293198 , n293199 , n2772 , n293201 , n293202 , n293203 , 
 n293204 , n2777 , n293206 , n293207 , n293208 , n293209 , n293210 , n293211 , n2784 , n293213 , 
 n293214 , n2787 , n293216 , n2789 , n293218 , n293219 , n2792 , n293221 , n293222 , n293223 , 
 n293224 , n2797 , n293226 , n293227 , n293228 , n293229 , n293230 , n293231 , n293232 , n293233 , 
 n2806 , n2807 , n293236 , n2809 , n293238 , n293239 , n293240 , n293241 , n2814 , n293243 , 
 n293244 , n293245 , n293246 , n2819 , n293248 , n293249 , n293250 , n2823 , n293252 , n293253 , 
 n2826 , n293255 , n293256 , n2829 , n293258 , n293259 , n2832 , n293261 , n293262 , n2835 , 
 n293264 , n293265 , n293266 , n293267 , n293268 , n293269 , n2842 , n293271 , n293272 , n2845 , 
 n293274 , n2847 , n2848 , n293277 , n293278 , n2851 , n293280 , n293281 , n293282 , n293283 , 
 n2856 , n293285 , n293286 , n293287 , n293288 , n293289 , n2862 , n293291 , n2864 , n2865 , 
 n293294 , n293295 , n2868 , n293297 , n293298 , n2871 , n293300 , n2873 , n2874 , n293303 , 
 n293304 , n2877 , n293306 , n293307 , n2880 , n293309 , n293310 , n293311 , n293312 , n293313 , 
 n293314 , n293315 , n293316 , n293317 , n293318 , n293319 , n2892 , n2893 , n293322 , n2895 , 
 n2896 , n293325 , n293326 , n293327 , n293328 , n293329 , n293330 , n293331 , n293332 , n293333 , 
 n293334 , n293335 , n2908 , n293337 , n293338 , n293339 , n293340 , n293341 , n293342 , n293343 , 
 n293344 , n293345 , n293346 , n293347 , n293348 , n293349 , n293350 , n293351 , n293352 , n293353 , 
 n293354 , n293355 , n2928 , n2929 , n2930 , n293359 , n293360 , n293361 , n293362 , n293363 , 
 n293364 , n293365 , n2938 , n293367 , n2940 , n2941 , n293370 , n293371 , n2944 , n293373 , 
 n293374 , n293375 , n293376 , n293377 , n2950 , n293379 , n293380 , n2953 , n293382 , n293383 , 
 n2956 , n293385 , n2958 , n293387 , n293388 , n293389 , n293390 , n293391 , n293392 , n2965 , 
 n293394 , n2967 , n2968 , n2969 , n293398 , n293399 , n2972 , n293401 , n293402 , n2975 , 
 n293404 , n293405 , n293406 , n293407 , n2980 , n293409 , n293410 , n293411 , n293412 , n293413 , 
 n293414 , n293415 , n2988 , n2989 , n293418 , n2991 , n293420 , n293421 , n2994 , n293423 , 
 n2996 , n2997 , n2998 , n2999 , n293428 , n3001 , n3002 , n293431 , n3004 , n293433 , 
 n293434 , n293435 , n3008 , n293437 , n3010 , n293439 , n293440 , n3013 , n293442 , n293443 , 
 n3016 , n3017 , n293446 , n3019 , n293448 , n293449 , n293450 , n3023 , n293452 , n3025 , 
 n293454 , n293455 , n3028 , n293457 , n3030 , n293459 , n293460 , n3033 , n293462 , n293463 , 
 n3036 , n293465 , n293466 , n293467 , n293468 , n3041 , n3042 , n293471 , n3044 , n3045 , 
 n293474 , n293475 , n3048 , n293477 , n293478 , n293479 , n3052 , n3053 , n293482 , n3055 , 
 n293484 , n293485 , n293486 , n293487 , n3060 , n293489 , n293490 , n3063 , n293492 , n293493 , 
 n3066 , n293495 , n3068 , n293497 , n3070 , n293499 , n3072 , n293501 , n3074 , n293503 , 
 n293504 , n293505 , n293506 , n3079 , n3080 , n293509 , n293510 , n293511 , n293512 , n293513 , 
 n293514 , n3087 , n293516 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n293523 , 
 n3096 , n293525 , n293526 , n293527 , n293528 , n293529 , n293530 , n293531 , n293532 , n293533 , 
 n293534 , n293535 , n3108 , n293537 , n293538 , n3111 , n3112 , n293541 , n3114 , n293543 , 
 n293544 , n293545 , n293546 , n3119 , n293548 , n293549 , n3122 , n3123 , n3124 , n3125 , 
 n3126 , n293555 , n293556 , n3129 , n293558 , n293559 , n3132 , n3133 , n3134 , n293563 , 
 n293564 , n3137 , n3138 , n3139 , n3140 , n293569 , n293570 , n293571 , n293572 , n293573 , 
 n293574 , n293575 , n293576 , n3149 , n3150 , n293579 , n293580 , n293581 , n3154 , n3155 , 
 n293584 , n293585 , n3158 , n293587 , n3160 , n293589 , n3162 , n293591 , n293592 , n293593 , 
 n293594 , n3167 , n293596 , n293597 , n293598 , n293599 , n3172 , n293601 , n293602 , n3175 , 
 n293604 , n3177 , n293606 , n293607 , n3180 , n3181 , n3182 , n293611 , n3184 , n293613 , 
 n293614 , n293615 , n293616 , n293617 , n293618 , n293619 , n3192 , n293621 , n293622 , n293623 , 
 n293624 , n3197 , n293626 , n293627 , n293628 , n293629 , n3202 , n293631 , n293632 , n293633 , 
 n293634 , n293635 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n293642 , n293643 , 
 n293644 , n293645 , n293646 , n293647 , n293648 , n293649 , n3222 , n3223 , n293652 , n3225 , 
 n293654 , n293655 , n3228 , n3229 , n3230 , n293659 , n293660 , n3233 , n3234 , n3235 , 
 n293664 , n293665 , n293666 , n293667 , n3240 , n293669 , n293670 , n3243 , n3244 , n3245 , 
 n3246 , n3247 , n3248 , n3249 , n293678 , n293679 , n293680 , n293681 , n293682 , n293683 , 
 n293684 , n293685 , n293686 , n293687 , n293688 , n293689 , n293690 , n293691 , n293692 , n293693 , 
 n293694 , n293695 , n3268 , n293697 , n293698 , n3271 , n293700 , n293701 , n293702 , n293703 , 
 n293704 , n293705 , n293706 , n293707 , n293708 , n3281 , n293710 , n293711 , n293712 , n293713 , 
 n293714 , n293715 , n293716 , n293717 , n293718 , n293719 , n3292 , n3293 , n3294 , n3295 , 
 n293724 , n293725 , n3298 , n3299 , n293728 , n293729 , n3302 , n293731 , n293732 , n3305 , 
 n293734 , n293735 , n3308 , n3309 , n3310 , n3311 , n3312 , n293741 , n3314 , n293743 , 
 n293744 , n3317 , n293746 , n293747 , n293748 , n293749 , n3322 , n293751 , n293752 , n293753 , 
 n293754 , n3327 , n293756 , n293757 , n3330 , n3331 , n293760 , n293761 , n3334 , n293763 , 
 n293764 , n3337 , n293766 , n293767 , n293768 , n3341 , n293770 , n293771 , n3344 , n293773 , 
 n293774 , n293775 , n293776 , n293777 , n293778 , n293779 , n293780 , n293781 , n3354 , n293783 , 
 n293784 , n293785 , n293786 , n293787 , n293788 , n293789 , n293790 , n293791 , n3364 , n293793 , 
 n3366 , n293795 , n293796 , n3369 , n293798 , n3371 , n293800 , n293801 , n293802 , n293803 , 
 n293804 , n293805 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , 
 n3386 , n3387 , n3388 , n3389 , n3390 , n293819 , n3392 , n293821 , n3394 , n3395 , 
 n293824 , n293825 , n293826 , n293827 , n293828 , n293829 , n293830 , n293831 , n293832 , n293833 , 
 n293834 , n293835 , n3408 , n293837 , n3410 , n293839 , n293840 , n293841 , n3414 , n293843 , 
 n3416 , n293845 , n293846 , n293847 , n293848 , n293849 , n293850 , n293851 , n293852 , n3425 , 
 n293854 , n3427 , n293856 , n293857 , n293858 , n293859 , n3432 , n293861 , n293862 , n293863 , 
 n293864 , n293865 , n293866 , n293867 , n293868 , n3441 , n3442 , n293871 , n293872 , n293873 , 
 n3446 , n3447 , n293876 , n293877 , n293878 , n293879 , n293880 , n293881 , n293882 , n293883 , 
 n293884 , n3457 , n3458 , n293887 , n293888 , n293889 , n293890 , n3463 , n293892 , n3465 , 
 n293894 , n3467 , n293896 , n3469 , n293898 , n3471 , n3472 , n293901 , n293902 , n293903 , 
 n293904 , n293905 , n293906 , n293907 , n293908 , n293909 , n3482 , n3483 , n293912 , n3485 , 
 n293914 , n293915 , n293916 , n293917 , n293918 , n293919 , n293920 , n3493 , n293922 , n3495 , 
 n293924 , n293925 , n293926 , n293927 , n3500 , n293929 , n3502 , n293931 , n293932 , n293933 , 
 n293934 , n293935 , n293936 , n293937 , n3510 , n293939 , n293940 , n3513 , n293942 , n293943 , 
 n3516 , n293945 , n293946 , n293947 , n3520 , n293949 , n3522 , n293951 , n293952 , n293953 , 
 n3526 , n293955 , n293956 , n293957 , n3530 , n293959 , n293960 , n3533 , n293962 , n293963 , 
 n293964 , n3537 , n3538 , n3539 , n293968 , n3541 , n3542 , n293971 , n293972 , n3545 , 
 n293974 , n293975 , n293976 , n3549 , n293978 , n293979 , n3552 , n293981 , n293982 , n3555 , 
 n293984 , n3557 , n293986 , n293987 , n3560 , n293989 , n293990 , n293991 , n3564 , n293993 , 
 n293994 , n3567 , n293996 , n293997 , n3570 , n293999 , n294000 , n3573 , n294002 , n294003 , 
 n3576 , n294005 , n3578 , n3579 , n294008 , n294009 , n294010 , n3583 , n294012 , n294013 , 
 n294014 , n294015 , n3588 , n294017 , n294018 , n3591 , n294020 , n294021 , n3594 , n294023 , 
 n294024 , n294025 , n294026 , n294027 , n3600 , n294029 , n3602 , n294031 , n294032 , n294033 , 
 n294034 , n294035 , n294036 , n294037 , n294038 , n294039 , n294040 , n294041 , n3614 , n294043 , 
 n294044 , n294045 , n294046 , n3619 , n294048 , n294049 , n294050 , n294051 , n294052 , n294053 , 
 n3626 , n3627 , n294056 , n294057 , n294058 , n294059 , n294060 , n294061 , n294062 , n294063 , 
 n3636 , n3637 , n3638 , n3639 , n294068 , n294069 , n3642 , n3643 , n294072 , n294073 , 
 n294074 , n3647 , n294076 , n294077 , n3650 , n294079 , n294080 , n3653 , n294082 , n3655 , 
 n3656 , n294085 , n3658 , n294087 , n294088 , n3661 , n294090 , n3663 , n294092 , n294093 , 
 n294094 , n294095 , n294096 , n3669 , n3670 , n294099 , n294100 , n294101 , n294102 , n294103 , 
 n294104 , n294105 , n3678 , n294107 , n294108 , n294109 , n3682 , n3683 , n294112 , n294113 , 
 n294114 , n3687 , n294116 , n294117 , n3690 , n294119 , n294120 , n3693 , n294122 , n294123 , 
 n294124 , n294125 , n294126 , n3699 , n3700 , n294129 , n3702 , n294131 , n3704 , n3705 , 
 n294134 , n294135 , n294136 , n294137 , n294138 , n294139 , n3712 , n294141 , n294142 , n294143 , 
 n294144 , n294145 , n3718 , n3719 , n294148 , n3721 , n294150 , n294151 , n294152 , n294153 , 
 n3726 , n294155 , n294156 , n294157 , n294158 , n294159 , n294160 , n294161 , n3734 , n294163 , 
 n3736 , n294165 , n294166 , n294167 , n294168 , n294169 , n294170 , n294171 , n3744 , n294173 , 
 n294174 , n294175 , n294176 , n294177 , n294178 , n294179 , n294180 , n294181 , n294182 , n294183 , 
 n294184 , n3757 , n294186 , n3759 , n294188 , n294189 , n3762 , n294191 , n3764 , n3765 , 
 n294194 , n3767 , n294196 , n3769 , n294198 , n294199 , n294200 , n294201 , n294202 , n294203 , 
 n294204 , n3777 , n294206 , n294207 , n294208 , n294209 , n294210 , n294211 , n294212 , n3785 , 
 n294214 , n294215 , n294216 , n294217 , n294218 , n294219 , n3792 , n294221 , n294222 , n294223 , 
 n294224 , n294225 , n3798 , n294227 , n294228 , n294229 , n294230 , n294231 , n3804 , n294233 , 
 n294234 , n294235 , n294236 , n3809 , n294238 , n294239 , n3812 , n294241 , n294242 , n294243 , 
 n294244 , n294245 , n294246 , n3819 , n294248 , n3821 , n294250 , n294251 , n294252 , n294253 , 
 n294254 , n294255 , n294256 , n294257 , n294258 , n3831 , n294260 , n294261 , n3834 , n294263 , 
 n294264 , n294265 , n294266 , n294267 , n3840 , n3841 , n294270 , n294271 , n3844 , n3845 , 
 n294274 , n294275 , n294276 , n294277 , n294278 , n294279 , n3852 , n294281 , n294282 , n294283 , 
 n294284 , n294285 , n3858 , n294287 , n294288 , n294289 , n3862 , n294291 , n3864 , n3865 , 
 n294294 , n294295 , n3868 , n294297 , n3870 , n294299 , n294300 , n294301 , n294302 , n294303 , 
 n3876 , n294305 , n294306 , n3879 , n3880 , n294309 , n294310 , n3883 , n294312 , n294313 , 
 n3886 , n294315 , n294316 , n3889 , n294318 , n294319 , n3892 , n294321 , n294322 , n294323 , 
 n3896 , n294325 , n294326 , n294327 , n3900 , n294329 , n294330 , n3903 , n294332 , n3905 , 
 n294334 , n294335 , n294336 , n294337 , n294338 , n294339 , n294340 , n294341 , n294342 , n294343 , 
 n294344 , n3917 , n3918 , n294347 , n294348 , n294349 , n3922 , n294351 , n294352 , n294353 , 
 n3926 , n294355 , n294356 , n294357 , n3930 , n294359 , n294360 , n294361 , n294362 , n294363 , 
 n3936 , n3937 , n294366 , n294367 , n294368 , n294369 , n294370 , n3943 , n294372 , n294373 , 
 n294374 , n294375 , n294376 , n294377 , n294378 , n294379 , n294380 , n3953 , n294382 , n3955 , 
 n294384 , n294385 , n294386 , n294387 , n294388 , n294389 , n294390 , n3963 , n294392 , n294393 , 
 n3966 , n3967 , n294396 , n3969 , n294398 , n294399 , n3972 , n3973 , n294402 , n3975 , 
 n3976 , n3977 , n294406 , n294407 , n3980 , n294409 , n3982 , n294411 , n294412 , n294413 , 
 n294414 , n294415 , n294416 , n294417 , n3990 , n294419 , n294420 , n294421 , n3994 , n294423 , 
 n294424 , n294425 , n294426 , n294427 , n4000 , n4001 , n4002 , n294431 , n4004 , n294433 , 
 n294434 , n4007 , n294436 , n294437 , n4010 , n294439 , n294440 , n294441 , n4014 , n294443 , 
 n294444 , n294445 , n294446 , n4019 , n4020 , n294449 , n294450 , n294451 , n294452 , n294453 , 
 n294454 , n294455 , n294456 , n294457 , n4030 , n4031 , n294460 , n4033 , n294462 , n4035 , 
 n294464 , n294465 , n294466 , n294467 , n4040 , n294469 , n4042 , n4043 , n294472 , n294473 , 
 n294474 , n4047 , n294476 , n4049 , n294478 , n294479 , n294480 , n294481 , n294482 , n294483 , 
 n294484 , n294485 , n294486 , n294487 , n4060 , n294489 , n294490 , n294491 , n4064 , n294493 , 
 n294494 , n4067 , n294496 , n294497 , n294498 , n294499 , n294500 , n4073 , n4074 , n4075 , 
 n294504 , n4077 , n4078 , n294507 , n4080 , n294509 , n4082 , n294511 , n4084 , n4085 , 
 n294514 , n294515 , n294516 , n294517 , n294518 , n294519 , n4092 , n294521 , n294522 , n294523 , 
 n294524 , n294525 , n294526 , n294527 , n294528 , n294529 , n294530 , n294531 , n294532 , n294533 , 
 n294534 , n4107 , n294536 , n294537 , n294538 , n294539 , n294540 , n294541 , n4114 , n294543 , 
 n294544 , n4117 , n294546 , n294547 , n294548 , n294549 , n294550 , n4123 , n294552 , n294553 , 
 n294554 , n294555 , n4128 , n294557 , n294558 , n294559 , n294560 , n294561 , n294562 , n294563 , 
 n4136 , n294565 , n294566 , n294567 , n294568 , n294569 , n4142 , n294571 , n294572 , n4145 , 
 n294574 , n4147 , n4148 , n294577 , n4150 , n4151 , n294580 , n294581 , n4154 , n294583 , 
 n4156 , n294585 , n4158 , n294587 , n4160 , n4161 , n4162 , n294591 , n294592 , n294593 , 
 n294594 , n294595 , n4168 , n294597 , n294598 , n294599 , n294600 , n4173 , n4174 , n294603 , 
 n294604 , n294605 , n294606 , n294607 , n294608 , n294609 , n4182 , n294611 , n4184 , n4185 , 
 n294614 , n294615 , n294616 , n4189 , n294618 , n294619 , n4192 , n294621 , n294622 , n4195 , 
 n4196 , n294625 , n4198 , n294627 , n294628 , n4201 , n294630 , n294631 , n294632 , n4205 , 
 n294634 , n294635 , n4208 , n294637 , n294638 , n4211 , n294640 , n294641 , n294642 , n4215 , 
 n294644 , n294645 , n294646 , n294647 , n4220 , n294649 , n294650 , n294651 , n294652 , n4225 , 
 n294654 , n4227 , n294656 , n4229 , n294658 , n294659 , n4232 , n294661 , n294662 , n294663 , 
 n4236 , n294665 , n294666 , n294667 , n4240 , n294669 , n4242 , n4243 , n4244 , n294673 , 
 n4246 , n294675 , n294676 , n294677 , n4250 , n294679 , n294680 , n4253 , n294682 , n294683 , 
 n294684 , n4257 , n294686 , n294687 , n4260 , n294689 , n294690 , n4263 , n294692 , n294693 , 
 n4266 , n294695 , n294696 , n294697 , n4270 , n294699 , n294700 , n294701 , n294702 , n294703 , 
 n294704 , n294705 , n294706 , n294707 , n294708 , n294709 , n294710 , n294711 , n4284 , n294713 , 
 n294714 , n294715 , n4288 , n294717 , n294718 , n294719 , n294720 , n4293 , n294722 , n294723 , 
 n4296 , n294725 , n294726 , n294727 , n4300 , n294729 , n294730 , n294731 , n294732 , n294733 , 
 n294734 , n294735 , n294736 , n4309 , n294738 , n4311 , n294740 , n4313 , n294742 , n4315 , 
 n294744 , n294745 , n294746 , n294747 , n294748 , n294749 , n294750 , n294751 , n294752 , n294753 , 
 n294754 , n294755 , n294756 , n294757 , n294758 , n4331 , n294760 , n294761 , n4334 , n294763 , 
 n294764 , n294765 , n294766 , n294767 , n294768 , n294769 , n294770 , n294771 , n294772 , n4345 , 
 n294774 , n294775 , n294776 , n294777 , n294778 , n294779 , n294780 , n294781 , n294782 , n294783 , 
 n294784 , n4357 , n294786 , n294787 , n294788 , n294789 , n294790 , n4363 , n294792 , n294793 , 
 n294794 , n294795 , n4368 , n294797 , n294798 , n4371 , n294800 , n4373 , n4374 , n294803 , 
 n4376 , n294805 , n4378 , n294807 , n294808 , n4381 , n294810 , n294811 , n294812 , n4385 , 
 n294814 , n294815 , n294816 , n4389 , n294818 , n294819 , n294820 , n294821 , n4394 , n294823 , 
 n294824 , n294825 , n4398 , n4399 , n294828 , n294829 , n4402 , n294831 , n294832 , n294833 , 
 n294834 , n294835 , n294836 , n294837 , n294838 , n294839 , n294840 , n294841 , n294842 , n4415 , 
 n294844 , n294845 , n294846 , n4419 , n294848 , n294849 , n294850 , n294851 , n294852 , n294853 , 
 n4426 , n294855 , n4428 , n4429 , n4430 , n4431 , n4432 , n294861 , n294862 , n294863 , 
 n4436 , n294865 , n4438 , n294867 , n4440 , n294869 , n294870 , n294871 , n294872 , n294873 , 
 n4446 , n4447 , n294876 , n4449 , n4450 , n294879 , n294880 , n294881 , n4454 , n294883 , 
 n294884 , n294885 , n294886 , n4459 , n294888 , n294889 , n294890 , n294891 , n4464 , n294893 , 
 n294894 , n294895 , n294896 , n4469 , n294898 , n294899 , n294900 , n294901 , n294902 , n4475 , 
 n294904 , n294905 , n4478 , n294907 , n4480 , n294909 , n294910 , n294911 , n294912 , n294913 , 
 n294914 , n4487 , n294916 , n294917 , n294918 , n294919 , n294920 , n294921 , n294922 , n294923 , 
 n4496 , n294925 , n294926 , n4499 , n4500 , n4501 , n4502 , n4503 , n294932 , n4505 , 
 n294934 , n294935 , n4508 , n4509 , n4510 , n4511 , n4512 , n294941 , n4514 , n294943 , 
 n294944 , n4517 , n294946 , n294947 , n294948 , n294949 , n294950 , n4523 , n294952 , n294953 , 
 n294954 , n4527 , n294956 , n294957 , n294958 , n4531 , n4532 , n294961 , n294962 , n294963 , 
 n294964 , n294965 , n4538 , n294967 , n294968 , n294969 , n4542 , n294971 , n4544 , n4545 , 
 n294974 , n294975 , n4548 , n294977 , n294978 , n4551 , n294980 , n294981 , n4554 , n294983 , 
 n294984 , n4557 , n294986 , n4559 , n294988 , n294989 , n294990 , n294991 , n294992 , n4565 , 
 n294994 , n294995 , n294996 , n294997 , n294998 , n294999 , n4572 , n4573 , n295002 , n295003 , 
 n4576 , n295005 , n295006 , n4579 , n295008 , n4581 , n4582 , n295011 , n295012 , n4585 , 
 n295014 , n4587 , n295016 , n295017 , n295018 , n295019 , n295020 , n295021 , n295022 , n295023 , 
 n295024 , n295025 , n295026 , n295027 , n295028 , n295029 , n295030 , n4603 , n295032 , n295033 , 
 n295034 , n295035 , n295036 , n295037 , n4610 , n295039 , n295040 , n295041 , n295042 , n295043 , 
 n295044 , n295045 , n295046 , n295047 , n295048 , n295049 , n4622 , n295051 , n295052 , n4625 , 
 n295054 , n295055 , n295056 , n295057 , n4630 , n295059 , n295060 , n295061 , n295062 , n295063 , 
 n295064 , n4637 , n295066 , n295067 , n4640 , n4641 , n295070 , n295071 , n295072 , n295073 , 
 n295074 , n4647 , n295076 , n295077 , n295078 , n295079 , n4652 , n295081 , n295082 , n295083 , 
 n295084 , n295085 , n295086 , n4659 , n295088 , n295089 , n295090 , n295091 , n295092 , n295093 , 
 n295094 , n295095 , n295096 , n295097 , n295098 , n295099 , n295100 , n295101 , n295102 , n295103 , 
 n4676 , n295105 , n295106 , n295107 , n295108 , n295109 , n295110 , n295111 , n295112 , n295113 , 
 n295114 , n4687 , n295116 , n295117 , n295118 , n295119 , n4692 , n4693 , n295122 , n295123 , 
 n4696 , n295125 , n295126 , n4699 , n295128 , n295129 , n4702 , n4703 , n295132 , n4705 , 
 n295134 , n295135 , n295136 , n295137 , n4710 , n295139 , n295140 , n4713 , n295142 , n4715 , 
 n295144 , n4717 , n295146 , n4719 , n295148 , n4721 , n295150 , n295151 , n295152 , n295153 , 
 n4726 , n295155 , n295156 , n4729 , n295158 , n295159 , n295160 , n4733 , n295162 , n295163 , 
 n295164 , n295165 , n295166 , n4739 , n4740 , n295169 , n4742 , n295171 , n4744 , n295173 , 
 n4746 , n295175 , n295176 , n295177 , n4750 , n4751 , n295180 , n295181 , n295182 , n4755 , 
 n295184 , n4757 , n295186 , n295187 , n4760 , n295189 , n4762 , n295191 , n4764 , n295193 , 
 n4766 , n4767 , n4768 , n295197 , n4770 , n4771 , n4772 , n4773 , n4774 , n295203 , 
 n4776 , n295205 , n295206 , n4779 , n295208 , n4781 , n295210 , n4783 , n295212 , n4785 , 
 n4786 , n4787 , n4788 , n4789 , n295218 , n295219 , n4792 , n295221 , n295222 , n4795 , 
 n295224 , n4797 , n4798 , n295227 , n295228 , n4801 , n295230 , n4803 , n295232 , n295233 , 
 n295234 , n295235 , n295236 , n295237 , n295238 , n295239 , n295240 , n295241 , n4814 , n295243 , 
 n4816 , n4817 , n295246 , n4819 , n295248 , n4821 , n295250 , n295251 , n295252 , n295253 , 
 n295254 , n295255 , n295256 , n295257 , n4830 , n295259 , n295260 , n295261 , n295262 , n4835 , 
 n295264 , n295265 , n4838 , n295267 , n295268 , n4841 , n4842 , n295271 , n295272 , n4845 , 
 n4846 , n295275 , n4848 , n4849 , n4850 , n4851 , n295280 , n4853 , n295282 , n4855 , 
 n295284 , n295285 , n295286 , n295287 , n4860 , n295289 , n295290 , n4863 , n295292 , n295293 , 
 n4866 , n295295 , n4868 , n295297 , n295298 , n295299 , n295300 , n295301 , n295302 , n295303 , 
 n4876 , n295305 , n295306 , n295307 , n295308 , n4881 , n295310 , n4883 , n295312 , n4885 , 
 n4886 , n295315 , n295316 , n4889 , n4890 , n295319 , n295320 , n4893 , n295322 , n4895 , 
 n295324 , n295325 , n4898 , n295327 , n4900 , n295329 , n295330 , n295331 , n295332 , n295333 , 
 n295334 , n295335 , n295336 , n4909 , n295338 , n4911 , n295340 , n295341 , n295342 , n4915 , 
 n295344 , n295345 , n4918 , n295347 , n4920 , n295349 , n295350 , n295351 , n295352 , n295353 , 
 n295354 , n4927 , n295356 , n295357 , n295358 , n295359 , n4932 , n295361 , n295362 , n295363 , 
 n295364 , n295365 , n295366 , n295367 , n295368 , n4941 , n295370 , n295371 , n295372 , n295373 , 
 n295374 , n295375 , n4948 , n295377 , n4950 , n295379 , n4952 , n295381 , n4954 , n295383 , 
 n295384 , n295385 , n295386 , n4959 , n4960 , n4961 , n295390 , n295391 , n295392 , n295393 , 
 n295394 , n295395 , n295396 , n4969 , n295398 , n4971 , n4972 , n295401 , n295402 , n4975 , 
 n295404 , n295405 , n4978 , n295407 , n295408 , n4981 , n295410 , n4983 , n295412 , n4985 , 
 n295414 , n4987 , n4988 , n4989 , n4990 , n295419 , n4992 , n4993 , n295422 , n295423 , 
 n295424 , n295425 , n4998 , n295427 , n295428 , n5001 , n295430 , n5003 , n5004 , n295433 , 
 n295434 , n5007 , n295436 , n295437 , n295438 , n295439 , n295440 , n5013 , n295442 , n295443 , 
 n295444 , n295445 , n5018 , n295447 , n5020 , n295449 , n295450 , n5023 , n295452 , n295453 , 
 n295454 , n295455 , n295456 , n295457 , n295458 , n295459 , n295460 , n5033 , n5034 , n295463 , 
 n5036 , n295465 , n5038 , n295467 , n295468 , n295469 , n295470 , n295471 , n295472 , n295473 , 
 n295474 , n295475 , n5048 , n5049 , n295478 , n5051 , n295480 , n5053 , n295482 , n295483 , 
 n295484 , n295485 , n295486 , n295487 , n295488 , n295489 , n295490 , n5063 , n5064 , n5065 , 
 n295494 , n295495 , n295496 , n295497 , n295498 , n295499 , n295500 , n295501 , n295502 , n295503 , 
 n295504 , n295505 , n295506 , n295507 , n295508 , n295509 , n5082 , n5083 , n295512 , n295513 , 
 n295514 , n5087 , n295516 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n295523 , 
 n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n295533 , 
 n5106 , n295535 , n5108 , n295537 , n295538 , n295539 , n295540 , n5113 , n295542 , n295543 , 
 n5116 , n295545 , n295546 , n295547 , n295548 , n5121 , n5122 , n5123 , n295552 , n295553 , 
 n5126 , n295555 , n5128 , n5129 , n295558 , n5131 , n5132 , n5133 , n295562 , n295563 , 
 n5136 , n5137 , n5138 , n295567 , n5140 , n5141 , n295570 , n5143 , n5144 , n295573 , 
 n5146 , n295575 , n295576 , n295577 , n295578 , n295579 , n295580 , n295581 , n295582 , n295583 , 
 n295584 , n5157 , n295586 , n295587 , n295588 , n295589 , n295590 , n295591 , n5164 , n295593 , 
 n295594 , n295595 , n295596 , n295597 , n295598 , n5171 , n295600 , n295601 , n295602 , n295603 , 
 n295604 , n5177 , n295606 , n5179 , n295608 , n295609 , n295610 , n295611 , n295612 , n295613 , 
 n295614 , n295615 , n295616 , n295617 , n295618 , n295619 , n295620 , n295621 , n295622 , n5195 , 
 n5196 , n295625 , n5198 , n295627 , n5200 , n295629 , n295630 , n295631 , n295632 , n295633 , 
 n295634 , n5207 , n295636 , n295637 , n295638 , n295639 , n295640 , n295641 , n5214 , n295643 , 
 n295644 , n295645 , n295646 , n295647 , n295648 , n295649 , n295650 , n5223 , n295652 , n295653 , 
 n5226 , n295655 , n5228 , n295657 , n295658 , n5231 , n295660 , n5233 , n5234 , n5235 , 
 n5236 , n5237 , n5238 , n295667 , n5240 , n295669 , n295670 , n295671 , n295672 , n295673 , 
 n295674 , n5247 , n295676 , n295677 , n295678 , n295679 , n5252 , n295681 , n5254 , n5255 , 
 n295684 , n295685 , n5258 , n5259 , n295688 , n5261 , n295690 , n295691 , n5264 , n295693 , 
 n5266 , n295695 , n5268 , n5269 , n295698 , n5271 , n295700 , n295701 , n295702 , n295703 , 
 n295704 , n295705 , n295706 , n295707 , n5280 , n5281 , n295710 , n295711 , n5284 , n295713 , 
 n295714 , n5287 , n295716 , n295717 , n5290 , n295719 , n295720 , n5293 , n295722 , n295723 , 
 n5296 , n5297 , n295726 , n295727 , n295728 , n5301 , n5302 , n5303 , n295732 , n295733 , 
 n295734 , n5307 , n295736 , n295737 , n5310 , n5311 , n295740 , n295741 , n295742 , n5315 , 
 n5316 , n295745 , n295746 , n5319 , n5320 , n295749 , n295750 , n295751 , n295752 , n5325 , 
 n295754 , n295755 , n295756 , n5329 , n5330 , n5331 , n295760 , n295761 , n5334 , n295763 , 
 n5336 , n295765 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n295772 , n5345 , 
 n295774 , n295775 , n5348 , n295777 , n295778 , n295779 , n295780 , n295781 , n295782 , n295783 , 
 n295784 , n295785 , n295786 , n5359 , n295788 , n295789 , n5362 , n295791 , n295792 , n5365 , 
 n295794 , n295795 , n5368 , n5369 , n295798 , n5371 , n295800 , n295801 , n5374 , n295803 , 
 n295804 , n295805 , n5378 , n295807 , n295808 , n5381 , n295810 , n5383 , n5384 , n295813 , 
 n295814 , n5387 , n295816 , n295817 , n5390 , n295819 , n295820 , n295821 , n295822 , n5395 , 
 n295824 , n5397 , n295826 , n295827 , n295828 , n5401 , n295830 , n295831 , n5404 , n295833 , 
 n295834 , n5407 , n295836 , n295837 , n5410 , n295839 , n295840 , n5413 , n295842 , n5415 , 
 n5416 , n5417 , n295846 , n295847 , n295848 , n295849 , n5422 , n295851 , n295852 , n5425 , 
 n295854 , n295855 , n295856 , n5429 , n295858 , n295859 , n295860 , n295861 , n5434 , n5435 , 
 n5436 , n5437 , n295866 , n5439 , n5440 , n5441 , n295870 , n5443 , n5444 , n295873 , 
 n295874 , n5447 , n5448 , n5449 , n295878 , n5451 , n295880 , n295881 , n5454 , n295883 , 
 n5456 , n5457 , n5458 , n5459 , n295888 , n295889 , n5462 , n295891 , n5464 , n295893 , 
 n5466 , n5467 , n5468 , n295897 , n295898 , n5471 , n5472 , n5473 , n5474 , n5475 , 
 n5476 , n5477 , n5478 , n5479 , n295908 , n5481 , n295910 , n295911 , n295912 , n5485 , 
 n5486 , n295915 , n5488 , n5489 , n295918 , n295919 , n295920 , n295921 , n295922 , n295923 , 
 n5496 , n295925 , n295926 , n5499 , n295928 , n295929 , n295930 , n295931 , n295932 , n5505 , 
 n295934 , n295935 , n5508 , n295937 , n295938 , n295939 , n5512 , n295941 , n295942 , n5515 , 
 n295944 , n295945 , n295946 , n295947 , n295948 , n295949 , n5522 , n295951 , n295952 , n295953 , 
 n295954 , n295955 , n295956 , n5529 , n295958 , n295959 , n295960 , n295961 , n5534 , n295963 , 
 n295964 , n5537 , n295966 , n5539 , n5540 , n295969 , n295970 , n5543 , n295972 , n295973 , 
 n295974 , n295975 , n295976 , n295977 , n295978 , n295979 , n295980 , n295981 , n5554 , n295983 , 
 n295984 , n5557 , n295986 , n295987 , n295988 , n295989 , n295990 , n295991 , n295992 , n295993 , 
 n295994 , n295995 , n295996 , n295997 , n295998 , n5571 , n296000 , n296001 , n296002 , n5575 , 
 n296004 , n5577 , n296006 , n296007 , n296008 , n296009 , n296010 , n296011 , n296012 , n296013 , 
 n296014 , n296015 , n296016 , n296017 , n5590 , n296019 , n5592 , n296021 , n296022 , n5595 , 
 n5596 , n5597 , n5598 , n296027 , n296028 , n296029 , n296030 , n5603 , n296032 , n296033 , 
 n5606 , n296035 , n296036 , n296037 , n296038 , n296039 , n296040 , n296041 , n5614 , n5615 , 
 n5616 , n5617 , n5618 , n5619 , n296048 , n5621 , n296050 , n296051 , n5624 , n296053 , 
 n5626 , n5627 , n5628 , n5629 , n296058 , n296059 , n296060 , n5633 , n296062 , n296063 , 
 n5636 , n296065 , n5638 , n5639 , n296068 , n296069 , n5642 , n296071 , n296072 , n5645 , 
 n296074 , n296075 , n5648 , n5649 , n296078 , n5651 , n296080 , n5653 , n5654 , n296083 , 
 n296084 , n5657 , n296086 , n296087 , n5660 , n296089 , n296090 , n5663 , n5664 , n5665 , 
 n296094 , n5667 , n5668 , n296097 , n296098 , n5671 , n296100 , n296101 , n5674 , n296103 , 
 n5676 , n296105 , n296106 , n296107 , n5680 , n296109 , n296110 , n296111 , n296112 , n296113 , 
 n296114 , n296115 , n296116 , n296117 , n5690 , n296119 , n5692 , n296121 , n296122 , n296123 , 
 n296124 , n5697 , n296126 , n296127 , n5700 , n296129 , n5702 , n5703 , n296132 , n296133 , 
 n296134 , n296135 , n296136 , n5709 , n296138 , n5711 , n296140 , n296141 , n296142 , n5715 , 
 n296144 , n296145 , n5718 , n296147 , n296148 , n5721 , n296150 , n296151 , n296152 , n296153 , 
 n5726 , n296155 , n296156 , n5729 , n296158 , n296159 , n5732 , n5733 , n5734 , n296163 , 
 n296164 , n5737 , n5738 , n5739 , n296168 , n296169 , n5742 , n296171 , n5744 , n296173 , 
 n296174 , n5747 , n5748 , n296177 , n296178 , n5751 , n5752 , n296181 , n296182 , n296183 , 
 n5756 , n5757 , n296186 , n5759 , n296188 , n296189 , n296190 , n296191 , n296192 , n296193 , 
 n296194 , n296195 , n5768 , n296197 , n296198 , n296199 , n5772 , n296201 , n296202 , n5775 , 
 n296204 , n296205 , n296206 , n296207 , n296208 , n296209 , n296210 , n296211 , n296212 , n296213 , 
 n5786 , n296215 , n296216 , n296217 , n296218 , n5791 , n296220 , n296221 , n296222 , n296223 , 
 n296224 , n296225 , n296226 , n296227 , n296228 , n296229 , n296230 , n5803 , n296232 , n5805 , 
 n296234 , n296235 , n296236 , n296237 , n296238 , n296239 , n5812 , n296241 , n296242 , n5815 , 
 n296244 , n296245 , n296246 , n5819 , n296248 , n296249 , n296250 , n296251 , n5824 , n296253 , 
 n296254 , n296255 , n296256 , n5829 , n296258 , n296259 , n296260 , n5833 , n5834 , n296263 , 
 n5836 , n296265 , n5838 , n5839 , n5840 , n5841 , n296270 , n5843 , n296272 , n5845 , 
 n296274 , n5847 , n5848 , n5849 , n296278 , n296279 , n5852 , n5853 , n5854 , n296283 , 
 n296284 , n5857 , n5858 , n5859 , n296288 , n296289 , n5862 , n5863 , n5864 , n296293 , 
 n296294 , n5867 , n296296 , n5869 , n296298 , n5871 , n5872 , n296301 , n296302 , n296303 , 
 n296304 , n296305 , n296306 , n296307 , n5880 , n5881 , n296310 , n296311 , n296312 , n296313 , 
 n296314 , n296315 , n296316 , n5889 , n296318 , n296319 , n5892 , n296321 , n5894 , n296323 , 
 n296324 , n5897 , n296326 , n5899 , n296328 , n296329 , n5902 , n296331 , n5904 , n296333 , 
 n296334 , n5907 , n296336 , n296337 , n296338 , n296339 , n296340 , n296341 , n296342 , n296343 , 
 n5916 , n296345 , n296346 , n296347 , n296348 , n5921 , n296350 , n296351 , n296352 , n296353 , 
 n296354 , n296355 , n296356 , n296357 , n5930 , n296359 , n296360 , n296361 , n296362 , n296363 , 
 n296364 , n296365 , n296366 , n5939 , n296368 , n296369 , n296370 , n296371 , n5944 , n296373 , 
 n5946 , n296375 , n296376 , n5949 , n296378 , n296379 , n5952 , n296381 , n296382 , n296383 , 
 n296384 , n5957 , n296386 , n5959 , n296388 , n296389 , n5962 , n296391 , n296392 , n296393 , 
 n296394 , n296395 , n296396 , n296397 , n5970 , n5971 , n296400 , n296401 , n296402 , n5975 , 
 n296404 , n296405 , n5978 , n296407 , n5980 , n296409 , n5982 , n296411 , n296412 , n5985 , 
 n296414 , n296415 , n5988 , n5989 , n296418 , n296419 , n296420 , n5993 , n296422 , n296423 , 
 n296424 , n296425 , n5998 , n296427 , n296428 , n6001 , n296430 , n6003 , n296432 , n296433 , 
 n296434 , n296435 , n296436 , n296437 , n6010 , n296439 , n296440 , n296441 , n296442 , n296443 , 
 n296444 , n6017 , n296446 , n6019 , n6020 , n6021 , n6022 , n6023 , n296452 , n6025 , 
 n296454 , n296455 , n6028 , n296457 , n6030 , n6031 , n296460 , n296461 , n6034 , n296463 , 
 n296464 , n6037 , n296466 , n296467 , n6040 , n296469 , n296470 , n6043 , n296472 , n296473 , 
 n6046 , n296475 , n6048 , n6049 , n296478 , n6051 , n296480 , n296481 , n296482 , n6055 , 
 n6056 , n6057 , n296486 , n6059 , n296488 , n6061 , n296490 , n296491 , n6064 , n296493 , 
 n296494 , n296495 , n296496 , n6069 , n296498 , n296499 , n296500 , n296501 , n296502 , n6075 , 
 n6076 , n296505 , n6078 , n6079 , n296508 , n296509 , n6082 , n6083 , n296512 , n6085 , 
 n296514 , n296515 , n296516 , n296517 , n296518 , n296519 , n296520 , n296521 , n296522 , n6095 , 
 n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n296531 , n296532 , n296533 , 
 n296534 , n296535 , n296536 , n296537 , n296538 , n296539 , n296540 , n296541 , n296542 , n6115 , 
 n6116 , n296545 , n296546 , n296547 , n296548 , n296549 , n6122 , n296551 , n296552 , n6125 , 
 n296554 , n6127 , n296556 , n296557 , n296558 , n296559 , n296560 , n296561 , n6134 , n6135 , 
 n296564 , n296565 , n6138 , n6139 , n296568 , n296569 , n6142 , n296571 , n6144 , n6145 , 
 n6146 , n296575 , n296576 , n296577 , n6150 , n296579 , n296580 , n6153 , n296582 , n6155 , 
 n6156 , n6157 , n6158 , n296587 , n6160 , n296589 , n6162 , n6163 , n296592 , n6165 , 
 n296594 , n6167 , n296596 , n296597 , n6170 , n296599 , n6172 , n296601 , n296602 , n6175 , 
 n6176 , n296605 , n296606 , n296607 , n296608 , n296609 , n296610 , n296611 , n296612 , n296613 , 
 n6186 , n296615 , n296616 , n296617 , n296618 , n6191 , n6192 , n296621 , n296622 , n296623 , 
 n296624 , n296625 , n296626 , n6199 , n296628 , n296629 , n6202 , n296631 , n296632 , n6205 , 
 n6206 , n296635 , n296636 , n6209 , n296638 , n296639 , n6212 , n296641 , n296642 , n296643 , 
 n296644 , n296645 , n296646 , n296647 , n296648 , n296649 , n296650 , n296651 , n296652 , n296653 , 
 n6226 , n296655 , n296656 , n296657 , n296658 , n6231 , n296660 , n6233 , n6234 , n296663 , 
 n296664 , n296665 , n296666 , n6239 , n296668 , n296669 , n296670 , n296671 , n296672 , n296673 , 
 n296674 , n296675 , n296676 , n296677 , n296678 , n296679 , n6252 , n296681 , n296682 , n296683 , 
 n296684 , n296685 , n296686 , n296687 , n296688 , n296689 , n296690 , n296691 , n296692 , n296693 , 
 n296694 , n296695 , n296696 , n296697 , n6270 , n296699 , n296700 , n6273 , n296702 , n296703 , 
 n6276 , n296705 , n296706 , n296707 , n296708 , n6281 , n296710 , n296711 , n296712 , n296713 , 
 n6286 , n296715 , n296716 , n296717 , n296718 , n6291 , n6292 , n296721 , n296722 , n296723 , 
 n296724 , n6297 , n296726 , n296727 , n6300 , n6301 , n296730 , n296731 , n6304 , n6305 , 
 n296734 , n296735 , n296736 , n296737 , n296738 , n6311 , n296740 , n296741 , n296742 , n6315 , 
 n296744 , n6317 , n296746 , n296747 , n6320 , n296749 , n296750 , n296751 , n6324 , n6325 , 
 n6326 , n296755 , n6328 , n6329 , n296758 , n6331 , n296760 , n296761 , n296762 , n6335 , 
 n6336 , n296765 , n296766 , n296767 , n6340 , n296769 , n296770 , n296771 , n296772 , n296773 , 
 n296774 , n296775 , n296776 , n296777 , n296778 , n6351 , n296780 , n296781 , n6354 , n296783 , 
 n6356 , n296785 , n296786 , n296787 , n296788 , n6361 , n296790 , n296791 , n296792 , n296793 , 
 n296794 , n296795 , n296796 , n296797 , n6370 , n296799 , n296800 , n6373 , n296802 , n6375 , 
 n6376 , n296805 , n6378 , n296807 , n296808 , n6381 , n296810 , n296811 , n296812 , n6385 , 
 n296814 , n296815 , n296816 , n296817 , n296818 , n296819 , n296820 , n6393 , n296822 , n296823 , 
 n296824 , n296825 , n296826 , n296827 , n6400 , n296829 , n296830 , n296831 , n296832 , n296833 , 
 n296834 , n6407 , n296836 , n296837 , n296838 , n296839 , n296840 , n296841 , n296842 , n6415 , 
 n296844 , n296845 , n296846 , n6419 , n296848 , n296849 , n296850 , n296851 , n296852 , n296853 , 
 n296854 , n296855 , n6428 , n296857 , n296858 , n6431 , n296860 , n296861 , n6434 , n296863 , 
 n296864 , n296865 , n296866 , n296867 , n296868 , n296869 , n296870 , n296871 , n296872 , n6445 , 
 n296874 , n296875 , n296876 , n296877 , n296878 , n296879 , n296880 , n296881 , n6454 , n6455 , 
 n296884 , n296885 , n296886 , n296887 , n296888 , n296889 , n296890 , n296891 , n296892 , n296893 , 
 n296894 , n6467 , n6468 , n296897 , n6470 , n296899 , n296900 , n296901 , n296902 , n296903 , 
 n6476 , n296905 , n296906 , n6479 , n296908 , n296909 , n296910 , n296911 , n6484 , n296913 , 
 n296914 , n6487 , n6488 , n296917 , n296918 , n6491 , n296920 , n296921 , n6494 , n296923 , 
 n296924 , n6497 , n296926 , n296927 , n6500 , n296929 , n6502 , n296931 , n296932 , n296933 , 
 n296934 , n296935 , n296936 , n6509 , n296938 , n296939 , n296940 , n296941 , n6514 , n296943 , 
 n296944 , n296945 , n296946 , n6519 , n296948 , n296949 , n296950 , n296951 , n296952 , n296953 , 
 n296954 , n296955 , n296956 , n6529 , n296958 , n296959 , n296960 , n296961 , n296962 , n6535 , 
 n296964 , n296965 , n296966 , n296967 , n296968 , n6541 , n296970 , n296971 , n296972 , n296973 , 
 n296974 , n6547 , n296976 , n6549 , n6550 , n6551 , n6552 , n296981 , n6554 , n296983 , 
 n296984 , n6557 , n296986 , n296987 , n6560 , n296989 , n296990 , n296991 , n296992 , n296993 , 
 n6566 , n296995 , n6568 , n296997 , n296998 , n296999 , n297000 , n6573 , n297002 , n297003 , 
 n6576 , n6577 , n297006 , n6579 , n297008 , n297009 , n297010 , n6583 , n6584 , n297013 , 
 n297014 , n297015 , n297016 , n297017 , n6590 , n297019 , n6592 , n6593 , n297022 , n297023 , 
 n297024 , n6597 , n297026 , n297027 , n6600 , n297029 , n297030 , n297031 , n297032 , n6605 , 
 n297034 , n297035 , n297036 , n297037 , n297038 , n297039 , n297040 , n297041 , n297042 , n6615 , 
 n297044 , n297045 , n6618 , n297047 , n297048 , n6621 , n297050 , n297051 , n6624 , n297053 , 
 n6626 , n297055 , n297056 , n6629 , n297058 , n297059 , n297060 , n297061 , n6634 , n297063 , 
 n297064 , n297065 , n297066 , n297067 , n297068 , n297069 , n297070 , n6643 , n297072 , n297073 , 
 n297074 , n297075 , n6648 , n297077 , n6650 , n6651 , n6652 , n297081 , n6654 , n297083 , 
 n6656 , n6657 , n297086 , n297087 , n6660 , n297089 , n297090 , n6663 , n297092 , n6665 , 
 n6666 , n297095 , n297096 , n297097 , n297098 , n297099 , n297100 , n6673 , n297102 , n297103 , 
 n297104 , n6677 , n6678 , n6679 , n297108 , n297109 , n297110 , n297111 , n297112 , n6685 , 
 n297114 , n297115 , n6688 , n6689 , n6690 , n6691 , n297120 , n6693 , n297122 , n6695 , 
 n6696 , n297125 , n297126 , n297127 , n297128 , n297129 , n6702 , n297131 , n6704 , n6705 , 
 n6706 , n297135 , n297136 , n297137 , n6710 , n297139 , n297140 , n297141 , n6714 , n6715 , 
 n297144 , n297145 , n297146 , n6719 , n297148 , n297149 , n6722 , n297151 , n297152 , n6725 , 
 n297154 , n297155 , n297156 , n297157 , n297158 , n297159 , n297160 , n297161 , n6734 , n6735 , 
 n297164 , n297165 , n297166 , n297167 , n297168 , n6741 , n297170 , n297171 , n6744 , n297173 , 
 n6746 , n297175 , n297176 , n6749 , n6750 , n297179 , n297180 , n297181 , n297182 , n297183 , 
 n6756 , n297185 , n297186 , n6759 , n6760 , n6761 , n297190 , n297191 , n6764 , n297193 , 
 n6766 , n297195 , n6768 , n6769 , n6770 , n6771 , n297200 , n6773 , n297202 , n297203 , 
 n297204 , n297205 , n297206 , n297207 , n297208 , n297209 , n6782 , n297211 , n6784 , n6785 , 
 n6786 , n6787 , n297216 , n6789 , n297218 , n297219 , n297220 , n297221 , n297222 , n297223 , 
 n6796 , n6797 , n297226 , n6799 , n6800 , n297229 , n297230 , n297231 , n6804 , n6805 , 
 n297234 , n6807 , n6808 , n297237 , n297238 , n6811 , n6812 , n6813 , n297242 , n297243 , 
 n297244 , n297245 , n6818 , n297247 , n6820 , n297249 , n6822 , n297251 , n297252 , n6825 , 
 n297254 , n297255 , n297256 , n6829 , n297258 , n297259 , n297260 , n6833 , n6834 , n297263 , 
 n297264 , n297265 , n6838 , n6839 , n6840 , n297269 , n297270 , n6843 , n297272 , n297273 , 
 n297274 , n297275 , n297276 , n6849 , n6850 , n297279 , n297280 , n297281 , n297282 , n297283 , 
 n6856 , n297285 , n297286 , n297287 , n297288 , n297289 , n6862 , n297291 , n297292 , n297293 , 
 n297294 , n297295 , n297296 , n297297 , n297298 , n6871 , n297300 , n297301 , n297302 , n6875 , 
 n6876 , n297305 , n6878 , n297307 , n297308 , n297309 , n6882 , n297311 , n6884 , n297313 , 
 n6886 , n297315 , n6888 , n6889 , n297318 , n6891 , n297320 , n6893 , n297322 , n297323 , 
 n297324 , n297325 , n297326 , n6899 , n297328 , n6901 , n297330 , n297331 , n297332 , n297333 , 
 n6906 , n297335 , n6908 , n6909 , n6910 , n297339 , n297340 , n297341 , n297342 , n297343 , 
 n297344 , n297345 , n6918 , n297347 , n6920 , n6921 , n297350 , n297351 , n6924 , n297353 , 
 n297354 , n6927 , n297356 , n297357 , n6930 , n297359 , n6932 , n6933 , n297362 , n297363 , 
 n297364 , n6937 , n297366 , n297367 , n297368 , n297369 , n297370 , n297371 , n297372 , n297373 , 
 n297374 , n6947 , n297376 , n6949 , n297378 , n297379 , n297380 , n297381 , n6954 , n6955 , 
 n297384 , n297385 , n297386 , n6959 , n6960 , n6961 , n297390 , n6963 , n297392 , n297393 , 
 n6966 , n297395 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n297402 , n6975 , 
 n297404 , n297405 , n297406 , n6979 , n297408 , n297409 , n297410 , n297411 , n297412 , n297413 , 
 n297414 , n297415 , n297416 , n297417 , n297418 , n297419 , n297420 , n297421 , n6994 , n297423 , 
 n297424 , n6997 , n297426 , n297427 , n7000 , n297429 , n7002 , n297431 , n297432 , n297433 , 
 n297434 , n297435 , n297436 , n297437 , n297438 , n297439 , n7012 , n297441 , n297442 , n7015 , 
 n297444 , n297445 , n7018 , n7019 , n297448 , n297449 , n297450 , n297451 , n7024 , n297453 , 
 n297454 , n7027 , n297456 , n297457 , n297458 , n297459 , n7032 , n297461 , n7034 , n297463 , 
 n297464 , n297465 , n297466 , n7039 , n7040 , n297469 , n297470 , n297471 , n297472 , n297473 , 
 n297474 , n7047 , n297476 , n297477 , n7050 , n297479 , n297480 , n7053 , n7054 , n297483 , 
 n7056 , n297485 , n297486 , n297487 , n297488 , n297489 , n297490 , n7063 , n297492 , n7065 , 
 n7066 , n297495 , n297496 , n297497 , n7070 , n297499 , n297500 , n297501 , n297502 , n7075 , 
 n297504 , n297505 , n7078 , n297507 , n297508 , n297509 , n297510 , n297511 , n297512 , n297513 , 
 n7086 , n7087 , n297516 , n297517 , n297518 , n7091 , n7092 , n297521 , n297522 , n297523 , 
 n7096 , n297525 , n297526 , n7099 , n297528 , n7101 , n7102 , n7103 , n7104 , n297533 , 
 n7106 , n7107 , n7108 , n297537 , n7110 , n7111 , n7112 , n297541 , n297542 , n7115 , 
 n7116 , n297545 , n297546 , n297547 , n297548 , n7121 , n297550 , n297551 , n297552 , n297553 , 
 n7126 , n7127 , n297556 , n7129 , n7130 , n297559 , n297560 , n297561 , n297562 , n297563 , 
 n297564 , n7137 , n297566 , n7139 , n7140 , n297569 , n297570 , n7143 , n297572 , n297573 , 
 n297574 , n297575 , n7148 , n297577 , n297578 , n297579 , n297580 , n297581 , n297582 , n7155 , 
 n297584 , n297585 , n297586 , n297587 , n297588 , n297589 , n297590 , n297591 , n297592 , n7165 , 
 n297594 , n297595 , n297596 , n297597 , n297598 , n297599 , n297600 , n297601 , n297602 , n297603 , 
 n7176 , n297605 , n7178 , n7179 , n297608 , n297609 , n7182 , n297611 , n297612 , n297613 , 
 n297614 , n297615 , n297616 , n297617 , n297618 , n7191 , n7192 , n297621 , n297622 , n297623 , 
 n297624 , n297625 , n297626 , n297627 , n297628 , n297629 , n7202 , n297631 , n297632 , n7205 , 
 n297634 , n297635 , n7208 , n7209 , n7210 , n7211 , n297640 , n297641 , n297642 , n297643 , 
 n7216 , n7217 , n7218 , n297647 , n297648 , n297649 , n297650 , n7223 , n297652 , n297653 , 
 n297654 , n297655 , n297656 , n297657 , n297658 , n7231 , n297660 , n297661 , n297662 , n297663 , 
 n297664 , n297665 , n7238 , n297667 , n297668 , n7241 , n297670 , n7243 , n297672 , n297673 , 
 n7246 , n297675 , n7248 , n297677 , n7250 , n297679 , n297680 , n297681 , n297682 , n297683 , 
 n297684 , n7257 , n297686 , n7259 , n297688 , n297689 , n297690 , n297691 , n297692 , n297693 , 
 n297694 , n297695 , n297696 , n7269 , n297698 , n297699 , n297700 , n297701 , n297702 , n297703 , 
 n297704 , n297705 , n297706 , n297707 , n7280 , n297709 , n297710 , n7283 , n297712 , n297713 , 
 n7286 , n297715 , n297716 , n7289 , n297718 , n297719 , n7292 , n297721 , n297722 , n297723 , 
 n297724 , n297725 , n297726 , n297727 , n297728 , n7301 , n297730 , n297731 , n7304 , n297733 , 
 n297734 , n7307 , n297736 , n297737 , n297738 , n297739 , n297740 , n297741 , n297742 , n7315 , 
 n297744 , n297745 , n297746 , n297747 , n297748 , n297749 , n297750 , n297751 , n297752 , n297753 , 
 n297754 , n7327 , n297756 , n297757 , n297758 , n297759 , n7332 , n297761 , n297762 , n7335 , 
 n297764 , n297765 , n7338 , n297767 , n7340 , n7341 , n297770 , n297771 , n297772 , n297773 , 
 n297774 , n297775 , n297776 , n297777 , n7350 , n7351 , n297780 , n7353 , n297782 , n297783 , 
 n297784 , n297785 , n7358 , n297787 , n297788 , n7361 , n297790 , n7363 , n297792 , n297793 , 
 n7366 , n297795 , n7368 , n297797 , n297798 , n297799 , n7372 , n297801 , n297802 , n7375 , 
 n297804 , n297805 , n7378 , n297807 , n7380 , n297809 , n7382 , n7383 , n297812 , n297813 , 
 n7386 , n7387 , n297816 , n297817 , n7390 , n297819 , n297820 , n297821 , n297822 , n297823 , 
 n297824 , n7397 , n297826 , n297827 , n7400 , n297829 , n7402 , n7403 , n297832 , n297833 , 
 n297834 , n297835 , n297836 , n7409 , n297838 , n297839 , n7412 , n297841 , n297842 , n7415 , 
 n297844 , n7417 , n7418 , n297847 , n297848 , n7421 , n297850 , n7423 , n297852 , n7425 , 
 n297854 , n297855 , n7428 , n297857 , n7430 , n297859 , n7432 , n7433 , n7434 , n297863 , 
 n297864 , n7437 , n7438 , n7439 , n297868 , n297869 , n7442 , n297871 , n7444 , n7445 , 
 n7446 , n297875 , n7448 , n7449 , n297878 , n297879 , n297880 , n7453 , n297882 , n297883 , 
 n297884 , n297885 , n297886 , n297887 , n7460 , n297889 , n7462 , n297891 , n297892 , n297893 , 
 n297894 , n7467 , n297896 , n297897 , n297898 , n297899 , n297900 , n297901 , n7474 , n297903 , 
 n297904 , n7477 , n297906 , n297907 , n297908 , n7481 , n297910 , n7483 , n297912 , n297913 , 
 n7486 , n297915 , n297916 , n7489 , n297918 , n297919 , n297920 , n297921 , n297922 , n297923 , 
 n7496 , n297925 , n7498 , n7499 , n297928 , n7501 , n7502 , n7503 , n297932 , n7505 , 
 n7506 , n297935 , n7508 , n297937 , n297938 , n297939 , n7512 , n297941 , n297942 , n297943 , 
 n7516 , n7517 , n7518 , n297947 , n7520 , n7521 , n297950 , n7523 , n297952 , n297953 , 
 n7526 , n297955 , n297956 , n7529 , n297958 , n7531 , n7532 , n297961 , n297962 , n7535 , 
 n297964 , n297965 , n297966 , n297967 , n297968 , n297969 , n297970 , n297971 , n7544 , n297973 , 
 n297974 , n297975 , n297976 , n297977 , n297978 , n7551 , n297980 , n297981 , n7554 , n297983 , 
 n297984 , n7557 , n297986 , n297987 , n7560 , n297989 , n7562 , n297991 , n297992 , n297993 , 
 n297994 , n297995 , n297996 , n297997 , n297998 , n297999 , n298000 , n298001 , n298002 , n298003 , 
 n298004 , n298005 , n298006 , n7579 , n298008 , n298009 , n298010 , n298011 , n298012 , n298013 , 
 n298014 , n298015 , n7588 , n298017 , n298018 , n298019 , n298020 , n298021 , n298022 , n298023 , 
 n298024 , n298025 , n298026 , n7599 , n298028 , n298029 , n298030 , n298031 , n298032 , n298033 , 
 n298034 , n298035 , n298036 , n298037 , n298038 , n7611 , n298040 , n298041 , n298042 , n7615 , 
 n7616 , n298045 , n7618 , n298047 , n298048 , n298049 , n298050 , n298051 , n298052 , n298053 , 
 n7626 , n298055 , n298056 , n298057 , n298058 , n7631 , n298060 , n298061 , n7634 , n298063 , 
 n298064 , n298065 , n298066 , n298067 , n298068 , n298069 , n298070 , n298071 , n7644 , n298073 , 
 n298074 , n298075 , n298076 , n7649 , n298078 , n298079 , n298080 , n298081 , n298082 , n7655 , 
 n298084 , n298085 , n7658 , n298087 , n7660 , n298089 , n7662 , n7663 , n7664 , n7665 , 
 n7666 , n7667 , n7668 , n298097 , n7670 , n298099 , n298100 , n7673 , n298102 , n7675 , 
 n7676 , n7677 , n7678 , n298107 , n298108 , n298109 , n7682 , n298111 , n298112 , n298113 , 
 n298114 , n298115 , n7688 , n298117 , n298118 , n298119 , n298120 , n7693 , n7694 , n7695 , 
 n298124 , n7697 , n7698 , n7699 , n7700 , n7701 , n298130 , n298131 , n298132 , n7705 , 
 n298134 , n298135 , n7708 , n298137 , n7710 , n7711 , n298140 , n298141 , n298142 , n7715 , 
 n298144 , n298145 , n7718 , n298147 , n298148 , n298149 , n298150 , n298151 , n298152 , n298153 , 
 n298154 , n298155 , n298156 , n298157 , n7730 , n298159 , n298160 , n7733 , n298162 , n7735 , 
 n298164 , n298165 , n298166 , n298167 , n7740 , n7741 , n298170 , n298171 , n7744 , n298173 , 
 n7746 , n298175 , n298176 , n298177 , n298178 , n7751 , n298180 , n298181 , n298182 , n298183 , 
 n298184 , n298185 , n298186 , n298187 , n298188 , n298189 , n298190 , n298191 , n298192 , n7765 , 
 n298194 , n298195 , n298196 , n7769 , n298198 , n298199 , n298200 , n298201 , n298202 , n7775 , 
 n298204 , n298205 , n298206 , n7779 , n298208 , n298209 , n7782 , n298211 , n298212 , n298213 , 
 n298214 , n298215 , n7788 , n298217 , n298218 , n7791 , n298220 , n7793 , n7794 , n7795 , 
 n7796 , n7797 , n298226 , n298227 , n7800 , n298229 , n7802 , n7803 , n7804 , n7805 , 
 n7806 , n7807 , n298236 , n298237 , n7810 , n298239 , n298240 , n7813 , n298242 , n7815 , 
 n7816 , n298245 , n7818 , n7819 , n298248 , n298249 , n7822 , n298251 , n298252 , n7825 , 
 n7826 , n298255 , n298256 , n7829 , n298258 , n298259 , n7832 , n298261 , n7834 , n298263 , 
 n298264 , n298265 , n298266 , n298267 , n298268 , n7841 , n298270 , n298271 , n7844 , n7845 , 
 n7846 , n7847 , n298276 , n298277 , n7850 , n7851 , n298280 , n298281 , n298282 , n298283 , 
 n298284 , n7857 , n298286 , n298287 , n7860 , n298289 , n7862 , n7863 , n298292 , n298293 , 
 n7866 , n298295 , n298296 , n7869 , n298298 , n298299 , n7872 , n298301 , n298302 , n298303 , 
 n298304 , n7877 , n298306 , n298307 , n7880 , n298309 , n7882 , n7883 , n7884 , n298313 , 
 n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n298322 , n7895 , 
 n7896 , n298325 , n7898 , n298327 , n7900 , n298329 , n298330 , n7903 , n7904 , n7905 , 
 n298334 , n7907 , n7908 , n7909 , n298338 , n298339 , n298340 , n7913 , n7914 , n7915 , 
 n7916 , n298345 , n298346 , n7919 , n7920 , n7921 , n7922 , n298351 , n7924 , n7925 , 
 n298354 , n298355 , n298356 , n7929 , n298358 , n298359 , n7932 , n7933 , n298362 , n298363 , 
 n7936 , n298365 , n298366 , n7939 , n298368 , n298369 , n7942 , n298371 , n7944 , n7945 , 
 n7946 , n298375 , n7948 , n7949 , n298378 , n7951 , n298380 , n298381 , n7954 , n7955 , 
 n298384 , n7957 , n7958 , n7959 , n7960 , n298389 , n298390 , n7963 , n298392 , n7965 , 
 n298394 , n298395 , n298396 , n7969 , n7970 , n298399 , n298400 , n298401 , n298402 , n7975 , 
 n7976 , n298405 , n7978 , n7979 , n298408 , n298409 , n298410 , n298411 , n7984 , n298413 , 
 n298414 , n7987 , n298416 , n7989 , n298418 , n298419 , n298420 , n298421 , n298422 , n298423 , 
 n7996 , n298425 , n298426 , n7999 , n298428 , n298429 , n298430 , n8003 , n8004 , n8005 , 
 n8006 , n298435 , n298436 , n298437 , n8010 , n298439 , n298440 , n8013 , n298442 , n8015 , 
 n8016 , n298445 , n298446 , n298447 , n298448 , n298449 , n298450 , n298451 , n298452 , n8025 , 
 n298454 , n298455 , n298456 , n298457 , n298458 , n298459 , n298460 , n8033 , n298462 , n298463 , 
 n298464 , n298465 , n298466 , n298467 , n8040 , n298469 , n298470 , n298471 , n8044 , n8045 , 
 n298474 , n298475 , n298476 , n8049 , n298478 , n298479 , n298480 , n298481 , n298482 , n298483 , 
 n298484 , n8057 , n298486 , n298487 , n298488 , n8061 , n8062 , n298491 , n298492 , n298493 , 
 n8066 , n8067 , n298496 , n8069 , n298498 , n298499 , n298500 , n298501 , n8074 , n298503 , 
 n298504 , n298505 , n298506 , n298507 , n298508 , n8081 , n298510 , n298511 , n8084 , n298513 , 
 n298514 , n8087 , n298516 , n8089 , n298518 , n298519 , n298520 , n8093 , n298522 , n298523 , 
 n8096 , n298525 , n298526 , n298527 , n298528 , n298529 , n8102 , n298531 , n298532 , n8105 , 
 n298534 , n298535 , n298536 , n298537 , n298538 , n298539 , n298540 , n8113 , n298542 , n298543 , 
 n298544 , n298545 , n8118 , n298547 , n298548 , n8121 , n298550 , n8123 , n298552 , n298553 , 
 n8126 , n298555 , n298556 , n298557 , n298558 , n298559 , n298560 , n298561 , n298562 , n8135 , 
 n298564 , n298565 , n298566 , n298567 , n298568 , n298569 , n8142 , n8143 , n298572 , n298573 , 
 n298574 , n298575 , n298576 , n8149 , n298578 , n298579 , n8152 , n8153 , n298582 , n298583 , 
 n298584 , n298585 , n8158 , n298587 , n298588 , n8161 , n8162 , n298591 , n298592 , n298593 , 
 n298594 , n298595 , n298596 , n8169 , n298598 , n298599 , n8172 , n8173 , n8174 , n8175 , 
 n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n298611 , n298612 , n298613 , 
 n298614 , n298615 , n298616 , n298617 , n298618 , n298619 , n298620 , n298621 , n8194 , n298623 , 
 n298624 , n298625 , n298626 , n298627 , n298628 , n298629 , n298630 , n8203 , n298632 , n8205 , 
 n298634 , n298635 , n298636 , n298637 , n298638 , n298639 , n298640 , n298641 , n298642 , n298643 , 
 n8216 , n8217 , n298646 , n298647 , n8220 , n298649 , n298650 , n298651 , n298652 , n298653 , 
 n298654 , n298655 , n298656 , n298657 , n298658 , n298659 , n298660 , n298661 , n298662 , n298663 , 
 n298664 , n298665 , n298666 , n298667 , n298668 , n298669 , n298670 , n298671 , n298672 , n298673 , 
 n8246 , n8247 , n298676 , n8249 , n298678 , n298679 , n8252 , n8253 , n298682 , n8255 , 
 n298684 , n298685 , n298686 , n8259 , n298688 , n298689 , n298690 , n298691 , n8264 , n298693 , 
 n298694 , n298695 , n298696 , n298697 , n8270 , n298699 , n298700 , n298701 , n8274 , n298703 , 
 n298704 , n8277 , n298706 , n298707 , n8280 , n8281 , n298710 , n8283 , n298712 , n8285 , 
 n298714 , n298715 , n298716 , n298717 , n298718 , n298719 , n8292 , n298721 , n298722 , n8295 , 
 n8296 , n298725 , n298726 , n8299 , n298728 , n298729 , n8302 , n298731 , n298732 , n298733 , 
 n298734 , n298735 , n298736 , n298737 , n298738 , n298739 , n298740 , n298741 , n298742 , n298743 , 
 n298744 , n8317 , n298746 , n298747 , n298748 , n298749 , n8322 , n298751 , n298752 , n8325 , 
 n298754 , n298755 , n8328 , n298757 , n298758 , n298759 , n298760 , n8333 , n298762 , n298763 , 
 n298764 , n8337 , n298766 , n298767 , n8340 , n298769 , n8342 , n298771 , n298772 , n8345 , 
 n298774 , n298775 , n8348 , n298777 , n8350 , n8351 , n298780 , n8353 , n8354 , n298783 , 
 n298784 , n298785 , n298786 , n298787 , n8360 , n298789 , n298790 , n8363 , n8364 , n298793 , 
 n298794 , n8367 , n298796 , n298797 , n298798 , n298799 , n298800 , n8373 , n298802 , n298803 , 
 n298804 , n298805 , n298806 , n8379 , n8380 , n298809 , n8382 , n298811 , n8384 , n8385 , 
 n8386 , n298815 , n8388 , n8389 , n298818 , n298819 , n298820 , n298821 , n8394 , n8395 , 
 n298824 , n298825 , n8398 , n298827 , n8400 , n298829 , n298830 , n298831 , n8404 , n298833 , 
 n298834 , n298835 , n298836 , n298837 , n298838 , n298839 , n298840 , n8413 , n298842 , n298843 , 
 n298844 , n8417 , n298846 , n298847 , n298848 , n298849 , n298850 , n298851 , n298852 , n8425 , 
 n298854 , n8427 , n298856 , n298857 , n8430 , n8431 , n298860 , n298861 , n8434 , n298863 , 
 n8436 , n8437 , n8438 , n8439 , n298868 , n8441 , n8442 , n8443 , n8444 , n8445 , 
 n8446 , n298875 , n298876 , n8449 , n298878 , n298879 , n8452 , n298881 , n8454 , n8455 , 
 n298884 , n298885 , n8458 , n298887 , n298888 , n8461 , n298890 , n298891 , n298892 , n298893 , 
 n8466 , n298895 , n298896 , n8469 , n298898 , n298899 , n8472 , n298901 , n8474 , n298903 , 
 n298904 , n298905 , n298906 , n8479 , n298908 , n298909 , n8482 , n298911 , n298912 , n8485 , 
 n298914 , n298915 , n298916 , n298917 , n298918 , n298919 , n8492 , n298921 , n298922 , n298923 , 
 n8496 , n8497 , n8498 , n8499 , n8500 , n298929 , n8502 , n298931 , n8504 , n8505 , 
 n298934 , n298935 , n298936 , n298937 , n8510 , n298939 , n8512 , n8513 , n8514 , n8515 , 
 n298944 , n298945 , n298946 , n298947 , n298948 , n298949 , n298950 , n298951 , n298952 , n298953 , 
 n8526 , n298955 , n298956 , n298957 , n298958 , n8531 , n8532 , n298961 , n298962 , n298963 , 
 n8536 , n298965 , n298966 , n8539 , n298968 , n298969 , n8542 , n298971 , n298972 , n298973 , 
 n298974 , n298975 , n298976 , n298977 , n298978 , n8551 , n298980 , n298981 , n8554 , n298983 , 
 n298984 , n298985 , n298986 , n298987 , n298988 , n8561 , n298990 , n298991 , n8564 , n298993 , 
 n298994 , n298995 , n298996 , n8569 , n298998 , n298999 , n8572 , n299001 , n299002 , n299003 , 
 n299004 , n8577 , n8578 , n299007 , n299008 , n8581 , n299010 , n299011 , n299012 , n299013 , 
 n299014 , n8587 , n299016 , n299017 , n8590 , n8591 , n299020 , n299021 , n8594 , n299023 , 
 n299024 , n299025 , n299026 , n299027 , n299028 , n299029 , n8602 , n299031 , n299032 , n8605 , 
 n299034 , n299035 , n299036 , n299037 , n8610 , n299039 , n299040 , n299041 , n8614 , n299043 , 
 n8616 , n299045 , n299046 , n8619 , n8620 , n8621 , n299050 , n8623 , n299052 , n299053 , 
 n8626 , n299055 , n8628 , n299057 , n8630 , n8631 , n299060 , n299061 , n8634 , n299063 , 
 n299064 , n8637 , n299066 , n299067 , n8640 , n8641 , n8642 , n299071 , n299072 , n8645 , 
 n299074 , n299075 , n299076 , n8649 , n299078 , n299079 , n299080 , n299081 , n299082 , n299083 , 
 n8656 , n8657 , n299086 , n299087 , n299088 , n299089 , n299090 , n299091 , n299092 , n299093 , 
 n299094 , n8667 , n299096 , n299097 , n8670 , n299099 , n299100 , n8673 , n299102 , n299103 , 
 n299104 , n299105 , n299106 , n299107 , n8680 , n299109 , n299110 , n299111 , n8684 , n299113 , 
 n299114 , n299115 , n299116 , n299117 , n299118 , n299119 , n8692 , n299121 , n299122 , n8695 , 
 n8696 , n8697 , n299126 , n299127 , n8700 , n299129 , n299130 , n8703 , n299132 , n299133 , 
 n299134 , n299135 , n299136 , n299137 , n8710 , n299139 , n299140 , n8713 , n299142 , n299143 , 
 n299144 , n299145 , n8718 , n299147 , n8720 , n8721 , n299150 , n299151 , n299152 , n299153 , 
 n299154 , n299155 , n8728 , n299157 , n299158 , n299159 , n299160 , n299161 , n8734 , n299163 , 
 n299164 , n299165 , n299166 , n299167 , n8740 , n299169 , n299170 , n299171 , n8744 , n299173 , 
 n299174 , n299175 , n299176 , n299177 , n8750 , n8751 , n8752 , n299181 , n299182 , n8755 , 
 n8756 , n8757 , n8758 , n299187 , n299188 , n8761 , n299190 , n299191 , n299192 , n8765 , 
 n299194 , n299195 , n8768 , n299197 , n299198 , n8771 , n299200 , n299201 , n8774 , n299203 , 
 n299204 , n299205 , n299206 , n299207 , n8780 , n299209 , n299210 , n299211 , n299212 , n299213 , 
 n299214 , n299215 , n299216 , n299217 , n299218 , n299219 , n299220 , n8793 , n299222 , n299223 , 
 n299224 , n299225 , n299226 , n299227 , n8800 , n299229 , n299230 , n299231 , n299232 , n299233 , 
 n299234 , n299235 , n8808 , n8809 , n299238 , n299239 , n8812 , n299241 , n299242 , n8815 , 
 n299244 , n299245 , n8818 , n299247 , n8820 , n299249 , n8822 , n299251 , n299252 , n8825 , 
 n299254 , n299255 , n299256 , n299257 , n8830 , n299259 , n299260 , n8833 , n299262 , n299263 , 
 n8836 , n299265 , n299266 , n299267 , n299268 , n8841 , n299270 , n299271 , n299272 , n299273 , 
 n299274 , n299275 , n299276 , n299277 , n299278 , n299279 , n299280 , n8853 , n299282 , n8855 , 
 n299284 , n299285 , n299286 , n299287 , n8860 , n299289 , n8862 , n299291 , n8864 , n299293 , 
 n8866 , n8867 , n299296 , n8869 , n299298 , n299299 , n299300 , n299301 , n8874 , n299303 , 
 n299304 , n299305 , n8878 , n299307 , n299308 , n299309 , n299310 , n299311 , n8884 , n299313 , 
 n299314 , n8887 , n299316 , n299317 , n299318 , n299319 , n299320 , n299321 , n299322 , n299323 , 
 n299324 , n299325 , n299326 , n299327 , n8900 , n299329 , n299330 , n299331 , n8904 , n299333 , 
 n299334 , n299335 , n299336 , n299337 , n8910 , n299339 , n299340 , n8913 , n299342 , n299343 , 
 n299344 , n299345 , n299346 , n299347 , n299348 , n299349 , n299350 , n8923 , n299352 , n299353 , 
 n299354 , n299355 , n299356 , n299357 , n299358 , n299359 , n299360 , n299361 , n8934 , n299363 , 
 n299364 , n299365 , n299366 , n8939 , n299368 , n299369 , n299370 , n299371 , n299372 , n299373 , 
 n299374 , n299375 , n299376 , n299377 , n299378 , n8951 , n299380 , n299381 , n8954 , n299383 , 
 n299384 , n299385 , n8958 , n299387 , n299388 , n8961 , n299390 , n8963 , n299392 , n299393 , 
 n299394 , n299395 , n8968 , n299397 , n299398 , n299399 , n8972 , n299401 , n299402 , n299403 , 
 n299404 , n8977 , n299406 , n299407 , n8980 , n299409 , n8982 , n299411 , n299412 , n299413 , 
 n299414 , n8987 , n299416 , n8989 , n8990 , n8991 , n299420 , n8993 , n299422 , n299423 , 
 n8996 , n299425 , n8998 , n299427 , n299428 , n299429 , n299430 , n299431 , n9004 , n299433 , 
 n9006 , n299435 , n299436 , n299437 , n299438 , n299439 , n299440 , n299441 , n9014 , n299443 , 
 n299444 , n299445 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n299453 , 
 n299454 , n299455 , n299456 , n299457 , n9030 , n299459 , n299460 , n9033 , n299462 , n299463 , 
 n9036 , n299465 , n299466 , n9039 , n299468 , n299469 , n9042 , n299471 , n299472 , n299473 , 
 n299474 , n299475 , n299476 , n299477 , n299478 , n299479 , n9052 , n299481 , n299482 , n9055 , 
 n299484 , n299485 , n299486 , n299487 , n299488 , n299489 , n299490 , n299491 , n299492 , n299493 , 
 n9066 , n299495 , n299496 , n299497 , n299498 , n299499 , n299500 , n299501 , n299502 , n299503 , 
 n299504 , n299505 , n299506 , n299507 , n299508 , n299509 , n299510 , n299511 , n299512 , n9085 , 
 n299514 , n299515 , n299516 , n299517 , n9090 , n299519 , n299520 , n299521 , n299522 , n299523 , 
 n299524 , n299525 , n299526 , n299527 , n9100 , n299529 , n299530 , n299531 , n299532 , n299533 , 
 n9106 , n9107 , n299536 , n299537 , n9110 , n9111 , n9112 , n299541 , n299542 , n299543 , 
 n299544 , n9117 , n299546 , n299547 , n9120 , n9121 , n9122 , n299551 , n299552 , n9125 , 
 n9126 , n299555 , n299556 , n299557 , n9130 , n299559 , n299560 , n299561 , n299562 , n299563 , 
 n299564 , n299565 , n299566 , n299567 , n299568 , n299569 , n299570 , n299571 , n299572 , n9145 , 
 n9146 , n299575 , n299576 , n299577 , n9150 , n9151 , n9152 , n9153 , n299582 , n299583 , 
 n299584 , n299585 , n9158 , n299587 , n299588 , n299589 , n299590 , n299591 , n9164 , n299593 , 
 n299594 , n9167 , n299596 , n299597 , n9170 , n299599 , n9172 , n299601 , n299602 , n299603 , 
 n299604 , n299605 , n299606 , n299607 , n299608 , n9181 , n9182 , n299611 , n9184 , n299613 , 
 n299614 , n299615 , n299616 , n299617 , n299618 , n9191 , n299620 , n299621 , n9194 , n299623 , 
 n299624 , n299625 , n299626 , n299627 , n9200 , n299629 , n299630 , n9203 , n299632 , n299633 , 
 n9206 , n9207 , n299636 , n299637 , n299638 , n299639 , n299640 , n9213 , n299642 , n299643 , 
 n9216 , n299645 , n299646 , n9219 , n9220 , n299649 , n9222 , n299651 , n9224 , n9225 , 
 n9226 , n9227 , n9228 , n9229 , n299658 , n9231 , n299660 , n9233 , n299662 , n299663 , 
 n299664 , n9237 , n299666 , n299667 , n9240 , n299669 , n9242 , n299671 , n299672 , n299673 , 
 n9246 , n299675 , n299676 , n299677 , n9250 , n299679 , n9252 , n299681 , n299682 , n299683 , 
 n9256 , n299685 , n299686 , n9259 , n299688 , n299689 , n9262 , n299691 , n299692 , n299693 , 
 n299694 , n299695 , n299696 , n299697 , n299698 , n299699 , n9272 , n299701 , n299702 , n9275 , 
 n299704 , n9277 , n299706 , n299707 , n299708 , n9281 , n299710 , n299711 , n9284 , n299713 , 
 n299714 , n299715 , n299716 , n299717 , n299718 , n299719 , n9292 , n299721 , n299722 , n299723 , 
 n299724 , n299725 , n299726 , n299727 , n9300 , n299729 , n299730 , n299731 , n299732 , n299733 , 
 n299734 , n299735 , n299736 , n299737 , n9310 , n299739 , n299740 , n299741 , n9314 , n299743 , 
 n299744 , n299745 , n9318 , n299747 , n299748 , n299749 , n299750 , n299751 , n299752 , n9325 , 
 n299754 , n299755 , n299756 , n299757 , n299758 , n299759 , n299760 , n299761 , n9334 , n299763 , 
 n299764 , n9337 , n299766 , n299767 , n299768 , n299769 , n9342 , n299771 , n299772 , n299773 , 
 n9346 , n9347 , n9348 , n299777 , n299778 , n9351 , n9352 , n9353 , n9354 , n299783 , 
 n9356 , n9357 , n9358 , n299787 , n299788 , n299789 , n299790 , n9363 , n299792 , n299793 , 
 n9366 , n299795 , n299796 , n299797 , n299798 , n299799 , n299800 , n299801 , n9374 , n299803 , 
 n299804 , n299805 , n299806 , n299807 , n299808 , n299809 , n299810 , n9383 , n299812 , n299813 , 
 n9386 , n299815 , n299816 , n9389 , n299818 , n299819 , n9392 , n299821 , n299822 , n9395 , 
 n299824 , n299825 , n299826 , n299827 , n9400 , n299829 , n9402 , n299831 , n299832 , n299833 , 
 n299834 , n9407 , n299836 , n299837 , n299838 , n9411 , n299840 , n299841 , n9414 , n299843 , 
 n299844 , n299845 , n299846 , n299847 , n9420 , n299849 , n299850 , n9423 , n299852 , n299853 , 
 n9426 , n299855 , n299856 , n9429 , n299858 , n299859 , n9432 , n299861 , n299862 , n9435 , 
 n9436 , n299865 , n299866 , n299867 , n299868 , n9441 , n299870 , n299871 , n299872 , n299873 , 
 n299874 , n299875 , n299876 , n299877 , n9450 , n299879 , n299880 , n9453 , n9454 , n299883 , 
 n9456 , n299885 , n299886 , n299887 , n299888 , n299889 , n299890 , n299891 , n299892 , n299893 , 
 n9466 , n9467 , n299896 , n299897 , n9470 , n299899 , n299900 , n299901 , n9474 , n9475 , 
 n9476 , n299905 , n9478 , n299907 , n299908 , n9481 , n299910 , n299911 , n299912 , n299913 , 
 n299914 , n9487 , n299916 , n299917 , n299918 , n299919 , n299920 , n299921 , n9494 , n9495 , 
 n299924 , n299925 , n299926 , n299927 , n9500 , n299929 , n299930 , n299931 , n9504 , n299933 , 
 n299934 , n299935 , n299936 , n9509 , n299938 , n9511 , n299940 , n299941 , n299942 , n299943 , 
 n299944 , n299945 , n9518 , n299947 , n299948 , n299949 , n9522 , n299951 , n299952 , n299953 , 
 n299954 , n9527 , n299956 , n9529 , n299958 , n299959 , n9532 , n9533 , n299962 , n299963 , 
 n9536 , n9537 , n299966 , n299967 , n9540 , n9541 , n299970 , n299971 , n299972 , n299973 , 
 n299974 , n299975 , n299976 , n299977 , n299978 , n299979 , n9552 , n299981 , n299982 , n299983 , 
 n299984 , n299985 , n299986 , n299987 , n299988 , n299989 , n299990 , n299991 , n299992 , n299993 , 
 n299994 , n299995 , n299996 , n9569 , n299998 , n299999 , n300000 , n300001 , n300002 , n300003 , 
 n300004 , n300005 , n300006 , n300007 , n300008 , n300009 , n300010 , n300011 , n300012 , n300013 , 
 n300014 , n9587 , n300016 , n300017 , n300018 , n300019 , n300020 , n300021 , n300022 , n300023 , 
 n300024 , n300025 , n9598 , n300027 , n300028 , n9601 , n300030 , n300031 , n300032 , n9605 , 
 n9606 , n9607 , n9608 , n9609 , n300038 , n9611 , n300040 , n9613 , n300042 , n300043 , 
 n300044 , n9617 , n300046 , n300047 , n300048 , n300049 , n300050 , n300051 , n300052 , n300053 , 
 n300054 , n300055 , n300056 , n9629 , n300058 , n9631 , n300060 , n300061 , n300062 , n300063 , 
 n300064 , n300065 , n9638 , n300067 , n300068 , n9641 , n9642 , n300071 , n300072 , n300073 , 
 n300074 , n300075 , n300076 , n300077 , n300078 , n300079 , n300080 , n300081 , n300082 , n300083 , 
 n300084 , n300085 , n300086 , n300087 , n9660 , n9661 , n300090 , n300091 , n300092 , n300093 , 
 n300094 , n300095 , n9668 , n9669 , n9670 , n300099 , n300100 , n300101 , n300102 , n300103 , 
 n300104 , n300105 , n300106 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , 
 n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n300123 , 
 n9696 , n300125 , n300126 , n9699 , n9700 , n300129 , n9702 , n300131 , n300132 , n9705 , 
 n300134 , n300135 , n300136 , n300137 , n300138 , n300139 , n300140 , n300141 , n300142 , n300143 , 
 n9716 , n300145 , n300146 , n9719 , n300148 , n9721 , n9722 , n300151 , n300152 , n300153 , 
 n300154 , n9727 , n9728 , n9729 , n300158 , n300159 , n9732 , n300161 , n300162 , n300163 , 
 n300164 , n300165 , n300166 , n300167 , n9740 , n300169 , n300170 , n300171 , n300172 , n300173 , 
 n300174 , n300175 , n300176 , n300177 , n300178 , n9751 , n9752 , n300181 , n9754 , n300183 , 
 n300184 , n300185 , n300186 , n300187 , n300188 , n9761 , n300190 , n300191 , n9764 , n300193 , 
 n300194 , n9767 , n300196 , n300197 , n9770 , n300199 , n300200 , n300201 , n300202 , n300203 , 
 n9776 , n300205 , n300206 , n300207 , n9780 , n300209 , n300210 , n300211 , n300212 , n9785 , 
 n9786 , n300215 , n300216 , n300217 , n300218 , n300219 , n9792 , n300221 , n9794 , n300223 , 
 n9796 , n9797 , n9798 , n9799 , n300228 , n300229 , n300230 , n9803 , n9804 , n300233 , 
 n9806 , n300235 , n300236 , n300237 , n300238 , n9811 , n300240 , n300241 , n9814 , n300243 , 
 n300244 , n9817 , n300246 , n300247 , n9820 , n300249 , n9822 , n300251 , n9824 , n9825 , 
 n300254 , n9827 , n300256 , n300257 , n300258 , n9831 , n300260 , n9833 , n300262 , n300263 , 
 n300264 , n300265 , n300266 , n300267 , n300268 , n300269 , n300270 , n300271 , n9844 , n300273 , 
 n9846 , n300275 , n9848 , n300277 , n300278 , n9851 , n300280 , n9853 , n300282 , n300283 , 
 n9856 , n300285 , n300286 , n9859 , n9860 , n300289 , n300290 , n9863 , n9864 , n9865 , 
 n9866 , n300295 , n300296 , n300297 , n300298 , n300299 , n300300 , n9873 , n300302 , n300303 , 
 n300304 , n300305 , n9878 , n9879 , n300308 , n300309 , n300310 , n300311 , n300312 , n9885 , 
 n300314 , n300315 , n300316 , n300317 , n300318 , n300319 , n9892 , n9893 , n9894 , n9895 , 
 n300324 , n9897 , n300326 , n300327 , n9900 , n300329 , n300330 , n9903 , n300332 , n300333 , 
 n9906 , n300335 , n300336 , n9909 , n9910 , n9911 , n300340 , n300341 , n300342 , n9915 , 
 n9916 , n300345 , n300346 , n300347 , n9920 , n300349 , n9922 , n9923 , n9924 , n300353 , 
 n9926 , n300355 , n300356 , n300357 , n300358 , n300359 , n300360 , n300361 , n300362 , n300363 , 
 n9936 , n300365 , n300366 , n9939 , n300368 , n300369 , n9942 , n9943 , n300372 , n300373 , 
 n300374 , n9947 , n300376 , n300377 , n9950 , n300379 , n9952 , n300381 , n300382 , n300383 , 
 n300384 , n300385 , n300386 , n300387 , n9960 , n9961 , n300390 , n9963 , n300392 , n300393 , 
 n300394 , n300395 , n300396 , n300397 , n9970 , n300399 , n300400 , n9973 , n300402 , n300403 , 
 n9976 , n300405 , n300406 , n300407 , n300408 , n300409 , n9982 , n300411 , n9984 , n300413 , 
 n9986 , n9987 , n9988 , n300417 , n300418 , n9991 , n9992 , n9993 , n300422 , n300423 , 
 n9996 , n300425 , n300426 , n9999 , n300428 , n300429 , n10002 , n300431 , n300432 , n10005 , 
 n300434 , n300435 , n10008 , n300437 , n300438 , n300439 , n300440 , n300441 , n10014 , n300443 , 
 n300444 , n300445 , n300446 , n300447 , n300448 , n10021 , n300450 , n300451 , n300452 , n300453 , 
 n300454 , n10027 , n10028 , n300457 , n300458 , n300459 , n10032 , n300461 , n300462 , n300463 , 
 n300464 , n300465 , n300466 , n10039 , n300468 , n300469 , n300470 , n10043 , n300472 , n300473 , 
 n300474 , n300475 , n300476 , n300477 , n300478 , n300479 , n300480 , n10053 , n300482 , n300483 , 
 n300484 , n300485 , n10058 , n300487 , n300488 , n10061 , n300490 , n300491 , n300492 , n300493 , 
 n300494 , n300495 , n300496 , n10069 , n300498 , n300499 , n300500 , n300501 , n300502 , n300503 , 
 n300504 , n300505 , n300506 , n300507 , n10080 , n300509 , n300510 , n300511 , n300512 , n300513 , 
 n300514 , n10087 , n300516 , n300517 , n10090 , n300519 , n10092 , n300521 , n300522 , n10095 , 
 n300524 , n300525 , n300526 , n300527 , n300528 , n300529 , n300530 , n300531 , n300532 , n300533 , 
 n300534 , n300535 , n300536 , n300537 , n300538 , n300539 , n300540 , n300541 , n10114 , n300543 , 
 n300544 , n300545 , n300546 , n10119 , n300548 , n10121 , n10122 , n10123 , n300552 , n10125 , 
 n300554 , n300555 , n300556 , n300557 , n300558 , n300559 , n300560 , n300561 , n300562 , n300563 , 
 n10136 , n300565 , n300566 , n300567 , n300568 , n300569 , n300570 , n300571 , n300572 , n300573 , 
 n300574 , n300575 , n300576 , n300577 , n300578 , n10151 , n300580 , n300581 , n300582 , n300583 , 
 n10156 , n300585 , n300586 , n10159 , n300588 , n300589 , n300590 , n300591 , n10164 , n300593 , 
 n10166 , n10167 , n300596 , n300597 , n300598 , n300599 , n300600 , n300601 , n300602 , n300603 , 
 n300604 , n300605 , n300606 , n300607 , n300608 , n300609 , n10182 , n300611 , n300612 , n10185 , 
 n300614 , n300615 , n10188 , n10189 , n300618 , n300619 , n300620 , n300621 , n300622 , n300623 , 
 n300624 , n10197 , n300626 , n10199 , n10200 , n300629 , n300630 , n10203 , n300632 , n300633 , 
 n10206 , n10207 , n300636 , n300637 , n300638 , n300639 , n300640 , n300641 , n300642 , n300643 , 
 n10216 , n300645 , n10218 , n10219 , n300648 , n300649 , n10222 , n300651 , n300652 , n300653 , 
 n300654 , n300655 , n300656 , n300657 , n300658 , n10231 , n300660 , n300661 , n300662 , n300663 , 
 n300664 , n10237 , n10238 , n10239 , n300668 , n10241 , n300670 , n300671 , n300672 , n10245 , 
 n300674 , n300675 , n10248 , n300677 , n300678 , n10251 , n300680 , n300681 , n300682 , n300683 , 
 n300684 , n300685 , n300686 , n300687 , n10260 , n300689 , n300690 , n300691 , n300692 , n300693 , 
 n300694 , n300695 , n300696 , n300697 , n300698 , n300699 , n300700 , n300701 , n10274 , n300703 , 
 n300704 , n300705 , n300706 , n300707 , n300708 , n300709 , n300710 , n300711 , n300712 , n300713 , 
 n300714 , n10287 , n10288 , n300717 , n10290 , n300719 , n300720 , n300721 , n300722 , n300723 , 
 n300724 , n300725 , n300726 , n10299 , n10300 , n300729 , n10302 , n10303 , n300732 , n10305 , 
 n10306 , n300735 , n300736 , n300737 , n300738 , n300739 , n300740 , n10313 , n300742 , n300743 , 
 n300744 , n300745 , n10318 , n300747 , n300748 , n10321 , n300750 , n300751 , n10324 , n300753 , 
 n300754 , n10327 , n300756 , n300757 , n300758 , n10331 , n300760 , n300761 , n10334 , n300763 , 
 n300764 , n300765 , n10338 , n300767 , n300768 , n300769 , n300770 , n300771 , n300772 , n300773 , 
 n300774 , n300775 , n300776 , n300777 , n10350 , n300779 , n300780 , n10353 , n300782 , n10355 , 
 n10356 , n300785 , n10358 , n300787 , n300788 , n10361 , n10362 , n300791 , n10364 , n300793 , 
 n10366 , n300795 , n10368 , n300797 , n300798 , n10371 , n300800 , n300801 , n300802 , n300803 , 
 n300804 , n300805 , n300806 , n300807 , n300808 , n300809 , n300810 , n300811 , n300812 , n300813 , 
 n10386 , n300815 , n10388 , n10389 , n300818 , n300819 , n10392 , n300821 , n300822 , n10395 , 
 n300824 , n10397 , n300826 , n300827 , n10400 , n300829 , n300830 , n10403 , n300832 , n10405 , 
 n10406 , n10407 , n10408 , n300837 , n300838 , n300839 , n300840 , n10413 , n300842 , n300843 , 
 n10416 , n300845 , n300846 , n300847 , n300848 , n300849 , n300850 , n300851 , n300852 , n300853 , 
 n300854 , n300855 , n300856 , n10429 , n300858 , n300859 , n300860 , n10433 , n10434 , n300863 , 
 n10436 , n300865 , n300866 , n10439 , n300868 , n10441 , n300870 , n300871 , n300872 , n300873 , 
 n300874 , n300875 , n300876 , n10449 , n300878 , n300879 , n10452 , n300881 , n10454 , n300883 , 
 n300884 , n300885 , n300886 , n300887 , n300888 , n300889 , n300890 , n300891 , n300892 , n300893 , 
 n300894 , n300895 , n10468 , n300897 , n300898 , n300899 , n300900 , n300901 , n300902 , n300903 , 
 n300904 , n300905 , n300906 , n300907 , n300908 , n10481 , n300910 , n300911 , n300912 , n300913 , 
 n10486 , n300915 , n300916 , n10489 , n300918 , n300919 , n10492 , n300921 , n300922 , n10495 , 
 n300924 , n300925 , n10498 , n300927 , n300928 , n300929 , n300930 , n300931 , n300932 , n300933 , 
 n300934 , n300935 , n300936 , n300937 , n300938 , n10511 , n300940 , n300941 , n300942 , n300943 , 
 n300944 , n300945 , n300946 , n300947 , n300948 , n300949 , n300950 , n300951 , n10524 , n300953 , 
 n10526 , n300955 , n300956 , n10529 , n300958 , n300959 , n300960 , n300961 , n10534 , n300963 , 
 n300964 , n300965 , n300966 , n300967 , n300968 , n300969 , n300970 , n300971 , n300972 , n300973 , 
 n300974 , n300975 , n10548 , n300977 , n300978 , n300979 , n300980 , n300981 , n300982 , n300983 , 
 n300984 , n300985 , n300986 , n300987 , n300988 , n300989 , n300990 , n300991 , n300992 , n300993 , 
 n300994 , n300995 , n300996 , n300997 , n300998 , n300999 , n10572 , n301001 , n301002 , n10575 , 
 n301004 , n301005 , n301006 , n301007 , n10580 , n301009 , n301010 , n301011 , n301012 , n301013 , 
 n301014 , n301015 , n10588 , n10589 , n301018 , n301019 , n301020 , n301021 , n301022 , n301023 , 
 n301024 , n301025 , n301026 , n10599 , n301028 , n301029 , n10602 , n301031 , n301032 , n10605 , 
 n10606 , n301035 , n301036 , n301037 , n301038 , n10611 , n10612 , n301041 , n10614 , n10615 , 
 n301044 , n301045 , n301046 , n301047 , n10620 , n10621 , n301050 , n301051 , n301052 , n301053 , 
 n10626 , n301055 , n10628 , n301057 , n301058 , n10631 , n301060 , n301061 , n301062 , n301063 , 
 n301064 , n10637 , n301066 , n301067 , n10640 , n301069 , n301070 , n10643 , n301072 , n301073 , 
 n301074 , n301075 , n301076 , n301077 , n301078 , n301079 , n301080 , n301081 , n10654 , n301083 , 
 n301084 , n301085 , n301086 , n301087 , n301088 , n301089 , n301090 , n301091 , n301092 , n301093 , 
 n301094 , n10667 , n10668 , n301097 , n301098 , n10671 , n10672 , n301101 , n301102 , n301103 , 
 n301104 , n10677 , n301106 , n301107 , n301108 , n301109 , n301110 , n301111 , n301112 , n301113 , 
 n301114 , n10687 , n301116 , n10689 , n301118 , n301119 , n10692 , n301121 , n301122 , n10695 , 
 n301124 , n301125 , n10698 , n301127 , n301128 , n301129 , n301130 , n301131 , n301132 , n301133 , 
 n301134 , n301135 , n301136 , n301137 , n10710 , n301139 , n301140 , n301141 , n301142 , n10715 , 
 n301144 , n301145 , n301146 , n301147 , n10720 , n301149 , n301150 , n10723 , n301152 , n301153 , 
 n301154 , n301155 , n301156 , n301157 , n301158 , n301159 , n301160 , n10733 , n301162 , n301163 , 
 n301164 , n301165 , n301166 , n301167 , n301168 , n301169 , n301170 , n301171 , n301172 , n301173 , 
 n301174 , n301175 , n301176 , n301177 , n301178 , n10751 , n301180 , n10753 , n10754 , n10755 , 
 n10756 , n10757 , n10758 , n10759 , n10760 , n301189 , n301190 , n10763 , n301192 , n301193 , 
 n10766 , n301195 , n301196 , n10769 , n301198 , n301199 , n301200 , n301201 , n301202 , n301203 , 
 n10776 , n301205 , n301206 , n301207 , n10780 , n10781 , n301210 , n301211 , n10784 , n301213 , 
 n301214 , n301215 , n301216 , n301217 , n301218 , n301219 , n301220 , n301221 , n301222 , n10795 , 
 n301224 , n301225 , n301226 , n301227 , n301228 , n301229 , n10802 , n301231 , n10804 , n301233 , 
 n10806 , n301235 , n10808 , n10809 , n301238 , n301239 , n301240 , n301241 , n301242 , n301243 , 
 n301244 , n301245 , n301246 , n301247 , n301248 , n301249 , n301250 , n301251 , n10824 , n301253 , 
 n10826 , n301255 , n10828 , n301257 , n301258 , n10831 , n301260 , n10833 , n10834 , n301263 , 
 n301264 , n301265 , n301266 , n301267 , n10840 , n301269 , n301270 , n10843 , n301272 , n301273 , 
 n10846 , n301275 , n301276 , n301277 , n10850 , n301279 , n301280 , n10853 , n301282 , n10855 , 
 n10856 , n301285 , n10858 , n301287 , n10860 , n301289 , n301290 , n301291 , n301292 , n301293 , 
 n301294 , n301295 , n301296 , n301297 , n301298 , n301299 , n301300 , n10873 , n301302 , n301303 , 
 n301304 , n10877 , n301306 , n301307 , n10880 , n301309 , n301310 , n301311 , n301312 , n301313 , 
 n301314 , n301315 , n301316 , n301317 , n301318 , n301319 , n10892 , n301321 , n301322 , n10895 , 
 n10896 , n301325 , n10898 , n301327 , n301328 , n10901 , n301330 , n301331 , n301332 , n301333 , 
 n301334 , n301335 , n301336 , n301337 , n301338 , n10911 , n301340 , n301341 , n301342 , n301343 , 
 n301344 , n301345 , n301346 , n301347 , n301348 , n301349 , n301350 , n10923 , n10924 , n10925 , 
 n10926 , n301355 , n10928 , n10929 , n10930 , n301359 , n10932 , n10933 , n301362 , n10935 , 
 n301364 , n301365 , n301366 , n301367 , n301368 , n301369 , n301370 , n10943 , n301372 , n301373 , 
 n301374 , n301375 , n301376 , n301377 , n301378 , n301379 , n301380 , n301381 , n301382 , n10955 , 
 n301384 , n10957 , n10958 , n301387 , n301388 , n301389 , n301390 , n10963 , n301392 , n301393 , 
 n301394 , n301395 , n301396 , n301397 , n301398 , n10971 , n301400 , n301401 , n10974 , n10975 , 
 n301404 , n10977 , n301406 , n10979 , n301408 , n301409 , n301410 , n301411 , n301412 , n301413 , 
 n10986 , n10987 , n301416 , n301417 , n301418 , n301419 , n301420 , n301421 , n301422 , n301423 , 
 n301424 , n10997 , n301426 , n10999 , n11000 , n11001 , n301430 , n11003 , n301432 , n11005 , 
 n301434 , n301435 , n11008 , n301437 , n301438 , n301439 , n301440 , n11013 , n301442 , n301443 , 
 n301444 , n301445 , n301446 , n301447 , n301448 , n301449 , n301450 , n301451 , n301452 , n301453 , 
 n301454 , n301455 , n11028 , n301457 , n301458 , n301459 , n301460 , n301461 , n301462 , n11035 , 
 n301464 , n11037 , n11038 , n301467 , n11040 , n301469 , n301470 , n301471 , n301472 , n301473 , 
 n301474 , n301475 , n301476 , n11049 , n301478 , n301479 , n11052 , n301481 , n301482 , n11055 , 
 n301484 , n301485 , n301486 , n301487 , n11060 , n301489 , n301490 , n301491 , n301492 , n11065 , 
 n301494 , n301495 , n301496 , n301497 , n301498 , n11071 , n301500 , n301501 , n11074 , n301503 , 
 n301504 , n301505 , n301506 , n301507 , n301508 , n11081 , n11082 , n301511 , n301512 , n301513 , 
 n301514 , n11087 , n301516 , n11089 , n11090 , n11091 , n11092 , n301521 , n11094 , n11095 , 
 n301524 , n11097 , n301526 , n301527 , n301528 , n11101 , n11102 , n301531 , n301532 , n11105 , 
 n301534 , n301535 , n301536 , n301537 , n301538 , n11111 , n301540 , n11113 , n301542 , n301543 , 
 n301544 , n301545 , n11118 , n301547 , n301548 , n11121 , n301550 , n301551 , n11124 , n301553 , 
 n301554 , n301555 , n11128 , n301557 , n301558 , n301559 , n11132 , n301561 , n301562 , n301563 , 
 n301564 , n301565 , n301566 , n11139 , n301568 , n301569 , n301570 , n301571 , n11144 , n11145 , 
 n11146 , n11147 , n11148 , n11149 , n301578 , n301579 , n301580 , n301581 , n301582 , n301583 , 
 n301584 , n301585 , n11158 , n301587 , n301588 , n301589 , n11162 , n11163 , n301592 , n301593 , 
 n301594 , n11167 , n301596 , n301597 , n301598 , n301599 , n11172 , n11173 , n301602 , n301603 , 
 n301604 , n11177 , n301606 , n301607 , n301608 , n301609 , n301610 , n301611 , n301612 , n11185 , 
 n301614 , n11187 , n11188 , n301617 , n301618 , n11191 , n301620 , n11193 , n11194 , n11195 , 
 n301624 , n301625 , n11198 , n301627 , n301628 , n11201 , n301630 , n301631 , n301632 , n301633 , 
 n301634 , n11207 , n11208 , n301637 , n11210 , n301639 , n11212 , n301641 , n301642 , n11215 , 
 n301644 , n301645 , n11218 , n301647 , n11220 , n301649 , n301650 , n11223 , n301652 , n301653 , 
 n301654 , n301655 , n301656 , n301657 , n301658 , n301659 , n301660 , n301661 , n301662 , n301663 , 
 n301664 , n301665 , n301666 , n301667 , n301668 , n301669 , n301670 , n301671 , n11244 , n301673 , 
 n301674 , n11247 , n11248 , n301677 , n11250 , n301679 , n301680 , n11253 , n301682 , n301683 , 
 n301684 , n11257 , n301686 , n301687 , n11260 , n301689 , n301690 , n11263 , n11264 , n301693 , 
 n11266 , n301695 , n11268 , n301697 , n301698 , n301699 , n11272 , n301701 , n301702 , n301703 , 
 n301704 , n301705 , n11278 , n301707 , n301708 , n11281 , n301710 , n301711 , n11284 , n11285 , 
 n11286 , n301715 , n11288 , n301717 , n301718 , n11291 , n11292 , n11293 , n301722 , n301723 , 
 n11296 , n11297 , n301726 , n11299 , n301728 , n301729 , n301730 , n301731 , n301732 , n11305 , 
 n301734 , n11307 , n11308 , n301737 , n301738 , n301739 , n301740 , n301741 , n11314 , n301743 , 
 n301744 , n301745 , n301746 , n11319 , n301748 , n301749 , n11322 , n301751 , n301752 , n11325 , 
 n11326 , n301755 , n301756 , n301757 , n301758 , n11331 , n301760 , n301761 , n301762 , n301763 , 
 n301764 , n301765 , n301766 , n301767 , n301768 , n301769 , n11342 , n11343 , n301772 , n11345 , 
 n301774 , n11347 , n11348 , n301777 , n301778 , n301779 , n301780 , n301781 , n301782 , n301783 , 
 n301784 , n301785 , n11358 , n301787 , n11360 , n301789 , n301790 , n11363 , n301792 , n301793 , 
 n11366 , n301795 , n301796 , n301797 , n301798 , n301799 , n301800 , n11373 , n301802 , n301803 , 
 n11376 , n301805 , n301806 , n301807 , n301808 , n301809 , n301810 , n11383 , n11384 , n301813 , 
 n301814 , n301815 , n11388 , n301817 , n301818 , n11391 , n301820 , n301821 , n301822 , n301823 , 
 n301824 , n301825 , n301826 , n301827 , n301828 , n301829 , n11402 , n301831 , n301832 , n301833 , 
 n301834 , n301835 , n301836 , n301837 , n301838 , n301839 , n301840 , n11413 , n301842 , n301843 , 
 n301844 , n301845 , n301846 , n301847 , n301848 , n301849 , n301850 , n11423 , n11424 , n11425 , 
 n11426 , n11427 , n11428 , n301857 , n301858 , n301859 , n301860 , n301861 , n301862 , n301863 , 
 n301864 , n301865 , n301866 , n301867 , n301868 , n11441 , n301870 , n11443 , n301872 , n301873 , 
 n301874 , n301875 , n11448 , n301877 , n301878 , n301879 , n301880 , n301881 , n11454 , n301883 , 
 n301884 , n301885 , n301886 , n11459 , n301888 , n11461 , n11462 , n301891 , n11464 , n11465 , 
 n11466 , n11467 , n301896 , n11469 , n301898 , n301899 , n11472 , n301901 , n301902 , n11475 , 
 n301904 , n301905 , n11478 , n301907 , n301908 , n301909 , n301910 , n301911 , n301912 , n11485 , 
 n301914 , n301915 , n301916 , n11489 , n301918 , n301919 , n301920 , n11493 , n301922 , n301923 , 
 n11496 , n11497 , n11498 , n301927 , n301928 , n11501 , n11502 , n301931 , n301932 , n11505 , 
 n11506 , n11507 , n301936 , n301937 , n11510 , n301939 , n301940 , n301941 , n301942 , n301943 , 
 n11516 , n301945 , n301946 , n11519 , n11520 , n11521 , n301950 , n11523 , n11524 , n11525 , 
 n301954 , n301955 , n301956 , n11529 , n301958 , n301959 , n11532 , n301961 , n301962 , n301963 , 
 n11536 , n301965 , n301966 , n301967 , n301968 , n301969 , n301970 , n301971 , n301972 , n301973 , 
 n11546 , n301975 , n301976 , n11549 , n301978 , n301979 , n11552 , n301981 , n301982 , n301983 , 
 n301984 , n301985 , n301986 , n301987 , n301988 , n301989 , n11562 , n301991 , n301992 , n301993 , 
 n301994 , n301995 , n301996 , n301997 , n301998 , n11571 , n302000 , n302001 , n11574 , n302003 , 
 n11576 , n302005 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n302012 , n11585 , 
 n302014 , n302015 , n11588 , n302017 , n302018 , n302019 , n302020 , n302021 , n11594 , n302023 , 
 n11596 , n302025 , n302026 , n302027 , n302028 , n302029 , n302030 , n302031 , n302032 , n302033 , 
 n302034 , n11607 , n11608 , n302037 , n11610 , n11611 , n302040 , n302041 , n302042 , n302043 , 
 n302044 , n11617 , n11618 , n11619 , n11620 , n302049 , n11622 , n302051 , n302052 , n302053 , 
 n302054 , n302055 , n11628 , n302057 , n302058 , n302059 , n302060 , n302061 , n302062 , n302063 , 
 n302064 , n302065 , n302066 , n302067 , n11640 , n302069 , n11642 , n302071 , n302072 , n302073 , 
 n302074 , n302075 , n302076 , n11649 , n11650 , n11651 , n302080 , n302081 , n302082 , n302083 , 
 n11656 , n302085 , n302086 , n302087 , n302088 , n11661 , n302090 , n302091 , n302092 , n302093 , 
 n302094 , n11667 , n302096 , n302097 , n11670 , n302099 , n11672 , n302101 , n302102 , n302103 , 
 n11676 , n11677 , n302106 , n302107 , n11680 , n302109 , n302110 , n302111 , n302112 , n11685 , 
 n11686 , n11687 , n302116 , n302117 , n302118 , n11691 , n11692 , n302121 , n302122 , n302123 , 
 n302124 , n302125 , n11698 , n302127 , n302128 , n302129 , n302130 , n11703 , n302132 , n302133 , 
 n302134 , n11707 , n11708 , n302137 , n11710 , n302139 , n302140 , n302141 , n302142 , n11715 , 
 n302144 , n302145 , n302146 , n11719 , n302148 , n302149 , n11722 , n302151 , n302152 , n302153 , 
 n302154 , n302155 , n302156 , n302157 , n302158 , n302159 , n302160 , n11733 , n302162 , n302163 , 
 n11736 , n302165 , n302166 , n11739 , n302168 , n302169 , n302170 , n302171 , n302172 , n302173 , 
 n302174 , n11747 , n302176 , n302177 , n11750 , n302179 , n302180 , n302181 , n302182 , n302183 , 
 n302184 , n302185 , n11758 , n302187 , n302188 , n11761 , n11762 , n302191 , n302192 , n302193 , 
 n11766 , n302195 , n302196 , n302197 , n302198 , n11771 , n302200 , n11773 , n11774 , n302203 , 
 n302204 , n11777 , n11778 , n302207 , n302208 , n11781 , n302210 , n11783 , n302212 , n11785 , 
 n302214 , n302215 , n302216 , n11789 , n11790 , n11791 , n302220 , n302221 , n302222 , n11795 , 
 n302224 , n302225 , n302226 , n302227 , n302228 , n302229 , n302230 , n302231 , n302232 , n302233 , 
 n11806 , n302235 , n302236 , n302237 , n302238 , n11811 , n302240 , n302241 , n302242 , n302243 , 
 n302244 , n302245 , n302246 , n302247 , n302248 , n11821 , n302250 , n302251 , n302252 , n302253 , 
 n11826 , n302255 , n302256 , n302257 , n302258 , n302259 , n302260 , n302261 , n302262 , n302263 , 
 n11836 , n302265 , n11838 , n11839 , n302268 , n11841 , n302270 , n11843 , n302272 , n302273 , 
 n302274 , n302275 , n11848 , n302277 , n302278 , n302279 , n11852 , n302281 , n302282 , n11855 , 
 n302284 , n11857 , n302286 , n11859 , n302288 , n11861 , n302290 , n302291 , n302292 , n302293 , 
 n11866 , n302295 , n302296 , n302297 , n302298 , n302299 , n302300 , n302301 , n302302 , n11875 , 
 n11876 , n11877 , n11878 , n11879 , n11880 , n302309 , n302310 , n302311 , n302312 , n302313 , 
 n302314 , n11887 , n302316 , n302317 , n302318 , n302319 , n302320 , n302321 , n302322 , n302323 , 
 n302324 , n302325 , n302326 , n302327 , n302328 , n302329 , n302330 , n302331 , n302332 , n302333 , 
 n302334 , n302335 , n302336 , n11909 , n11910 , n302339 , n302340 , n302341 , n302342 , n302343 , 
 n11916 , n302345 , n302346 , n302347 , n302348 , n302349 , n302350 , n302351 , n302352 , n11925 , 
 n302354 , n302355 , n11928 , n302357 , n302358 , n11931 , n302360 , n302361 , n11934 , n302363 , 
 n302364 , n302365 , n11938 , n302367 , n302368 , n11941 , n302370 , n302371 , n302372 , n11945 , 
 n302374 , n302375 , n11948 , n302377 , n302378 , n11951 , n302380 , n302381 , n302382 , n302383 , 
 n11956 , n302385 , n302386 , n11959 , n302388 , n11961 , n302390 , n302391 , n11964 , n302393 , 
 n302394 , n302395 , n11968 , n302397 , n302398 , n302399 , n11972 , n302401 , n302402 , n302403 , 
 n302404 , n302405 , n302406 , n302407 , n11980 , n302409 , n302410 , n11983 , n302412 , n302413 , 
 n11986 , n302415 , n302416 , n302417 , n302418 , n302419 , n302420 , n302421 , n302422 , n302423 , 
 n11996 , n11997 , n302426 , n302427 , n12000 , n302429 , n302430 , n302431 , n302432 , n302433 , 
 n12006 , n302435 , n302436 , n12009 , n302438 , n302439 , n12012 , n302441 , n302442 , n12015 , 
 n302444 , n302445 , n302446 , n302447 , n302448 , n12021 , n302450 , n302451 , n302452 , n12025 , 
 n302454 , n302455 , n302456 , n302457 , n302458 , n302459 , n302460 , n302461 , n302462 , n12035 , 
 n302464 , n302465 , n302466 , n302467 , n302468 , n302469 , n302470 , n302471 , n302472 , n302473 , 
 n302474 , n12047 , n302476 , n302477 , n12050 , n302479 , n302480 , n302481 , n302482 , n302483 , 
 n12056 , n302485 , n12058 , n302487 , n302488 , n302489 , n12062 , n302491 , n302492 , n302493 , 
 n302494 , n302495 , n302496 , n302497 , n302498 , n302499 , n302500 , n12073 , n12074 , n302503 , 
 n302504 , n302505 , n12078 , n302507 , n302508 , n302509 , n12082 , n302511 , n12084 , n302513 , 
 n302514 , n302515 , n12088 , n302517 , n302518 , n12091 , n302520 , n302521 , n12094 , n12095 , 
 n302524 , n302525 , n12098 , n302527 , n302528 , n302529 , n12102 , n12103 , n12104 , n12105 , 
 n12106 , n12107 , n12108 , n302537 , n12110 , n302539 , n302540 , n302541 , n302542 , n302543 , 
 n12116 , n302545 , n302546 , n302547 , n302548 , n302549 , n302550 , n302551 , n302552 , n12125 , 
 n12126 , n12127 , n12128 , n302557 , n12130 , n302559 , n302560 , n12133 , n302562 , n302563 , 
 n12136 , n302565 , n12138 , n302567 , n302568 , n302569 , n302570 , n302571 , n302572 , n12145 , 
 n12146 , n12147 , n302576 , n302577 , n302578 , n302579 , n12152 , n302581 , n302582 , n302583 , 
 n12156 , n302585 , n302586 , n302587 , n12160 , n302589 , n302590 , n302591 , n302592 , n302593 , 
 n12166 , n302595 , n12168 , n302597 , n12170 , n12171 , n12172 , n302601 , n302602 , n302603 , 
 n302604 , n302605 , n12178 , n12179 , n302608 , n302609 , n12182 , n12183 , n302612 , n302613 , 
 n12186 , n12187 , n302616 , n302617 , n12190 , n302619 , n302620 , n302621 , n12194 , n302623 , 
 n302624 , n12197 , n302626 , n12199 , n302628 , n12201 , n302630 , n302631 , n302632 , n302633 , 
 n12206 , n302635 , n302636 , n302637 , n12210 , n302639 , n302640 , n302641 , n12214 , n302643 , 
 n12216 , n302645 , n12218 , n12219 , n302648 , n302649 , n12222 , n302651 , n302652 , n302653 , 
 n302654 , n302655 , n302656 , n302657 , n302658 , n302659 , n302660 , n302661 , n12234 , n302663 , 
 n302664 , n302665 , n12238 , n302667 , n302668 , n302669 , n302670 , n302671 , n302672 , n12245 , 
 n302674 , n302675 , n12248 , n302677 , n12250 , n302679 , n12252 , n302681 , n12254 , n12255 , 
 n12256 , n302685 , n302686 , n302687 , n12260 , n302689 , n302690 , n302691 , n12264 , n302693 , 
 n302694 , n302695 , n302696 , n302697 , n302698 , n302699 , n302700 , n302701 , n302702 , n302703 , 
 n302704 , n302705 , n302706 , n302707 , n302708 , n12281 , n302710 , n302711 , n302712 , n302713 , 
 n302714 , n302715 , n302716 , n302717 , n302718 , n302719 , n12292 , n302721 , n302722 , n12295 , 
 n302724 , n302725 , n302726 , n302727 , n12300 , n12301 , n12302 , n302731 , n302732 , n302733 , 
 n12306 , n302735 , n302736 , n302737 , n302738 , n12311 , n302740 , n302741 , n302742 , n302743 , 
 n302744 , n12317 , n302746 , n302747 , n12320 , n302749 , n302750 , n302751 , n302752 , n12325 , 
 n302754 , n302755 , n302756 , n12329 , n302758 , n302759 , n12332 , n302761 , n302762 , n302763 , 
 n12336 , n302765 , n302766 , n12339 , n12340 , n302769 , n302770 , n302771 , n12344 , n302773 , 
 n302774 , n302775 , n302776 , n302777 , n12350 , n12351 , n12352 , n302781 , n302782 , n12355 , 
 n12356 , n12357 , n302786 , n12359 , n302788 , n302789 , n302790 , n302791 , n302792 , n302793 , 
 n12366 , n302795 , n12368 , n302797 , n302798 , n302799 , n302800 , n302801 , n302802 , n302803 , 
 n302804 , n302805 , n12378 , n302807 , n302808 , n302809 , n302810 , n302811 , n302812 , n302813 , 
 n302814 , n302815 , n12388 , n302817 , n12390 , n12391 , n302820 , n302821 , n302822 , n302823 , 
 n302824 , n302825 , n302826 , n302827 , n302828 , n302829 , n302830 , n302831 , n12404 , n302833 , 
 n302834 , n302835 , n12408 , n12409 , n302838 , n12411 , n302840 , n302841 , n12414 , n302843 , 
 n12416 , n302845 , n302846 , n12419 , n302848 , n302849 , n302850 , n12423 , n12424 , n302853 , 
 n302854 , n302855 , n302856 , n302857 , n12430 , n302859 , n302860 , n302861 , n302862 , n12435 , 
 n302864 , n302865 , n302866 , n12439 , n302868 , n302869 , n12442 , n302871 , n302872 , n302873 , 
 n302874 , n302875 , n12448 , n302877 , n12450 , n12451 , n302880 , n302881 , n302882 , n302883 , 
 n302884 , n302885 , n302886 , n302887 , n302888 , n302889 , n302890 , n12463 , n302892 , n12465 , 
 n302894 , n302895 , n12468 , n12469 , n302898 , n302899 , n302900 , n12473 , n302902 , n12475 , 
 n12476 , n302905 , n302906 , n302907 , n12480 , n302909 , n302910 , n12483 , n302912 , n12485 , 
 n302914 , n302915 , n302916 , n302917 , n12490 , n302919 , n302920 , n12493 , n302922 , n12495 , 
 n302924 , n12497 , n302926 , n12499 , n12500 , n302929 , n302930 , n302931 , n302932 , n302933 , 
 n302934 , n302935 , n302936 , n302937 , n12510 , n302939 , n302940 , n302941 , n12514 , n12515 , 
 n12516 , n302945 , n302946 , n302947 , n12520 , n302949 , n302950 , n302951 , n302952 , n12525 , 
 n12526 , n302955 , n302956 , n302957 , n302958 , n302959 , n302960 , n302961 , n302962 , n302963 , 
 n12536 , n302965 , n302966 , n12539 , n302968 , n12541 , n302970 , n302971 , n302972 , n302973 , 
 n12546 , n302975 , n302976 , n302977 , n302978 , n12551 , n302980 , n302981 , n302982 , n302983 , 
 n302984 , n302985 , n12558 , n302987 , n302988 , n12561 , n12562 , n12563 , n12564 , n302993 , 
 n302994 , n12567 , n12568 , n12569 , n302998 , n12571 , n12572 , n12573 , n303002 , n303003 , 
 n12576 , n12577 , n12578 , n303007 , n303008 , n303009 , n303010 , n303011 , n12584 , n303013 , 
 n303014 , n12587 , n12588 , n303017 , n303018 , n303019 , n303020 , n12593 , n12594 , n12595 , 
 n12596 , n12597 , n12598 , n303027 , n303028 , n12601 , n12602 , n303031 , n12604 , n303033 , 
 n303034 , n303035 , n12608 , n12609 , n12610 , n303039 , n12612 , n303041 , n303042 , n12615 , 
 n12616 , n12617 , n12618 , n303047 , n303048 , n12621 , n303050 , n12623 , n303052 , n303053 , 
 n303054 , n303055 , n303056 , n303057 , n303058 , n12631 , n303060 , n12633 , n303062 , n12635 , 
 n12636 , n303065 , n12638 , n303067 , n12640 , n303069 , n303070 , n303071 , n12644 , n303073 , 
 n303074 , n303075 , n12648 , n12649 , n12650 , n303079 , n12652 , n303081 , n12654 , n303083 , 
 n303084 , n303085 , n303086 , n12659 , n303088 , n303089 , n12662 , n303091 , n303092 , n303093 , 
 n303094 , n12667 , n303096 , n303097 , n12670 , n303099 , n12672 , n303101 , n303102 , n12675 , 
 n303104 , n303105 , n303106 , n303107 , n303108 , n303109 , n12682 , n303111 , n303112 , n12685 , 
 n303114 , n303115 , n303116 , n12689 , n303118 , n12691 , n12692 , n303121 , n303122 , n12695 , 
 n303124 , n12697 , n12698 , n12699 , n303128 , n303129 , n12702 , n12703 , n303132 , n303133 , 
 n12706 , n303135 , n303136 , n12709 , n303138 , n12711 , n12712 , n303141 , n12714 , n303143 , 
 n12716 , n12717 , n303146 , n303147 , n303148 , n303149 , n303150 , n12723 , n12724 , n303153 , 
 n12726 , n303155 , n303156 , n303157 , n12730 , n12731 , n12732 , n12733 , n303162 , n303163 , 
 n303164 , n303165 , n12738 , n303167 , n303168 , n303169 , n12742 , n303171 , n12744 , n303173 , 
 n303174 , n303175 , n12748 , n12749 , n303178 , n303179 , n12752 , n303181 , n303182 , n12755 , 
 n12756 , n12757 , n12758 , n303187 , n303188 , n303189 , n303190 , n12763 , n303192 , n303193 , 
 n303194 , n303195 , n12768 , n303197 , n12770 , n303199 , n303200 , n12773 , n303202 , n303203 , 
 n303204 , n303205 , n12778 , n12779 , n303208 , n12781 , n12782 , n12783 , n12784 , n12785 , 
 n12786 , n303215 , n303216 , n303217 , n303218 , n303219 , n303220 , n303221 , n303222 , n303223 , 
 n303224 , n303225 , n12798 , n303227 , n303228 , n303229 , n303230 , n303231 , n303232 , n303233 , 
 n303234 , n303235 , n12808 , n303237 , n303238 , n12811 , n303240 , n303241 , n12814 , n303243 , 
 n303244 , n12817 , n303246 , n303247 , n303248 , n303249 , n303250 , n303251 , n303252 , n303253 , 
 n303254 , n303255 , n12828 , n303257 , n303258 , n12831 , n303260 , n303261 , n12834 , n303263 , 
 n303264 , n12837 , n12838 , n12839 , n303268 , n303269 , n12842 , n303271 , n303272 , n12845 , 
 n303274 , n303275 , n12848 , n303277 , n303278 , n303279 , n303280 , n303281 , n303282 , n303283 , 
 n303284 , n303285 , n303286 , n303287 , n303288 , n12861 , n303290 , n303291 , n12864 , n303293 , 
 n303294 , n303295 , n303296 , n303297 , n303298 , n12871 , n303300 , n303301 , n303302 , n303303 , 
 n303304 , n303305 , n303306 , n303307 , n303308 , n303309 , n303310 , n303311 , n303312 , n303313 , 
 n12886 , n12887 , n303316 , n303317 , n303318 , n303319 , n303320 , n303321 , n303322 , n303323 , 
 n12896 , n12897 , n303326 , n12899 , n303328 , n303329 , n303330 , n303331 , n303332 , n303333 , 
 n303334 , n303335 , n303336 , n303337 , n303338 , n303339 , n303340 , n303341 , n303342 , n303343 , 
 n303344 , n303345 , n12918 , n303347 , n12920 , n303349 , n12922 , n303351 , n303352 , n12925 , 
 n303354 , n303355 , n12928 , n12929 , n303358 , n12931 , n303360 , n303361 , n303362 , n303363 , 
 n303364 , n12937 , n12938 , n12939 , n12940 , n303369 , n12942 , n303371 , n12944 , n303373 , 
 n303374 , n303375 , n303376 , n303377 , n303378 , n303379 , n303380 , n303381 , n303382 , n303383 , 
 n303384 , n303385 , n12958 , n303387 , n12960 , n303389 , n303390 , n12963 , n303392 , n303393 , 
 n12966 , n303395 , n303396 , n12969 , n303398 , n303399 , n12972 , n303401 , n303402 , n12975 , 
 n303404 , n303405 , n303406 , n303407 , n12980 , n303409 , n12982 , n12983 , n303412 , n303413 , 
 n303414 , n303415 , n12988 , n12989 , n12990 , n303419 , n12992 , n303421 , n12994 , n303423 , 
 n303424 , n303425 , n303426 , n12999 , n303428 , n303429 , n13002 , n303431 , n303432 , n303433 , 
 n303434 , n303435 , n303436 , n303437 , n303438 , n303439 , n303440 , n303441 , n303442 , n303443 , 
 n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n303450 , n13023 , n303452 , n13025 , 
 n303454 , n303455 , n303456 , n303457 , n13030 , n303459 , n303460 , n13033 , n13034 , n303463 , 
 n303464 , n303465 , n13038 , n13039 , n303468 , n303469 , n303470 , n13043 , n303472 , n303473 , 
 n303474 , n303475 , n303476 , n303477 , n13050 , n303479 , n303480 , n303481 , n13054 , n303483 , 
 n303484 , n303485 , n303486 , n13059 , n303488 , n303489 , n303490 , n303491 , n303492 , n303493 , 
 n303494 , n303495 , n303496 , n13069 , n303498 , n13071 , n303500 , n303501 , n303502 , n303503 , 
 n13076 , n303505 , n303506 , n13079 , n303508 , n303509 , n13082 , n303511 , n303512 , n13085 , 
 n303514 , n303515 , n303516 , n303517 , n13090 , n303519 , n303520 , n13093 , n303522 , n13095 , 
 n13096 , n303525 , n303526 , n303527 , n303528 , n13101 , n303530 , n303531 , n303532 , n303533 , 
 n13106 , n303535 , n13108 , n13109 , n303538 , n303539 , n303540 , n303541 , n303542 , n13115 , 
 n13116 , n303545 , n303546 , n13119 , n303548 , n13121 , n303550 , n303551 , n13124 , n303553 , 
 n303554 , n303555 , n303556 , n13129 , n303558 , n13131 , n303560 , n303561 , n303562 , n13135 , 
 n13136 , n13137 , n303566 , n303567 , n13140 , n303569 , n303570 , n13143 , n303572 , n303573 , 
 n303574 , n303575 , n13148 , n303577 , n13150 , n303579 , n303580 , n13153 , n303582 , n13155 , 
 n303584 , n13157 , n303586 , n303587 , n13160 , n303589 , n13162 , n303591 , n13164 , n303593 , 
 n303594 , n13167 , n13168 , n303597 , n13170 , n303599 , n303600 , n13173 , n303602 , n303603 , 
 n13176 , n13177 , n303606 , n303607 , n13180 , n303609 , n303610 , n303611 , n303612 , n303613 , 
 n303614 , n303615 , n303616 , n13189 , n303618 , n303619 , n303620 , n303621 , n303622 , n303623 , 
 n13196 , n13197 , n303626 , n303627 , n303628 , n303629 , n303630 , n303631 , n303632 , n13205 , 
 n303634 , n303635 , n303636 , n303637 , n303638 , n303639 , n13212 , n303641 , n13214 , n303643 , 
 n303644 , n13217 , n303646 , n303647 , n13220 , n303649 , n303650 , n13223 , n13224 , n303653 , 
 n13226 , n303655 , n303656 , n13229 , n303658 , n303659 , n13232 , n303661 , n303662 , n13235 , 
 n13236 , n303665 , n303666 , n13239 , n303668 , n303669 , n13242 , n13243 , n303672 , n303673 , 
 n303674 , n303675 , n303676 , n303677 , n303678 , n303679 , n303680 , n303681 , n303682 , n303683 , 
 n303684 , n303685 , n13258 , n303687 , n303688 , n303689 , n303690 , n13263 , n303692 , n303693 , 
 n13266 , n303695 , n303696 , n13269 , n13270 , n303699 , n13272 , n303701 , n303702 , n13275 , 
 n13276 , n303705 , n13278 , n303707 , n13280 , n13281 , n303710 , n303711 , n13284 , n303713 , 
 n303714 , n13287 , n303716 , n303717 , n13290 , n303719 , n303720 , n303721 , n303722 , n13295 , 
 n303724 , n13297 , n303726 , n13299 , n13300 , n13301 , n13302 , n303731 , n303732 , n13305 , 
 n303734 , n13307 , n303736 , n13309 , n303738 , n13311 , n303740 , n303741 , n13314 , n303743 , 
 n303744 , n303745 , n303746 , n303747 , n303748 , n303749 , n303750 , n303751 , n303752 , n303753 , 
 n303754 , n303755 , n303756 , n303757 , n303758 , n303759 , n303760 , n303761 , n303762 , n13335 , 
 n303764 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n303771 , n13344 , n303773 , 
 n303774 , n303775 , n303776 , n303777 , n13350 , n303779 , n303780 , n303781 , n303782 , n303783 , 
 n303784 , n303785 , n303786 , n303787 , n13360 , n303789 , n303790 , n13363 , n13364 , n303793 , 
 n303794 , n13367 , n13368 , n303797 , n303798 , n303799 , n13372 , n303801 , n13374 , n13375 , 
 n303804 , n13377 , n13378 , n13379 , n13380 , n303809 , n13382 , n303811 , n303812 , n13385 , 
 n13386 , n303815 , n303816 , n303817 , n303818 , n13391 , n303820 , n303821 , n303822 , n303823 , 
 n303824 , n303825 , n303826 , n303827 , n303828 , n303829 , n303830 , n303831 , n303832 , n303833 , 
 n13406 , n303835 , n13408 , n13409 , n303838 , n13411 , n303840 , n13413 , n303842 , n13415 , 
 n303844 , n13417 , n303846 , n303847 , n13420 , n303849 , n303850 , n303851 , n303852 , n303853 , 
 n13426 , n303855 , n303856 , n303857 , n303858 , n303859 , n303860 , n303861 , n303862 , n303863 , 
 n303864 , n303865 , n303866 , n303867 , n303868 , n13441 , n303870 , n13443 , n303872 , n303873 , 
 n303874 , n303875 , n303876 , n303877 , n13450 , n303879 , n303880 , n13453 , n303882 , n303883 , 
 n303884 , n13457 , n303886 , n13459 , n13460 , n13461 , n303890 , n13463 , n303892 , n303893 , 
 n303894 , n13467 , n303896 , n303897 , n13470 , n303899 , n303900 , n303901 , n13474 , n303903 , 
 n303904 , n13477 , n303906 , n303907 , n303908 , n303909 , n303910 , n303911 , n303912 , n303913 , 
 n303914 , n13487 , n303916 , n303917 , n303918 , n303919 , n13492 , n303921 , n303922 , n13495 , 
 n303924 , n13497 , n303926 , n13499 , n13500 , n303929 , n303930 , n303931 , n13504 , n303933 , 
 n303934 , n303935 , n303936 , n303937 , n13510 , n303939 , n303940 , n13513 , n13514 , n303943 , 
 n13516 , n303945 , n13518 , n303947 , n13520 , n303949 , n13522 , n303951 , n303952 , n303953 , 
 n13526 , n303955 , n303956 , n13529 , n303958 , n303959 , n303960 , n13533 , n303962 , n303963 , 
 n13536 , n303965 , n303966 , n13539 , n303968 , n303969 , n13542 , n303971 , n13544 , n303973 , 
 n13546 , n303975 , n13548 , n303977 , n303978 , n303979 , n13552 , n303981 , n303982 , n303983 , 
 n13556 , n303985 , n13558 , n303987 , n13560 , n303989 , n303990 , n303991 , n303992 , n303993 , 
 n303994 , n303995 , n13568 , n303997 , n303998 , n303999 , n304000 , n304001 , n13574 , n304003 , 
 n304004 , n304005 , n13578 , n304007 , n304008 , n304009 , n304010 , n304011 , n13584 , n304013 , 
 n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n304020 , n304021 , n13594 , n13595 , 
 n304024 , n13597 , n304026 , n304027 , n304028 , n13601 , n304030 , n13603 , n304032 , n304033 , 
 n13606 , n304035 , n304036 , n304037 , n304038 , n304039 , n13612 , n304041 , n13614 , n304043 , 
 n304044 , n304045 , n13618 , n304047 , n304048 , n304049 , n304050 , n304051 , n304052 , n304053 , 
 n13626 , n13627 , n304056 , n304057 , n304058 , n304059 , n304060 , n304061 , n304062 , n304063 , 
 n304064 , n13637 , n304066 , n304067 , n13640 , n304069 , n304070 , n13643 , n304072 , n304073 , 
 n13646 , n304075 , n304076 , n13649 , n304078 , n304079 , n304080 , n304081 , n304082 , n304083 , 
 n304084 , n304085 , n304086 , n304087 , n13660 , n13661 , n304090 , n304091 , n13664 , n304093 , 
 n304094 , n13667 , n304096 , n304097 , n13670 , n13671 , n304100 , n13673 , n13674 , n13675 , 
 n13676 , n304105 , n304106 , n13679 , n304108 , n304109 , n13682 , n13683 , n13684 , n13685 , 
 n13686 , n13687 , n13688 , n13689 , n13690 , n304119 , n13692 , n304121 , n13694 , n13695 , 
 n304124 , n13697 , n304126 , n304127 , n13700 , n304129 , n304130 , n304131 , n304132 , n13705 , 
 n13706 , n13707 , n13708 , n13709 , n13710 , n304139 , n13712 , n13713 , n13714 , n13715 , 
 n13716 , n304145 , n13718 , n304147 , n304148 , n13721 , n304150 , n13723 , n304152 , n304153 , 
 n13726 , n304155 , n304156 , n13729 , n304158 , n304159 , n304160 , n304161 , n304162 , n13735 , 
 n304164 , n304165 , n13738 , n304167 , n304168 , n13741 , n304170 , n304171 , n304172 , n13745 , 
 n304174 , n304175 , n304176 , n304177 , n13750 , n13751 , n13752 , n304181 , n304182 , n304183 , 
 n13756 , n304185 , n304186 , n304187 , n304188 , n304189 , n304190 , n304191 , n13764 , n304193 , 
 n304194 , n13767 , n304196 , n304197 , n13770 , n13771 , n304200 , n13773 , n304202 , n304203 , 
 n304204 , n304205 , n304206 , n13779 , n13780 , n304209 , n304210 , n304211 , n304212 , n304213 , 
 n13786 , n304215 , n304216 , n304217 , n304218 , n304219 , n304220 , n13793 , n304222 , n304223 , 
 n304224 , n304225 , n304226 , n304227 , n13800 , n304229 , n304230 , n304231 , n304232 , n304233 , 
 n304234 , n304235 , n304236 , n304237 , n304238 , n13811 , n304240 , n304241 , n13814 , n304243 , 
 n13816 , n304245 , n304246 , n304247 , n304248 , n304249 , n304250 , n304251 , n304252 , n304253 , 
 n304254 , n304255 , n304256 , n304257 , n304258 , n13831 , n304260 , n13833 , n13834 , n13835 , 
 n304264 , n13837 , n304266 , n304267 , n304268 , n304269 , n304270 , n304271 , n304272 , n304273 , 
 n13846 , n304275 , n304276 , n13849 , n304278 , n304279 , n13852 , n13853 , n304282 , n13855 , 
 n304284 , n304285 , n13858 , n304287 , n304288 , n304289 , n304290 , n304291 , n304292 , n304293 , 
 n304294 , n304295 , n304296 , n304297 , n304298 , n304299 , n304300 , n13873 , n304302 , n304303 , 
 n304304 , n13877 , n13878 , n304307 , n13880 , n304309 , n304310 , n304311 , n304312 , n13885 , 
 n304314 , n304315 , n304316 , n13889 , n304318 , n304319 , n13892 , n304321 , n304322 , n304323 , 
 n304324 , n304325 , n13898 , n304327 , n13900 , n13901 , n13902 , n304331 , n304332 , n304333 , 
 n304334 , n304335 , n13908 , n304337 , n304338 , n13911 , n304340 , n13913 , n304342 , n304343 , 
 n304344 , n13917 , n304346 , n304347 , n13920 , n304349 , n13922 , n304351 , n304352 , n304353 , 
 n304354 , n304355 , n304356 , n13929 , n304358 , n304359 , n13932 , n13933 , n13934 , n13935 , 
 n304364 , n304365 , n304366 , n304367 , n13940 , n304369 , n13942 , n304371 , n304372 , n13945 , 
 n304374 , n13947 , n13948 , n304377 , n13950 , n13951 , n304380 , n304381 , n304382 , n304383 , 
 n13956 , n304385 , n304386 , n304387 , n13960 , n304389 , n304390 , n13963 , n304392 , n304393 , 
 n13966 , n304395 , n304396 , n13969 , n304398 , n304399 , n13972 , n13973 , n13974 , n13975 , 
 n304404 , n304405 , n13978 , n13979 , n13980 , n13981 , n13982 , n304411 , n304412 , n13985 , 
 n304414 , n304415 , n13988 , n304417 , n304418 , n13991 , n304420 , n13993 , n304422 , n13995 , 
 n304424 , n304425 , n13998 , n304427 , n304428 , n14001 , n304430 , n304431 , n304432 , n304433 , 
 n14006 , n304435 , n304436 , n304437 , n14010 , n304439 , n14012 , n304441 , n14014 , n14015 , 
 n14016 , n14017 , n14018 , n304447 , n304448 , n304449 , n304450 , n304451 , n304452 , n304453 , 
 n14026 , n304455 , n304456 , n304457 , n14030 , n304459 , n14032 , n14033 , n304462 , n304463 , 
 n304464 , n304465 , n304466 , n304467 , n14040 , n304469 , n304470 , n304471 , n304472 , n304473 , 
 n14046 , n304475 , n14048 , n304477 , n304478 , n14051 , n304480 , n304481 , n304482 , n14055 , 
 n304484 , n304485 , n304486 , n304487 , n304488 , n304489 , n304490 , n304491 , n14064 , n304493 , 
 n304494 , n304495 , n304496 , n304497 , n304498 , n14071 , n304500 , n304501 , n14074 , n14075 , 
 n304504 , n304505 , n304506 , n14079 , n14080 , n304509 , n304510 , n304511 , n304512 , n304513 , 
 n304514 , n14087 , n304516 , n304517 , n304518 , n304519 , n304520 , n304521 , n14094 , n14095 , 
 n304524 , n14097 , n304526 , n304527 , n14100 , n304529 , n14102 , n304531 , n14104 , n304533 , 
 n304534 , n14107 , n304536 , n304537 , n14110 , n304539 , n14112 , n304541 , n14114 , n14115 , 
 n14116 , n14117 , n304546 , n304547 , n304548 , n304549 , n14122 , n14123 , n14124 , n304553 , 
 n304554 , n14127 , n14128 , n304557 , n14130 , n304559 , n304560 , n304561 , n304562 , n304563 , 
 n304564 , n304565 , n304566 , n14139 , n14140 , n304569 , n304570 , n304571 , n304572 , n304573 , 
 n304574 , n304575 , n304576 , n304577 , n14150 , n304579 , n14152 , n304581 , n14154 , n14155 , 
 n304584 , n304585 , n304586 , n304587 , n304588 , n304589 , n14162 , n304591 , n304592 , n304593 , 
 n304594 , n14167 , n304596 , n304597 , n304598 , n304599 , n304600 , n304601 , n304602 , n304603 , 
 n304604 , n304605 , n304606 , n14179 , n304608 , n304609 , n304610 , n304611 , n14184 , n14185 , 
 n304614 , n304615 , n14188 , n304617 , n304618 , n304619 , n14192 , n304621 , n304622 , n14195 , 
 n304624 , n304625 , n14198 , n304627 , n14200 , n304629 , n304630 , n304631 , n14204 , n304633 , 
 n304634 , n304635 , n14208 , n304637 , n14210 , n304639 , n14212 , n304641 , n14214 , n304643 , 
 n304644 , n304645 , n304646 , n304647 , n304648 , n304649 , n304650 , n304651 , n304652 , n304653 , 
 n14226 , n304655 , n304656 , n304657 , n304658 , n304659 , n304660 , n304661 , n304662 , n14235 , 
 n14236 , n14237 , n14238 , n304667 , n304668 , n14241 , n304670 , n304671 , n304672 , n304673 , 
 n304674 , n304675 , n14248 , n304677 , n304678 , n304679 , n304680 , n304681 , n304682 , n304683 , 
 n304684 , n304685 , n304686 , n304687 , n304688 , n304689 , n304690 , n304691 , n304692 , n304693 , 
 n304694 , n304695 , n304696 , n304697 , n304698 , n14271 , n14272 , n304701 , n304702 , n14275 , 
 n304704 , n14277 , n304706 , n304707 , n304708 , n304709 , n304710 , n14283 , n304712 , n304713 , 
 n304714 , n14287 , n14288 , n14289 , n304718 , n14291 , n304720 , n304721 , n304722 , n304723 , 
 n304724 , n304725 , n304726 , n14299 , n304728 , n304729 , n14302 , n304731 , n304732 , n304733 , 
 n304734 , n304735 , n304736 , n14309 , n304738 , n304739 , n304740 , n304741 , n304742 , n304743 , 
 n304744 , n14317 , n14318 , n304747 , n14320 , n304749 , n14322 , n14323 , n304752 , n14325 , 
 n304754 , n304755 , n304756 , n14329 , n304758 , n14331 , n304760 , n14333 , n304762 , n304763 , 
 n304764 , n304765 , n304766 , n304767 , n304768 , n304769 , n304770 , n304771 , n304772 , n304773 , 
 n304774 , n304775 , n304776 , n14349 , n304778 , n304779 , n14352 , n304781 , n304782 , n304783 , 
 n304784 , n14357 , n304786 , n304787 , n14360 , n304789 , n304790 , n14363 , n304792 , n304793 , 
 n304794 , n304795 , n304796 , n14369 , n14370 , n304799 , n304800 , n14373 , n304802 , n14375 , 
 n304804 , n304805 , n304806 , n304807 , n304808 , n304809 , n304810 , n304811 , n304812 , n304813 , 
 n304814 , n304815 , n304816 , n304817 , n14390 , n304819 , n304820 , n304821 , n304822 , n304823 , 
 n304824 , n304825 , n14398 , n304827 , n304828 , n14401 , n14402 , n14403 , n304832 , n14405 , 
 n304834 , n304835 , n14408 , n304837 , n304838 , n14411 , n304840 , n304841 , n304842 , n304843 , 
 n304844 , n304845 , n304846 , n14419 , n14420 , n14421 , n14422 , n304851 , n304852 , n14425 , 
 n304854 , n304855 , n304856 , n304857 , n304858 , n304859 , n304860 , n14433 , n304862 , n14435 , 
 n304864 , n304865 , n14438 , n14439 , n304868 , n304869 , n304870 , n304871 , n14444 , n304873 , 
 n14446 , n14447 , n14448 , n304877 , n304878 , n304879 , n304880 , n304881 , n304882 , n304883 , 
 n304884 , n14457 , n304886 , n304887 , n14460 , n304889 , n304890 , n304891 , n304892 , n304893 , 
 n304894 , n304895 , n304896 , n14469 , n304898 , n304899 , n304900 , n304901 , n304902 , n304903 , 
 n304904 , n14477 , n304906 , n304907 , n14480 , n304909 , n304910 , n14483 , n304912 , n304913 , 
 n14486 , n14487 , n304916 , n304917 , n14490 , n304919 , n304920 , n14493 , n304922 , n14495 , 
 n304924 , n304925 , n304926 , n304927 , n304928 , n14501 , n304930 , n304931 , n304932 , n304933 , 
 n14506 , n14507 , n304936 , n14509 , n304938 , n304939 , n14512 , n304941 , n304942 , n304943 , 
 n304944 , n304945 , n304946 , n304947 , n304948 , n304949 , n14522 , n14523 , n304952 , n304953 , 
 n304954 , n14527 , n304956 , n304957 , n14530 , n14531 , n14532 , n14533 , n304962 , n304963 , 
 n304964 , n14537 , n304966 , n304967 , n304968 , n304969 , n14542 , n304971 , n304972 , n304973 , 
 n304974 , n304975 , n304976 , n304977 , n14550 , n304979 , n304980 , n304981 , n304982 , n14555 , 
 n304984 , n14557 , n304986 , n304987 , n304988 , n304989 , n14562 , n14563 , n14564 , n304993 , 
 n14566 , n304995 , n304996 , n304997 , n304998 , n14571 , n305000 , n305001 , n305002 , n305003 , 
 n305004 , n305005 , n305006 , n305007 , n305008 , n305009 , n14582 , n305011 , n305012 , n305013 , 
 n14586 , n305015 , n305016 , n14589 , n305018 , n305019 , n305020 , n305021 , n305022 , n305023 , 
 n14596 , n305025 , n305026 , n305027 , n305028 , n305029 , n305030 , n305031 , n305032 , n305033 , 
 n14606 , n305035 , n305036 , n305037 , n305038 , n305039 , n305040 , n305041 , n305042 , n305043 , 
 n305044 , n305045 , n305046 , n305047 , n305048 , n305049 , n305050 , n14623 , n305052 , n305053 , 
 n305054 , n305055 , n305056 , n305057 , n305058 , n305059 , n305060 , n305061 , n305062 , n305063 , 
 n305064 , n305065 , n305066 , n305067 , n305068 , n14641 , n305070 , n305071 , n14644 , n305073 , 
 n305074 , n305075 , n14648 , n305077 , n305078 , n305079 , n305080 , n305081 , n305082 , n305083 , 
 n305084 , n305085 , n305086 , n305087 , n305088 , n305089 , n305090 , n305091 , n305092 , n305093 , 
 n14666 , n305095 , n305096 , n305097 , n305098 , n305099 , n305100 , n14673 , n305102 , n305103 , 
 n305104 , n305105 , n305106 , n305107 , n14680 , n14681 , n305110 , n305111 , n305112 , n305113 , 
 n14686 , n305115 , n305116 , n305117 , n305118 , n14691 , n14692 , n305121 , n305122 , n305123 , 
 n305124 , n305125 , n305126 , n305127 , n305128 , n14701 , n305130 , n305131 , n305132 , n305133 , 
 n305134 , n305135 , n305136 , n305137 , n305138 , n305139 , n14712 , n14713 , n14714 , n305143 , 
 n305144 , n305145 , n14718 , n305147 , n14720 , n305149 , n305150 , n14723 , n305152 , n305153 , 
 n305154 , n305155 , n305156 , n305157 , n305158 , n305159 , n305160 , n305161 , n305162 , n14735 , 
 n14736 , n305165 , n305166 , n305167 , n305168 , n305169 , n305170 , n305171 , n305172 , n305173 , 
 n305174 , n305175 , n305176 , n305177 , n14750 , n305179 , n305180 , n14753 , n305182 , n305183 , 
 n14756 , n305185 , n305186 , n14759 , n14760 , n305189 , n14762 , n305191 , n305192 , n305193 , 
 n14766 , n305195 , n305196 , n305197 , n305198 , n305199 , n305200 , n14773 , n305202 , n305203 , 
 n14776 , n305205 , n14778 , n305207 , n305208 , n305209 , n305210 , n305211 , n305212 , n305213 , 
 n305214 , n305215 , n14788 , n305217 , n14790 , n305219 , n305220 , n14793 , n305222 , n305223 , 
 n305224 , n305225 , n305226 , n305227 , n305228 , n305229 , n305230 , n305231 , n305232 , n14805 , 
 n305234 , n305235 , n305236 , n14809 , n14810 , n305239 , n305240 , n305241 , n305242 , n305243 , 
 n305244 , n305245 , n305246 , n305247 , n305248 , n305249 , n14822 , n305251 , n305252 , n14825 , 
 n305254 , n305255 , n305256 , n305257 , n305258 , n305259 , n14832 , n305261 , n14834 , n14835 , 
 n14836 , n305265 , n14838 , n14839 , n305268 , n305269 , n305270 , n305271 , n305272 , n305273 , 
 n305274 , n305275 , n305276 , n14849 , n305278 , n305279 , n305280 , n14853 , n305282 , n305283 , 
 n305284 , n305285 , n305286 , n305287 , n14860 , n305289 , n305290 , n305291 , n305292 , n305293 , 
 n305294 , n305295 , n305296 , n305297 , n305298 , n14871 , n305300 , n305301 , n305302 , n305303 , 
 n305304 , n305305 , n305306 , n305307 , n305308 , n305309 , n305310 , n305311 , n305312 , n305313 , 
 n14886 , n14887 , n14888 , n305317 , n14890 , n305319 , n305320 , n305321 , n14894 , n305323 , 
 n305324 , n14897 , n305326 , n305327 , n14900 , n14901 , n305330 , n305331 , n305332 , n305333 , 
 n305334 , n305335 , n14908 , n305337 , n305338 , n305339 , n305340 , n305341 , n305342 , n305343 , 
 n305344 , n305345 , n14918 , n305347 , n305348 , n305349 , n305350 , n305351 , n305352 , n305353 , 
 n305354 , n305355 , n305356 , n305357 , n305358 , n305359 , n305360 , n305361 , n305362 , n305363 , 
 n305364 , n305365 , n305366 , n14939 , n305368 , n305369 , n305370 , n14943 , n14944 , n305373 , 
 n14946 , n305375 , n14948 , n305377 , n305378 , n305379 , n305380 , n305381 , n305382 , n305383 , 
 n305384 , n305385 , n14958 , n14959 , n14960 , n14961 , n305390 , n305391 , n305392 , n305393 , 
 n305394 , n14967 , n305396 , n14969 , n305398 , n305399 , n14972 , n305401 , n305402 , n305403 , 
 n305404 , n305405 , n305406 , n305407 , n305408 , n305409 , n305410 , n14983 , n305412 , n305413 , 
 n305414 , n305415 , n14988 , n14989 , n305418 , n14991 , n14992 , n305421 , n14994 , n305423 , 
 n305424 , n305425 , n14998 , n305427 , n15000 , n305429 , n305430 , n305431 , n305432 , n305433 , 
 n15006 , n305435 , n305436 , n305437 , n305438 , n305439 , n305440 , n305441 , n305442 , n15015 , 
 n305444 , n305445 , n15018 , n15019 , n305448 , n305449 , n305450 , n305451 , n305452 , n305453 , 
 n305454 , n305455 , n305456 , n15029 , n305458 , n305459 , n305460 , n305461 , n305462 , n15035 , 
 n305464 , n305465 , n305466 , n305467 , n305468 , n305469 , n305470 , n305471 , n305472 , n305473 , 
 n305474 , n305475 , n15048 , n305477 , n305478 , n305479 , n305480 , n305481 , n305482 , n305483 , 
 n15056 , n15057 , n305486 , n305487 , n305488 , n305489 , n305490 , n305491 , n15064 , n15065 , 
 n305494 , n15067 , n15068 , n305497 , n305498 , n15071 , n305500 , n305501 , n305502 , n305503 , 
 n305504 , n305505 , n305506 , n15079 , n305508 , n15081 , n305510 , n15083 , n305512 , n305513 , 
 n305514 , n305515 , n305516 , n305517 , n305518 , n305519 , n305520 , n305521 , n305522 , n305523 , 
 n305524 , n305525 , n305526 , n305527 , n305528 , n15101 , n305530 , n305531 , n305532 , n305533 , 
 n305534 , n15107 , n15108 , n305537 , n305538 , n305539 , n15112 , n305541 , n305542 , n305543 , 
 n305544 , n15117 , n305546 , n305547 , n305548 , n305549 , n305550 , n305551 , n15124 , n305553 , 
 n305554 , n305555 , n15128 , n15129 , n305558 , n305559 , n305560 , n305561 , n305562 , n305563 , 
 n305564 , n15137 , n305566 , n305567 , n305568 , n15141 , n305570 , n305571 , n15144 , n15145 , 
 n305574 , n15147 , n305576 , n305577 , n305578 , n15151 , n305580 , n305581 , n15154 , n305583 , 
 n305584 , n15157 , n15158 , n305587 , n15160 , n15161 , n305590 , n305591 , n15164 , n305593 , 
 n305594 , n305595 , n305596 , n305597 , n305598 , n15171 , n305600 , n305601 , n15174 , n305603 , 
 n305604 , n15177 , n305606 , n305607 , n305608 , n15181 , n305610 , n305611 , n15184 , n15185 , 
 n305614 , n15187 , n305616 , n305617 , n305618 , n305619 , n15192 , n305621 , n305622 , n305623 , 
 n305624 , n305625 , n15198 , n305627 , n305628 , n15201 , n305630 , n15203 , n305632 , n305633 , 
 n15206 , n15207 , n305636 , n305637 , n305638 , n305639 , n305640 , n15213 , n305642 , n305643 , 
 n305644 , n305645 , n305646 , n15219 , n15220 , n305649 , n305650 , n305651 , n305652 , n15225 , 
 n15226 , n305655 , n305656 , n15229 , n305658 , n305659 , n305660 , n15233 , n305662 , n15235 , 
 n305664 , n305665 , n305666 , n305667 , n305668 , n15241 , n305670 , n305671 , n15244 , n15245 , 
 n305674 , n15247 , n305676 , n305677 , n305678 , n15251 , n15252 , n305681 , n305682 , n305683 , 
 n305684 , n305685 , n15258 , n305687 , n305688 , n305689 , n305690 , n305691 , n305692 , n305693 , 
 n305694 , n305695 , n305696 , n305697 , n15270 , n305699 , n305700 , n305701 , n305702 , n305703 , 
 n305704 , n15277 , n15278 , n305707 , n305708 , n305709 , n15282 , n305711 , n305712 , n305713 , 
 n305714 , n15287 , n15288 , n305717 , n305718 , n305719 , n305720 , n305721 , n305722 , n305723 , 
 n305724 , n305725 , n15298 , n305727 , n305728 , n15301 , n305730 , n305731 , n305732 , n305733 , 
 n305734 , n305735 , n15308 , n15309 , n305738 , n305739 , n305740 , n305741 , n305742 , n305743 , 
 n305744 , n305745 , n305746 , n305747 , n305748 , n305749 , n305750 , n305751 , n305752 , n305753 , 
 n305754 , n15327 , n15328 , n305757 , n15330 , n15331 , n305760 , n305761 , n305762 , n305763 , 
 n305764 , n305765 , n305766 , n305767 , n15340 , n15341 , n305770 , n305771 , n15344 , n15345 , 
 n15346 , n305775 , n15348 , n15349 , n305778 , n15351 , n305780 , n305781 , n15354 , n305783 , 
 n305784 , n15357 , n305786 , n305787 , n305788 , n305789 , n305790 , n305791 , n15364 , n305793 , 
 n15366 , n305795 , n305796 , n305797 , n305798 , n305799 , n305800 , n15373 , n15374 , n15375 , 
 n305804 , n15377 , n15378 , n305807 , n15380 , n305809 , n15382 , n305811 , n305812 , n15385 , 
 n305814 , n305815 , n305816 , n15389 , n305818 , n305819 , n305820 , n305821 , n305822 , n305823 , 
 n305824 , n305825 , n305826 , n305827 , n305828 , n305829 , n305830 , n15403 , n305832 , n305833 , 
 n305834 , n305835 , n305836 , n305837 , n305838 , n305839 , n305840 , n305841 , n305842 , n305843 , 
 n305844 , n305845 , n15418 , n305847 , n305848 , n305849 , n305850 , n305851 , n305852 , n15425 , 
 n15426 , n15427 , n15428 , n305857 , n305858 , n15431 , n305860 , n305861 , n15434 , n305863 , 
 n305864 , n305865 , n15438 , n305867 , n305868 , n305869 , n305870 , n305871 , n305872 , n305873 , 
 n305874 , n305875 , n305876 , n15449 , n305878 , n305879 , n15452 , n305881 , n305882 , n305883 , 
 n305884 , n305885 , n305886 , n305887 , n305888 , n305889 , n305890 , n15463 , n305892 , n305893 , 
 n15466 , n15467 , n15468 , n15469 , n305898 , n305899 , n305900 , n305901 , n305902 , n305903 , 
 n15476 , n305905 , n305906 , n305907 , n305908 , n305909 , n15482 , n15483 , n15484 , n305913 , 
 n305914 , n305915 , n15488 , n15489 , n305918 , n305919 , n305920 , n305921 , n305922 , n305923 , 
 n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n305930 , n15503 , n305932 , n305933 , 
 n305934 , n305935 , n305936 , n15509 , n15510 , n305939 , n305940 , n15513 , n305942 , n305943 , 
 n15516 , n305945 , n305946 , n305947 , n15520 , n15521 , n305950 , n305951 , n305952 , n305953 , 
 n305954 , n305955 , n305956 , n305957 , n15530 , n305959 , n305960 , n305961 , n305962 , n305963 , 
 n15536 , n305965 , n305966 , n305967 , n305968 , n15541 , n305970 , n305971 , n15544 , n305973 , 
 n305974 , n15547 , n305976 , n305977 , n15550 , n305979 , n305980 , n305981 , n305982 , n305983 , 
 n305984 , n15557 , n15558 , n305987 , n305988 , n15561 , n15562 , n305991 , n305992 , n305993 , 
 n305994 , n15567 , n305996 , n305997 , n15570 , n15571 , n15572 , n306001 , n15574 , n15575 , 
 n306004 , n306005 , n306006 , n306007 , n306008 , n15581 , n15582 , n306011 , n306012 , n306013 , 
 n306014 , n306015 , n306016 , n306017 , n306018 , n306019 , n306020 , n306021 , n15594 , n15595 , 
 n306024 , n306025 , n306026 , n306027 , n306028 , n306029 , n306030 , n306031 , n306032 , n15605 , 
 n15606 , n306035 , n306036 , n306037 , n306038 , n306039 , n306040 , n15613 , n306042 , n306043 , 
 n306044 , n306045 , n306046 , n15619 , n306048 , n306049 , n306050 , n306051 , n15624 , n15625 , 
 n306054 , n15627 , n306056 , n306057 , n15630 , n306059 , n306060 , n15633 , n306062 , n306063 , 
 n306064 , n306065 , n306066 , n306067 , n306068 , n306069 , n306070 , n306071 , n15644 , n306073 , 
 n15646 , n15647 , n306076 , n306077 , n306078 , n306079 , n306080 , n15653 , n306082 , n306083 , 
 n15656 , n306085 , n15658 , n306087 , n15660 , n306089 , n306090 , n306091 , n306092 , n306093 , 
 n15666 , n15667 , n306096 , n306097 , n306098 , n306099 , n15672 , n306101 , n306102 , n15675 , 
 n306104 , n306105 , n306106 , n306107 , n306108 , n306109 , n306110 , n15683 , n306112 , n306113 , 
 n15686 , n306115 , n306116 , n306117 , n306118 , n306119 , n306120 , n306121 , n15694 , n306123 , 
 n15696 , n15697 , n306126 , n306127 , n15700 , n306129 , n306130 , n306131 , n306132 , n306133 , 
 n306134 , n15707 , n306136 , n306137 , n15710 , n306139 , n306140 , n306141 , n306142 , n15715 , 
 n306144 , n15717 , n15718 , n306147 , n306148 , n15721 , n306150 , n306151 , n306152 , n306153 , 
 n306154 , n306155 , n306156 , n15729 , n306158 , n15731 , n306160 , n306161 , n15734 , n306163 , 
 n15736 , n306165 , n15738 , n306167 , n15740 , n15741 , n15742 , n306171 , n306172 , n306173 , 
 n15746 , n15747 , n306176 , n306177 , n306178 , n306179 , n306180 , n15753 , n15754 , n15755 , 
 n15756 , n15757 , n306186 , n15759 , n306188 , n306189 , n15762 , n306191 , n306192 , n306193 , 
 n306194 , n306195 , n306196 , n15769 , n306198 , n15771 , n306200 , n306201 , n306202 , n306203 , 
 n306204 , n306205 , n306206 , n306207 , n306208 , n306209 , n306210 , n306211 , n306212 , n306213 , 
 n306214 , n306215 , n306216 , n306217 , n306218 , n306219 , n306220 , n15793 , n306222 , n306223 , 
 n306224 , n306225 , n306226 , n306227 , n306228 , n306229 , n306230 , n15803 , n15804 , n306233 , 
 n306234 , n306235 , n15808 , n15809 , n306238 , n306239 , n306240 , n306241 , n306242 , n306243 , 
 n306244 , n306245 , n306246 , n306247 , n306248 , n306249 , n306250 , n306251 , n306252 , n306253 , 
 n306254 , n306255 , n15828 , n306257 , n306258 , n306259 , n306260 , n306261 , n306262 , n306263 , 
 n15836 , n306265 , n306266 , n306267 , n306268 , n15841 , n306270 , n306271 , n306272 , n306273 , 
 n306274 , n306275 , n306276 , n15849 , n306278 , n306279 , n306280 , n306281 , n306282 , n306283 , 
 n306284 , n306285 , n306286 , n306287 , n15860 , n15861 , n306290 , n306291 , n306292 , n306293 , 
 n306294 , n306295 , n306296 , n306297 , n306298 , n306299 , n306300 , n306301 , n15874 , n15875 , 
 n15876 , n15877 , n306306 , n306307 , n306308 , n306309 , n306310 , n306311 , n306312 , n306313 , 
 n15886 , n15887 , n306316 , n15889 , n306318 , n15891 , n306320 , n306321 , n306322 , n306323 , 
 n306324 , n306325 , n15898 , n306327 , n306328 , n306329 , n306330 , n306331 , n306332 , n306333 , 
 n306334 , n306335 , n306336 , n306337 , n306338 , n306339 , n306340 , n306341 , n306342 , n306343 , 
 n306344 , n306345 , n306346 , n306347 , n306348 , n306349 , n15922 , n306351 , n306352 , n15925 , 
 n15926 , n306355 , n15928 , n15929 , n15930 , n306359 , n15932 , n306361 , n306362 , n306363 , 
 n306364 , n306365 , n306366 , n306367 , n306368 , n306369 , n15942 , n15943 , n15944 , n306373 , 
 n306374 , n306375 , n15948 , n306377 , n15950 , n306379 , n306380 , n306381 , n15954 , n15955 , 
 n306384 , n15957 , n306386 , n306387 , n15960 , n306389 , n306390 , n306391 , n15964 , n306393 , 
 n306394 , n15967 , n306396 , n306397 , n306398 , n15971 , n306400 , n306401 , n306402 , n306403 , 
 n306404 , n15977 , n306406 , n306407 , n306408 , n306409 , n306410 , n15983 , n15984 , n306413 , 
 n306414 , n15987 , n15988 , n306417 , n306418 , n15991 , n306420 , n306421 , n306422 , n306423 , 
 n306424 , n15997 , n306426 , n306427 , n306428 , n306429 , n306430 , n16003 , n306432 , n306433 , 
 n306434 , n306435 , n306436 , n306437 , n306438 , n306439 , n306440 , n306441 , n306442 , n306443 , 
 n16016 , n306445 , n306446 , n306447 , n16020 , n16021 , n306450 , n16023 , n306452 , n16025 , 
 n16026 , n306455 , n306456 , n306457 , n306458 , n306459 , n306460 , n306461 , n306462 , n306463 , 
 n306464 , n306465 , n306466 , n306467 , n16040 , n306469 , n306470 , n16043 , n306472 , n306473 , 
 n16046 , n306475 , n16048 , n16049 , n306478 , n16051 , n306480 , n306481 , n16054 , n306483 , 
 n306484 , n306485 , n306486 , n306487 , n306488 , n16061 , n306490 , n306491 , n306492 , n306493 , 
 n306494 , n16067 , n306496 , n306497 , n306498 , n306499 , n306500 , n16073 , n306502 , n16075 , 
 n16076 , n306505 , n306506 , n16079 , n306508 , n306509 , n16082 , n306511 , n306512 , n16085 , 
 n306514 , n16087 , n16088 , n306517 , n306518 , n16091 , n306520 , n16093 , n306522 , n306523 , 
 n16096 , n306525 , n306526 , n306527 , n16100 , n16101 , n16102 , n306531 , n306532 , n306533 , 
 n16106 , n16107 , n306536 , n306537 , n16110 , n306539 , n306540 , n16113 , n306542 , n306543 , 
 n306544 , n16117 , n306546 , n306547 , n16120 , n306549 , n16122 , n306551 , n16124 , n16125 , 
 n306554 , n306555 , n16128 , n306557 , n306558 , n306559 , n306560 , n306561 , n306562 , n306563 , 
 n306564 , n306565 , n306566 , n306567 , n306568 , n306569 , n306570 , n306571 , n306572 , n306573 , 
 n306574 , n16147 , n16148 , n306577 , n306578 , n306579 , n16152 , n306581 , n306582 , n16155 , 
 n306584 , n306585 , n16158 , n306587 , n306588 , n16161 , n306590 , n306591 , n306592 , n16165 , 
 n16166 , n306595 , n306596 , n306597 , n306598 , n306599 , n306600 , n16173 , n306602 , n306603 , 
 n16176 , n306605 , n306606 , n306607 , n306608 , n306609 , n16182 , n306611 , n306612 , n16185 , 
 n16186 , n306615 , n306616 , n306617 , n306618 , n306619 , n16192 , n16193 , n306622 , n306623 , 
 n306624 , n306625 , n306626 , n306627 , n16200 , n16201 , n16202 , n306631 , n306632 , n16205 , 
 n306634 , n16207 , n16208 , n306637 , n306638 , n16211 , n16212 , n306641 , n306642 , n306643 , 
 n306644 , n16217 , n306646 , n16219 , n306648 , n306649 , n306650 , n306651 , n306652 , n306653 , 
 n306654 , n306655 , n16228 , n306657 , n306658 , n16231 , n306660 , n306661 , n16234 , n306663 , 
 n16236 , n306665 , n306666 , n16239 , n306668 , n306669 , n306670 , n306671 , n306672 , n16245 , 
 n306674 , n306675 , n16248 , n16249 , n306678 , n16251 , n306680 , n16253 , n16254 , n306683 , 
 n306684 , n306685 , n16258 , n16259 , n306688 , n16261 , n306690 , n16263 , n306692 , n16265 , 
 n306694 , n16267 , n306696 , n306697 , n306698 , n306699 , n306700 , n16273 , n16274 , n306703 , 
 n306704 , n306705 , n306706 , n306707 , n306708 , n306709 , n306710 , n306711 , n16284 , n306713 , 
 n306714 , n306715 , n306716 , n16289 , n306718 , n306719 , n306720 , n16293 , n16294 , n306723 , 
 n306724 , n16297 , n16298 , n16299 , n16300 , n16301 , n306730 , n306731 , n306732 , n306733 , 
 n306734 , n306735 , n16308 , n306737 , n306738 , n16311 , n16312 , n16313 , n306742 , n16315 , 
 n306744 , n16317 , n16318 , n306747 , n306748 , n306749 , n306750 , n306751 , n306752 , n16325 , 
 n306754 , n306755 , n16328 , n306757 , n16330 , n16331 , n16332 , n16333 , n306762 , n306763 , 
 n306764 , n16337 , n306766 , n306767 , n16340 , n306769 , n306770 , n306771 , n16344 , n306773 , 
 n306774 , n306775 , n306776 , n306777 , n306778 , n306779 , n306780 , n306781 , n16354 , n306783 , 
 n16356 , n16357 , n16358 , n16359 , n306788 , n306789 , n306790 , n306791 , n16364 , n306793 , 
 n306794 , n306795 , n306796 , n16369 , n306798 , n306799 , n306800 , n306801 , n16374 , n306803 , 
 n306804 , n16377 , n306806 , n306807 , n16380 , n306809 , n306810 , n306811 , n16384 , n306813 , 
 n306814 , n16387 , n306816 , n306817 , n16390 , n306819 , n306820 , n16393 , n306822 , n306823 , 
 n16396 , n16397 , n306826 , n306827 , n306828 , n306829 , n306830 , n306831 , n306832 , n16405 , 
 n306834 , n16407 , n306836 , n306837 , n16410 , n306839 , n306840 , n16413 , n306842 , n306843 , 
 n306844 , n306845 , n16418 , n306847 , n306848 , n16421 , n306850 , n16423 , n306852 , n16425 , 
 n16426 , n306855 , n306856 , n16429 , n306858 , n306859 , n16432 , n306861 , n16434 , n16435 , 
 n306864 , n16437 , n16438 , n16439 , n16440 , n306869 , n306870 , n16443 , n16444 , n16445 , 
 n16446 , n306875 , n306876 , n306877 , n16450 , n16451 , n306880 , n306881 , n306882 , n306883 , 
 n16456 , n306885 , n306886 , n16459 , n306888 , n306889 , n306890 , n16463 , n306892 , n16465 , 
 n16466 , n306895 , n306896 , n306897 , n16470 , n306899 , n306900 , n16473 , n306902 , n306903 , 
 n16476 , n306905 , n306906 , n306907 , n306908 , n16481 , n306910 , n16483 , n16484 , n306913 , 
 n306914 , n306915 , n306916 , n16489 , n306918 , n16491 , n16492 , n306921 , n306922 , n16495 , 
 n306924 , n306925 , n16498 , n306927 , n306928 , n16501 , n306930 , n306931 , n16504 , n306933 , 
 n306934 , n306935 , n306936 , n306937 , n16510 , n16511 , n306940 , n306941 , n306942 , n306943 , 
 n306944 , n306945 , n16518 , n306947 , n306948 , n16521 , n306950 , n306951 , n306952 , n16525 , 
 n306954 , n16527 , n16528 , n306957 , n306958 , n306959 , n16532 , n306961 , n306962 , n16535 , 
 n306964 , n306965 , n16538 , n306967 , n306968 , n16541 , n306970 , n16543 , n306972 , n16545 , 
 n16546 , n306975 , n306976 , n306977 , n16550 , n306979 , n306980 , n16553 , n306982 , n306983 , 
 n16556 , n306985 , n306986 , n16559 , n306988 , n306989 , n306990 , n16563 , n306992 , n16565 , 
 n16566 , n306995 , n306996 , n306997 , n16570 , n306999 , n307000 , n16573 , n307002 , n307003 , 
 n16576 , n307005 , n307006 , n307007 , n307008 , n16581 , n307010 , n307011 , n307012 , n307013 , 
 n16586 , n307015 , n307016 , n307017 , n16590 , n16591 , n307020 , n307021 , n307022 , n307023 , 
 n307024 , n307025 , n307026 , n307027 , n307028 , n16601 , n307030 , n307031 , n16604 , n307033 , 
 n307034 , n16607 , n307036 , n307037 , n16610 , n307039 , n307040 , n16613 , n307042 , n16615 , 
 n16616 , n307045 , n307046 , n307047 , n16620 , n307049 , n307050 , n16623 , n307052 , n307053 , 
 n16626 , n307055 , n307056 , n16629 , n307058 , n16631 , n16632 , n16633 , n307062 , n307063 , 
 n16636 , n307065 , n307066 , n16639 , n307068 , n307069 , n16642 , n307071 , n16644 , n16645 , 
 n307074 , n307075 , n16648 , n307077 , n307078 , n16651 , n307080 , n307081 , n16654 , n307083 , 
 n16656 , n307085 , n307086 , n307087 , n307088 , n307089 , n307090 , n307091 , n16664 , n307093 , 
 n307094 , n16667 , n307096 , n307097 , n16670 , n16671 , n16672 , n16673 , n16674 , n307103 , 
 n307104 , n16677 , n307106 , n307107 , n16680 , n16681 , n16682 , n16683 , n307112 , n307113 , 
 n16686 , n307115 , n307116 , n16689 , n307118 , n307119 , n16692 , n307121 , n307122 , n16695 , 
 n307124 , n307125 , n16698 , n307127 , n307128 , n16701 , n16702 , n307131 , n16704 , n307133 , 
 n307134 , n16707 , n16708 , n307137 , n16710 , n16711 , n16712 , n307141 , n16714 , n307143 , 
 n16716 , n16717 , n16718 , n16719 , n16720 , n307149 , n307150 , n307151 , n307152 , n307153 , 
 n16726 , n307155 , n307156 , n307157 , n307158 , n16731 , n307160 , n307161 , n307162 , n16735 , 
 n16736 , n307165 , n307166 , n16739 , n307168 , n16741 , n307170 , n307171 , n16744 , n307173 , 
 n307174 , n16747 , n307176 , n307177 , n307178 , n307179 , n307180 , n16753 , n307182 , n307183 , 
 n16756 , n307185 , n307186 , n307187 , n307188 , n307189 , n16762 , n307191 , n307192 , n16765 , 
 n307194 , n307195 , n16768 , n16769 , n307198 , n16771 , n307200 , n307201 , n16774 , n307203 , 
 n307204 , n16777 , n307206 , n307207 , n16780 , n307209 , n307210 , n16783 , n307212 , n307213 , 
 n16786 , n307215 , n307216 , n307217 , n307218 , n307219 , n16792 , n16793 , n16794 , n307223 , 
 n307224 , n16797 , n16798 , n16799 , n307228 , n307229 , n307230 , n16803 , n16804 , n307233 , 
 n16806 , n307235 , n307236 , n307237 , n307238 , n16811 , n16812 , n16813 , n307242 , n307243 , 
 n16816 , n307245 , n16818 , n307247 , n16820 , n307249 , n307250 , n16823 , n307252 , n307253 , 
 n16826 , n307255 , n16828 , n16829 , n307258 , n16831 , n307260 , n307261 , n307262 , n307263 , 
 n307264 , n16837 , n307266 , n307267 , n16840 , n307269 , n307270 , n16843 , n307272 , n307273 , 
 n307274 , n307275 , n307276 , n307277 , n307278 , n307279 , n16852 , n16853 , n16854 , n16855 , 
 n16856 , n16857 , n16858 , n307287 , n16860 , n307289 , n307290 , n307291 , n16864 , n307293 , 
 n307294 , n307295 , n307296 , n307297 , n307298 , n16871 , n16872 , n307301 , n307302 , n307303 , 
 n16876 , n307305 , n307306 , n307307 , n307308 , n307309 , n307310 , n307311 , n307312 , n307313 , 
 n307314 , n307315 , n307316 , n16889 , n16890 , n307319 , n307320 , n16893 , n307322 , n307323 , 
 n16896 , n307325 , n307326 , n307327 , n307328 , n307329 , n307330 , n307331 , n307332 , n307333 , 
 n307334 , n307335 , n307336 , n307337 , n307338 , n16911 , n307340 , n16913 , n16914 , n16915 , 
 n307344 , n16917 , n16918 , n307347 , n307348 , n307349 , n307350 , n307351 , n307352 , n307353 , 
 n16926 , n307355 , n307356 , n307357 , n307358 , n307359 , n307360 , n307361 , n307362 , n16935 , 
 n307364 , n307365 , n307366 , n307367 , n307368 , n16941 , n307370 , n16943 , n307372 , n16945 , 
 n16946 , n307375 , n16948 , n307377 , n16950 , n307379 , n16952 , n16953 , n307382 , n307383 , 
 n307384 , n307385 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n307392 , n307393 , 
 n16966 , n307395 , n307396 , n307397 , n307398 , n307399 , n307400 , n307401 , n307402 , n307403 , 
 n307404 , n307405 , n307406 , n16979 , n307408 , n16981 , n307410 , n307411 , n16984 , n307413 , 
 n307414 , n16987 , n307416 , n307417 , n16990 , n16991 , n16992 , n307421 , n307422 , n16995 , 
 n307424 , n307425 , n16998 , n307427 , n307428 , n17001 , n307430 , n17003 , n17004 , n307433 , 
 n17006 , n307435 , n307436 , n307437 , n307438 , n17011 , n307440 , n307441 , n17014 , n307443 , 
 n17016 , n307445 , n307446 , n307447 , n307448 , n17021 , n17022 , n307451 , n17024 , n307453 , 
 n307454 , n17027 , n307456 , n17029 , n307458 , n307459 , n17032 , n17033 , n307462 , n17035 , 
 n17036 , n307465 , n307466 , n17039 , n307468 , n307469 , n307470 , n17043 , n307472 , n17045 , 
 n17046 , n307475 , n307476 , n17049 , n307478 , n307479 , n17052 , n307481 , n307482 , n307483 , 
 n17056 , n307485 , n307486 , n17059 , n307488 , n17061 , n17062 , n307491 , n307492 , n17065 , 
 n307494 , n307495 , n17068 , n307497 , n17070 , n17071 , n307500 , n307501 , n17074 , n307503 , 
 n307504 , n17077 , n307506 , n17079 , n17080 , n307509 , n307510 , n17083 , n307512 , n307513 , 
 n17086 , n307515 , n17088 , n17089 , n17090 , n17091 , n307520 , n307521 , n17094 , n307523 , 
 n307524 , n17097 , n307526 , n17099 , n17100 , n307529 , n307530 , n17103 , n307532 , n307533 , 
 n17106 , n307535 , n307536 , n307537 , n307538 , n17111 , n307540 , n307541 , n17114 , n307543 , 
 n17116 , n17117 , n307546 , n307547 , n17120 , n307549 , n307550 , n17123 , n307552 , n307553 , 
 n17126 , n17127 , n307556 , n17129 , n307558 , n17131 , n17132 , n307561 , n307562 , n307563 , 
 n17136 , n307565 , n307566 , n17139 , n307568 , n307569 , n17142 , n307571 , n307572 , n307573 , 
 n17146 , n17147 , n307576 , n17149 , n17150 , n307579 , n307580 , n17153 , n307582 , n307583 , 
 n307584 , n307585 , n307586 , n307587 , n307588 , n17161 , n307590 , n17163 , n17164 , n307593 , 
 n17166 , n17167 , n307596 , n307597 , n307598 , n307599 , n307600 , n17173 , n307602 , n307603 , 
 n17176 , n307605 , n17178 , n17179 , n307608 , n307609 , n307610 , n17183 , n307612 , n307613 , 
 n17186 , n307615 , n307616 , n17189 , n307618 , n307619 , n17192 , n17193 , n17194 , n307623 , 
 n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n307630 , n307631 , n17204 , n17205 , 
 n17206 , n307635 , n307636 , n17209 , n17210 , n307639 , n307640 , n307641 , n307642 , n307643 , 
 n307644 , n17217 , n307646 , n307647 , n307648 , n307649 , n307650 , n17223 , n17224 , n307653 , 
 n307654 , n307655 , n307656 , n307657 , n307658 , n307659 , n307660 , n307661 , n307662 , n17235 , 
 n307664 , n17237 , n17238 , n307667 , n17240 , n307669 , n17242 , n307671 , n307672 , n17245 , 
 n307674 , n307675 , n17248 , n307677 , n307678 , n17251 , n17252 , n17253 , n307682 , n307683 , 
 n17256 , n307685 , n307686 , n17259 , n307688 , n307689 , n307690 , n17263 , n307692 , n17265 , 
 n17266 , n307695 , n307696 , n307697 , n17270 , n307699 , n307700 , n17273 , n307702 , n307703 , 
 n17276 , n17277 , n307706 , n17279 , n307708 , n17281 , n307710 , n17283 , n17284 , n307713 , 
 n17286 , n307715 , n17288 , n307717 , n307718 , n17291 , n307720 , n307721 , n17294 , n307723 , 
 n17296 , n307725 , n17298 , n17299 , n17300 , n307729 , n307730 , n17303 , n17304 , n307733 , 
 n307734 , n17307 , n307736 , n17309 , n307738 , n17311 , n17312 , n307741 , n17314 , n307743 , 
 n17316 , n307745 , n307746 , n17319 , n307748 , n307749 , n307750 , n17323 , n307752 , n17325 , 
 n17326 , n307755 , n307756 , n17329 , n307758 , n307759 , n17332 , n307761 , n307762 , n17335 , 
 n17336 , n17337 , n17338 , n17339 , n17340 , n307769 , n17342 , n17343 , n307772 , n307773 , 
 n17346 , n307775 , n17348 , n307777 , n17350 , n17351 , n307780 , n307781 , n17354 , n307783 , 
 n307784 , n17357 , n307786 , n307787 , n17360 , n307789 , n307790 , n17363 , n307792 , n307793 , 
 n17366 , n307795 , n307796 , n17369 , n307798 , n307799 , n307800 , n17373 , n307802 , n17375 , 
 n17376 , n307805 , n307806 , n17379 , n307808 , n307809 , n17382 , n307811 , n307812 , n17385 , 
 n307814 , n17387 , n307816 , n17389 , n17390 , n307819 , n307820 , n17393 , n307822 , n307823 , 
 n17396 , n307825 , n307826 , n17399 , n17400 , n17401 , n307830 , n307831 , n17404 , n17405 , 
 n17406 , n307835 , n307836 , n17409 , n17410 , n17411 , n307840 , n307841 , n17414 , n307843 , 
 n307844 , n17417 , n17418 , n17419 , n307848 , n307849 , n17422 , n17423 , n307852 , n307853 , 
 n17426 , n17427 , n307856 , n307857 , n17430 , n17431 , n307860 , n17433 , n17434 , n307863 , 
 n307864 , n17437 , n17438 , n17439 , n307868 , n307869 , n17442 , n17443 , n17444 , n17445 , 
 n17446 , n17447 , n17448 , n307877 , n17450 , n17451 , n17452 , n307881 , n307882 , n17455 , 
 n17456 , n17457 , n307886 , n307887 , n17460 , n307889 , n307890 , n307891 , n17464 , n307893 , 
 n17466 , n17467 , n307896 , n307897 , n17470 , n307899 , n307900 , n17473 , n307902 , n307903 , 
 n307904 , n17477 , n307906 , n17479 , n17480 , n307909 , n307910 , n17483 , n307912 , n307913 , 
 n17486 , n307915 , n307916 , n17489 , n307918 , n307919 , n307920 , n307921 , n17494 , n17495 , 
 n17496 , n307925 , n307926 , n17499 , n17500 , n17501 , n307930 , n17503 , n17504 , n17505 , 
 n17506 , n307935 , n307936 , n307937 , n307938 , n17511 , n17512 , n307941 , n307942 , n307943 , 
 n17516 , n307945 , n307946 , n17519 , n17520 , n307949 , n307950 , n307951 , n307952 , n17525 , 
 n307954 , n307955 , n17528 , n17529 , n17530 , n307959 , n307960 , n17533 , n17534 , n307963 , 
 n307964 , n17537 , n17538 , n307967 , n307968 , n307969 , n17542 , n307971 , n307972 , n17545 , 
 n17546 , n17547 , n307976 , n307977 , n17550 , n17551 , n307980 , n307981 , n307982 , n17555 , 
 n17556 , n307985 , n307986 , n17559 , n307988 , n307989 , n17562 , n307991 , n307992 , n307993 , 
 n307994 , n17567 , n17568 , n17569 , n307998 , n307999 , n17572 , n17573 , n17574 , n308003 , 
 n308004 , n17577 , n17578 , n17579 , n308008 , n308009 , n17582 , n17583 , n17584 , n308013 , 
 n308014 , n17587 , n17588 , n17589 , n308018 , n308019 , n17592 , n308021 , n308022 , n17595 , 
 n308024 , n308025 , n17598 , n17599 , n308028 , n308029 , n17602 , n17603 , n308032 , n308033 , 
 n17606 , n17607 , n17608 , n17609 , n308038 , n308039 , n17612 , n17613 , n308042 , n308043 , 
 n17616 , n17617 , n17618 , n17619 , n17620 , n308049 , n308050 , n17623 , n17624 , n308053 , 
 n308054 , n308055 , n17628 , n17629 , n17630 , n308059 , n308060 , n17633 , n17634 , n17635 , 
 n308064 , n308065 , n308066 , n308067 , n308068 , n17641 , n308070 , n308071 , n308072 , n308073 , 
 n308074 , n308075 , n17648 , n308077 , n308078 , n17651 , n308080 , n308081 , n308082 , n17655 , 
 n308084 , n308085 , n308086 , n308087 , n308088 , n17661 , n308090 , n308091 , n308092 , n308093 , 
 n308094 , n17667 , n17668 , n308097 , n308098 , n308099 , n308100 , n308101 , n308102 , n17675 , 
 n308104 , n308105 , n17678 , n17679 , n17680 , n17681 , n308110 , n308111 , n308112 , n308113 , 
 n308114 , n308115 , n17688 , n17689 , n17690 , n308119 , n308120 , n308121 , n308122 , n308123 , 
 n308124 , n17697 , n308126 , n308127 , n17700 , n17701 , n308130 , n308131 , n308132 , n308133 , 
 n308134 , n308135 , n308136 , n17709 , n308138 , n17711 , n308140 , n308141 , n308142 , n17715 , 
 n308144 , n308145 , n308146 , n308147 , n308148 , n308149 , n17722 , n308151 , n308152 , n17725 , 
 n308154 , n308155 , n308156 , n308157 , n308158 , n308159 , n308160 , n308161 , n308162 , n308163 , 
 n308164 , n17737 , n308166 , n17739 , n308168 , n308169 , n308170 , n17743 , n308172 , n17745 , 
 n17746 , n308175 , n308176 , n308177 , n308178 , n308179 , n17752 , n308181 , n308182 , n308183 , 
 n308184 , n308185 , n308186 , n17759 , n308188 , n308189 , n17762 , n308191 , n308192 , n308193 , 
 n308194 , n308195 , n308196 , n308197 , n308198 , n308199 , n308200 , n308201 , n308202 , n308203 , 
 n308204 , n308205 , n308206 , n308207 , n308208 , n308209 , n308210 , n308211 , n308212 , n308213 , 
 n308214 , n308215 , n17788 , n17789 , n17790 , n17791 , n308220 , n308221 , n17794 , n308223 , 
 n17796 , n308225 , n308226 , n308227 , n308228 , n308229 , n308230 , n308231 , n308232 , n17805 , 
 n308234 , n308235 , n308236 , n17809 , n308238 , n308239 , n308240 , n308241 , n308242 , n308243 , 
 n308244 , n308245 , n308246 , n308247 , n308248 , n17821 , n308250 , n308251 , n308252 , n308253 , 
 n308254 , n308255 , n17828 , n308257 , n308258 , n17831 , n308260 , n17833 , n308262 , n17835 , 
 n308264 , n308265 , n308266 , n308267 , n308268 , n17841 , n308270 , n308271 , n308272 , n308273 , 
 n308274 , n308275 , n17848 , n308277 , n308278 , n308279 , n308280 , n308281 , n308282 , n308283 , 
 n308284 , n308285 , n308286 , n308287 , n308288 , n308289 , n308290 , n17863 , n308292 , n17865 , 
 n308294 , n308295 , n308296 , n308297 , n308298 , n308299 , n308300 , n308301 , n308302 , n308303 , 
 n308304 , n308305 , n308306 , n308307 , n308308 , n308309 , n308310 , n17883 , n308312 , n308313 , 
 n308314 , n308315 , n17888 , n308317 , n308318 , n308319 , n308320 , n308321 , n308322 , n308323 , 
 n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n308330 , n17903 , n17904 , n308333 , 
 n308334 , n17907 , n17908 , n308337 , n308338 , n308339 , n17912 , n308341 , n308342 , n308343 , 
 n308344 , n308345 , n308346 , n308347 , n17920 , n308349 , n308350 , n17923 , n308352 , n308353 , 
 n17926 , n308355 , n308356 , n17929 , n308358 , n308359 , n17932 , n17933 , n308362 , n17935 , 
 n17936 , n17937 , n308366 , n308367 , n308368 , n308369 , n17942 , n17943 , n308372 , n308373 , 
 n17946 , n17947 , n308376 , n308377 , n17950 , n308379 , n308380 , n308381 , n308382 , n308383 , 
 n308384 , n17957 , n308386 , n17959 , n17960 , n308389 , n308390 , n308391 , n308392 , n17965 , 
 n308394 , n17967 , n308396 , n17969 , n17970 , n308399 , n308400 , n308401 , n17974 , n308403 , 
 n308404 , n308405 , n308406 , n308407 , n308408 , n308409 , n308410 , n308411 , n308412 , n308413 , 
 n17986 , n308415 , n17988 , n308417 , n17990 , n308419 , n308420 , n308421 , n17994 , n17995 , 
 n308424 , n308425 , n17998 , n308427 , n308428 , n308429 , n308430 , n308431 , n308432 , n18005 , 
 n308434 , n18007 , n18008 , n308437 , n308438 , n308439 , n18012 , n308441 , n308442 , n18015 , 
 n308444 , n308445 , n18018 , n308447 , n18020 , n18021 , n308450 , n18023 , n308452 , n18025 , 
 n18026 , n308455 , n308456 , n308457 , n18030 , n308459 , n308460 , n18033 , n308462 , n308463 , 
 n18036 , n308465 , n308466 , n18039 , n308468 , n308469 , n18042 , n308471 , n308472 , n18045 , 
 n308474 , n308475 , n308476 , n18049 , n18050 , n18051 , n308480 , n308481 , n308482 , n308483 , 
 n18056 , n308485 , n308486 , n308487 , n18060 , n308489 , n18062 , n308491 , n308492 , n18065 , 
 n308494 , n308495 , n18068 , n308497 , n308498 , n308499 , n308500 , n308501 , n308502 , n308503 , 
 n308504 , n18077 , n18078 , n18079 , n308508 , n308509 , n308510 , n308511 , n308512 , n18085 , 
 n18086 , n18087 , n18088 , n308517 , n308518 , n18091 , n18092 , n308521 , n308522 , n18095 , 
 n308524 , n308525 , n308526 , n308527 , n308528 , n18101 , n308530 , n308531 , n308532 , n308533 , 
 n308534 , n308535 , n308536 , n18109 , n18110 , n308539 , n308540 , n308541 , n308542 , n308543 , 
 n308544 , n308545 , n18118 , n308547 , n308548 , n308549 , n308550 , n308551 , n308552 , n308553 , 
 n308554 , n308555 , n308556 , n308557 , n308558 , n308559 , n308560 , n308561 , n308562 , n18135 , 
 n308564 , n18137 , n308566 , n308567 , n308568 , n308569 , n308570 , n308571 , n308572 , n308573 , 
 n308574 , n308575 , n308576 , n308577 , n308578 , n308579 , n18152 , n308581 , n18154 , n308583 , 
 n18156 , n18157 , n308586 , n308587 , n308588 , n18161 , n308590 , n308591 , n308592 , n308593 , 
 n308594 , n308595 , n18168 , n308597 , n308598 , n18171 , n18172 , n308601 , n308602 , n308603 , 
 n308604 , n308605 , n308606 , n308607 , n308608 , n308609 , n308610 , n18183 , n308612 , n308613 , 
 n18186 , n308615 , n308616 , n308617 , n308618 , n308619 , n308620 , n308621 , n308622 , n308623 , 
 n308624 , n308625 , n308626 , n308627 , n308628 , n308629 , n18202 , n308631 , n308632 , n18205 , 
 n308634 , n308635 , n18208 , n308637 , n308638 , n18211 , n308640 , n308641 , n18214 , n308643 , 
 n308644 , n18217 , n308646 , n18219 , n18220 , n308649 , n308650 , n18223 , n18224 , n18225 , 
 n18226 , n308655 , n308656 , n18229 , n18230 , n18231 , n18232 , n308661 , n308662 , n18235 , 
 n308664 , n18237 , n308666 , n18239 , n18240 , n308669 , n308670 , n308671 , n18244 , n308673 , 
 n308674 , n18247 , n308676 , n308677 , n18250 , n308679 , n308680 , n18253 , n308682 , n18255 , 
 n18256 , n308685 , n308686 , n18259 , n308688 , n308689 , n18262 , n308691 , n308692 , n308693 , 
 n18266 , n308695 , n18268 , n308697 , n18270 , n308699 , n308700 , n308701 , n308702 , n308703 , 
 n308704 , n308705 , n308706 , n18279 , n18280 , n308709 , n308710 , n308711 , n308712 , n308713 , 
 n308714 , n308715 , n308716 , n308717 , n308718 , n308719 , n18292 , n308721 , n18294 , n308723 , 
 n308724 , n308725 , n308726 , n308727 , n308728 , n308729 , n308730 , n308731 , n308732 , n308733 , 
 n308734 , n308735 , n308736 , n308737 , n18310 , n308739 , n18312 , n308741 , n308742 , n308743 , 
 n308744 , n308745 , n308746 , n308747 , n308748 , n308749 , n308750 , n308751 , n308752 , n308753 , 
 n308754 , n308755 , n18328 , n308757 , n18330 , n308759 , n308760 , n18333 , n308762 , n18335 , 
 n308764 , n308765 , n308766 , n308767 , n308768 , n308769 , n308770 , n18343 , n308772 , n18345 , 
 n308774 , n308775 , n308776 , n308777 , n18350 , n308779 , n308780 , n18353 , n18354 , n18355 , 
 n308784 , n308785 , n18358 , n18359 , n308788 , n18361 , n18362 , n18363 , n308792 , n18365 , 
 n18366 , n308795 , n308796 , n308797 , n308798 , n18371 , n308800 , n308801 , n18374 , n308803 , 
 n308804 , n308805 , n308806 , n308807 , n18380 , n308809 , n308810 , n308811 , n308812 , n18385 , 
 n308814 , n18387 , n18388 , n308817 , n308818 , n18391 , n308820 , n308821 , n18394 , n308823 , 
 n18396 , n308825 , n308826 , n308827 , n308828 , n308829 , n308830 , n308831 , n308832 , n18405 , 
 n308834 , n308835 , n308836 , n308837 , n308838 , n308839 , n308840 , n18413 , n308842 , n308843 , 
 n18416 , n18417 , n308846 , n18419 , n18420 , n308849 , n18422 , n308851 , n18424 , n18425 , 
 n18426 , n308855 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , 
 n308864 , n18437 , n308866 , n308867 , n18440 , n308869 , n308870 , n308871 , n308872 , n18445 , 
 n308874 , n308875 , n18448 , n18449 , n308878 , n18451 , n308880 , n308881 , n308882 , n18455 , 
 n308884 , n308885 , n308886 , n18459 , n308888 , n308889 , n18462 , n308891 , n18464 , n18465 , 
 n308894 , n18467 , n308896 , n308897 , n308898 , n308899 , n308900 , n18473 , n308902 , n308903 , 
 n308904 , n308905 , n308906 , n308907 , n18480 , n18481 , n308910 , n308911 , n308912 , n308913 , 
 n308914 , n18487 , n308916 , n18489 , n308918 , n18491 , n18492 , n18493 , n18494 , n18495 , 
 n308924 , n18497 , n18498 , n308927 , n18500 , n308929 , n18502 , n308931 , n18504 , n308933 , 
 n308934 , n308935 , n18508 , n18509 , n308938 , n18511 , n308940 , n308941 , n308942 , n308943 , 
 n18516 , n18517 , n308946 , n18519 , n308948 , n308949 , n308950 , n308951 , n308952 , n308953 , 
 n308954 , n308955 , n308956 , n308957 , n18530 , n308959 , n308960 , n308961 , n18534 , n308963 , 
 n308964 , n308965 , n308966 , n18539 , n308968 , n18541 , n308970 , n308971 , n308972 , n308973 , 
 n308974 , n308975 , n308976 , n18549 , n308978 , n308979 , n18552 , n308981 , n308982 , n18555 , 
 n18556 , n18557 , n18558 , n308987 , n308988 , n308989 , n308990 , n18563 , n308992 , n308993 , 
 n308994 , n308995 , n308996 , n308997 , n308998 , n308999 , n309000 , n309001 , n309002 , n18575 , 
 n309004 , n309005 , n18578 , n309007 , n309008 , n309009 , n309010 , n309011 , n18584 , n18585 , 
 n18586 , n309015 , n309016 , n309017 , n309018 , n309019 , n309020 , n309021 , n309022 , n18595 , 
 n309024 , n18597 , n18598 , n309027 , n309028 , n18601 , n18602 , n309031 , n18604 , n309033 , 
 n309034 , n309035 , n309036 , n18609 , n309038 , n18611 , n309040 , n309041 , n309042 , n309043 , 
 n309044 , n309045 , n309046 , n309047 , n18620 , n309049 , n309050 , n309051 , n309052 , n309053 , 
 n309054 , n309055 , n18628 , n309057 , n18630 , n309059 , n309060 , n309061 , n309062 , n309063 , 
 n18636 , n309065 , n309066 , n309067 , n309068 , n309069 , n18642 , n309071 , n18644 , n309073 , 
 n309074 , n309075 , n309076 , n18649 , n18650 , n309079 , n18652 , n18653 , n309082 , n18655 , 
 n309084 , n18657 , n18658 , n309087 , n309088 , n309089 , n309090 , n309091 , n18664 , n18665 , 
 n309094 , n309095 , n18668 , n18669 , n309098 , n309099 , n18672 , n18673 , n309102 , n309103 , 
 n18676 , n309105 , n309106 , n309107 , n309108 , n309109 , n18682 , n309111 , n18684 , n18685 , 
 n309114 , n309115 , n18688 , n18689 , n309118 , n18691 , n309120 , n18693 , n309122 , n309123 , 
 n18696 , n309125 , n309126 , n18699 , n309128 , n309129 , n309130 , n309131 , n309132 , n18705 , 
 n309134 , n309135 , n309136 , n309137 , n309138 , n309139 , n309140 , n309141 , n309142 , n309143 , 
 n309144 , n309145 , n309146 , n309147 , n18720 , n309149 , n309150 , n18723 , n309152 , n309153 , 
 n18726 , n309155 , n309156 , n18729 , n309158 , n18731 , n309160 , n309161 , n309162 , n309163 , 
 n309164 , n309165 , n309166 , n309167 , n18740 , n309169 , n309170 , n18743 , n309172 , n309173 , 
 n18746 , n309175 , n309176 , n18749 , n309178 , n309179 , n18752 , n309181 , n309182 , n309183 , 
 n309184 , n309185 , n18758 , n309187 , n309188 , n309189 , n18762 , n309191 , n18764 , n309193 , 
 n309194 , n309195 , n18768 , n309197 , n309198 , n18771 , n309200 , n18773 , n18774 , n309203 , 
 n309204 , n18777 , n309206 , n18779 , n309208 , n309209 , n18782 , n309211 , n309212 , n309213 , 
 n309214 , n309215 , n309216 , n18789 , n309218 , n18791 , n18792 , n18793 , n18794 , n309223 , 
 n18796 , n18797 , n309226 , n309227 , n309228 , n18801 , n18802 , n309231 , n309232 , n309233 , 
 n18806 , n309235 , n309236 , n18809 , n309238 , n309239 , n309240 , n18813 , n309242 , n309243 , 
 n309244 , n18817 , n309246 , n18819 , n309248 , n309249 , n309250 , n309251 , n309252 , n309253 , 
 n309254 , n309255 , n18828 , n18829 , n18830 , n309259 , n18832 , n18833 , n309262 , n309263 , 
 n309264 , n309265 , n309266 , n309267 , n309268 , n309269 , n18842 , n309271 , n309272 , n18845 , 
 n18846 , n309275 , n18848 , n18849 , n309278 , n309279 , n18852 , n309281 , n18854 , n309283 , 
 n309284 , n18857 , n309286 , n309287 , n18860 , n309289 , n309290 , n309291 , n309292 , n309293 , 
 n18866 , n309295 , n309296 , n309297 , n309298 , n309299 , n309300 , n309301 , n309302 , n309303 , 
 n18876 , n309305 , n309306 , n309307 , n18880 , n309309 , n309310 , n18883 , n309312 , n309313 , 
 n18886 , n309315 , n309316 , n18889 , n309318 , n309319 , n18892 , n309321 , n309322 , n309323 , 
 n309324 , n18897 , n309326 , n18899 , n309328 , n309329 , n309330 , n309331 , n309332 , n309333 , 
 n309334 , n309335 , n309336 , n309337 , n309338 , n18911 , n18912 , n309341 , n309342 , n309343 , 
 n309344 , n18917 , n309346 , n18919 , n309348 , n309349 , n309350 , n18923 , n309352 , n309353 , 
 n309354 , n309355 , n309356 , n309357 , n18930 , n309359 , n309360 , n309361 , n18934 , n309363 , 
 n309364 , n18937 , n309366 , n309367 , n18940 , n309369 , n309370 , n18943 , n309372 , n309373 , 
 n309374 , n309375 , n18948 , n309377 , n309378 , n18951 , n309380 , n309381 , n18954 , n309383 , 
 n309384 , n309385 , n309386 , n18959 , n309388 , n309389 , n309390 , n309391 , n18964 , n309393 , 
 n18966 , n18967 , n309396 , n309397 , n18970 , n18971 , n18972 , n309401 , n18974 , n309403 , 
 n309404 , n309405 , n309406 , n309407 , n309408 , n18981 , n309410 , n309411 , n309412 , n309413 , 
 n309414 , n309415 , n309416 , n309417 , n309418 , n309419 , n309420 , n309421 , n18994 , n309423 , 
 n309424 , n18997 , n309426 , n309427 , n19000 , n309429 , n309430 , n309431 , n19004 , n309433 , 
 n309434 , n19007 , n19008 , n309437 , n309438 , n19011 , n19012 , n309441 , n309442 , n19015 , 
 n309444 , n309445 , n309446 , n309447 , n19020 , n309449 , n309450 , n19023 , n309452 , n309453 , 
 n309454 , n309455 , n309456 , n19029 , n309458 , n309459 , n19032 , n309461 , n309462 , n309463 , 
 n309464 , n19037 , n309466 , n309467 , n309468 , n309469 , n309470 , n19043 , n19044 , n309473 , 
 n309474 , n309475 , n19048 , n309477 , n309478 , n309479 , n309480 , n309481 , n309482 , n309483 , 
 n309484 , n309485 , n309486 , n19059 , n309488 , n309489 , n309490 , n309491 , n19064 , n309493 , 
 n309494 , n19067 , n19068 , n19069 , n19070 , n309499 , n309500 , n19073 , n19074 , n19075 , 
 n19076 , n19077 , n309506 , n309507 , n19080 , n19081 , n19082 , n309511 , n19084 , n309513 , 
 n309514 , n309515 , n309516 , n19089 , n309518 , n309519 , n19092 , n309521 , n309522 , n19095 , 
 n309524 , n19097 , n19098 , n309527 , n309528 , n19101 , n309530 , n309531 , n19104 , n309533 , 
 n19106 , n19107 , n19108 , n309537 , n19110 , n309539 , n309540 , n309541 , n19114 , n309543 , 
 n19116 , n309545 , n309546 , n309547 , n309548 , n19121 , n309550 , n309551 , n19124 , n309553 , 
 n309554 , n309555 , n19128 , n309557 , n19130 , n309559 , n309560 , n19133 , n309562 , n309563 , 
 n309564 , n309565 , n19138 , n309567 , n309568 , n19141 , n309570 , n309571 , n19144 , n309573 , 
 n19146 , n309575 , n309576 , n19149 , n309578 , n309579 , n309580 , n309581 , n309582 , n309583 , 
 n19156 , n309585 , n309586 , n309587 , n309588 , n19161 , n309590 , n309591 , n19164 , n309593 , 
 n309594 , n19167 , n309596 , n309597 , n309598 , n309599 , n309600 , n19173 , n309602 , n309603 , 
 n309604 , n309605 , n309606 , n309607 , n309608 , n309609 , n309610 , n19183 , n19184 , n309613 , 
 n19186 , n309615 , n309616 , n19189 , n309618 , n309619 , n19192 , n309621 , n19194 , n19195 , 
 n309624 , n309625 , n19198 , n309627 , n309628 , n19201 , n309630 , n19203 , n309632 , n19205 , 
 n309634 , n19207 , n309636 , n19209 , n309638 , n309639 , n309640 , n19213 , n309642 , n309643 , 
 n309644 , n19217 , n309646 , n309647 , n19220 , n309649 , n309650 , n19223 , n309652 , n309653 , 
 n309654 , n309655 , n309656 , n309657 , n309658 , n309659 , n309660 , n19233 , n309662 , n309663 , 
 n309664 , n309665 , n309666 , n19239 , n309668 , n309669 , n309670 , n309671 , n309672 , n309673 , 
 n309674 , n19247 , n309676 , n309677 , n19250 , n309679 , n309680 , n309681 , n19254 , n309683 , 
 n309684 , n309685 , n309686 , n309687 , n309688 , n19261 , n19262 , n309691 , n309692 , n309693 , 
 n309694 , n309695 , n309696 , n19269 , n309698 , n309699 , n19272 , n309701 , n309702 , n19275 , 
 n309704 , n19277 , n309706 , n309707 , n19280 , n309709 , n19282 , n309711 , n309712 , n309713 , 
 n19286 , n309715 , n19288 , n19289 , n309718 , n309719 , n19292 , n309721 , n19294 , n309723 , 
 n309724 , n19297 , n309726 , n309727 , n309728 , n19301 , n309730 , n19303 , n19304 , n309733 , 
 n19306 , n19307 , n19308 , n19309 , n309738 , n309739 , n309740 , n309741 , n309742 , n309743 , 
 n309744 , n19317 , n309746 , n19319 , n19320 , n309749 , n19322 , n19323 , n19324 , n309753 , 
 n309754 , n19327 , n309756 , n309757 , n19330 , n309759 , n19332 , n19333 , n309762 , n309763 , 
 n309764 , n309765 , n309766 , n309767 , n19340 , n309769 , n309770 , n19343 , n19344 , n19345 , 
 n309774 , n309775 , n19348 , n309777 , n19350 , n309779 , n19352 , n19353 , n309782 , n309783 , 
 n309784 , n19357 , n309786 , n309787 , n19360 , n309789 , n309790 , n19363 , n309792 , n309793 , 
 n309794 , n309795 , n19368 , n309797 , n19370 , n309799 , n309800 , n19373 , n309802 , n19375 , 
 n309804 , n19377 , n19378 , n309807 , n309808 , n309809 , n19382 , n309811 , n309812 , n19385 , 
 n309814 , n309815 , n19388 , n309817 , n309818 , n19391 , n19392 , n19393 , n309822 , n309823 , 
 n19396 , n309825 , n309826 , n19399 , n309828 , n309829 , n309830 , n309831 , n19404 , n309833 , 
 n309834 , n309835 , n19408 , n309837 , n19410 , n19411 , n309840 , n19413 , n309842 , n19415 , 
 n309844 , n309845 , n19418 , n309847 , n309848 , n19421 , n309850 , n19423 , n309852 , n19425 , 
 n19426 , n309855 , n19428 , n309857 , n19430 , n309859 , n309860 , n19433 , n309862 , n309863 , 
 n19436 , n309865 , n309866 , n309867 , n19440 , n309869 , n19442 , n19443 , n309872 , n309873 , 
 n309874 , n19447 , n309876 , n309877 , n19450 , n309879 , n309880 , n19453 , n309882 , n309883 , 
 n309884 , n19457 , n309886 , n19459 , n19460 , n19461 , n309890 , n309891 , n309892 , n19465 , 
 n309894 , n309895 , n19468 , n309897 , n309898 , n19471 , n309900 , n309901 , n19474 , n309903 , 
 n19476 , n309905 , n19478 , n309907 , n309908 , n19481 , n19482 , n309911 , n309912 , n19485 , 
 n309914 , n309915 , n19488 , n309917 , n309918 , n19491 , n309920 , n309921 , n19494 , n309923 , 
 n309924 , n19497 , n309926 , n19499 , n309928 , n19501 , n19502 , n309931 , n19504 , n309933 , 
 n19506 , n309935 , n309936 , n19509 , n309938 , n309939 , n309940 , n19513 , n309942 , n19515 , 
 n19516 , n309945 , n19518 , n309947 , n19520 , n309949 , n309950 , n309951 , n309952 , n19525 , 
 n19526 , n309955 , n19528 , n309957 , n19530 , n309959 , n19532 , n309961 , n309962 , n309963 , 
 n309964 , n309965 , n19538 , n309967 , n309968 , n309969 , n309970 , n309971 , n309972 , n309973 , 
 n19546 , n309975 , n19548 , n309977 , n309978 , n19551 , n309980 , n309981 , n309982 , n19555 , 
 n19556 , n19557 , n309986 , n309987 , n19560 , n309989 , n19562 , n309991 , n309992 , n309993 , 
 n309994 , n309995 , n309996 , n19569 , n19570 , n19571 , n310000 , n19573 , n19574 , n310003 , 
 n19576 , n310005 , n310006 , n19579 , n310008 , n19581 , n19582 , n310011 , n310012 , n19585 , 
 n310014 , n310015 , n19588 , n310017 , n19590 , n19591 , n19592 , n19593 , n310022 , n310023 , 
 n310024 , n310025 , n19598 , n19599 , n310028 , n310029 , n310030 , n310031 , n310032 , n310033 , 
 n310034 , n19607 , n19608 , n310037 , n310038 , n310039 , n310040 , n19613 , n19614 , n310043 , 
 n310044 , n310045 , n310046 , n310047 , n19620 , n310049 , n310050 , n310051 , n310052 , n310053 , 
 n19626 , n310055 , n310056 , n310057 , n310058 , n19631 , n310060 , n310061 , n19634 , n19635 , 
 n310064 , n310065 , n19638 , n310067 , n310068 , n19641 , n310070 , n310071 , n310072 , n310073 , 
 n310074 , n19647 , n310076 , n310077 , n19650 , n310079 , n310080 , n19653 , n310082 , n310083 , 
 n19656 , n310085 , n19658 , n19659 , n310088 , n310089 , n310090 , n310091 , n310092 , n19665 , 
 n310094 , n310095 , n19668 , n19669 , n310098 , n310099 , n310100 , n310101 , n310102 , n19675 , 
 n310104 , n310105 , n310106 , n19679 , n310108 , n310109 , n310110 , n19683 , n310112 , n310113 , 
 n19686 , n310115 , n310116 , n19689 , n310118 , n310119 , n310120 , n310121 , n310122 , n19695 , 
 n310124 , n310125 , n19698 , n310127 , n310128 , n19701 , n310130 , n310131 , n19704 , n310133 , 
 n19706 , n310135 , n310136 , n310137 , n19710 , n310139 , n310140 , n19713 , n310142 , n310143 , 
 n310144 , n310145 , n310146 , n310147 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , 
 n19726 , n310155 , n310156 , n19729 , n310158 , n310159 , n310160 , n310161 , n310162 , n19735 , 
 n310164 , n19737 , n310166 , n19739 , n19740 , n310169 , n19742 , n19743 , n310172 , n310173 , 
 n19746 , n310175 , n310176 , n310177 , n19750 , n310179 , n310180 , n310181 , n310182 , n310183 , 
 n19756 , n19757 , n310186 , n19759 , n310188 , n19761 , n19762 , n310191 , n310192 , n310193 , 
 n310194 , n19767 , n19768 , n310197 , n19770 , n19771 , n310200 , n19773 , n310202 , n310203 , 
 n310204 , n19777 , n19778 , n310207 , n310208 , n19781 , n19782 , n19783 , n310212 , n310213 , 
 n310214 , n310215 , n310216 , n310217 , n310218 , n310219 , n19792 , n310221 , n310222 , n19795 , 
 n19796 , n310225 , n310226 , n310227 , n310228 , n310229 , n19802 , n310231 , n19804 , n310233 , 
 n310234 , n310235 , n310236 , n310237 , n19810 , n310239 , n310240 , n310241 , n310242 , n19815 , 
 n19816 , n310245 , n310246 , n310247 , n310248 , n310249 , n19822 , n310251 , n19824 , n310253 , 
 n19826 , n19827 , n19828 , n310257 , n310258 , n310259 , n310260 , n310261 , n19834 , n310263 , 
 n19836 , n310265 , n19838 , n310267 , n19840 , n310269 , n19842 , n310271 , n310272 , n310273 , 
 n310274 , n310275 , n19848 , n310277 , n19850 , n310279 , n19852 , n19853 , n19854 , n310283 , 
 n310284 , n310285 , n19860 , n310287 , n19862 , n310289 , n310290 , n310291 , n310292 , n310293 , 
 n19868 , n310295 , n310296 , n310297 , n310298 , n310299 , n310300 , n310301 , n310302 , n310303 , 
 n310304 , n310305 , n310306 , n310307 , n310308 , n310309 , n310310 , n310311 , n310312 , n310313 , 
 n310314 , n310315 , n19890 , n310317 , n310318 , n310319 , n310320 , n310321 , n19896 , n310323 , 
 n310324 , n19899 , n310326 , n19901 , n310328 , n19903 , n310330 , n19905 , n19906 , n310333 , 
 n19908 , n310335 , n19910 , n310337 , n310338 , n19913 , n19914 , n310341 , n19916 , n310343 , 
 n310344 , n310345 , n310346 , n19921 , n310348 , n310349 , n310350 , n310351 , n310352 , n310353 , 
 n310354 , n310355 , n310356 , n310357 , n310358 , n310359 , n310360 , n310361 , n310362 , n310363 , 
 n310364 , n310365 , n310366 , n310367 , n310368 , n310369 , n19944 , n310371 , n310372 , n310373 , 
 n19948 , n310375 , n310376 , n310377 , n310378 , n310379 , n19954 , n19955 , n310382 , n310383 , 
 n310384 , n19959 , n310386 , n310387 , n19962 , n310389 , n310390 , n310391 , n310392 , n310393 , 
 n310394 , n310395 , n310396 , n310397 , n310398 , n310399 , n310400 , n310401 , n310402 , n310403 , 
 n310404 , n310405 , n310406 , n19981 , n19982 , n310409 , n19984 , n19985 , n19986 , n310413 , 
 n19988 , n310415 , n310416 , n310417 , n310418 , n310419 , n19994 , n310421 , n19996 , n19997 , 
 n19998 , n310425 , n20000 , n310427 , n310428 , n310429 , n310430 , n20005 , n310432 , n310433 , 
 n310434 , n310435 , n310436 , n20011 , n310438 , n310439 , n310440 , n310441 , n310442 , n20017 , 
 n310444 , n310445 , n310446 , n310447 , n310448 , n20023 , n310450 , n310451 , n310452 , n20027 , 
 n20028 , n310455 , n310456 , n20031 , n310458 , n310459 , n310460 , n310461 , n20036 , n310463 , 
 n310464 , n20039 , n310466 , n310467 , n20042 , n310469 , n310470 , n310471 , n310472 , n310473 , 
 n20048 , n310475 , n20050 , n310477 , n310478 , n20053 , n310480 , n310481 , n310482 , n310483 , 
 n310484 , n310485 , n310486 , n310487 , n310488 , n310489 , n20064 , n20065 , n310492 , n310493 , 
 n310494 , n310495 , n310496 , n310497 , n20072 , n310499 , n310500 , n20075 , n310502 , n310503 , 
 n310504 , n310505 , n310506 , n310507 , n310508 , n310509 , n310510 , n310511 , n310512 , n310513 , 
 n310514 , n310515 , n310516 , n20091 , n310518 , n310519 , n20094 , n310521 , n310522 , n310523 , 
 n310524 , n310525 , n310526 , n310527 , n310528 , n20103 , n310530 , n310531 , n310532 , n310533 , 
 n310534 , n310535 , n310536 , n310537 , n310538 , n310539 , n310540 , n310541 , n310542 , n310543 , 
 n310544 , n310545 , n310546 , n310547 , n310548 , n310549 , n310550 , n310551 , n310552 , n20127 , 
 n20128 , n310555 , n310556 , n310557 , n310558 , n20133 , n310560 , n310561 , n310562 , n20137 , 
 n20138 , n310565 , n310566 , n20141 , n310568 , n310569 , n310570 , n310571 , n20146 , n310573 , 
 n310574 , n20149 , n310576 , n310577 , n20152 , n20153 , n310580 , n20155 , n310582 , n20157 , 
 n310584 , n310585 , n310586 , n310587 , n310588 , n20163 , n310590 , n310591 , n20166 , n20167 , 
 n310594 , n20169 , n310596 , n310597 , n310598 , n310599 , n310600 , n310601 , n310602 , n20177 , 
 n310604 , n20179 , n310606 , n310607 , n310608 , n20183 , n310610 , n310611 , n310612 , n20187 , 
 n20188 , n310615 , n310616 , n310617 , n310618 , n310619 , n310620 , n310621 , n310622 , n310623 , 
 n20198 , n310625 , n20200 , n310627 , n310628 , n310629 , n310630 , n310631 , n310632 , n20207 , 
 n310634 , n310635 , n20210 , n310637 , n310638 , n310639 , n310640 , n20215 , n310642 , n20217 , 
 n310644 , n310645 , n310646 , n20221 , n310648 , n310649 , n20224 , n20225 , n310652 , n310653 , 
 n310654 , n310655 , n310656 , n310657 , n310658 , n310659 , n20234 , n20235 , n310662 , n20237 , 
 n20238 , n310665 , n310666 , n20241 , n310668 , n310669 , n20244 , n310671 , n310672 , n310673 , 
 n20248 , n310675 , n310676 , n310677 , n310678 , n310679 , n20254 , n20255 , n310682 , n20257 , 
 n20258 , n310685 , n310686 , n20261 , n310688 , n310689 , n20264 , n310691 , n310692 , n20267 , 
 n310694 , n310695 , n310696 , n20271 , n310698 , n310699 , n310700 , n310701 , n310702 , n310703 , 
 n310704 , n310705 , n310706 , n310707 , n310708 , n310709 , n310710 , n310711 , n310712 , n20287 , 
 n310714 , n310715 , n20290 , n310717 , n310718 , n20293 , n310720 , n310721 , n310722 , n310723 , 
 n310724 , n310725 , n310726 , n310727 , n310728 , n310729 , n20304 , n310731 , n310732 , n20307 , 
 n20308 , n310735 , n310736 , n310737 , n310738 , n310739 , n310740 , n310741 , n310742 , n310743 , 
 n20318 , n310745 , n310746 , n310747 , n310748 , n310749 , n310750 , n20325 , n20326 , n310753 , 
 n310754 , n310755 , n310756 , n310757 , n20332 , n310759 , n310760 , n20335 , n310762 , n20337 , 
 n310764 , n310765 , n310766 , n310767 , n20342 , n310769 , n310770 , n20345 , n20346 , n310773 , 
 n310774 , n310775 , n20350 , n310777 , n310778 , n20353 , n20354 , n310781 , n20356 , n20357 , 
 n310784 , n310785 , n20360 , n310787 , n310788 , n20363 , n310790 , n20365 , n310792 , n310793 , 
 n310794 , n310795 , n20370 , n310797 , n310798 , n20373 , n20374 , n20375 , n310802 , n310803 , 
 n310804 , n310805 , n310806 , n310807 , n310808 , n20383 , n310810 , n310811 , n20386 , n310813 , 
 n310814 , n310815 , n310816 , n310817 , n20392 , n310819 , n310820 , n310821 , n310822 , n20397 , 
 n310824 , n310825 , n310826 , n310827 , n310828 , n310829 , n20404 , n310831 , n310832 , n20407 , 
 n310834 , n310835 , n310836 , n20411 , n20412 , n310839 , n20414 , n310841 , n310842 , n310843 , 
 n310844 , n20419 , n20420 , n20421 , n20422 , n310849 , n310850 , n20425 , n310852 , n20427 , 
 n20428 , n310855 , n310856 , n310857 , n20432 , n310859 , n310860 , n20435 , n310862 , n310863 , 
 n310864 , n310865 , n310866 , n310867 , n310868 , n20443 , n310870 , n310871 , n310872 , n20447 , 
 n310874 , n20449 , n310876 , n310877 , n310878 , n310879 , n310880 , n20455 , n310882 , n310883 , 
 n20458 , n310885 , n310886 , n310887 , n310888 , n310889 , n310890 , n20465 , n20466 , n310893 , 
 n310894 , n310895 , n310896 , n310897 , n310898 , n20473 , n310900 , n310901 , n310902 , n310903 , 
 n310904 , n310905 , n20480 , n310907 , n310908 , n310909 , n310910 , n310911 , n20486 , n310913 , 
 n310914 , n310915 , n310916 , n310917 , n310918 , n310919 , n310920 , n310921 , n20496 , n310923 , 
 n310924 , n310925 , n310926 , n310927 , n310928 , n20503 , n310930 , n310931 , n20506 , n310933 , 
 n310934 , n20509 , n310936 , n20511 , n310938 , n20513 , n20514 , n20515 , n310942 , n310943 , 
 n310944 , n310945 , n20520 , n20521 , n310948 , n310949 , n20524 , n20525 , n310952 , n310953 , 
 n310954 , n20529 , n310956 , n310957 , n310958 , n310959 , n310960 , n20535 , n310962 , n20537 , 
 n310964 , n310965 , n20540 , n310967 , n310968 , n310969 , n310970 , n310971 , n310972 , n20547 , 
 n20548 , n310975 , n310976 , n20551 , n20552 , n310979 , n310980 , n310981 , n310982 , n20557 , 
 n310984 , n310985 , n310986 , n310987 , n20562 , n310989 , n310990 , n310991 , n310992 , n310993 , 
 n310994 , n310995 , n310996 , n310997 , n310998 , n20573 , n20574 , n311001 , n311002 , n311003 , 
 n20578 , n311005 , n311006 , n20581 , n311008 , n20583 , n311010 , n311011 , n311012 , n311013 , 
 n311014 , n311015 , n311016 , n311017 , n311018 , n311019 , n311020 , n311021 , n311022 , n311023 , 
 n311024 , n311025 , n20600 , n20601 , n311028 , n311029 , n311030 , n311031 , n311032 , n20607 , 
 n311034 , n311035 , n20610 , n311037 , n311038 , n311039 , n311040 , n311041 , n20616 , n311043 , 
 n311044 , n20619 , n20620 , n20621 , n311048 , n20623 , n311050 , n311051 , n311052 , n20627 , 
 n20628 , n20629 , n311056 , n20631 , n311058 , n311059 , n311060 , n20635 , n311062 , n311063 , 
 n20638 , n311065 , n311066 , n311067 , n20642 , n311069 , n20644 , n20645 , n20646 , n311073 , 
 n20648 , n311075 , n20650 , n311077 , n20652 , n311079 , n20654 , n311081 , n311082 , n311083 , 
 n311084 , n311085 , n311086 , n311087 , n20662 , n311089 , n311090 , n20665 , n311092 , n311093 , 
 n311094 , n311095 , n311096 , n311097 , n311098 , n311099 , n20674 , n20675 , n311102 , n311103 , 
 n20678 , n311105 , n20680 , n311107 , n20682 , n311109 , n311110 , n20685 , n311112 , n20687 , 
 n20688 , n20689 , n311116 , n20691 , n311118 , n311119 , n311120 , n311121 , n20696 , n20697 , 
 n20698 , n20699 , n20700 , n20701 , n311128 , n20703 , n20704 , n311131 , n20706 , n311133 , 
 n20708 , n311135 , n311136 , n311137 , n311138 , n311139 , n311140 , n311141 , n311142 , n311143 , 
 n311144 , n311145 , n311146 , n311147 , n311148 , n311149 , n311150 , n311151 , n20726 , n20727 , 
 n311154 , n20729 , n311156 , n311157 , n311158 , n311159 , n311160 , n311161 , n20736 , n311163 , 
 n311164 , n311165 , n311166 , n311167 , n311168 , n311169 , n311170 , n20745 , n311172 , n311173 , 
 n311174 , n311175 , n311176 , n20751 , n311178 , n311179 , n20754 , n20755 , n20756 , n311183 , 
 n311184 , n311185 , n20760 , n20761 , n311188 , n311189 , n20764 , n311191 , n311192 , n311193 , 
 n311194 , n311195 , n311196 , n311197 , n311198 , n20773 , n20774 , n311201 , n311202 , n20777 , 
 n311204 , n311205 , n311206 , n311207 , n311208 , n311209 , n20784 , n311211 , n20786 , n311213 , 
 n20788 , n20789 , n20790 , n20791 , n311218 , n20793 , n20794 , n311221 , n20796 , n20797 , 
 n311224 , n311225 , n311226 , n311227 , n311228 , n311229 , n311230 , n311231 , n311232 , n20807 , 
 n311234 , n311235 , n20810 , n311237 , n311238 , n20813 , n20814 , n311241 , n311242 , n20817 , 
 n311244 , n20819 , n311246 , n311247 , n311248 , n311249 , n20824 , n311251 , n311252 , n20827 , 
 n20828 , n311255 , n311256 , n311257 , n20832 , n20833 , n311260 , n20835 , n311262 , n311263 , 
 n311264 , n311265 , n20840 , n311267 , n311268 , n311269 , n20844 , n311271 , n20846 , n311273 , 
 n311274 , n311275 , n311276 , n20851 , n311278 , n311279 , n20854 , n20855 , n311282 , n311283 , 
 n311284 , n311285 , n311286 , n20861 , n311288 , n311289 , n311290 , n311291 , n311292 , n311293 , 
 n311294 , n20869 , n311296 , n311297 , n20872 , n20873 , n311300 , n311301 , n311302 , n311303 , 
 n20878 , n311305 , n20880 , n311307 , n311308 , n311309 , n311310 , n311311 , n311312 , n311313 , 
 n20888 , n311315 , n311316 , n20891 , n311318 , n311319 , n20894 , n20895 , n311322 , n311323 , 
 n20898 , n311325 , n311326 , n311327 , n20902 , n311329 , n311330 , n311331 , n311332 , n311333 , 
 n311334 , n311335 , n20910 , n311337 , n311338 , n311339 , n311340 , n311341 , n20916 , n311343 , 
 n311344 , n20919 , n311346 , n311347 , n311348 , n311349 , n311350 , n20925 , n311352 , n311353 , 
 n311354 , n311355 , n311356 , n20931 , n311358 , n20933 , n20934 , n20935 , n20936 , n311363 , 
 n20938 , n311365 , n311366 , n20941 , n311368 , n311369 , n20944 , n311371 , n311372 , n311373 , 
 n311374 , n311375 , n311376 , n311377 , n311378 , n311379 , n311380 , n20955 , n20956 , n311383 , 
 n311384 , n20959 , n20960 , n20961 , n311388 , n311389 , n20964 , n311391 , n311392 , n311393 , 
 n311394 , n311395 , n311396 , n311397 , n311398 , n20973 , n311400 , n311401 , n311402 , n20977 , 
 n311404 , n311405 , n311406 , n311407 , n20982 , n20983 , n311410 , n311411 , n311412 , n311413 , 
 n20988 , n311415 , n311416 , n311417 , n311418 , n311419 , n311420 , n311421 , n311422 , n311423 , 
 n20998 , n311425 , n311426 , n21001 , n311428 , n21003 , n21004 , n311431 , n311432 , n21007 , 
 n21008 , n21009 , n21010 , n21011 , n311438 , n311439 , n21014 , n311441 , n311442 , n21017 , 
 n21018 , n21019 , n311446 , n311447 , n21022 , n311449 , n21024 , n311451 , n311452 , n311453 , 
 n311454 , n21029 , n311456 , n21031 , n311458 , n311459 , n311460 , n311461 , n311462 , n311463 , 
 n21038 , n311465 , n311466 , n311467 , n21042 , n311469 , n311470 , n21045 , n311472 , n311473 , 
 n311474 , n311475 , n311476 , n21051 , n311478 , n311479 , n21054 , n311481 , n21056 , n311483 , 
 n311484 , n21059 , n311486 , n21061 , n311488 , n21063 , n311490 , n311491 , n311492 , n311493 , 
 n311494 , n311495 , n311496 , n311497 , n311498 , n311499 , n311500 , n311501 , n311502 , n311503 , 
 n311504 , n311505 , n311506 , n21081 , n21082 , n21083 , n311510 , n311511 , n21086 , n311513 , 
 n21088 , n311515 , n311516 , n311517 , n311518 , n311519 , n311520 , n311521 , n311522 , n21097 , 
 n311524 , n311525 , n311526 , n311527 , n311528 , n311529 , n21104 , n311531 , n21106 , n21107 , 
 n21108 , n21109 , n21110 , n21111 , n311538 , n21113 , n311540 , n311541 , n21116 , n311543 , 
 n311544 , n21119 , n21120 , n21121 , n311548 , n21123 , n311550 , n21125 , n311552 , n311553 , 
 n21128 , n311555 , n311556 , n21131 , n311558 , n311559 , n311560 , n311561 , n311562 , n311563 , 
 n21138 , n21139 , n21140 , n311567 , n311568 , n311569 , n311570 , n311571 , n21146 , n311573 , 
 n311574 , n311575 , n21150 , n21151 , n21152 , n311579 , n311580 , n21155 , n311582 , n311583 , 
 n311584 , n21159 , n21160 , n311587 , n311588 , n21163 , n311590 , n21165 , n311592 , n21167 , 
 n21168 , n311595 , n311596 , n21171 , n311598 , n311599 , n21174 , n21175 , n311602 , n311603 , 
 n311604 , n311605 , n311606 , n311607 , n21182 , n311609 , n311610 , n311611 , n21186 , n311613 , 
 n21188 , n311615 , n311616 , n311617 , n311618 , n21193 , n311620 , n311621 , n311622 , n311623 , 
 n311624 , n21199 , n311626 , n311627 , n311628 , n311629 , n311630 , n311631 , n311632 , n311633 , 
 n311634 , n21209 , n311636 , n311637 , n311638 , n311639 , n21214 , n311641 , n311642 , n21217 , 
 n311644 , n311645 , n311646 , n311647 , n311648 , n311649 , n21224 , n311651 , n311652 , n21227 , 
 n21228 , n311655 , n311656 , n21231 , n21232 , n311659 , n311660 , n311661 , n311662 , n311663 , 
 n311664 , n311665 , n311666 , n311667 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , 
 n311674 , n311675 , n311676 , n311677 , n21252 , n21253 , n311680 , n311681 , n311682 , n311683 , 
 n311684 , n311685 , n21260 , n21261 , n311688 , n21263 , n311690 , n311691 , n311692 , n311693 , 
 n311694 , n311695 , n311696 , n311697 , n311698 , n311699 , n311700 , n311701 , n311702 , n311703 , 
 n311704 , n21279 , n21280 , n21281 , n311708 , n311709 , n311710 , n311711 , n311712 , n311713 , 
 n311714 , n21289 , n311716 , n311717 , n311718 , n311719 , n311720 , n21295 , n21296 , n311723 , 
 n311724 , n21299 , n311726 , n311727 , n311728 , n311729 , n311730 , n311731 , n311732 , n311733 , 
 n311734 , n311735 , n311736 , n311737 , n311738 , n311739 , n311740 , n311741 , n311742 , n311743 , 
 n21318 , n311745 , n311746 , n21321 , n311748 , n311749 , n21324 , n311751 , n311752 , n311753 , 
 n311754 , n311755 , n311756 , n311757 , n311758 , n311759 , n311760 , n311761 , n311762 , n21337 , 
 n311764 , n311765 , n311766 , n311767 , n311768 , n311769 , n311770 , n311771 , n311772 , n311773 , 
 n311774 , n21349 , n21350 , n311777 , n311778 , n311779 , n311780 , n311781 , n21356 , n311783 , 
 n311784 , n21359 , n311786 , n311787 , n311788 , n311789 , n311790 , n21365 , n311792 , n311793 , 
 n311794 , n21369 , n311796 , n21371 , n311798 , n311799 , n311800 , n311801 , n311802 , n311803 , 
 n311804 , n311805 , n311806 , n311807 , n311808 , n311809 , n311810 , n311811 , n311812 , n311813 , 
 n311814 , n311815 , n21390 , n311817 , n311818 , n311819 , n311820 , n311821 , n311822 , n311823 , 
 n311824 , n311825 , n311826 , n311827 , n21402 , n311829 , n21404 , n311831 , n311832 , n311833 , 
 n311834 , n21409 , n21410 , n311837 , n311838 , n311839 , n21414 , n311841 , n311842 , n21417 , 
 n21418 , n311845 , n311846 , n21421 , n21422 , n311849 , n311850 , n311851 , n311852 , n21427 , 
 n21428 , n311855 , n311856 , n311857 , n311858 , n21433 , n21434 , n311861 , n311862 , n21437 , 
 n21438 , n311865 , n311866 , n311867 , n21442 , n311869 , n311870 , n311871 , n311872 , n311873 , 
 n311874 , n311875 , n21450 , n311877 , n311878 , n21453 , n311880 , n311881 , n311882 , n311883 , 
 n21458 , n311885 , n311886 , n311887 , n311888 , n311889 , n311890 , n311891 , n311892 , n21467 , 
 n311894 , n311895 , n311896 , n311897 , n311898 , n311899 , n311900 , n311901 , n21476 , n21477 , 
 n311904 , n21479 , n311906 , n311907 , n311908 , n311909 , n21484 , n311911 , n21486 , n21487 , 
 n311914 , n311915 , n21490 , n311917 , n311918 , n21493 , n311920 , n311921 , n21496 , n311923 , 
 n311924 , n311925 , n21500 , n21501 , n311928 , n311929 , n311930 , n311931 , n311932 , n21507 , 
 n311934 , n311935 , n21510 , n311937 , n311938 , n311939 , n311940 , n311941 , n311942 , n311943 , 
 n311944 , n311945 , n21520 , n311947 , n311948 , n311949 , n311950 , n21525 , n311952 , n311953 , 
 n21528 , n311955 , n311956 , n311957 , n311958 , n21533 , n311960 , n311961 , n21536 , n311963 , 
 n311964 , n21539 , n21540 , n21541 , n311968 , n311969 , n21544 , n21545 , n311972 , n311973 , 
 n21548 , n311975 , n311976 , n21551 , n311978 , n311979 , n21554 , n311981 , n311982 , n21557 , 
 n311984 , n311985 , n311986 , n311987 , n311988 , n311989 , n311990 , n311991 , n21566 , n311993 , 
 n21568 , n311995 , n311996 , n311997 , n311998 , n311999 , n312000 , n21575 , n312002 , n312003 , 
 n21578 , n312005 , n312006 , n21581 , n312008 , n312009 , n312010 , n312011 , n21586 , n312013 , 
 n21588 , n21589 , n21590 , n312017 , n312018 , n312019 , n312020 , n21595 , n21596 , n312023 , 
 n21598 , n312025 , n312026 , n21601 , n21602 , n312029 , n21604 , n21605 , n312032 , n312033 , 
 n21608 , n312035 , n21610 , n21611 , n312038 , n21613 , n312040 , n21615 , n312042 , n312043 , 
 n21618 , n312045 , n312046 , n21621 , n21622 , n21623 , n312050 , n312051 , n21626 , n312053 , 
 n312054 , n312055 , n312056 , n312057 , n312058 , n312059 , n21634 , n21635 , n312062 , n312063 , 
 n312064 , n312065 , n312066 , n312067 , n312068 , n312069 , n312070 , n312071 , n21646 , n21647 , 
 n21648 , n312075 , n21650 , n21651 , n312078 , n21653 , n312080 , n312081 , n21656 , n312083 , 
 n312084 , n312085 , n312086 , n312087 , n312088 , n312089 , n312090 , n312091 , n312092 , n312093 , 
 n312094 , n312095 , n21670 , n312097 , n312098 , n21673 , n21674 , n312101 , n21676 , n312103 , 
 n312104 , n21679 , n312106 , n312107 , n312108 , n21683 , n21684 , n312111 , n21686 , n312113 , 
 n21688 , n312115 , n312116 , n312117 , n21692 , n312119 , n312120 , n312121 , n312122 , n312123 , 
 n21698 , n312125 , n312126 , n21701 , n21702 , n312129 , n21704 , n21705 , n312132 , n312133 , 
 n312134 , n312135 , n312136 , n312137 , n312138 , n21713 , n312140 , n21715 , n312142 , n312143 , 
 n21718 , n312145 , n21720 , n312147 , n312148 , n312149 , n312150 , n312151 , n312152 , n312153 , 
 n312154 , n312155 , n312156 , n312157 , n21732 , n312159 , n21734 , n21735 , n312162 , n312163 , 
 n21738 , n312165 , n21740 , n312167 , n312168 , n312169 , n312170 , n312171 , n312172 , n21747 , 
 n312174 , n21749 , n312176 , n312177 , n21752 , n312179 , n21754 , n312181 , n21756 , n312183 , 
 n21758 , n21759 , n312186 , n312187 , n21762 , n21763 , n312190 , n312191 , n312192 , n312193 , 
 n21768 , n312195 , n312196 , n312197 , n21772 , n312199 , n312200 , n312201 , n312202 , n312203 , 
 n312204 , n312205 , n312206 , n312207 , n312208 , n312209 , n312210 , n21785 , n312212 , n312213 , 
 n312214 , n312215 , n312216 , n312217 , n21792 , n312219 , n312220 , n312221 , n21796 , n312223 , 
 n312224 , n21799 , n21800 , n312227 , n21802 , n312229 , n312230 , n21805 , n312232 , n312233 , 
 n312234 , n312235 , n21810 , n312237 , n312238 , n312239 , n312240 , n312241 , n21816 , n312243 , 
 n312244 , n21819 , n21820 , n312247 , n312248 , n21823 , n312250 , n312251 , n312252 , n312253 , 
 n312254 , n21829 , n312256 , n312257 , n312258 , n21833 , n312260 , n312261 , n312262 , n312263 , 
 n312264 , n21839 , n312266 , n312267 , n21842 , n312269 , n312270 , n312271 , n312272 , n312273 , 
 n21848 , n312275 , n312276 , n21851 , n312278 , n312279 , n312280 , n312281 , n312282 , n21857 , 
 n312284 , n312285 , n312286 , n312287 , n21862 , n312289 , n312290 , n21865 , n312292 , n312293 , 
 n21868 , n312295 , n312296 , n21871 , n312298 , n312299 , n312300 , n21875 , n312302 , n312303 , 
 n312304 , n312305 , n312306 , n312307 , n312308 , n312309 , n312310 , n312311 , n312312 , n21887 , 
 n312314 , n21889 , n312316 , n312317 , n312318 , n312319 , n312320 , n312321 , n312322 , n312323 , 
 n312324 , n312325 , n21900 , n312327 , n312328 , n312329 , n312330 , n312331 , n312332 , n312333 , 
 n312334 , n312335 , n312336 , n312337 , n312338 , n21913 , n312340 , n312341 , n312342 , n312343 , 
 n312344 , n312345 , n312346 , n21921 , n312348 , n312349 , n21924 , n312351 , n312352 , n312353 , 
 n312354 , n312355 , n312356 , n312357 , n312358 , n312359 , n312360 , n312361 , n21936 , n312363 , 
 n312364 , n312365 , n312366 , n312367 , n312368 , n21943 , n312370 , n312371 , n312372 , n312373 , 
 n312374 , n312375 , n312376 , n312377 , n21952 , n312379 , n312380 , n21955 , n312382 , n312383 , 
 n312384 , n312385 , n312386 , n312387 , n21962 , n312389 , n312390 , n312391 , n312392 , n312393 , 
 n312394 , n312395 , n312396 , n312397 , n21972 , n312399 , n21974 , n21975 , n312402 , n312403 , 
 n312404 , n312405 , n312406 , n312407 , n312408 , n312409 , n312410 , n21985 , n312412 , n312413 , 
 n21988 , n312415 , n312416 , n312417 , n312418 , n21993 , n21994 , n21995 , n312422 , n21997 , 
 n21998 , n312425 , n22000 , n312427 , n312428 , n22003 , n312430 , n312431 , n312432 , n312433 , 
 n312434 , n312435 , n312436 , n22011 , n22012 , n312439 , n22014 , n312441 , n312442 , n312443 , 
 n312444 , n312445 , n312446 , n312447 , n312448 , n22023 , n312450 , n312451 , n312452 , n312453 , 
 n312454 , n312455 , n312456 , n312457 , n312458 , n312459 , n312460 , n312461 , n312462 , n312463 , 
 n312464 , n312465 , n22040 , n312467 , n312468 , n22043 , n22044 , n312471 , n312472 , n22047 , 
 n312474 , n312475 , n312476 , n22051 , n22052 , n312479 , n312480 , n22055 , n312482 , n312483 , 
 n22058 , n312485 , n312486 , n312487 , n312488 , n22063 , n312490 , n312491 , n22066 , n22067 , 
 n312494 , n312495 , n22070 , n312497 , n22072 , n22073 , n312500 , n312501 , n312502 , n312503 , 
 n312504 , n312505 , n22080 , n312507 , n22082 , n22083 , n22084 , n22085 , n312512 , n312513 , 
 n22088 , n312515 , n22090 , n22091 , n312518 , n312519 , n312520 , n22095 , n312522 , n312523 , 
 n312524 , n22099 , n312526 , n312527 , n312528 , n312529 , n312530 , n312531 , n312532 , n312533 , 
 n312534 , n312535 , n312536 , n312537 , n312538 , n312539 , n312540 , n312541 , n22116 , n312543 , 
 n312544 , n22119 , n312546 , n312547 , n22122 , n312549 , n312550 , n312551 , n22126 , n312553 , 
 n312554 , n312555 , n312556 , n312557 , n22132 , n312559 , n22134 , n312561 , n312562 , n312563 , 
 n22138 , n22139 , n312566 , n312567 , n312568 , n312569 , n312570 , n312571 , n22146 , n312573 , 
 n312574 , n22149 , n312576 , n312577 , n312578 , n22153 , n312580 , n312581 , n312582 , n312583 , 
 n312584 , n312585 , n312586 , n312587 , n22162 , n312589 , n22164 , n312591 , n22166 , n312593 , 
 n22168 , n312595 , n312596 , n22171 , n312598 , n22173 , n312600 , n312601 , n312602 , n22177 , 
 n312604 , n312605 , n312606 , n312607 , n312608 , n312609 , n312610 , n312611 , n312612 , n312613 , 
 n312614 , n312615 , n22190 , n312617 , n312618 , n312619 , n22194 , n22195 , n312622 , n312623 , 
 n22198 , n312625 , n22200 , n312627 , n22202 , n312629 , n312630 , n22205 , n312632 , n312633 , 
 n22208 , n22209 , n312636 , n312637 , n312638 , n312639 , n312640 , n22215 , n312642 , n312643 , 
 n312644 , n312645 , n22220 , n312647 , n22222 , n312649 , n22224 , n312651 , n312652 , n312653 , 
 n312654 , n312655 , n312656 , n312657 , n312658 , n312659 , n312660 , n312661 , n312662 , n312663 , 
 n312664 , n312665 , n312666 , n312667 , n22242 , n312669 , n312670 , n312671 , n22246 , n312673 , 
 n312674 , n312675 , n312676 , n312677 , n312678 , n312679 , n312680 , n312681 , n312682 , n22257 , 
 n312684 , n312685 , n312686 , n22261 , n312688 , n22263 , n312690 , n312691 , n312692 , n312693 , 
 n312694 , n312695 , n312696 , n22271 , n312698 , n312699 , n312700 , n312701 , n312702 , n312703 , 
 n312704 , n312705 , n312706 , n312707 , n312708 , n312709 , n22284 , n312711 , n312712 , n22287 , 
 n312714 , n312715 , n312716 , n22291 , n22292 , n312719 , n22294 , n312721 , n22296 , n312723 , 
 n22298 , n312725 , n312726 , n22301 , n22302 , n312729 , n312730 , n22305 , n312732 , n312733 , 
 n312734 , n312735 , n312736 , n312737 , n22312 , n312739 , n22314 , n22315 , n312742 , n312743 , 
 n22318 , n312745 , n312746 , n312747 , n312748 , n22323 , n312750 , n312751 , n312752 , n312753 , 
 n312754 , n312755 , n312756 , n312757 , n22332 , n312759 , n312760 , n312761 , n22336 , n312763 , 
 n312764 , n312765 , n312766 , n312767 , n22342 , n312769 , n312770 , n312771 , n312772 , n312773 , 
 n22348 , n22349 , n22350 , n312777 , n312778 , n312779 , n312780 , n22355 , n312782 , n22357 , 
 n312784 , n312785 , n312786 , n312787 , n22362 , n312789 , n312790 , n312791 , n312792 , n312793 , 
 n312794 , n312795 , n312796 , n312797 , n312798 , n312799 , n312800 , n312801 , n312802 , n312803 , 
 n312804 , n22379 , n312806 , n312807 , n22382 , n312809 , n312810 , n312811 , n312812 , n312813 , 
 n22388 , n312815 , n312816 , n312817 , n22392 , n312819 , n22394 , n22395 , n22396 , n22397 , 
 n22398 , n22399 , n22400 , n22401 , n312828 , n312829 , n312830 , n22405 , n22406 , n22407 , 
 n312834 , n312835 , n312836 , n312837 , n312838 , n22413 , n312840 , n312841 , n312842 , n312843 , 
 n312844 , n22419 , n312846 , n22421 , n22422 , n22423 , n312850 , n22425 , n22426 , n312853 , 
 n312854 , n312855 , n312856 , n22431 , n312858 , n312859 , n22434 , n312861 , n312862 , n312863 , 
 n312864 , n312865 , n312866 , n312867 , n312868 , n312869 , n312870 , n312871 , n312872 , n312873 , 
 n312874 , n312875 , n22450 , n312877 , n312878 , n312879 , n312880 , n312881 , n312882 , n22457 , 
 n312884 , n312885 , n22460 , n312887 , n312888 , n312889 , n312890 , n312891 , n22466 , n312893 , 
 n312894 , n312895 , n312896 , n312897 , n22472 , n312899 , n312900 , n22475 , n312902 , n312903 , 
 n312904 , n312905 , n312906 , n22481 , n312908 , n22483 , n312910 , n22485 , n22486 , n312913 , 
 n22488 , n312915 , n22490 , n312917 , n312918 , n22493 , n312920 , n22495 , n312922 , n312923 , 
 n22498 , n22499 , n312926 , n22501 , n312928 , n312929 , n22504 , n312931 , n22506 , n312933 , 
 n22508 , n22509 , n312936 , n312937 , n22512 , n312939 , n22514 , n22515 , n22516 , n312943 , 
 n312944 , n22519 , n312946 , n312947 , n312948 , n312949 , n312950 , n312951 , n312952 , n312953 , 
 n22528 , n312955 , n312956 , n312957 , n312958 , n312959 , n312960 , n312961 , n312962 , n312963 , 
 n312964 , n22539 , n312966 , n22541 , n22542 , n312969 , n312970 , n22545 , n22546 , n312973 , 
 n312974 , n22549 , n22550 , n22551 , n22552 , n312979 , n312980 , n312981 , n22556 , n22557 , 
 n312984 , n312985 , n22560 , n22561 , n22562 , n312989 , n312990 , n22565 , n22566 , n22567 , 
 n312994 , n312995 , n22570 , n312997 , n312998 , n22573 , n313000 , n313001 , n313002 , n22577 , 
 n22578 , n313005 , n22580 , n22581 , n313008 , n313009 , n313010 , n313011 , n22586 , n22587 , 
 n313014 , n313015 , n313016 , n313017 , n313018 , n313019 , n313020 , n313021 , n313022 , n313023 , 
 n313024 , n313025 , n313026 , n313027 , n313028 , n313029 , n313030 , n313031 , n313032 , n313033 , 
 n313034 , n313035 , n313036 , n313037 , n313038 , n22613 , n313040 , n313041 , n22616 , n313043 , 
 n22618 , n22619 , n313046 , n313047 , n313048 , n313049 , n313050 , n313051 , n313052 , n313053 , 
 n313054 , n313055 , n313056 , n313057 , n313058 , n313059 , n313060 , n313061 , n313062 , n313063 , 
 n313064 , n313065 , n313066 , n313067 , n313068 , n313069 , n22644 , n22645 , n313072 , n313073 , 
 n313074 , n313075 , n313076 , n313077 , n313078 , n313079 , n313080 , n313081 , n313082 , n313083 , 
 n313084 , n313085 , n22660 , n22661 , n313088 , n22663 , n313090 , n22665 , n313092 , n313093 , 
 n22668 , n313095 , n22670 , n22671 , n313098 , n313099 , n313100 , n313101 , n22676 , n313103 , 
 n313104 , n313105 , n313106 , n313107 , n313108 , n313109 , n313110 , n22685 , n313112 , n22687 , 
 n22688 , n313115 , n313116 , n313117 , n313118 , n22693 , n313120 , n313121 , n313122 , n313123 , 
 n313124 , n313125 , n313126 , n313127 , n313128 , n22703 , n313130 , n313131 , n22706 , n22707 , 
 n22708 , n22709 , n22710 , n313137 , n22712 , n313139 , n313140 , n22715 , n313142 , n313143 , 
 n22718 , n22719 , n313146 , n22721 , n313148 , n313149 , n22724 , n22725 , n313152 , n22727 , 
 n22728 , n313155 , n313156 , n22731 , n313158 , n313159 , n22734 , n313161 , n313162 , n22737 , 
 n22738 , n313165 , n313166 , n22741 , n22742 , n22743 , n22744 , n313171 , n22746 , n22747 , 
 n313174 , n22749 , n22750 , n313177 , n313178 , n313179 , n313180 , n313181 , n313182 , n313183 , 
 n22758 , n313185 , n313186 , n313187 , n313188 , n22763 , n313190 , n313191 , n313192 , n22767 , 
 n313194 , n313195 , n313196 , n313197 , n313198 , n313199 , n313200 , n22775 , n22776 , n313203 , 
 n313204 , n22779 , n313206 , n313207 , n22782 , n313209 , n313210 , n313211 , n313212 , n313213 , 
 n22788 , n313215 , n313216 , n22791 , n313218 , n313219 , n313220 , n313221 , n313222 , n313223 , 
 n313224 , n313225 , n22800 , n22801 , n22802 , n22803 , n313230 , n22805 , n22806 , n313233 , 
 n22808 , n313235 , n313236 , n313237 , n313238 , n313239 , n313240 , n22815 , n313242 , n22817 , 
 n313244 , n313245 , n313246 , n313247 , n313248 , n313249 , n313250 , n22825 , n22826 , n22827 , 
 n22828 , n313255 , n313256 , n22831 , n22832 , n22833 , n22834 , n22835 , n313262 , n313263 , 
 n22838 , n313265 , n313266 , n22841 , n313268 , n313269 , n313270 , n313271 , n313272 , n22847 , 
 n22848 , n22849 , n22850 , n313277 , n313278 , n22853 , n22854 , n313281 , n313282 , n22857 , 
 n313284 , n313285 , n313286 , n313287 , n22862 , n313289 , n22864 , n313291 , n313292 , n313293 , 
 n313294 , n313295 , n313296 , n22871 , n22872 , n22873 , n22874 , n313301 , n313302 , n22877 , 
 n313304 , n22879 , n22880 , n313307 , n313308 , n22883 , n313310 , n313311 , n313312 , n313313 , 
 n313314 , n313315 , n313316 , n313317 , n313318 , n313319 , n313320 , n313321 , n22896 , n313323 , 
 n313324 , n313325 , n22900 , n313327 , n313328 , n22903 , n313330 , n22905 , n313332 , n313333 , 
 n313334 , n313335 , n313336 , n313337 , n313338 , n313339 , n22914 , n313341 , n313342 , n313343 , 
 n313344 , n313345 , n313346 , n313347 , n22922 , n313349 , n313350 , n22925 , n313352 , n313353 , 
 n313354 , n22929 , n313356 , n313357 , n22932 , n313359 , n313360 , n22935 , n313362 , n22937 , 
 n313364 , n313365 , n313366 , n313367 , n22942 , n22943 , n22944 , n22945 , n313372 , n22947 , 
 n313374 , n313375 , n313376 , n313377 , n313378 , n313379 , n313380 , n313381 , n313382 , n313383 , 
 n313384 , n313385 , n313386 , n22961 , n22962 , n313389 , n22964 , n313391 , n313392 , n313393 , 
 n313394 , n313395 , n313396 , n22971 , n22972 , n313399 , n22974 , n22975 , n22976 , n313403 , 
 n313404 , n313405 , n313406 , n313407 , n313408 , n313409 , n313410 , n22985 , n313412 , n22987 , 
 n313414 , n313415 , n313416 , n22991 , n313418 , n313419 , n313420 , n313421 , n313422 , n313423 , 
 n313424 , n313425 , n23000 , n313427 , n313428 , n23003 , n23004 , n23005 , n313432 , n313433 , 
 n313434 , n313435 , n23010 , n313437 , n23012 , n23013 , n313440 , n313441 , n313442 , n313443 , 
 n23018 , n313445 , n313446 , n313447 , n313448 , n313449 , n313450 , n313451 , n313452 , n313453 , 
 n313454 , n23029 , n313456 , n313457 , n313458 , n313459 , n313460 , n313461 , n313462 , n313463 , 
 n313464 , n313465 , n313466 , n313467 , n313468 , n313469 , n313470 , n313471 , n313472 , n313473 , 
 n313474 , n23049 , n313476 , n313477 , n313478 , n313479 , n313480 , n313481 , n313482 , n313483 , 
 n313484 , n313485 , n313486 , n313487 , n313488 , n313489 , n313490 , n23065 , n313492 , n313493 , 
 n313494 , n313495 , n23070 , n23071 , n313498 , n23073 , n313500 , n313501 , n313502 , n313503 , 
 n313504 , n313505 , n313506 , n313507 , n313508 , n23083 , n313510 , n313511 , n313512 , n313513 , 
 n313514 , n313515 , n313516 , n313517 , n313518 , n23093 , n23094 , n23095 , n313522 , n23097 , 
 n23098 , n313525 , n23100 , n23101 , n313528 , n313529 , n313530 , n313531 , n313532 , n313533 , 
 n313534 , n313535 , n313536 , n313537 , n313538 , n313539 , n313540 , n313541 , n313542 , n313543 , 
 n23118 , n313545 , n23120 , n23121 , n313548 , n313549 , n23124 , n313551 , n313552 , n313553 , 
 n313554 , n313555 , n313556 , n313557 , n313558 , n313559 , n23134 , n313561 , n313562 , n313563 , 
 n23138 , n313565 , n313566 , n313567 , n313568 , n23143 , n313570 , n313571 , n23146 , n313573 , 
 n313574 , n313575 , n313576 , n313577 , n313578 , n313579 , n313580 , n313581 , n313582 , n313583 , 
 n313584 , n313585 , n313586 , n313587 , n313588 , n313589 , n313590 , n313591 , n313592 , n313593 , 
 n313594 , n313595 , n313596 , n313597 , n313598 , n313599 , n23174 , n23175 , n313602 , n23177 , 
 n313604 , n313605 , n313606 , n313607 , n313608 , n23183 , n313610 , n23185 , n23186 , n313613 , 
 n23188 , n313615 , n313616 , n313617 , n313618 , n313619 , n313620 , n313621 , n313622 , n23197 , 
 n313624 , n313625 , n313626 , n313627 , n313628 , n313629 , n23204 , n313631 , n23206 , n313633 , 
 n313634 , n313635 , n313636 , n313637 , n313638 , n313639 , n313640 , n313641 , n23216 , n313643 , 
 n313644 , n23219 , n313646 , n23221 , n313648 , n313649 , n23224 , n313651 , n313652 , n313653 , 
 n313654 , n313655 , n313656 , n313657 , n23232 , n313659 , n313660 , n313661 , n313662 , n23237 , 
 n313664 , n313665 , n23240 , n23241 , n313668 , n313669 , n313670 , n313671 , n313672 , n313673 , 
 n313674 , n313675 , n23250 , n23251 , n313678 , n313679 , n313680 , n313681 , n313682 , n313683 , 
 n313684 , n313685 , n313686 , n23261 , n23262 , n313689 , n23264 , n313691 , n313692 , n313693 , 
 n313694 , n23269 , n313696 , n23271 , n313698 , n23273 , n23274 , n313701 , n23276 , n313703 , 
 n313704 , n23279 , n313706 , n313707 , n23282 , n313709 , n313710 , n23285 , n313712 , n23287 , 
 n313714 , n313715 , n23290 , n313717 , n313718 , n313719 , n313720 , n313721 , n313722 , n313723 , 
 n313724 , n313725 , n313726 , n23301 , n313728 , n23303 , n313730 , n313731 , n313732 , n313733 , 
 n313734 , n313735 , n313736 , n313737 , n313738 , n313739 , n23314 , n313741 , n313742 , n313743 , 
 n313744 , n23319 , n313746 , n313747 , n313748 , n313749 , n313750 , n313751 , n23326 , n313753 , 
 n313754 , n313755 , n23330 , n313757 , n313758 , n313759 , n23334 , n313761 , n313762 , n23337 , 
 n313764 , n313765 , n313766 , n313767 , n313768 , n313769 , n313770 , n313771 , n313772 , n313773 , 
 n23348 , n313775 , n313776 , n313777 , n313778 , n313779 , n313780 , n313781 , n313782 , n313783 , 
 n313784 , n313785 , n313786 , n313787 , n313788 , n313789 , n313790 , n313791 , n23366 , n313793 , 
 n313794 , n313795 , n313796 , n313797 , n313798 , n313799 , n313800 , n313801 , n313802 , n313803 , 
 n313804 , n23379 , n313806 , n313807 , n23382 , n313809 , n23384 , n313811 , n313812 , n313813 , 
 n23388 , n23389 , n23390 , n313817 , n313818 , n23393 , n23394 , n313821 , n313822 , n313823 , 
 n23398 , n313825 , n23400 , n313827 , n313828 , n313829 , n313830 , n23405 , n313832 , n313833 , 
 n23408 , n313835 , n313836 , n23411 , n313838 , n313839 , n23414 , n313841 , n23416 , n313843 , 
 n23418 , n313845 , n313846 , n313847 , n313848 , n313849 , n313850 , n313851 , n313852 , n313853 , 
 n313854 , n313855 , n313856 , n313857 , n313858 , n313859 , n313860 , n313861 , n313862 , n313863 , 
 n313864 , n313865 , n23440 , n23441 , n313868 , n23443 , n313870 , n313871 , n313872 , n313873 , 
 n23448 , n23449 , n313876 , n313877 , n313878 , n313879 , n23454 , n313881 , n23456 , n313883 , 
 n23458 , n313885 , n313886 , n313887 , n313888 , n313889 , n313890 , n313891 , n23466 , n313893 , 
 n313894 , n313895 , n313896 , n313897 , n313898 , n313899 , n313900 , n313901 , n313902 , n313903 , 
 n313904 , n313905 , n313906 , n313907 , n313908 , n313909 , n313910 , n313911 , n313912 , n313913 , 
 n313914 , n313915 , n313916 , n313917 , n313918 , n313919 , n313920 , n313921 , n23496 , n313923 , 
 n313924 , n23499 , n23500 , n313927 , n313928 , n23503 , n23504 , n313931 , n313932 , n23507 , 
 n313934 , n313935 , n313936 , n313937 , n313938 , n313939 , n313940 , n313941 , n313942 , n313943 , 
 n23518 , n313945 , n313946 , n313947 , n313948 , n313949 , n313950 , n313951 , n313952 , n313953 , 
 n313954 , n313955 , n313956 , n313957 , n23532 , n313959 , n313960 , n313961 , n313962 , n313963 , 
 n313964 , n23539 , n313966 , n313967 , n313968 , n313969 , n313970 , n23545 , n313972 , n313973 , 
 n23548 , n313975 , n313976 , n313977 , n23552 , n23553 , n313980 , n23555 , n313982 , n313983 , 
 n313984 , n23559 , n313986 , n313987 , n313988 , n23563 , n313990 , n313991 , n313992 , n313993 , 
 n313994 , n313995 , n313996 , n313997 , n313998 , n313999 , n23574 , n314001 , n314002 , n314003 , 
 n23578 , n23579 , n23580 , n23581 , n314008 , n314009 , n314010 , n23585 , n23586 , n23587 , 
 n23588 , n314015 , n314016 , n314017 , n314018 , n314019 , n314020 , n314021 , n314022 , n23597 , 
 n314024 , n314025 , n314026 , n23601 , n314028 , n314029 , n23604 , n314031 , n23606 , n314033 , 
 n23608 , n314035 , n314036 , n23611 , n314038 , n314039 , n314040 , n314041 , n314042 , n314043 , 
 n314044 , n314045 , n23620 , n314047 , n314048 , n23623 , n23624 , n314051 , n314052 , n23627 , 
 n23628 , n314055 , n314056 , n314057 , n23632 , n314059 , n314060 , n314061 , n314062 , n23637 , 
 n314064 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n314071 , n314072 , n314073 , 
 n314074 , n23649 , n314076 , n23651 , n23652 , n23653 , n23654 , n314081 , n23656 , n23657 , 
 n314084 , n23659 , n314086 , n314087 , n23662 , n314089 , n314090 , n23665 , n314092 , n314093 , 
 n314094 , n23669 , n314096 , n314097 , n314098 , n314099 , n23674 , n314101 , n314102 , n23677 , 
 n23678 , n23679 , n23680 , n23681 , n314108 , n314109 , n23684 , n23685 , n314112 , n314113 , 
 n23688 , n314115 , n314116 , n314117 , n314118 , n23693 , n23694 , n314121 , n314122 , n314123 , 
 n314124 , n314125 , n314126 , n23701 , n23702 , n314129 , n23704 , n314131 , n23706 , n314133 , 
 n314134 , n314135 , n314136 , n314137 , n314138 , n314139 , n314140 , n314141 , n314142 , n314143 , 
 n314144 , n23719 , n314146 , n314147 , n314148 , n314149 , n23724 , n314151 , n314152 , n314153 , 
 n23728 , n23729 , n314156 , n314157 , n314158 , n314159 , n23734 , n314161 , n314162 , n314163 , 
 n23738 , n314165 , n314166 , n314167 , n23742 , n314169 , n314170 , n314171 , n23746 , n314173 , 
 n23748 , n23749 , n314176 , n314177 , n314178 , n314179 , n314180 , n23755 , n314182 , n23757 , 
 n314184 , n314185 , n314186 , n314187 , n314188 , n23763 , n23764 , n314191 , n314192 , n23767 , 
 n314194 , n314195 , n314196 , n314197 , n314198 , n314199 , n314200 , n314201 , n314202 , n23777 , 
 n23778 , n23779 , n314206 , n23781 , n23782 , n314209 , n314210 , n23785 , n23786 , n314213 , 
 n314214 , n23789 , n314216 , n314217 , n23792 , n314219 , n314220 , n314221 , n314222 , n314223 , 
 n314224 , n314225 , n314226 , n314227 , n314228 , n23803 , n23804 , n23805 , n314232 , n314233 , 
 n314234 , n314235 , n314236 , n23811 , n23812 , n314239 , n23814 , n314241 , n314242 , n23817 , 
 n314244 , n23819 , n314246 , n23821 , n23822 , n314249 , n314250 , n314251 , n23826 , n314253 , 
 n314254 , n23829 , n314256 , n314257 , n23832 , n314259 , n314260 , n314261 , n314262 , n314263 , 
 n314264 , n314265 , n23840 , n23841 , n23842 , n23843 , n314270 , n314271 , n314272 , n23847 , 
 n314274 , n314275 , n314276 , n314277 , n23852 , n314279 , n23854 , n23855 , n314282 , n23857 , 
 n23858 , n23859 , n23860 , n314287 , n314288 , n314289 , n23864 , n314291 , n314292 , n23867 , 
 n314294 , n314295 , n23870 , n23871 , n314298 , n314299 , n314300 , n23875 , n23876 , n314303 , 
 n314304 , n314305 , n23880 , n314307 , n314308 , n314309 , n314310 , n314311 , n314312 , n314313 , 
 n314314 , n314315 , n314316 , n314317 , n23892 , n314319 , n314320 , n23895 , n23896 , n314323 , 
 n23898 , n314325 , n23900 , n314327 , n314328 , n314329 , n314330 , n314331 , n23906 , n314333 , 
 n314334 , n314335 , n314336 , n23911 , n314338 , n314339 , n314340 , n314341 , n23916 , n314343 , 
 n314344 , n314345 , n314346 , n314347 , n314348 , n314349 , n314350 , n314351 , n314352 , n314353 , 
 n314354 , n314355 , n23930 , n314357 , n314358 , n314359 , n23934 , n314361 , n314362 , n23937 , 
 n23938 , n314365 , n314366 , n314367 , n23942 , n314369 , n23944 , n314371 , n314372 , n314373 , 
 n314374 , n314375 , n314376 , n314377 , n23952 , n314379 , n314380 , n23955 , n314382 , n314383 , 
 n23958 , n314385 , n23960 , n23961 , n314388 , n23963 , n314390 , n23965 , n314392 , n23967 , 
 n23968 , n314395 , n314396 , n23971 , n314398 , n314399 , n314400 , n23975 , n314402 , n314403 , 
 n314404 , n314405 , n314406 , n314407 , n314408 , n314409 , n314410 , n23985 , n314412 , n314413 , 
 n314414 , n314415 , n23990 , n314417 , n23992 , n314419 , n314420 , n23995 , n23996 , n314423 , 
 n314424 , n23999 , n314426 , n314427 , n314428 , n314429 , n24004 , n24005 , n24006 , n314433 , 
 n314434 , n314435 , n24010 , n24011 , n24012 , n314439 , n314440 , n24015 , n24016 , n314443 , 
 n314444 , n24019 , n24020 , n24021 , n314448 , n24023 , n24024 , n24025 , n24026 , n24027 , 
 n24028 , n314455 , n314456 , n24031 , n24032 , n314459 , n24034 , n314461 , n314462 , n24037 , 
 n24038 , n314465 , n314466 , n24041 , n24042 , n314469 , n24044 , n24045 , n24046 , n314473 , 
 n314474 , n24049 , n314476 , n314477 , n314478 , n314479 , n314480 , n314481 , n314482 , n314483 , 
 n314484 , n314485 , n314486 , n24061 , n314488 , n314489 , n314490 , n314491 , n314492 , n314493 , 
 n314494 , n24069 , n314496 , n314497 , n24072 , n24073 , n314500 , n314501 , n314502 , n314503 , 
 n314504 , n24079 , n314506 , n314507 , n24082 , n314509 , n314510 , n24085 , n314512 , n24087 , 
 n24088 , n24089 , n24090 , n314517 , n24092 , n24093 , n24094 , n314521 , n314522 , n314523 , 
 n24098 , n314525 , n314526 , n314527 , n314528 , n24103 , n314530 , n314531 , n314532 , n314533 , 
 n314534 , n314535 , n314536 , n314537 , n24112 , n314539 , n314540 , n24115 , n24116 , n314543 , 
 n314544 , n314545 , n314546 , n24121 , n314548 , n314549 , n314550 , n314551 , n314552 , n314553 , 
 n314554 , n314555 , n24130 , n314557 , n314558 , n314559 , n314560 , n314561 , n314562 , n314563 , 
 n314564 , n314565 , n314566 , n314567 , n314568 , n24143 , n314570 , n314571 , n24146 , n314573 , 
 n314574 , n24149 , n314576 , n314577 , n314578 , n314579 , n24154 , n24155 , n314582 , n314583 , 
 n314584 , n314585 , n314586 , n314587 , n314588 , n24163 , n314590 , n314591 , n314592 , n314593 , 
 n24168 , n314595 , n314596 , n314597 , n314598 , n314599 , n314600 , n314601 , n314602 , n314603 , 
 n314604 , n24179 , n24180 , n24181 , n24182 , n314609 , n24184 , n314611 , n314612 , n24187 , 
 n314614 , n314615 , n314616 , n314617 , n314618 , n24193 , n314620 , n314621 , n24196 , n314623 , 
 n314624 , n314625 , n314626 , n314627 , n314628 , n24203 , n24204 , n24205 , n314632 , n314633 , 
 n314634 , n314635 , n314636 , n314637 , n314638 , n314639 , n314640 , n314641 , n24216 , n24217 , 
 n314644 , n314645 , n24220 , n314647 , n314648 , n314649 , n314650 , n314651 , n314652 , n24227 , 
 n314654 , n24229 , n314656 , n314657 , n314658 , n314659 , n24234 , n314661 , n314662 , n314663 , 
 n314664 , n314665 , n314666 , n314667 , n314668 , n314669 , n24244 , n314671 , n314672 , n24247 , 
 n314674 , n24249 , n24250 , n24251 , n24252 , n314679 , n24254 , n24255 , n314682 , n314683 , 
 n314684 , n314685 , n314686 , n314687 , n314688 , n314689 , n314690 , n24265 , n314692 , n314693 , 
 n314694 , n24269 , n24270 , n24271 , n314698 , n314699 , n24274 , n24275 , n314702 , n314703 , 
 n24278 , n314705 , n314706 , n24281 , n24282 , n314709 , n24284 , n24285 , n314712 , n314713 , 
 n314714 , n314715 , n314716 , n24291 , n24292 , n24293 , n24294 , n24295 , n314722 , n314723 , 
 n314724 , n314725 , n314726 , n314727 , n314728 , n314729 , n314730 , n314731 , n24306 , n314733 , 
 n314734 , n314735 , n24310 , n314737 , n24312 , n314739 , n314740 , n24315 , n314742 , n314743 , 
 n24318 , n314745 , n24320 , n314747 , n314748 , n314749 , n314750 , n24325 , n314752 , n314753 , 
 n24328 , n24329 , n314756 , n314757 , n24332 , n314759 , n314760 , n24335 , n314762 , n314763 , 
 n24338 , n314765 , n314766 , n314767 , n314768 , n24343 , n24344 , n314771 , n314772 , n24347 , 
 n314774 , n314775 , n24350 , n314777 , n24352 , n24353 , n24354 , n314781 , n314782 , n314783 , 
 n314784 , n314785 , n314786 , n314787 , n24362 , n24363 , n314790 , n314791 , n314792 , n314793 , 
 n314794 , n24369 , n314796 , n314797 , n24372 , n314799 , n314800 , n314801 , n314802 , n314803 , 
 n24378 , n314805 , n314806 , n24381 , n314808 , n314809 , n24384 , n314811 , n314812 , n24387 , 
 n314814 , n314815 , n314816 , n24391 , n314818 , n24393 , n314820 , n314821 , n24396 , n314823 , 
 n314824 , n24399 , n314826 , n314827 , n314828 , n314829 , n314830 , n314831 , n314832 , n314833 , 
 n314834 , n24409 , n314836 , n314837 , n314838 , n314839 , n314840 , n314841 , n24416 , n314843 , 
 n314844 , n314845 , n314846 , n314847 , n24422 , n314849 , n314850 , n24425 , n314852 , n314853 , 
 n314854 , n24429 , n314856 , n24431 , n24432 , n314859 , n24434 , n314861 , n314862 , n314863 , 
 n314864 , n314865 , n314866 , n314867 , n24442 , n314869 , n314870 , n24445 , n24446 , n314873 , 
 n314874 , n314875 , n24450 , n24451 , n314878 , n314879 , n24454 , n314881 , n314882 , n314883 , 
 n314884 , n314885 , n314886 , n314887 , n314888 , n314889 , n314890 , n314891 , n314892 , n314893 , 
 n314894 , n24469 , n314896 , n314897 , n314898 , n314899 , n314900 , n314901 , n314902 , n314903 , 
 n314904 , n314905 , n24480 , n314907 , n314908 , n314909 , n314910 , n314911 , n24486 , n314913 , 
 n24488 , n314915 , n314916 , n314917 , n314918 , n314919 , n314920 , n24495 , n314922 , n314923 , 
 n24498 , n314925 , n314926 , n24501 , n314928 , n314929 , n314930 , n24505 , n314932 , n314933 , 
 n24508 , n314935 , n314936 , n314937 , n314938 , n24513 , n314940 , n314941 , n314942 , n314943 , 
 n314944 , n314945 , n314946 , n314947 , n314948 , n24523 , n314950 , n314951 , n24526 , n314953 , 
 n314954 , n314955 , n314956 , n314957 , n314958 , n314959 , n24534 , n314961 , n314962 , n314963 , 
 n314964 , n314965 , n314966 , n24541 , n314968 , n314969 , n24544 , n314971 , n314972 , n314973 , 
 n314974 , n314975 , n314976 , n314977 , n314978 , n314979 , n314980 , n314981 , n314982 , n24557 , 
 n24558 , n314985 , n314986 , n314987 , n314988 , n314989 , n24564 , n314991 , n24566 , n314993 , 
 n314994 , n314995 , n314996 , n314997 , n314998 , n314999 , n24574 , n24575 , n315002 , n315003 , 
 n315004 , n315005 , n315006 , n315007 , n315008 , n315009 , n315010 , n315011 , n315012 , n315013 , 
 n315014 , n315015 , n315016 , n315017 , n315018 , n315019 , n315020 , n24595 , n315022 , n315023 , 
 n24598 , n315025 , n315026 , n24601 , n315028 , n315029 , n24604 , n315031 , n315032 , n24607 , 
 n315034 , n315035 , n315036 , n315037 , n315038 , n315039 , n24614 , n315041 , n315042 , n315043 , 
 n315044 , n24619 , n315046 , n315047 , n24622 , n315049 , n315050 , n24625 , n315052 , n24627 , 
 n315054 , n24629 , n315056 , n315057 , n315058 , n315059 , n315060 , n315061 , n315062 , n315063 , 
 n315064 , n315065 , n315066 , n315067 , n315068 , n315069 , n315070 , n315071 , n24646 , n315073 , 
 n315074 , n315075 , n315076 , n315077 , n315078 , n315079 , n315080 , n315081 , n315082 , n24657 , 
 n315084 , n315085 , n24660 , n315087 , n315088 , n24663 , n315090 , n315091 , n315092 , n24667 , 
 n315094 , n315095 , n24670 , n24671 , n315098 , n315099 , n315100 , n24675 , n315102 , n315103 , 
 n24678 , n315105 , n315106 , n315107 , n315108 , n315109 , n24684 , n315111 , n315112 , n24687 , 
 n315114 , n315115 , n24690 , n315117 , n315118 , n24693 , n315120 , n315121 , n315122 , n315123 , 
 n24698 , n315125 , n315126 , n315127 , n315128 , n315129 , n24704 , n315131 , n315132 , n315133 , 
 n315134 , n315135 , n24710 , n315137 , n315138 , n24713 , n24714 , n315141 , n24716 , n315143 , 
 n315144 , n315145 , n24720 , n315147 , n24722 , n315149 , n315150 , n24725 , n315152 , n315153 , 
 n24728 , n315155 , n315156 , n315157 , n315158 , n315159 , n24734 , n315161 , n315162 , n315163 , 
 n315164 , n315165 , n315166 , n315167 , n315168 , n315169 , n315170 , n315171 , n24746 , n24747 , 
 n315174 , n315175 , n24750 , n315177 , n315178 , n24753 , n315180 , n315181 , n24756 , n315183 , 
 n315184 , n24759 , n315186 , n315187 , n315188 , n315189 , n24764 , n315191 , n315192 , n315193 , 
 n315194 , n315195 , n24770 , n315197 , n315198 , n315199 , n24774 , n315201 , n315202 , n315203 , 
 n315204 , n315205 , n315206 , n24781 , n24782 , n315209 , n24784 , n315211 , n24786 , n24787 , 
 n315214 , n315215 , n24790 , n315217 , n315218 , n315219 , n315220 , n315221 , n24796 , n315223 , 
 n315224 , n315225 , n315226 , n315227 , n24802 , n24803 , n24804 , n315231 , n315232 , n315233 , 
 n24808 , n24809 , n315236 , n315237 , n24812 , n315239 , n315240 , n315241 , n24816 , n315243 , 
 n24818 , n315245 , n315246 , n315247 , n315248 , n315249 , n315250 , n315251 , n315252 , n24827 , 
 n24828 , n315255 , n315256 , n315257 , n24832 , n24833 , n315260 , n315261 , n315262 , n315263 , 
 n315264 , n24839 , n315266 , n24841 , n24842 , n315269 , n315270 , n24845 , n24846 , n315273 , 
 n315274 , n315275 , n315276 , n315277 , n315278 , n24853 , n315280 , n315281 , n315282 , n315283 , 
 n24858 , n315285 , n315286 , n315287 , n315288 , n24863 , n315290 , n315291 , n315292 , n315293 , 
 n24868 , n315295 , n315296 , n24871 , n315298 , n315299 , n24874 , n315301 , n315302 , n315303 , 
 n24878 , n315305 , n315306 , n315307 , n315308 , n24883 , n315310 , n315311 , n315312 , n315313 , 
 n315314 , n315315 , n315316 , n315317 , n315318 , n315319 , n24894 , n24895 , n315322 , n24897 , 
 n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n315332 , n315333 , 
 n24908 , n24909 , n24910 , n315337 , n24912 , n24913 , n315340 , n24915 , n315342 , n315343 , 
 n315344 , n315345 , n24920 , n315347 , n315348 , n315349 , n315350 , n315351 , n315352 , n315353 , 
 n315354 , n315355 , n24930 , n315357 , n315358 , n315359 , n315360 , n315361 , n315362 , n315363 , 
 n315364 , n24939 , n315366 , n315367 , n315368 , n315369 , n315370 , n24945 , n315372 , n315373 , 
 n24948 , n315375 , n315376 , n24951 , n315378 , n315379 , n315380 , n315381 , n315382 , n315383 , 
 n315384 , n315385 , n315386 , n24961 , n315388 , n315389 , n24964 , n315391 , n315392 , n315393 , 
 n315394 , n315395 , n315396 , n315397 , n24972 , n315399 , n315400 , n315401 , n315402 , n24977 , 
 n315404 , n24979 , n24980 , n315407 , n315408 , n315409 , n315410 , n315411 , n315412 , n315413 , 
 n315414 , n315415 , n24990 , n315417 , n315418 , n315419 , n315420 , n315421 , n24996 , n24997 , 
 n315424 , n315425 , n315426 , n315427 , n25002 , n25003 , n315430 , n315431 , n315432 , n315433 , 
 n315434 , n315435 , n315436 , n25011 , n315438 , n315439 , n315440 , n315441 , n315442 , n315443 , 
 n315444 , n315445 , n315446 , n25021 , n315448 , n315449 , n25024 , n315451 , n25026 , n315453 , 
 n25028 , n25029 , n315456 , n25031 , n315458 , n25033 , n25034 , n315461 , n315462 , n25037 , 
 n25038 , n25039 , n315466 , n315467 , n315468 , n315469 , n315470 , n315471 , n25046 , n315473 , 
 n315474 , n25049 , n315476 , n315477 , n315478 , n25053 , n315480 , n315481 , n315482 , n315483 , 
 n315484 , n315485 , n315486 , n315487 , n25062 , n315489 , n315490 , n315491 , n315492 , n315493 , 
 n25068 , n315495 , n315496 , n25071 , n315498 , n315499 , n315500 , n315501 , n315502 , n315503 , 
 n315504 , n315505 , n315506 , n315507 , n315508 , n315509 , n315510 , n315511 , n315512 , n315513 , 
 n315514 , n315515 , n315516 , n25091 , n315518 , n315519 , n315520 , n315521 , n315522 , n315523 , 
 n315524 , n315525 , n315526 , n315527 , n315528 , n315529 , n315530 , n315531 , n315532 , n25107 , 
 n315534 , n315535 , n315536 , n315537 , n315538 , n315539 , n315540 , n315541 , n315542 , n315543 , 
 n315544 , n315545 , n315546 , n315547 , n25122 , n315549 , n315550 , n315551 , n315552 , n315553 , 
 n315554 , n315555 , n25130 , n25131 , n315558 , n315559 , n315560 , n315561 , n315562 , n25137 , 
 n315564 , n315565 , n315566 , n315567 , n25142 , n315569 , n315570 , n315571 , n315572 , n25147 , 
 n25148 , n315575 , n315576 , n25151 , n315578 , n315579 , n25154 , n315581 , n315582 , n315583 , 
 n315584 , n315585 , n315586 , n315587 , n315588 , n315589 , n315590 , n315591 , n315592 , n315593 , 
 n315594 , n25169 , n315596 , n25171 , n315598 , n315599 , n315600 , n315601 , n25176 , n25177 , 
 n25178 , n25179 , n315606 , n315607 , n25182 , n315609 , n315610 , n315611 , n315612 , n25187 , 
 n315614 , n315615 , n315616 , n25191 , n315618 , n25193 , n25194 , n25195 , n25196 , n315623 , 
 n315624 , n315625 , n315626 , n315627 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , 
 n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n315642 , n25217 , 
 n315644 , n315645 , n315646 , n315647 , n315648 , n315649 , n315650 , n315651 , n315652 , n315653 , 
 n315654 , n315655 , n315656 , n315657 , n315658 , n25233 , n315660 , n315661 , n25236 , n315663 , 
 n315664 , n315665 , n315666 , n315667 , n25242 , n315669 , n315670 , n25245 , n315672 , n25247 , 
 n315674 , n315675 , n315676 , n25251 , n315678 , n315679 , n25254 , n315681 , n315682 , n25257 , 
 n315684 , n315685 , n25260 , n315687 , n25262 , n315689 , n315690 , n315691 , n25266 , n315693 , 
 n315694 , n315695 , n315696 , n315697 , n25272 , n315699 , n315700 , n315701 , n315702 , n315703 , 
 n25278 , n315705 , n315706 , n25281 , n315708 , n315709 , n25284 , n25285 , n315712 , n25287 , 
 n315714 , n25289 , n315716 , n315717 , n315718 , n315719 , n315720 , n315721 , n315722 , n315723 , 
 n315724 , n315725 , n315726 , n315727 , n315728 , n315729 , n315730 , n315731 , n25306 , n315733 , 
 n315734 , n25309 , n315736 , n315737 , n315738 , n315739 , n315740 , n315741 , n25316 , n315743 , 
 n315744 , n315745 , n315746 , n315747 , n315748 , n315749 , n315750 , n25325 , n315752 , n315753 , 
 n25328 , n315755 , n315756 , n25331 , n25332 , n25333 , n315760 , n25335 , n25336 , n315763 , 
 n25338 , n315765 , n315766 , n25341 , n315768 , n25343 , n315770 , n315771 , n25346 , n315773 , 
 n315774 , n315775 , n315776 , n315777 , n315778 , n25353 , n315780 , n315781 , n25356 , n25357 , 
 n25358 , n315785 , n25360 , n25361 , n315788 , n315789 , n25364 , n315791 , n315792 , n315793 , 
 n315794 , n315795 , n315796 , n25371 , n315798 , n25373 , n25374 , n25375 , n315802 , n315803 , 
 n315804 , n315805 , n315806 , n315807 , n315808 , n315809 , n25384 , n315811 , n315812 , n315813 , 
 n315814 , n315815 , n315816 , n315817 , n315818 , n315819 , n315820 , n315821 , n315822 , n315823 , 
 n315824 , n25399 , n25400 , n315827 , n315828 , n315829 , n25404 , n315831 , n315832 , n25407 , 
 n315834 , n315835 , n25410 , n315837 , n315838 , n315839 , n315840 , n315841 , n315842 , n315843 , 
 n315844 , n315845 , n315846 , n315847 , n315848 , n25423 , n315850 , n315851 , n315852 , n315853 , 
 n315854 , n315855 , n315856 , n25431 , n315858 , n315859 , n25434 , n315861 , n315862 , n25437 , 
 n315864 , n315865 , n315866 , n315867 , n315868 , n315869 , n315870 , n315871 , n315872 , n315873 , 
 n315874 , n315875 , n315876 , n315877 , n315878 , n25453 , n315880 , n315881 , n315882 , n315883 , 
 n315884 , n315885 , n25460 , n315887 , n25462 , n315889 , n315890 , n315891 , n25466 , n315893 , 
 n25468 , n315895 , n315896 , n315897 , n315898 , n315899 , n315900 , n315901 , n315902 , n315903 , 
 n25478 , n315905 , n315906 , n25481 , n315908 , n315909 , n315910 , n25485 , n315912 , n315913 , 
 n25488 , n315915 , n315916 , n315917 , n315918 , n315919 , n315920 , n25495 , n315922 , n315923 , 
 n315924 , n315925 , n315926 , n315927 , n25502 , n315929 , n315930 , n25505 , n315932 , n315933 , 
 n315934 , n315935 , n315936 , n315937 , n25512 , n315939 , n315940 , n25515 , n315942 , n315943 , 
 n25518 , n25519 , n25520 , n25521 , n315948 , n25523 , n315950 , n315951 , n315952 , n315953 , 
 n315954 , n315955 , n315956 , n315957 , n315958 , n315959 , n315960 , n315961 , n315962 , n315963 , 
 n315964 , n315965 , n315966 , n315967 , n25542 , n25543 , n315970 , n25545 , n315972 , n315973 , 
 n25548 , n315975 , n315976 , n315977 , n25552 , n315979 , n315980 , n25555 , n315982 , n315983 , 
 n315984 , n315985 , n315986 , n315987 , n315988 , n315989 , n315990 , n315991 , n315992 , n315993 , 
 n315994 , n315995 , n315996 , n315997 , n315998 , n25573 , n25574 , n316001 , n316002 , n25577 , 
 n316004 , n25579 , n316006 , n316007 , n316008 , n316009 , n25584 , n316011 , n316012 , n316013 , 
 n316014 , n316015 , n316016 , n25591 , n316018 , n316019 , n316020 , n316021 , n316022 , n316023 , 
 n25598 , n316025 , n316026 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , 
 n316034 , n316035 , n316036 , n316037 , n316038 , n316039 , n316040 , n316041 , n316042 , n316043 , 
 n316044 , n316045 , n316046 , n316047 , n316048 , n25623 , n316050 , n316051 , n25626 , n316053 , 
 n316054 , n316055 , n316056 , n25631 , n316058 , n316059 , n25634 , n316061 , n316062 , n316063 , 
 n316064 , n316065 , n316066 , n25641 , n25642 , n316069 , n316070 , n316071 , n316072 , n316073 , 
 n316074 , n316075 , n316076 , n316077 , n316078 , n316079 , n25654 , n316081 , n25656 , n316083 , 
 n316084 , n316085 , n316086 , n316087 , n25662 , n316089 , n316090 , n316091 , n25666 , n316093 , 
 n316094 , n316095 , n316096 , n316097 , n25672 , n25673 , n316100 , n316101 , n25676 , n316103 , 
 n25678 , n316105 , n316106 , n316107 , n316108 , n316109 , n316110 , n316111 , n25686 , n316113 , 
 n316114 , n316115 , n316116 , n316117 , n316118 , n25693 , n316120 , n316121 , n25696 , n316123 , 
 n25698 , n316125 , n316126 , n316127 , n316128 , n316129 , n316130 , n316131 , n316132 , n316133 , 
 n316134 , n316135 , n316136 , n25711 , n25712 , n316139 , n316140 , n25715 , n316142 , n316143 , 
 n316144 , n316145 , n25720 , n25721 , n25722 , n316149 , n316150 , n316151 , n316152 , n25727 , 
 n316154 , n316155 , n316156 , n316157 , n25732 , n25733 , n25734 , n316161 , n316162 , n316163 , 
 n316164 , n316165 , n316166 , n316167 , n316168 , n316169 , n316170 , n316171 , n316172 , n316173 , 
 n25748 , n316175 , n316176 , n25751 , n316178 , n316179 , n316180 , n25755 , n316182 , n316183 , 
 n25758 , n316185 , n316186 , n316187 , n316188 , n316189 , n316190 , n316191 , n316192 , n316193 , 
 n25768 , n316195 , n316196 , n316197 , n316198 , n316199 , n316200 , n316201 , n316202 , n316203 , 
 n316204 , n316205 , n316206 , n316207 , n316208 , n316209 , n316210 , n316211 , n316212 , n316213 , 
 n316214 , n316215 , n316216 , n316217 , n316218 , n316219 , n316220 , n316221 , n316222 , n316223 , 
 n25798 , n316225 , n316226 , n316227 , n316228 , n316229 , n316230 , n316231 , n316232 , n316233 , 
 n316234 , n316235 , n316236 , n316237 , n316238 , n316239 , n316240 , n316241 , n316242 , n316243 , 
 n316244 , n25819 , n316246 , n316247 , n25822 , n316249 , n316250 , n25825 , n25826 , n316253 , 
 n316254 , n25829 , n316256 , n316257 , n25832 , n316259 , n316260 , n25835 , n316262 , n316263 , 
 n25838 , n316265 , n316266 , n316267 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , 
 n25848 , n25849 , n316276 , n316277 , n316278 , n316279 , n25854 , n25855 , n25856 , n25857 , 
 n25858 , n316285 , n316286 , n316287 , n25862 , n25863 , n316290 , n316291 , n316292 , n25867 , 
 n25868 , n316295 , n316296 , n316297 , n25872 , n25873 , n316300 , n316301 , n316302 , n25877 , 
 n25878 , n316305 , n316306 , n316307 , n316308 , n316309 , n316310 , n316311 , n316312 , n316313 , 
 n316314 , n316315 , n316316 , n316317 , n316318 , n316319 , n316320 , n316321 , n316322 , n316323 , 
 n316324 , n316325 , n316326 , n316327 , n25902 , n316329 , n316330 , n316331 , n316332 , n316333 , 
 n316334 , n316335 , n316336 , n316337 , n316338 , n316339 , n316340 , n316341 , n316342 , n316343 , 
 n316344 , n316345 , n316346 , n316347 , n316348 , n316349 , n316350 , n316351 , n316352 , n316353 , 
 n316354 , n316355 , n316356 , n316357 , n316358 , n316359 , n316360 , n25935 , n316362 , n316363 , 
 n316364 , n316365 , n316366 , n316367 , n25942 , n316369 , n316370 , n25945 , n316372 , n316373 , 
 n25948 , n316375 , n316376 , n316377 , n316378 , n316379 , n25954 , n316381 , n25956 , n25957 , 
 n316384 , n316385 , n25960 , n316387 , n25962 , n25963 , n25964 , n316391 , n316392 , n316393 , 
 n316394 , n316395 , n316396 , n316397 , n316398 , n25973 , n316400 , n316401 , n25976 , n316403 , 
 n316404 , n25979 , n316406 , n316407 , n316408 , n316409 , n316410 , n316411 , n25986 , n316413 , 
 n316414 , n25989 , n25990 , n316417 , n316418 , n25993 , n316420 , n316421 , n25996 , n316423 , 
 n316424 , n316425 , n316426 , n316427 , n26002 , n26003 , n316430 , n316431 , n316432 , n26007 , 
 n316434 , n316435 , n26010 , n316437 , n316438 , n316439 , n316440 , n316441 , n26016 , n26017 , 
 n316444 , n26019 , n26020 , n26021 , n316448 , n26023 , n26024 , n316451 , n26026 , n316453 , 
 n26028 , n316455 , n316456 , n316457 , n316458 , n316459 , n26034 , n316461 , n26036 , n316463 , 
 n316464 , n316465 , n316466 , n316467 , n316468 , n26043 , n26044 , n316471 , n26046 , n316473 , 
 n316474 , n26049 , n316476 , n316477 , n26052 , n316479 , n316480 , n26055 , n316482 , n316483 , 
 n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n316490 , n316491 , n316492 , n316493 , 
 n316494 , n316495 , n316496 , n316497 , n26072 , n316499 , n316500 , n26075 , n316502 , n316503 , 
 n316504 , n316505 , n316506 , n26081 , n316508 , n316509 , n316510 , n26085 , n316512 , n316513 , 
 n26088 , n316515 , n316516 , n26091 , n316518 , n316519 , n316520 , n26095 , n316522 , n316523 , 
 n316524 , n316525 , n316526 , n316527 , n26102 , n316529 , n316530 , n26105 , n316532 , n26107 , 
 n316534 , n316535 , n316536 , n316537 , n316538 , n316539 , n26114 , n316541 , n26116 , n316543 , 
 n316544 , n316545 , n316546 , n26121 , n316548 , n316549 , n26124 , n316551 , n316552 , n316553 , 
 n316554 , n316555 , n316556 , n26131 , n316558 , n316559 , n316560 , n316561 , n316562 , n26137 , 
 n316564 , n316565 , n26140 , n316567 , n316568 , n26143 , n26144 , n316571 , n26146 , n26147 , 
 n316574 , n316575 , n26150 , n316577 , n316578 , n316579 , n26154 , n26155 , n316582 , n26157 , 
 n26158 , n26159 , n316586 , n26161 , n316588 , n316589 , n316590 , n316591 , n26166 , n316593 , 
 n26168 , n26169 , n316596 , n316597 , n26172 , n316599 , n316600 , n26175 , n316602 , n316603 , 
 n316604 , n316605 , n316606 , n316607 , n316608 , n316609 , n316610 , n316611 , n26186 , n316613 , 
 n316614 , n316615 , n316616 , n316617 , n26192 , n316619 , n316620 , n316621 , n316622 , n316623 , 
 n26198 , n316625 , n316626 , n26201 , n316628 , n316629 , n26204 , n26205 , n316632 , n316633 , 
 n26208 , n316635 , n316636 , n26211 , n316638 , n316639 , n26214 , n316641 , n316642 , n26217 , 
 n316644 , n316645 , n26220 , n316647 , n316648 , n316649 , n316650 , n26225 , n316652 , n26227 , 
 n26228 , n26229 , n26230 , n26231 , n26232 , n316659 , n316660 , n316661 , n316662 , n316663 , 
 n316664 , n316665 , n316666 , n316667 , n316668 , n316669 , n26244 , n26245 , n316672 , n316673 , 
 n316674 , n316675 , n26250 , n316677 , n26252 , n26253 , n26254 , n26255 , n316682 , n26257 , 
 n26258 , n316685 , n316686 , n316687 , n316688 , n26263 , n316690 , n316691 , n316692 , n316693 , 
 n316694 , n26269 , n316696 , n316697 , n316698 , n316699 , n316700 , n316701 , n316702 , n316703 , 
 n316704 , n316705 , n316706 , n316707 , n316708 , n316709 , n26284 , n316711 , n316712 , n26287 , 
 n316714 , n316715 , n316716 , n26291 , n316718 , n316719 , n26294 , n316721 , n316722 , n26297 , 
 n26298 , n316725 , n26300 , n316727 , n316728 , n316729 , n26304 , n26305 , n316732 , n316733 , 
 n316734 , n26309 , n316736 , n316737 , n316738 , n316739 , n316740 , n316741 , n316742 , n316743 , 
 n316744 , n316745 , n316746 , n316747 , n316748 , n316749 , n316750 , n26325 , n316752 , n316753 , 
 n26328 , n316755 , n26330 , n316757 , n316758 , n316759 , n316760 , n316761 , n316762 , n316763 , 
 n316764 , n316765 , n316766 , n316767 , n26342 , n26343 , n316770 , n316771 , n26346 , n26347 , 
 n316774 , n316775 , n316776 , n316777 , n316778 , n26353 , n316780 , n26355 , n316782 , n316783 , 
 n316784 , n316785 , n316786 , n316787 , n26362 , n316789 , n316790 , n316791 , n316792 , n26367 , 
 n316794 , n316795 , n26370 , n316797 , n316798 , n26373 , n26374 , n316801 , n316802 , n316803 , 
 n316804 , n26379 , n316806 , n316807 , n26382 , n26383 , n316810 , n316811 , n316812 , n316813 , 
 n26388 , n316815 , n316816 , n316817 , n26392 , n316819 , n316820 , n316821 , n316822 , n26397 , 
 n316824 , n316825 , n316826 , n316827 , n316828 , n316829 , n26404 , n316831 , n26406 , n316833 , 
 n316834 , n316835 , n316836 , n26411 , n316838 , n316839 , n316840 , n316841 , n316842 , n26417 , 
 n316844 , n316845 , n26420 , n316847 , n26422 , n316849 , n316850 , n26425 , n316852 , n316853 , 
 n26428 , n316855 , n316856 , n316857 , n316858 , n316859 , n316860 , n316861 , n316862 , n316863 , 
 n26438 , n316865 , n316866 , n316867 , n316868 , n316869 , n316870 , n316871 , n316872 , n26447 , 
 n26448 , n26449 , n316876 , n316877 , n316878 , n316879 , n316880 , n316881 , n26456 , n316883 , 
 n316884 , n316885 , n316886 , n316887 , n316888 , n316889 , n316890 , n316891 , n26466 , n316893 , 
 n316894 , n316895 , n316896 , n316897 , n316898 , n316899 , n316900 , n316901 , n26476 , n316903 , 
 n316904 , n26479 , n316906 , n316907 , n26482 , n316909 , n316910 , n316911 , n26486 , n316913 , 
 n316914 , n26489 , n316916 , n316917 , n316918 , n316919 , n316920 , n316921 , n316922 , n316923 , 
 n26498 , n26499 , n316926 , n316927 , n316928 , n316929 , n316930 , n316931 , n316932 , n316933 , 
 n316934 , n316935 , n316936 , n316937 , n316938 , n316939 , n26514 , n26515 , n316942 , n316943 , 
 n316944 , n26519 , n316946 , n316947 , n316948 , n316949 , n316950 , n316951 , n316952 , n26527 , 
 n316954 , n316955 , n316956 , n316957 , n316958 , n316959 , n26534 , n316961 , n316962 , n316963 , 
 n26538 , n316965 , n316966 , n316967 , n316968 , n316969 , n316970 , n26545 , n316972 , n316973 , 
 n26548 , n316975 , n316976 , n26551 , n316978 , n316979 , n26554 , n316981 , n316982 , n26557 , 
 n316984 , n316985 , n26560 , n316987 , n316988 , n316989 , n316990 , n316991 , n26566 , n316993 , 
 n316994 , n316995 , n316996 , n316997 , n316998 , n316999 , n317000 , n26575 , n317002 , n317003 , 
 n317004 , n317005 , n317006 , n317007 , n317008 , n317009 , n317010 , n317011 , n317012 , n317013 , 
 n317014 , n317015 , n317016 , n317017 , n317018 , n26593 , n317020 , n317021 , n26596 , n26597 , 
 n26598 , n317025 , n26600 , n317027 , n317028 , n317029 , n317030 , n317031 , n317032 , n317033 , 
 n317034 , n317035 , n317036 , n317037 , n317038 , n317039 , n317040 , n317041 , n317042 , n317043 , 
 n317044 , n317045 , n317046 , n26621 , n317048 , n317049 , n26624 , n317051 , n317052 , n317053 , 
 n26628 , n317055 , n317056 , n317057 , n317058 , n317059 , n26634 , n317061 , n317062 , n26637 , 
 n26638 , n26639 , n317066 , n317067 , n317068 , n26643 , n317070 , n26645 , n26646 , n317073 , 
 n26648 , n26649 , n317076 , n317077 , n26652 , n317079 , n317080 , n317081 , n317082 , n26657 , 
 n317084 , n26659 , n317086 , n317087 , n317088 , n317089 , n26664 , n317091 , n317092 , n317093 , 
 n317094 , n317095 , n317096 , n317097 , n317098 , n26673 , n26674 , n317101 , n317102 , n317103 , 
 n317104 , n26679 , n317106 , n317107 , n317108 , n317109 , n317110 , n317111 , n317112 , n317113 , 
 n317114 , n317115 , n317116 , n317117 , n317118 , n317119 , n317120 , n317121 , n317122 , n317123 , 
 n26698 , n317125 , n317126 , n317127 , n317128 , n317129 , n26704 , n317131 , n317132 , n26707 , 
 n317134 , n317135 , n317136 , n317137 , n317138 , n317139 , n317140 , n317141 , n26716 , n317143 , 
 n317144 , n317145 , n317146 , n317147 , n317148 , n317149 , n317150 , n317151 , n26726 , n317153 , 
 n317154 , n26729 , n317156 , n317157 , n317158 , n26733 , n26734 , n317161 , n317162 , n317163 , 
 n317164 , n317165 , n26740 , n26741 , n26742 , n317169 , n317170 , n317171 , n317172 , n26747 , 
 n317174 , n317175 , n317176 , n317177 , n26752 , n26753 , n317180 , n317181 , n26756 , n26757 , 
 n317184 , n317185 , n317186 , n317187 , n317188 , n317189 , n317190 , n317191 , n317192 , n317193 , 
 n317194 , n317195 , n317196 , n317197 , n317198 , n317199 , n26774 , n317201 , n317202 , n317203 , 
 n317204 , n26779 , n26780 , n26781 , n26782 , n317209 , n317210 , n26785 , n317212 , n317213 , 
 n317214 , n26789 , n317216 , n317217 , n26792 , n26793 , n317220 , n317221 , n317222 , n26797 , 
 n317224 , n317225 , n317226 , n317227 , n317228 , n317229 , n317230 , n317231 , n317232 , n317233 , 
 n317234 , n317235 , n26810 , n317237 , n317238 , n26813 , n26814 , n317241 , n26816 , n317243 , 
 n317244 , n317245 , n317246 , n317247 , n317248 , n317249 , n317250 , n26825 , n317252 , n317253 , 
 n317254 , n317255 , n317256 , n317257 , n317258 , n317259 , n317260 , n26835 , n317262 , n317263 , 
 n26838 , n317265 , n26840 , n26841 , n317268 , n317269 , n317270 , n317271 , n317272 , n317273 , 
 n317274 , n26849 , n317276 , n317277 , n26852 , n317279 , n317280 , n317281 , n317282 , n317283 , 
 n317284 , n317285 , n317286 , n26861 , n317288 , n26863 , n317290 , n317291 , n317292 , n317293 , 
 n26868 , n317295 , n317296 , n26871 , n26872 , n317299 , n317300 , n317301 , n317302 , n317303 , 
 n26878 , n317305 , n317306 , n317307 , n317308 , n26883 , n317310 , n317311 , n317312 , n317313 , 
 n26888 , n317315 , n317316 , n26891 , n317318 , n317319 , n26894 , n317321 , n317322 , n317323 , 
 n317324 , n317325 , n317326 , n317327 , n317328 , n317329 , n317330 , n317331 , n317332 , n317333 , 
 n317334 , n26909 , n317336 , n317337 , n317338 , n26913 , n26914 , n317341 , n26916 , n317343 , 
 n317344 , n317345 , n317346 , n317347 , n317348 , n317349 , n317350 , n317351 , n317352 , n26927 , 
 n317354 , n317355 , n317356 , n26931 , n317358 , n317359 , n317360 , n317361 , n317362 , n26937 , 
 n317364 , n317365 , n26940 , n317367 , n317368 , n26943 , n317370 , n317371 , n26946 , n317373 , 
 n317374 , n26949 , n317376 , n317377 , n26952 , n317379 , n317380 , n317381 , n317382 , n317383 , 
 n317384 , n317385 , n26960 , n317387 , n317388 , n317389 , n317390 , n317391 , n317392 , n317393 , 
 n26968 , n317395 , n26970 , n317397 , n317398 , n317399 , n317400 , n317401 , n317402 , n26977 , 
 n317404 , n317405 , n317406 , n317407 , n317408 , n317409 , n317410 , n317411 , n317412 , n317413 , 
 n317414 , n317415 , n317416 , n26991 , n317418 , n317419 , n26994 , n317421 , n26996 , n317423 , 
 n317424 , n317425 , n317426 , n317427 , n27002 , n317429 , n317430 , n317431 , n317432 , n27007 , 
 n317434 , n27009 , n317436 , n317437 , n317438 , n317439 , n317440 , n27015 , n317442 , n317443 , 
 n317444 , n317445 , n27020 , n27021 , n27022 , n317449 , n317450 , n27025 , n317452 , n317453 , 
 n27028 , n317455 , n317456 , n317457 , n317458 , n27033 , n317460 , n317461 , n317462 , n27037 , 
 n27038 , n317465 , n27040 , n27041 , n317468 , n317469 , n27044 , n27045 , n317472 , n317473 , 
 n317474 , n27049 , n317476 , n317477 , n317478 , n317479 , n317480 , n317481 , n27056 , n317483 , 
 n317484 , n317485 , n27060 , n317487 , n317488 , n27063 , n317490 , n317491 , n317492 , n317493 , 
 n317494 , n317495 , n317496 , n317497 , n317498 , n317499 , n317500 , n27075 , n317502 , n317503 , 
 n27078 , n317505 , n317506 , n317507 , n317508 , n317509 , n27084 , n317511 , n317512 , n317513 , 
 n317514 , n317515 , n317516 , n317517 , n317518 , n317519 , n317520 , n317521 , n27096 , n317523 , 
 n317524 , n317525 , n317526 , n317527 , n317528 , n317529 , n317530 , n317531 , n317532 , n317533 , 
 n317534 , n317535 , n317536 , n317537 , n317538 , n317539 , n317540 , n317541 , n317542 , n27117 , 
 n317544 , n317545 , n27120 , n317547 , n317548 , n317549 , n317550 , n27125 , n317552 , n317553 , 
 n317554 , n317555 , n317556 , n27131 , n317558 , n317559 , n317560 , n317561 , n27136 , n317563 , 
 n27138 , n317565 , n317566 , n317567 , n27142 , n317569 , n317570 , n317571 , n27146 , n317573 , 
 n317574 , n27149 , n317576 , n317577 , n27152 , n317579 , n317580 , n317581 , n317582 , n317583 , 
 n317584 , n317585 , n317586 , n317587 , n317588 , n27163 , n317590 , n317591 , n27166 , n27167 , 
 n317594 , n317595 , n317596 , n27171 , n317598 , n317599 , n317600 , n317601 , n27176 , n27177 , 
 n317604 , n317605 , n317606 , n27181 , n317608 , n27183 , n317610 , n27185 , n317612 , n317613 , 
 n27188 , n317615 , n27190 , n317617 , n27192 , n317619 , n317620 , n27195 , n317622 , n317623 , 
 n317624 , n27199 , n317626 , n27201 , n317628 , n317629 , n317630 , n27205 , n317632 , n317633 , 
 n27208 , n317635 , n27210 , n317637 , n317638 , n317639 , n27214 , n317641 , n317642 , n317643 , 
 n317644 , n317645 , n317646 , n27221 , n317648 , n317649 , n317650 , n317651 , n317652 , n27227 , 
 n27228 , n317655 , n27230 , n317657 , n317658 , n317659 , n317660 , n317661 , n317662 , n317663 , 
 n317664 , n317665 , n317666 , n317667 , n27242 , n317669 , n317670 , n317671 , n317672 , n317673 , 
 n317674 , n317675 , n317676 , n317677 , n317678 , n317679 , n27254 , n317681 , n317682 , n317683 , 
 n27258 , n317685 , n317686 , n317687 , n317688 , n317689 , n317690 , n317691 , n317692 , n317693 , 
 n317694 , n317695 , n317696 , n27271 , n317698 , n317699 , n27274 , n317701 , n317702 , n317703 , 
 n317704 , n317705 , n317706 , n317707 , n317708 , n317709 , n317710 , n317711 , n317712 , n317713 , 
 n317714 , n27289 , n317716 , n317717 , n27292 , n317719 , n317720 , n317721 , n317722 , n317723 , 
 n317724 , n317725 , n317726 , n317727 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , 
 n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n317740 , n317741 , n317742 , n317743 , 
 n27318 , n317745 , n317746 , n317747 , n27322 , n317749 , n317750 , n27325 , n317752 , n317753 , 
 n27328 , n317755 , n27330 , n317757 , n317758 , n27333 , n317760 , n317761 , n27336 , n317763 , 
 n317764 , n317765 , n317766 , n317767 , n317768 , n317769 , n317770 , n317771 , n27346 , n317773 , 
 n317774 , n27349 , n317776 , n317777 , n27352 , n317779 , n317780 , n317781 , n317782 , n317783 , 
 n317784 , n317785 , n317786 , n317787 , n27362 , n317789 , n317790 , n317791 , n317792 , n317793 , 
 n27368 , n317795 , n317796 , n27371 , n317798 , n27373 , n27374 , n317801 , n317802 , n27377 , 
 n317804 , n317805 , n317806 , n317807 , n317808 , n317809 , n27384 , n27385 , n317812 , n317813 , 
 n27388 , n317815 , n317816 , n317817 , n317818 , n317819 , n317820 , n27395 , n317822 , n317823 , 
 n317824 , n27399 , n317826 , n317827 , n317828 , n317829 , n317830 , n317831 , n27406 , n317833 , 
 n317834 , n27409 , n317836 , n317837 , n27412 , n317839 , n317840 , n27415 , n27416 , n317843 , 
 n27418 , n317845 , n317846 , n317847 , n317848 , n317849 , n317850 , n317851 , n317852 , n317853 , 
 n27428 , n317855 , n317856 , n317857 , n317858 , n317859 , n317860 , n317861 , n317862 , n317863 , 
 n317864 , n317865 , n27440 , n317867 , n27442 , n317869 , n27444 , n317871 , n317872 , n317873 , 
 n317874 , n317875 , n317876 , n317877 , n317878 , n317879 , n317880 , n317881 , n317882 , n27457 , 
 n317884 , n317885 , n317886 , n317887 , n27462 , n27463 , n27464 , n317891 , n317892 , n317893 , 
 n317894 , n317895 , n317896 , n27471 , n317898 , n317899 , n317900 , n317901 , n317902 , n317903 , 
 n317904 , n317905 , n317906 , n317907 , n317908 , n317909 , n317910 , n317911 , n317912 , n27487 , 
 n317914 , n317915 , n27490 , n317917 , n317918 , n27493 , n317920 , n317921 , n27496 , n317923 , 
 n317924 , n317925 , n27500 , n317927 , n317928 , n27503 , n317930 , n27505 , n27506 , n317933 , 
 n27508 , n27509 , n27510 , n317937 , n317938 , n317939 , n27514 , n27515 , n317942 , n317943 , 
 n317944 , n317945 , n317946 , n317947 , n317948 , n317949 , n27524 , n317951 , n317952 , n27527 , 
 n317954 , n317955 , n27530 , n317957 , n317958 , n317959 , n27534 , n317961 , n317962 , n27537 , 
 n317964 , n317965 , n317966 , n27541 , n27542 , n27543 , n317970 , n317971 , n317972 , n27547 , 
 n317974 , n317975 , n27550 , n317977 , n27552 , n27553 , n317980 , n317981 , n317982 , n27557 , 
 n317984 , n317985 , n27560 , n317987 , n317988 , n317989 , n27564 , n317991 , n317992 , n317993 , 
 n27568 , n317995 , n317996 , n317997 , n317998 , n27573 , n318000 , n318001 , n27576 , n318003 , 
 n318004 , n318005 , n27580 , n318007 , n27582 , n318009 , n318010 , n27585 , n318012 , n318013 , 
 n27588 , n27589 , n318016 , n318017 , n27592 , n27593 , n27594 , n318021 , n318022 , n27597 , 
 n318024 , n318025 , n27600 , n318027 , n318028 , n318029 , n318030 , n27605 , n318032 , n27607 , 
 n318034 , n318035 , n318036 , n318037 , n27612 , n318039 , n318040 , n318041 , n27616 , n318043 , 
 n318044 , n318045 , n27620 , n318047 , n318048 , n318049 , n27624 , n27625 , n318052 , n27627 , 
 n318054 , n27629 , n318056 , n318057 , n318058 , n318059 , n318060 , n27635 , n318062 , n318063 , 
 n27638 , n318065 , n318066 , n318067 , n318068 , n318069 , n27644 , n318071 , n318072 , n318073 , 
 n318074 , n27649 , n318076 , n27651 , n318078 , n318079 , n318080 , n318081 , n318082 , n27657 , 
 n318084 , n318085 , n318086 , n318087 , n27662 , n318089 , n318090 , n318091 , n318092 , n27667 , 
 n318094 , n318095 , n318096 , n318097 , n27672 , n318099 , n318100 , n318101 , n318102 , n27677 , 
 n318104 , n318105 , n318106 , n318107 , n27682 , n318109 , n318110 , n27685 , n318112 , n318113 , 
 n27688 , n318115 , n318116 , n318117 , n318118 , n27693 , n318120 , n318121 , n27696 , n27697 , 
 n318124 , n318125 , n318126 , n27701 , n318128 , n318129 , n27704 , n318131 , n318132 , n27707 , 
 n27708 , n318135 , n27710 , n318137 , n318138 , n318139 , n318140 , n318141 , n27716 , n318143 , 
 n318144 , n27719 , n318146 , n318147 , n318148 , n318149 , n318150 , n27725 , n318152 , n318153 , 
 n318154 , n318155 , n27730 , n318157 , n318158 , n27733 , n318160 , n318161 , n318162 , n318163 , 
 n318164 , n318165 , n318166 , n318167 , n318168 , n318169 , n318170 , n318171 , n318172 , n318173 , 
 n318174 , n318175 , n27750 , n318177 , n318178 , n27753 , n318180 , n318181 , n318182 , n318183 , 
 n27758 , n318185 , n318186 , n318187 , n318188 , n27763 , n318190 , n318191 , n318192 , n27767 , 
 n27768 , n318195 , n318196 , n318197 , n27772 , n318199 , n318200 , n27775 , n318202 , n27777 , 
 n318204 , n318205 , n27780 , n318207 , n318208 , n318209 , n318210 , n27785 , n27786 , n318213 , 
 n318214 , n318215 , n318216 , n318217 , n318218 , n27793 , n318220 , n318221 , n27796 , n318223 , 
 n318224 , n318225 , n318226 , n318227 , n27802 , n318229 , n318230 , n27805 , n318232 , n318233 , 
 n318234 , n318235 , n318236 , n318237 , n27812 , n318239 , n318240 , n27815 , n318242 , n318243 , 
 n27818 , n318245 , n318246 , n27821 , n27822 , n318249 , n318250 , n318251 , n27826 , n27827 , 
 n27828 , n27829 , n318256 , n27831 , n27832 , n318259 , n27834 , n318261 , n318262 , n27837 , 
 n318264 , n27839 , n27840 , n318267 , n27842 , n318269 , n318270 , n27845 , n318272 , n318273 , 
 n318274 , n27849 , n318276 , n318277 , n27852 , n318279 , n318280 , n27855 , n318282 , n318283 , 
 n318284 , n27859 , n318286 , n27861 , n27862 , n318289 , n318290 , n318291 , n27866 , n318293 , 
 n318294 , n27869 , n318296 , n318297 , n27872 , n318299 , n27874 , n318301 , n318302 , n318303 , 
 n318304 , n318305 , n318306 , n318307 , n318308 , n27883 , n318310 , n318311 , n318312 , n318313 , 
 n27888 , n318315 , n318316 , n318317 , n318318 , n318319 , n27894 , n318321 , n27896 , n318323 , 
 n318324 , n318325 , n318326 , n318327 , n318328 , n318329 , n318330 , n318331 , n318332 , n318333 , 
 n318334 , n27909 , n318336 , n318337 , n318338 , n318339 , n318340 , n318341 , n318342 , n27917 , 
 n318344 , n318345 , n318346 , n318347 , n318348 , n318349 , n318350 , n318351 , n318352 , n318353 , 
 n27928 , n318355 , n27930 , n318357 , n318358 , n318359 , n318360 , n318361 , n318362 , n318363 , 
 n318364 , n318365 , n27940 , n318367 , n318368 , n27943 , n318370 , n318371 , n318372 , n318373 , 
 n318374 , n318375 , n27950 , n318377 , n318378 , n27953 , n318380 , n318381 , n318382 , n318383 , 
 n318384 , n27959 , n318386 , n318387 , n318388 , n27963 , n318390 , n318391 , n318392 , n318393 , 
 n27968 , n318395 , n318396 , n318397 , n318398 , n318399 , n27974 , n318401 , n318402 , n318403 , 
 n318404 , n318405 , n318406 , n318407 , n318408 , n318409 , n318410 , n318411 , n27986 , n318413 , 
 n318414 , n27989 , n318416 , n318417 , n318418 , n318419 , n318420 , n318421 , n318422 , n318423 , 
 n318424 , n318425 , n318426 , n318427 , n28002 , n318429 , n318430 , n318431 , n318432 , n318433 , 
 n318434 , n318435 , n318436 , n28011 , n318438 , n28013 , n318440 , n318441 , n318442 , n318443 , 
 n318444 , n318445 , n318446 , n318447 , n318448 , n28023 , n318450 , n318451 , n318452 , n28027 , 
 n318454 , n28029 , n318456 , n318457 , n318458 , n318459 , n318460 , n318461 , n318462 , n318463 , 
 n318464 , n28039 , n318466 , n318467 , n28042 , n318469 , n318470 , n28045 , n318472 , n318473 , 
 n318474 , n28049 , n318476 , n28051 , n318478 , n318479 , n318480 , n318481 , n28056 , n318483 , 
 n318484 , n28059 , n318486 , n318487 , n28062 , n318489 , n318490 , n318491 , n28066 , n28067 , 
 n28068 , n318495 , n318496 , n318497 , n28072 , n318499 , n318500 , n318501 , n318502 , n28077 , 
 n28078 , n318505 , n28080 , n318507 , n318508 , n318509 , n318510 , n318511 , n318512 , n28087 , 
 n318514 , n318515 , n318516 , n318517 , n318518 , n318519 , n318520 , n318521 , n28096 , n318523 , 
 n318524 , n318525 , n318526 , n318527 , n28102 , n318529 , n318530 , n318531 , n318532 , n318533 , 
 n318534 , n318535 , n318536 , n318537 , n28112 , n28113 , n318540 , n318541 , n318542 , n318543 , 
 n318544 , n318545 , n318546 , n318547 , n318548 , n318549 , n318550 , n318551 , n318552 , n318553 , 
 n28128 , n318555 , n318556 , n28131 , n318558 , n28133 , n318560 , n318561 , n318562 , n318563 , 
 n318564 , n318565 , n318566 , n28141 , n318568 , n28143 , n318570 , n318571 , n318572 , n318573 , 
 n28148 , n318575 , n318576 , n28151 , n318578 , n318579 , n318580 , n318581 , n318582 , n318583 , 
 n318584 , n318585 , n318586 , n318587 , n28162 , n318589 , n318590 , n318591 , n318592 , n28167 , 
 n318594 , n318595 , n28170 , n318597 , n318598 , n318599 , n318600 , n318601 , n28176 , n28177 , 
 n318604 , n318605 , n318606 , n318607 , n318608 , n318609 , n318610 , n318611 , n318612 , n318613 , 
 n28188 , n318615 , n28190 , n28191 , n318618 , n318619 , n28194 , n318621 , n28196 , n28197 , 
 n318624 , n318625 , n318626 , n28201 , n318628 , n318629 , n318630 , n318631 , n318632 , n318633 , 
 n318634 , n28209 , n318636 , n318637 , n28212 , n318639 , n318640 , n28215 , n318642 , n318643 , 
 n28218 , n28219 , n318646 , n318647 , n318648 , n318649 , n28224 , n318651 , n318652 , n318653 , 
 n318654 , n318655 , n318656 , n318657 , n318658 , n318659 , n28234 , n318661 , n318662 , n318663 , 
 n318664 , n318665 , n318666 , n318667 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , 
 n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n318680 , n28255 , n318682 , n318683 , 
 n318684 , n28259 , n318686 , n318687 , n318688 , n28263 , n318690 , n318691 , n318692 , n318693 , 
 n28268 , n28269 , n318696 , n318697 , n318698 , n28273 , n28274 , n318701 , n318702 , n318703 , 
 n28278 , n318705 , n318706 , n318707 , n28282 , n28283 , n318710 , n318711 , n28286 , n318713 , 
 n318714 , n318715 , n28290 , n318717 , n28292 , n318719 , n318720 , n318721 , n318722 , n318723 , 
 n318724 , n318725 , n318726 , n318727 , n318728 , n318729 , n318730 , n28305 , n318732 , n318733 , 
 n318734 , n318735 , n318736 , n28311 , n318738 , n28313 , n318740 , n318741 , n318742 , n318743 , 
 n28318 , n318745 , n318746 , n28321 , n318748 , n318749 , n318750 , n28325 , n318752 , n318753 , 
 n28328 , n318755 , n318756 , n28331 , n318758 , n318759 , n318760 , n318761 , n28336 , n318763 , 
 n318764 , n318765 , n318766 , n318767 , n318768 , n28343 , n318770 , n318771 , n28346 , n318773 , 
 n318774 , n318775 , n318776 , n28351 , n318778 , n318779 , n318780 , n318781 , n318782 , n318783 , 
 n28358 , n28359 , n28360 , n28361 , n28362 , n318789 , n28364 , n28365 , n318792 , n318793 , 
 n318794 , n318795 , n28370 , n318797 , n318798 , n318799 , n318800 , n318801 , n318802 , n318803 , 
 n318804 , n318805 , n318806 , n318807 , n318808 , n318809 , n318810 , n318811 , n28386 , n318813 , 
 n318814 , n318815 , n318816 , n28391 , n318818 , n318819 , n318820 , n318821 , n318822 , n318823 , 
 n318824 , n318825 , n318826 , n28401 , n318828 , n28403 , n28404 , n318831 , n318832 , n318833 , 
 n318834 , n318835 , n318836 , n318837 , n318838 , n318839 , n28414 , n318841 , n318842 , n318843 , 
 n318844 , n318845 , n318846 , n318847 , n318848 , n318849 , n318850 , n318851 , n318852 , n318853 , 
 n28428 , n318855 , n318856 , n28431 , n318858 , n318859 , n28434 , n28435 , n318862 , n318863 , 
 n318864 , n318865 , n318866 , n318867 , n318868 , n318869 , n28444 , n318871 , n28446 , n28447 , 
 n318874 , n318875 , n318876 , n318877 , n318878 , n318879 , n318880 , n318881 , n318882 , n318883 , 
 n318884 , n318885 , n28460 , n28461 , n318888 , n28463 , n28464 , n28465 , n318892 , n28467 , 
 n318894 , n318895 , n28470 , n318897 , n28472 , n28473 , n318900 , n318901 , n28476 , n318903 , 
 n318904 , n28479 , n28480 , n28481 , n318908 , n28483 , n318910 , n318911 , n318912 , n28487 , 
 n28488 , n28489 , n318916 , n318917 , n318918 , n28493 , n28494 , n318921 , n318922 , n318923 , 
 n318924 , n28499 , n318926 , n318927 , n318928 , n28503 , n318930 , n318931 , n318932 , n28507 , 
 n318934 , n318935 , n318936 , n28511 , n318938 , n318939 , n28514 , n318941 , n318942 , n318943 , 
 n28518 , n318945 , n318946 , n318947 , n318948 , n318949 , n318950 , n318951 , n318952 , n318953 , 
 n318954 , n318955 , n318956 , n28531 , n318958 , n318959 , n318960 , n318961 , n28536 , n318963 , 
 n318964 , n318965 , n318966 , n318967 , n318968 , n318969 , n318970 , n318971 , n28546 , n318973 , 
 n318974 , n318975 , n318976 , n318977 , n318978 , n318979 , n318980 , n28555 , n318982 , n318983 , 
 n28558 , n28559 , n318986 , n318987 , n318988 , n318989 , n318990 , n318991 , n318992 , n318993 , 
 n28568 , n318995 , n318996 , n28571 , n318998 , n28573 , n319000 , n28575 , n319002 , n319003 , 
 n319004 , n319005 , n319006 , n319007 , n319008 , n319009 , n319010 , n319011 , n319012 , n319013 , 
 n319014 , n319015 , n319016 , n319017 , n319018 , n319019 , n319020 , n28595 , n319022 , n319023 , 
 n319024 , n319025 , n319026 , n319027 , n28602 , n319029 , n319030 , n319031 , n319032 , n28607 , 
 n319034 , n319035 , n319036 , n319037 , n319038 , n319039 , n319040 , n319041 , n319042 , n28617 , 
 n319044 , n319045 , n28620 , n319047 , n28622 , n319049 , n28624 , n28625 , n319052 , n28627 , 
 n319054 , n28629 , n319056 , n319057 , n319058 , n319059 , n319060 , n319061 , n319062 , n28637 , 
 n319064 , n28639 , n28640 , n319067 , n319068 , n28643 , n319070 , n319071 , n28646 , n319073 , 
 n319074 , n28649 , n319076 , n319077 , n319078 , n319079 , n319080 , n319081 , n319082 , n319083 , 
 n319084 , n319085 , n319086 , n28661 , n28662 , n319089 , n319090 , n319091 , n319092 , n319093 , 
 n319094 , n319095 , n319096 , n319097 , n319098 , n319099 , n319100 , n319101 , n319102 , n319103 , 
 n28678 , n319105 , n319106 , n319107 , n319108 , n319109 , n319110 , n319111 , n319112 , n319113 , 
 n319114 , n319115 , n319116 , n319117 , n319118 , n319119 , n319120 , n319121 , n319122 , n319123 , 
 n28698 , n319125 , n319126 , n319127 , n319128 , n28703 , n319130 , n319131 , n319132 , n319133 , 
 n319134 , n28709 , n28710 , n28711 , n319138 , n28713 , n28714 , n319141 , n28716 , n319143 , 
 n319144 , n28719 , n319146 , n319147 , n28722 , n319149 , n319150 , n319151 , n319152 , n319153 , 
 n319154 , n319155 , n319156 , n319157 , n319158 , n28733 , n28734 , n319161 , n28736 , n28737 , 
 n28738 , n319165 , n319166 , n319167 , n319168 , n319169 , n28744 , n319171 , n319172 , n319173 , 
 n28748 , n319175 , n319176 , n319177 , n319178 , n319179 , n28754 , n319181 , n319182 , n319183 , 
 n319184 , n28759 , n319186 , n319187 , n319188 , n28763 , n28764 , n319191 , n319192 , n28767 , 
 n28768 , n28769 , n319196 , n319197 , n319198 , n319199 , n319200 , n319201 , n319202 , n319203 , 
 n28778 , n319205 , n28780 , n319207 , n319208 , n319209 , n319210 , n319211 , n319212 , n319213 , 
 n319214 , n319215 , n319216 , n319217 , n28792 , n319219 , n319220 , n319221 , n319222 , n28797 , 
 n319224 , n319225 , n319226 , n319227 , n319228 , n319229 , n319230 , n28805 , n28806 , n319233 , 
 n319234 , n319235 , n319236 , n319237 , n319238 , n319239 , n28814 , n319241 , n28816 , n28817 , 
 n28818 , n28819 , n28820 , n319247 , n319248 , n319249 , n319250 , n319251 , n319252 , n319253 , 
 n319254 , n319255 , n319256 , n319257 , n319258 , n28833 , n319260 , n28835 , n319262 , n319263 , 
 n28838 , n319265 , n28840 , n28841 , n319268 , n319269 , n319270 , n319271 , n319272 , n319273 , 
 n319274 , n28849 , n28850 , n319277 , n319278 , n28853 , n319280 , n319281 , n319282 , n319283 , 
 n28858 , n28859 , n319286 , n319287 , n28862 , n319289 , n319290 , n319291 , n319292 , n319293 , 
 n28868 , n319295 , n319296 , n319297 , n319298 , n28873 , n319300 , n319301 , n28876 , n319303 , 
 n319304 , n319305 , n319306 , n319307 , n319308 , n319309 , n319310 , n319311 , n319312 , n319313 , 
 n28888 , n319315 , n319316 , n28891 , n319318 , n319319 , n319320 , n319321 , n319322 , n319323 , 
 n319324 , n319325 , n28900 , n319327 , n319328 , n319329 , n319330 , n319331 , n319332 , n28907 , 
 n28908 , n319335 , n319336 , n28911 , n28912 , n28913 , n319340 , n319341 , n28916 , n319343 , 
 n28918 , n319345 , n319346 , n28921 , n319348 , n319349 , n319350 , n319351 , n319352 , n319353 , 
 n319354 , n319355 , n319356 , n319357 , n319358 , n28933 , n319360 , n28935 , n28936 , n319363 , 
 n28938 , n28939 , n319366 , n319367 , n28942 , n319369 , n319370 , n319371 , n319372 , n319373 , 
 n28948 , n319375 , n28950 , n319377 , n319378 , n319379 , n28954 , n319381 , n319382 , n28957 , 
 n319384 , n319385 , n319386 , n319387 , n319388 , n319389 , n319390 , n319391 , n319392 , n319393 , 
 n319394 , n319395 , n319396 , n319397 , n319398 , n319399 , n319400 , n319401 , n28976 , n319403 , 
 n319404 , n319405 , n319406 , n319407 , n28982 , n28983 , n319410 , n319411 , n28986 , n28987 , 
 n319414 , n319415 , n319416 , n28991 , n319418 , n28993 , n28994 , n319421 , n319422 , n28997 , 
 n319424 , n319425 , n319426 , n29001 , n29002 , n319429 , n29004 , n319431 , n29006 , n319433 , 
 n319434 , n319435 , n29010 , n319437 , n319438 , n319439 , n319440 , n319441 , n319442 , n319443 , 
 n319444 , n319445 , n319446 , n319447 , n319448 , n319449 , n319450 , n319451 , n319452 , n29027 , 
 n29028 , n319455 , n319456 , n29031 , n319458 , n319459 , n319460 , n319461 , n319462 , n319463 , 
 n29038 , n29039 , n319466 , n29041 , n319468 , n319469 , n319470 , n319471 , n319472 , n319473 , 
 n319474 , n319475 , n29050 , n319477 , n319478 , n29053 , n319480 , n29055 , n319482 , n319483 , 
 n319484 , n319485 , n29060 , n319487 , n29062 , n29063 , n319490 , n319491 , n319492 , n319493 , 
 n319494 , n29069 , n29070 , n319497 , n319498 , n319499 , n29074 , n319501 , n29076 , n319503 , 
 n29078 , n29079 , n319506 , n319507 , n319508 , n29083 , n319510 , n319511 , n29086 , n319513 , 
 n319514 , n29089 , n319516 , n319517 , n319518 , n319519 , n29094 , n29095 , n319522 , n319523 , 
 n29098 , n319525 , n319526 , n29101 , n319528 , n319529 , n29104 , n319531 , n319532 , n29107 , 
 n319534 , n319535 , n29110 , n319537 , n319538 , n29113 , n319540 , n319541 , n319542 , n319543 , 
 n319544 , n319545 , n29120 , n319547 , n319548 , n29123 , n319550 , n29125 , n29126 , n319553 , 
 n319554 , n319555 , n319556 , n29131 , n319558 , n29133 , n319560 , n319561 , n319562 , n319563 , 
 n319564 , n319565 , n319566 , n319567 , n29142 , n319569 , n319570 , n319571 , n319572 , n319573 , 
 n319574 , n319575 , n319576 , n319577 , n319578 , n319579 , n319580 , n319581 , n319582 , n29157 , 
 n319584 , n319585 , n319586 , n29161 , n29162 , n319589 , n319590 , n319591 , n29166 , n319593 , 
 n319594 , n29169 , n319596 , n319597 , n319598 , n319599 , n319600 , n319601 , n29176 , n319603 , 
 n319604 , n319605 , n319606 , n319607 , n319608 , n319609 , n319610 , n319611 , n319612 , n319613 , 
 n319614 , n319615 , n319616 , n319617 , n319618 , n319619 , n319620 , n29195 , n319622 , n319623 , 
 n29198 , n319625 , n29200 , n319627 , n319628 , n319629 , n319630 , n319631 , n319632 , n319633 , 
 n29208 , n319635 , n319636 , n319637 , n319638 , n319639 , n319640 , n29215 , n319642 , n319643 , 
 n319644 , n319645 , n29220 , n29221 , n29222 , n29223 , n319650 , n319651 , n319652 , n319653 , 
 n319654 , n319655 , n319656 , n319657 , n319658 , n319659 , n319660 , n319661 , n319662 , n319663 , 
 n319664 , n319665 , n319666 , n319667 , n29242 , n29243 , n319670 , n29245 , n319672 , n319673 , 
 n319674 , n319675 , n319676 , n319677 , n319678 , n319679 , n319680 , n319681 , n319682 , n29257 , 
 n319684 , n319685 , n29260 , n319687 , n319688 , n319689 , n319690 , n319691 , n29266 , n319693 , 
 n319694 , n319695 , n319696 , n319697 , n29272 , n319699 , n319700 , n319701 , n29276 , n319703 , 
 n319704 , n319705 , n319706 , n319707 , n319708 , n319709 , n319710 , n29285 , n29286 , n29287 , 
 n319714 , n319715 , n319716 , n319717 , n319718 , n319719 , n29294 , n319721 , n319722 , n29297 , 
 n319724 , n319725 , n29300 , n319727 , n319728 , n319729 , n319730 , n319731 , n319732 , n319733 , 
 n29308 , n319735 , n319736 , n319737 , n319738 , n319739 , n319740 , n29315 , n29316 , n319743 , 
 n319744 , n319745 , n319746 , n319747 , n319748 , n319749 , n319750 , n319751 , n319752 , n319753 , 
 n319754 , n319755 , n319756 , n29331 , n319758 , n319759 , n319760 , n319761 , n319762 , n319763 , 
 n319764 , n319765 , n319766 , n319767 , n319768 , n319769 , n319770 , n319771 , n319772 , n319773 , 
 n319774 , n29349 , n319776 , n319777 , n319778 , n29353 , n29354 , n319781 , n29356 , n319783 , 
 n319784 , n319785 , n29360 , n29361 , n319788 , n319789 , n319790 , n29365 , n319792 , n319793 , 
 n29368 , n319795 , n319796 , n319797 , n319798 , n29373 , n319800 , n29375 , n319802 , n319803 , 
 n319804 , n319805 , n319806 , n319807 , n319808 , n319809 , n319810 , n319811 , n319812 , n319813 , 
 n319814 , n319815 , n319816 , n319817 , n29392 , n319819 , n319820 , n29395 , n319822 , n319823 , 
 n319824 , n319825 , n319826 , n319827 , n319828 , n319829 , n319830 , n319831 , n319832 , n319833 , 
 n319834 , n319835 , n319836 , n319837 , n319838 , n319839 , n319840 , n319841 , n319842 , n319843 , 
 n29418 , n29419 , n319846 , n319847 , n319848 , n319849 , n319850 , n29425 , n319852 , n319853 , 
 n319854 , n319855 , n319856 , n319857 , n319858 , n319859 , n319860 , n319861 , n29436 , n319863 , 
 n29438 , n29439 , n319866 , n319867 , n319868 , n319869 , n319870 , n29445 , n319872 , n319873 , 
 n29448 , n319875 , n319876 , n29451 , n319878 , n319879 , n29454 , n319881 , n319882 , n319883 , 
 n319884 , n319885 , n319886 , n319887 , n319888 , n29463 , n319890 , n319891 , n29466 , n319893 , 
 n29468 , n29469 , n319896 , n319897 , n319898 , n319899 , n319900 , n29475 , n319902 , n319903 , 
 n29478 , n319905 , n29480 , n319907 , n319908 , n29483 , n319910 , n29485 , n319912 , n319913 , 
 n29488 , n319915 , n319916 , n29491 , n319918 , n319919 , n319920 , n319921 , n29496 , n29497 , 
 n319924 , n319925 , n319926 , n319927 , n319928 , n319929 , n319930 , n319931 , n319932 , n319933 , 
 n319934 , n319935 , n319936 , n319937 , n319938 , n29513 , n29514 , n319941 , n319942 , n29517 , 
 n319944 , n319945 , n319946 , n319947 , n319948 , n29523 , n319950 , n319951 , n319952 , n29527 , 
 n29528 , n319955 , n319956 , n319957 , n319958 , n319959 , n319960 , n319961 , n319962 , n319963 , 
 n319964 , n319965 , n319966 , n319967 , n29542 , n319969 , n319970 , n29545 , n319972 , n319973 , 
 n319974 , n29549 , n319976 , n319977 , n319978 , n29553 , n319980 , n319981 , n29556 , n319983 , 
 n319984 , n29559 , n29560 , n319987 , n319988 , n319989 , n29564 , n29565 , n319992 , n319993 , 
 n319994 , n319995 , n319996 , n319997 , n319998 , n319999 , n320000 , n320001 , n29576 , n320003 , 
 n29578 , n320005 , n320006 , n320007 , n320008 , n29583 , n29584 , n320011 , n320012 , n320013 , 
 n320014 , n320015 , n320016 , n320017 , n320018 , n320019 , n320020 , n320021 , n320022 , n29597 , 
 n320024 , n320025 , n320026 , n320027 , n320028 , n320029 , n320030 , n320031 , n320032 , n29607 , 
 n320034 , n320035 , n320036 , n320037 , n320038 , n29613 , n29614 , n320041 , n320042 , n320043 , 
 n29618 , n320045 , n320046 , n320047 , n29622 , n29623 , n320050 , n320051 , n320052 , n320053 , 
 n29628 , n320055 , n29630 , n320057 , n320058 , n320059 , n29634 , n29635 , n29636 , n320063 , 
 n29638 , n29639 , n29640 , n320067 , n320068 , n320069 , n29644 , n320071 , n320072 , n320073 , 
 n320074 , n320075 , n320076 , n320077 , n320078 , n320079 , n320080 , n320081 , n320082 , n320083 , 
 n320084 , n320085 , n320086 , n29661 , n320088 , n320089 , n320090 , n320091 , n320092 , n320093 , 
 n320094 , n320095 , n320096 , n320097 , n29672 , n29673 , n320100 , n29675 , n320102 , n29677 , 
 n320104 , n320105 , n29680 , n320107 , n320108 , n320109 , n320110 , n320111 , n320112 , n29687 , 
 n320114 , n320115 , n29690 , n320117 , n320118 , n320119 , n320120 , n320121 , n29696 , n320123 , 
 n320124 , n320125 , n29700 , n320127 , n320128 , n320129 , n320130 , n29705 , n320132 , n320133 , 
 n29708 , n320135 , n320136 , n320137 , n320138 , n29713 , n320140 , n29715 , n320142 , n29717 , 
 n320144 , n320145 , n320146 , n320147 , n320148 , n320149 , n29724 , n320151 , n320152 , n320153 , 
 n320154 , n320155 , n29730 , n320157 , n29732 , n320159 , n320160 , n320161 , n320162 , n320163 , 
 n320164 , n320165 , n29740 , n29741 , n320168 , n320169 , n320170 , n320171 , n320172 , n29747 , 
 n320174 , n320175 , n29750 , n320177 , n320178 , n320179 , n320180 , n320181 , n29756 , n320183 , 
 n320184 , n320185 , n320186 , n320187 , n320188 , n320189 , n320190 , n320191 , n320192 , n320193 , 
 n320194 , n320195 , n29770 , n320197 , n320198 , n320199 , n320200 , n320201 , n320202 , n320203 , 
 n320204 , n320205 , n320206 , n320207 , n320208 , n320209 , n29784 , n320211 , n320212 , n320213 , 
 n29788 , n320215 , n320216 , n29791 , n320218 , n320219 , n29794 , n29795 , n320222 , n320223 , 
 n29798 , n29799 , n320226 , n29801 , n320228 , n320229 , n320230 , n29805 , n320232 , n320233 , 
 n320234 , n320235 , n320236 , n320237 , n29812 , n320239 , n320240 , n320241 , n320242 , n29817 , 
 n320244 , n320245 , n320246 , n320247 , n320248 , n320249 , n320250 , n320251 , n29826 , n320253 , 
 n29828 , n320255 , n29830 , n29831 , n320258 , n29833 , n320260 , n320261 , n29836 , n320263 , 
 n320264 , n320265 , n320266 , n320267 , n320268 , n320269 , n29844 , n320271 , n320272 , n320273 , 
 n320274 , n320275 , n320276 , n320277 , n320278 , n29853 , n29854 , n320281 , n320282 , n320283 , 
 n320284 , n29859 , n320286 , n320287 , n29862 , n29863 , n320290 , n29865 , n29866 , n320293 , 
 n320294 , n29869 , n29870 , n29871 , n320298 , n320299 , n29874 , n29875 , n320302 , n320303 , 
 n320304 , n29879 , n320306 , n320307 , n320308 , n320309 , n320310 , n320311 , n320312 , n29887 , 
 n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n320320 , n320321 , n320322 , n320323 , 
 n320324 , n320325 , n320326 , n29901 , n320328 , n29903 , n320330 , n320331 , n320332 , n320333 , 
 n320334 , n320335 , n320336 , n320337 , n320338 , n320339 , n29914 , n29915 , n29916 , n320343 , 
 n320344 , n320345 , n320346 , n320347 , n320348 , n320349 , n320350 , n29925 , n320352 , n320353 , 
 n320354 , n320355 , n320356 , n320357 , n320358 , n320359 , n320360 , n320361 , n320362 , n320363 , 
 n320364 , n320365 , n320366 , n29941 , n320368 , n29943 , n320370 , n29945 , n320372 , n320373 , 
 n320374 , n320375 , n320376 , n320377 , n320378 , n320379 , n320380 , n320381 , n320382 , n29957 , 
 n320384 , n320385 , n320386 , n320387 , n29962 , n320389 , n320390 , n29965 , n320392 , n320393 , 
 n320394 , n320395 , n320396 , n320397 , n320398 , n320399 , n320400 , n29975 , n320402 , n320403 , 
 n29978 , n320405 , n320406 , n320407 , n320408 , n320409 , n320410 , n29985 , n320412 , n320413 , 
 n320414 , n320415 , n320416 , n320417 , n320418 , n320419 , n320420 , n320421 , n29996 , n320423 , 
 n320424 , n320425 , n320426 , n320427 , n320428 , n320429 , n320430 , n320431 , n320432 , n320433 , 
 n320434 , n320435 , n30010 , n320437 , n320438 , n30013 , n30014 , n320441 , n320442 , n320443 , 
 n320444 , n30019 , n320446 , n320447 , n320448 , n30023 , n320450 , n320451 , n320452 , n320453 , 
 n320454 , n320455 , n30030 , n320457 , n320458 , n320459 , n320460 , n320461 , n320462 , n320463 , 
 n320464 , n320465 , n320466 , n30041 , n30042 , n320469 , n30044 , n320471 , n320472 , n320473 , 
 n320474 , n320475 , n30050 , n320477 , n320478 , n320479 , n320480 , n320481 , n30056 , n320483 , 
 n320484 , n320485 , n320486 , n30061 , n320488 , n320489 , n30064 , n320491 , n320492 , n320493 , 
 n320494 , n320495 , n320496 , n320497 , n320498 , n320499 , n30074 , n320501 , n320502 , n320503 , 
 n30078 , n320505 , n320506 , n30081 , n320508 , n320509 , n320510 , n30085 , n320512 , n320513 , 
 n30088 , n320515 , n320516 , n30091 , n320518 , n320519 , n30094 , n320521 , n30096 , n320523 , 
 n320524 , n320525 , n320526 , n320527 , n320528 , n320529 , n320530 , n320531 , n30106 , n320533 , 
 n320534 , n320535 , n320536 , n320537 , n320538 , n30113 , n320540 , n320541 , n30116 , n320543 , 
 n320544 , n320545 , n320546 , n320547 , n320548 , n320549 , n320550 , n320551 , n30126 , n320553 , 
 n320554 , n320555 , n320556 , n320557 , n320558 , n320559 , n320560 , n30135 , n320562 , n320563 , 
 n30138 , n30139 , n320566 , n320567 , n320568 , n320569 , n320570 , n320571 , n30146 , n320573 , 
 n320574 , n320575 , n30150 , n320577 , n320578 , n320579 , n320580 , n320581 , n320582 , n30157 , 
 n320584 , n320585 , n30160 , n30161 , n320588 , n320589 , n320590 , n320591 , n320592 , n320593 , 
 n30168 , n320595 , n320596 , n320597 , n320598 , n30173 , n30174 , n320601 , n320602 , n320603 , 
 n320604 , n320605 , n320606 , n320607 , n320608 , n320609 , n30184 , n320611 , n320612 , n320613 , 
 n320614 , n320615 , n320616 , n320617 , n320618 , n320619 , n320620 , n320621 , n320622 , n320623 , 
 n320624 , n320625 , n320626 , n320627 , n320628 , n320629 , n320630 , n320631 , n30206 , n320633 , 
 n320634 , n30209 , n30210 , n320637 , n320638 , n30213 , n320640 , n320641 , n320642 , n320643 , 
 n320644 , n320645 , n320646 , n320647 , n320648 , n320649 , n320650 , n320651 , n320652 , n320653 , 
 n320654 , n30229 , n320656 , n320657 , n320658 , n320659 , n320660 , n30235 , n30236 , n30237 , 
 n320664 , n320665 , n30240 , n320667 , n320668 , n30243 , n320670 , n320671 , n320672 , n320673 , 
 n30248 , n320675 , n320676 , n320677 , n320678 , n320679 , n320680 , n320681 , n30256 , n30257 , 
 n30258 , n30259 , n30260 , n320687 , n320688 , n320689 , n320690 , n30265 , n30266 , n320693 , 
 n320694 , n320695 , n30270 , n320697 , n30272 , n320699 , n320700 , n320701 , n320702 , n30277 , 
 n320704 , n320705 , n320706 , n320707 , n320708 , n30283 , n320710 , n320711 , n320712 , n30287 , 
 n320714 , n30289 , n320716 , n320717 , n320718 , n320719 , n320720 , n320721 , n320722 , n320723 , 
 n320724 , n320725 , n320726 , n30301 , n320728 , n320729 , n320730 , n320731 , n320732 , n30307 , 
 n320734 , n30309 , n320736 , n320737 , n30312 , n320739 , n320740 , n30315 , n320742 , n320743 , 
 n320744 , n320745 , n320746 , n320747 , n320748 , n320749 , n320750 , n320751 , n30326 , n320753 , 
 n320754 , n320755 , n320756 , n30331 , n30332 , n320759 , n320760 , n320761 , n320762 , n320763 , 
 n320764 , n30339 , n30340 , n320767 , n30342 , n30343 , n30344 , n320771 , n30346 , n320773 , 
 n320774 , n30349 , n320776 , n320777 , n30352 , n320779 , n320780 , n30355 , n320782 , n320783 , 
 n30358 , n320785 , n320786 , n320787 , n320788 , n320789 , n30364 , n320791 , n320792 , n30367 , 
 n320794 , n320795 , n320796 , n30371 , n30372 , n320799 , n30374 , n320801 , n320802 , n320803 , 
 n30378 , n320805 , n320806 , n30381 , n320808 , n320809 , n320810 , n320811 , n320812 , n320813 , 
 n320814 , n320815 , n320816 , n320817 , n320818 , n30393 , n320820 , n320821 , n320822 , n320823 , 
 n320824 , n30399 , n320826 , n320827 , n320828 , n320829 , n320830 , n30405 , n320832 , n320833 , 
 n320834 , n320835 , n320836 , n320837 , n30412 , n320839 , n320840 , n320841 , n30416 , n30417 , 
 n320844 , n30419 , n320846 , n320847 , n320848 , n320849 , n30424 , n320851 , n320852 , n320853 , 
 n320854 , n320855 , n320856 , n320857 , n320858 , n320859 , n320860 , n320861 , n30436 , n30437 , 
 n320864 , n30439 , n320866 , n320867 , n30442 , n320869 , n320870 , n320871 , n320872 , n30447 , 
 n320874 , n320875 , n320876 , n320877 , n320878 , n320879 , n320880 , n320881 , n320882 , n30457 , 
 n320884 , n320885 , n320886 , n30461 , n320888 , n30463 , n30464 , n320891 , n320892 , n320893 , 
 n320894 , n320895 , n320896 , n320897 , n320898 , n320899 , n320900 , n320901 , n320902 , n320903 , 
 n320904 , n320905 , n30480 , n320907 , n320908 , n320909 , n320910 , n320911 , n320912 , n30487 , 
 n320914 , n320915 , n320916 , n320917 , n320918 , n320919 , n320920 , n30495 , n320922 , n320923 , 
 n30498 , n320925 , n320926 , n320927 , n320928 , n320929 , n320930 , n320931 , n320932 , n30507 , 
 n320934 , n320935 , n30510 , n320937 , n30512 , n320939 , n320940 , n30515 , n320942 , n320943 , 
 n320944 , n320945 , n320946 , n30521 , n30522 , n320949 , n320950 , n30525 , n30526 , n320953 , 
 n30528 , n320955 , n30530 , n30531 , n320958 , n30533 , n320960 , n320961 , n320962 , n30537 , 
 n320964 , n320965 , n320966 , n320967 , n30542 , n320969 , n320970 , n320971 , n30546 , n320973 , 
 n320974 , n30549 , n320976 , n30551 , n30552 , n320979 , n30554 , n320981 , n30556 , n30557 , 
 n320984 , n30559 , n320986 , n320987 , n320988 , n320989 , n30564 , n320991 , n320992 , n320993 , 
 n320994 , n320995 , n30570 , n320997 , n320998 , n30573 , n30574 , n321001 , n30576 , n30577 , 
 n321004 , n321005 , n321006 , n30581 , n321008 , n321009 , n321010 , n30585 , n321012 , n321013 , 
 n30588 , n30589 , n321016 , n321017 , n30592 , n321019 , n30594 , n30595 , n321022 , n321023 , 
 n30598 , n321025 , n321026 , n321027 , n30602 , n321029 , n30604 , n321031 , n321032 , n30607 , 
 n321034 , n321035 , n30610 , n30611 , n321038 , n30613 , n321040 , n30615 , n321042 , n30617 , 
 n30618 , n321045 , n321046 , n321047 , n321048 , n321049 , n321050 , n321051 , n321052 , n321053 , 
 n321054 , n321055 , n321056 , n321057 , n30632 , n30633 , n321060 , n321061 , n30636 , n321063 , 
 n321064 , n321065 , n321066 , n321067 , n321068 , n321069 , n30644 , n321071 , n321072 , n321073 , 
 n321074 , n321075 , n321076 , n321077 , n30652 , n321079 , n321080 , n321081 , n30656 , n321083 , 
 n321084 , n321085 , n321086 , n321087 , n30662 , n321089 , n321090 , n321091 , n321092 , n30667 , 
 n30668 , n321095 , n321096 , n30671 , n30672 , n30673 , n30674 , n321101 , n321102 , n321103 , 
 n321104 , n321105 , n321106 , n321107 , n321108 , n30683 , n321110 , n321111 , n321112 , n321113 , 
 n30688 , n321115 , n321116 , n30691 , n321118 , n30693 , n321120 , n321121 , n321122 , n321123 , 
 n321124 , n321125 , n321126 , n321127 , n321128 , n321129 , n30704 , n321131 , n30706 , n321133 , 
 n321134 , n321135 , n30710 , n321137 , n321138 , n321139 , n321140 , n321141 , n321142 , n321143 , 
 n30718 , n321145 , n321146 , n321147 , n30722 , n321149 , n321150 , n30725 , n321152 , n321153 , 
 n321154 , n30729 , n321156 , n321157 , n321158 , n30733 , n321160 , n321161 , n321162 , n30737 , 
 n321164 , n321165 , n30740 , n321167 , n321168 , n321169 , n30744 , n321171 , n321172 , n321173 , 
 n321174 , n321175 , n321176 , n321177 , n30752 , n321179 , n321180 , n321181 , n321182 , n321183 , 
 n321184 , n321185 , n321186 , n321187 , n321188 , n321189 , n321190 , n321191 , n321192 , n321193 , 
 n321194 , n30769 , n321196 , n321197 , n321198 , n30773 , n30774 , n321201 , n30776 , n321203 , 
 n321204 , n30779 , n321206 , n321207 , n321208 , n321209 , n321210 , n321211 , n321212 , n321213 , 
 n321214 , n321215 , n321216 , n321217 , n321218 , n321219 , n321220 , n321221 , n321222 , n321223 , 
 n321224 , n321225 , n321226 , n321227 , n321228 , n321229 , n321230 , n321231 , n321232 , n321233 , 
 n321234 , n321235 , n321236 , n321237 , n321238 , n321239 , n321240 , n321241 , n321242 , n321243 , 
 n321244 , n30819 , n321246 , n321247 , n30822 , n30823 , n321250 , n321251 , n321252 , n321253 , 
 n321254 , n321255 , n321256 , n321257 , n321258 , n321259 , n321260 , n321261 , n321262 , n321263 , 
 n30838 , n321265 , n30840 , n321267 , n321268 , n321269 , n321270 , n321271 , n321272 , n321273 , 
 n30848 , n321275 , n321276 , n321277 , n321278 , n321279 , n30854 , n321281 , n321282 , n321283 , 
 n321284 , n321285 , n321286 , n30861 , n321288 , n321289 , n30864 , n321291 , n30866 , n321293 , 
 n321294 , n321295 , n321296 , n30871 , n30872 , n321299 , n30874 , n321301 , n321302 , n321303 , 
 n30878 , n321305 , n321306 , n30881 , n30882 , n321309 , n321310 , n321311 , n321312 , n321313 , 
 n321314 , n321315 , n321316 , n30891 , n30892 , n321319 , n321320 , n321321 , n321322 , n321323 , 
 n30898 , n321325 , n321326 , n321327 , n321328 , n321329 , n321330 , n321331 , n321332 , n321333 , 
 n321334 , n30909 , n321336 , n321337 , n321338 , n321339 , n321340 , n321341 , n321342 , n321343 , 
 n321344 , n30919 , n321346 , n321347 , n321348 , n321349 , n30924 , n30925 , n321352 , n30927 , 
 n30928 , n321355 , n321356 , n321357 , n321358 , n321359 , n321360 , n321361 , n30936 , n321363 , 
 n321364 , n30939 , n321366 , n30941 , n30942 , n321369 , n30944 , n30945 , n321372 , n30947 , 
 n321374 , n321375 , n321376 , n321377 , n321378 , n321379 , n30954 , n30955 , n30956 , n321383 , 
 n30958 , n321385 , n321386 , n30961 , n30962 , n321389 , n321390 , n30965 , n321392 , n30967 , 
 n321394 , n321395 , n321396 , n321397 , n30972 , n30973 , n321400 , n321401 , n321402 , n321403 , 
 n321404 , n321405 , n321406 , n30981 , n30982 , n30983 , n321410 , n321411 , n321412 , n321413 , 
 n321414 , n321415 , n321416 , n30991 , n321418 , n321419 , n30994 , n321421 , n321422 , n30997 , 
 n321424 , n321425 , n321426 , n321427 , n321428 , n321429 , n321430 , n321431 , n321432 , n31007 , 
 n31008 , n321435 , n321436 , n31011 , n321438 , n321439 , n321440 , n321441 , n321442 , n321443 , 
 n321444 , n31019 , n31020 , n31021 , n321448 , n321449 , n321450 , n321451 , n31026 , n321453 , 
 n321454 , n321455 , n31030 , n321457 , n31032 , n321459 , n321460 , n31035 , n31036 , n321463 , 
 n31038 , n321465 , n321466 , n321467 , n321468 , n321469 , n321470 , n31045 , n31046 , n321473 , 
 n321474 , n321475 , n321476 , n321477 , n321478 , n31053 , n321480 , n321481 , n31056 , n321483 , 
 n321484 , n321485 , n321486 , n321487 , n321488 , n321489 , n31064 , n321491 , n321492 , n321493 , 
 n321494 , n321495 , n321496 , n31071 , n321498 , n321499 , n321500 , n31075 , n321502 , n321503 , 
 n321504 , n321505 , n31080 , n321507 , n31082 , n321509 , n321510 , n321511 , n321512 , n321513 , 
 n321514 , n321515 , n321516 , n31091 , n31092 , n321519 , n321520 , n321521 , n321522 , n31097 , 
 n321524 , n321525 , n321526 , n31101 , n321528 , n321529 , n31104 , n31105 , n321532 , n321533 , 
 n321534 , n321535 , n31110 , n31111 , n321538 , n321539 , n31114 , n321541 , n321542 , n321543 , 
 n31118 , n321545 , n321546 , n321547 , n31122 , n31123 , n321550 , n321551 , n31126 , n321553 , 
 n321554 , n31129 , n321556 , n321557 , n31132 , n321559 , n321560 , n321561 , n321562 , n321563 , 
 n321564 , n321565 , n321566 , n31141 , n321568 , n321569 , n31144 , n321571 , n31146 , n321573 , 
 n31148 , n321575 , n321576 , n31151 , n321578 , n321579 , n31154 , n321581 , n321582 , n321583 , 
 n321584 , n321585 , n321586 , n321587 , n321588 , n321589 , n321590 , n31165 , n321592 , n31167 , 
 n321594 , n321595 , n31170 , n321597 , n321598 , n31173 , n31174 , n321601 , n31176 , n321603 , 
 n321604 , n31179 , n321606 , n321607 , n31182 , n31183 , n321610 , n31185 , n321612 , n321613 , 
 n31188 , n321615 , n31190 , n321617 , n321618 , n321619 , n321620 , n321621 , n321622 , n31197 , 
 n31198 , n31199 , n31200 , n31201 , n31202 , n321629 , n321630 , n321631 , n31206 , n321633 , 
 n321634 , n321635 , n321636 , n31211 , n321638 , n321639 , n321640 , n321641 , n321642 , n321643 , 
 n321644 , n321645 , n321646 , n31221 , n31222 , n321649 , n31224 , n321651 , n321652 , n321653 , 
 n321654 , n321655 , n321656 , n31231 , n321658 , n321659 , n321660 , n31235 , n321662 , n321663 , 
 n321664 , n31239 , n31240 , n31241 , n321668 , n321669 , n321670 , n321671 , n321672 , n321673 , 
 n321674 , n321675 , n321676 , n321677 , n321678 , n321679 , n321680 , n321681 , n321682 , n321683 , 
 n321684 , n321685 , n321686 , n321687 , n31262 , n31263 , n321690 , n321691 , n31266 , n321693 , 
 n321694 , n321695 , n321696 , n321697 , n31272 , n321699 , n321700 , n321701 , n321702 , n321703 , 
 n31278 , n321705 , n321706 , n31281 , n321708 , n321709 , n321710 , n31285 , n321712 , n321713 , 
 n321714 , n321715 , n321716 , n321717 , n31292 , n31293 , n321720 , n321721 , n321722 , n31297 , 
 n31298 , n31299 , n321726 , n321727 , n321728 , n321729 , n31304 , n321731 , n321732 , n31307 , 
 n321734 , n321735 , n31310 , n321737 , n321738 , n321739 , n321740 , n321741 , n321742 , n321743 , 
 n321744 , n321745 , n321746 , n321747 , n321748 , n321749 , n31324 , n31325 , n31326 , n31327 , 
 n31328 , n31329 , n321756 , n321757 , n321758 , n321759 , n321760 , n321761 , n321762 , n321763 , 
 n321764 , n31339 , n321766 , n321767 , n31342 , n321769 , n321770 , n321771 , n321772 , n321773 , 
 n321774 , n321775 , n321776 , n321777 , n321778 , n31353 , n31354 , n321781 , n321782 , n321783 , 
 n321784 , n321785 , n321786 , n321787 , n31362 , n321789 , n321790 , n31365 , n321792 , n321793 , 
 n321794 , n321795 , n321796 , n321797 , n31372 , n321799 , n321800 , n31375 , n321802 , n321803 , 
 n321804 , n321805 , n31380 , n321807 , n321808 , n31383 , n321810 , n321811 , n31386 , n321813 , 
 n321814 , n31389 , n31390 , n321817 , n321818 , n321819 , n321820 , n321821 , n321822 , n321823 , 
 n321824 , n321825 , n31400 , n321827 , n321828 , n31403 , n321830 , n321831 , n321832 , n31407 , 
 n321834 , n321835 , n321836 , n321837 , n321838 , n321839 , n321840 , n321841 , n321842 , n321843 , 
 n321844 , n31419 , n321846 , n321847 , n31422 , n321849 , n321850 , n321851 , n31426 , n321853 , 
 n321854 , n321855 , n321856 , n321857 , n321858 , n321859 , n31434 , n321861 , n321862 , n321863 , 
 n321864 , n31439 , n321866 , n321867 , n321868 , n321869 , n321870 , n31445 , n321872 , n321873 , 
 n321874 , n31449 , n321876 , n321877 , n31452 , n321879 , n321880 , n321881 , n321882 , n321883 , 
 n321884 , n321885 , n321886 , n321887 , n321888 , n31463 , n321890 , n321891 , n31466 , n321893 , 
 n321894 , n321895 , n31470 , n321897 , n321898 , n31473 , n321900 , n321901 , n31476 , n31477 , 
 n321904 , n321905 , n321906 , n321907 , n321908 , n321909 , n31484 , n321911 , n321912 , n321913 , 
 n321914 , n321915 , n321916 , n321917 , n321918 , n321919 , n321920 , n321921 , n321922 , n321923 , 
 n321924 , n321925 , n31500 , n321927 , n321928 , n31503 , n321930 , n321931 , n321932 , n321933 , 
 n321934 , n321935 , n321936 , n31511 , n31512 , n321939 , n31514 , n321941 , n321942 , n321943 , 
 n321944 , n31519 , n321946 , n321947 , n321948 , n321949 , n321950 , n31525 , n321952 , n321953 , 
 n321954 , n321955 , n321956 , n321957 , n321958 , n321959 , n321960 , n31535 , n31536 , n321963 , 
 n321964 , n321965 , n321966 , n31541 , n31542 , n321969 , n321970 , n321971 , n321972 , n31547 , 
 n321974 , n321975 , n31550 , n321977 , n321978 , n321979 , n321980 , n321981 , n321982 , n321983 , 
 n321984 , n321985 , n321986 , n321987 , n321988 , n321989 , n321990 , n31565 , n31566 , n321993 , 
 n321994 , n31569 , n321996 , n321997 , n321998 , n321999 , n322000 , n322001 , n322002 , n31577 , 
 n322004 , n322005 , n31580 , n322007 , n322008 , n322009 , n322010 , n31585 , n31586 , n322013 , 
 n31588 , n322015 , n31590 , n322017 , n322018 , n31593 , n322020 , n322021 , n31596 , n322023 , 
 n322024 , n31599 , n322026 , n322027 , n31602 , n31603 , n322030 , n322031 , n31606 , n322033 , 
 n322034 , n322035 , n322036 , n322037 , n322038 , n322039 , n322040 , n322041 , n322042 , n322043 , 
 n322044 , n322045 , n31620 , n322047 , n322048 , n31623 , n322050 , n322051 , n322052 , n322053 , 
 n31628 , n322055 , n322056 , n31631 , n322058 , n322059 , n322060 , n31635 , n322062 , n322063 , 
 n322064 , n322065 , n322066 , n322067 , n322068 , n322069 , n322070 , n31645 , n322072 , n322073 , 
 n322074 , n322075 , n322076 , n31651 , n322078 , n322079 , n322080 , n322081 , n322082 , n322083 , 
 n322084 , n322085 , n322086 , n322087 , n322088 , n322089 , n322090 , n322091 , n322092 , n322093 , 
 n322094 , n322095 , n322096 , n322097 , n31672 , n322099 , n322100 , n322101 , n322102 , n31677 , 
 n322104 , n322105 , n31680 , n322107 , n322108 , n322109 , n322110 , n322111 , n322112 , n322113 , 
 n322114 , n31689 , n322116 , n322117 , n31692 , n322119 , n322120 , n322121 , n322122 , n31697 , 
 n322124 , n322125 , n322126 , n322127 , n322128 , n322129 , n322130 , n322131 , n322132 , n31707 , 
 n322134 , n322135 , n322136 , n322137 , n322138 , n322139 , n31714 , n31715 , n322142 , n322143 , 
 n322144 , n322145 , n322146 , n322147 , n322148 , n31723 , n322150 , n322151 , n31726 , n322153 , 
 n322154 , n322155 , n31730 , n322157 , n322158 , n31733 , n322160 , n322161 , n322162 , n31737 , 
 n322164 , n322165 , n31740 , n322167 , n322168 , n322169 , n322170 , n322171 , n31746 , n31747 , 
 n322174 , n322175 , n31750 , n322177 , n322178 , n322179 , n322180 , n322181 , n31756 , n322183 , 
 n322184 , n322185 , n322186 , n322187 , n322188 , n322189 , n31764 , n31765 , n322192 , n322193 , 
 n31768 , n31769 , n322196 , n31771 , n31772 , n322199 , n31774 , n322201 , n322202 , n31777 , 
 n322204 , n322205 , n31780 , n322207 , n322208 , n31783 , n322210 , n322211 , n31786 , n31787 , 
 n322214 , n322215 , n322216 , n322217 , n322218 , n322219 , n31794 , n322221 , n322222 , n322223 , 
 n31798 , n322225 , n322226 , n322227 , n322228 , n322229 , n322230 , n322231 , n322232 , n31807 , 
 n322234 , n322235 , n31810 , n322237 , n322238 , n322239 , n31814 , n31815 , n322242 , n322243 , 
 n31818 , n322245 , n322246 , n31821 , n322248 , n322249 , n31824 , n322251 , n322252 , n322253 , 
 n322254 , n322255 , n322256 , n31831 , n322258 , n322259 , n322260 , n322261 , n322262 , n31837 , 
 n322264 , n322265 , n31840 , n31841 , n31842 , n322269 , n31844 , n31845 , n322272 , n322273 , 
 n322274 , n31849 , n322276 , n322277 , n31852 , n31853 , n31854 , n31855 , n322282 , n322283 , 
 n31858 , n322285 , n322286 , n31861 , n322288 , n31863 , n31864 , n322291 , n31866 , n31867 , 
 n31868 , n31869 , n322296 , n31871 , n322298 , n31873 , n322300 , n322301 , n322302 , n322303 , 
 n31878 , n322305 , n322306 , n31881 , n322308 , n322309 , n322310 , n322311 , n322312 , n322313 , 
 n322314 , n322315 , n31890 , n322317 , n322318 , n322319 , n322320 , n31895 , n322322 , n31897 , 
 n31898 , n31899 , n322326 , n31901 , n31902 , n31903 , n31904 , n322331 , n322332 , n31907 , 
 n322334 , n322335 , n31910 , n31911 , n322338 , n322339 , n31914 , n322341 , n322342 , n322343 , 
 n322344 , n322345 , n31920 , n322347 , n322348 , n31923 , n322350 , n322351 , n31926 , n322353 , 
 n322354 , n31929 , n31930 , n322357 , n322358 , n322359 , n322360 , n322361 , n322362 , n322363 , 
 n322364 , n322365 , n31940 , n31941 , n322368 , n322369 , n322370 , n322371 , n322372 , n322373 , 
 n322374 , n322375 , n322376 , n322377 , n322378 , n322379 , n31954 , n322381 , n322382 , n31957 , 
 n322384 , n322385 , n31960 , n322387 , n322388 , n322389 , n31964 , n31965 , n322392 , n31967 , 
 n322394 , n322395 , n31970 , n322397 , n31972 , n322399 , n322400 , n322401 , n322402 , n31977 , 
 n322404 , n322405 , n322406 , n31981 , n322408 , n31983 , n322410 , n322411 , n322412 , n322413 , 
 n322414 , n322415 , n322416 , n322417 , n31992 , n322419 , n31994 , n31995 , n322422 , n322423 , 
 n322424 , n322425 , n322426 , n322427 , n322428 , n322429 , n32004 , n322431 , n322432 , n32007 , 
 n322434 , n322435 , n32010 , n322437 , n32012 , n322439 , n322440 , n32015 , n322442 , n322443 , 
 n322444 , n322445 , n32020 , n322447 , n322448 , n32023 , n322450 , n322451 , n32026 , n322453 , 
 n322454 , n32029 , n322456 , n322457 , n32032 , n322459 , n322460 , n322461 , n322462 , n322463 , 
 n322464 , n322465 , n322466 , n322467 , n322468 , n322469 , n322470 , n322471 , n322472 , n32047 , 
 n322474 , n322475 , n322476 , n322477 , n322478 , n322479 , n322480 , n322481 , n32056 , n322483 , 
 n322484 , n32059 , n322486 , n322487 , n32062 , n322489 , n322490 , n32065 , n322492 , n322493 , 
 n322494 , n322495 , n322496 , n322497 , n322498 , n322499 , n32074 , n322501 , n322502 , n322503 , 
 n322504 , n32079 , n322506 , n322507 , n32082 , n322509 , n322510 , n322511 , n322512 , n32087 , 
 n32088 , n322515 , n32090 , n322517 , n322518 , n322519 , n322520 , n322521 , n322522 , n322523 , 
 n322524 , n322525 , n322526 , n322527 , n322528 , n322529 , n322530 , n322531 , n322532 , n322533 , 
 n32108 , n322535 , n322536 , n322537 , n32112 , n322539 , n32114 , n322541 , n322542 , n322543 , 
 n322544 , n32119 , n322546 , n322547 , n32122 , n32123 , n322550 , n322551 , n322552 , n32127 , 
 n322554 , n322555 , n322556 , n322557 , n322558 , n322559 , n32134 , n322561 , n322562 , n322563 , 
 n322564 , n32139 , n322566 , n32141 , n32142 , n322569 , n322570 , n322571 , n322572 , n322573 , 
 n32148 , n322575 , n322576 , n322577 , n32152 , n322579 , n322580 , n32155 , n322582 , n32157 , 
 n322584 , n322585 , n322586 , n32161 , n322588 , n322589 , n322590 , n322591 , n32166 , n322593 , 
 n32168 , n32169 , n322596 , n322597 , n322598 , n322599 , n322600 , n322601 , n322602 , n322603 , 
 n322604 , n322605 , n322606 , n322607 , n322608 , n32183 , n322610 , n322611 , n32186 , n322613 , 
 n322614 , n322615 , n32190 , n322617 , n322618 , n322619 , n322620 , n322621 , n322622 , n322623 , 
 n32198 , n322625 , n322626 , n32201 , n32202 , n322629 , n322630 , n32205 , n32206 , n322633 , 
 n322634 , n322635 , n322636 , n322637 , n322638 , n322639 , n322640 , n322641 , n32216 , n32217 , 
 n322644 , n322645 , n32220 , n322647 , n322648 , n322649 , n322650 , n322651 , n322652 , n322653 , 
 n322654 , n322655 , n322656 , n322657 , n322658 , n322659 , n32234 , n322661 , n322662 , n322663 , 
 n32238 , n322665 , n322666 , n32241 , n322668 , n322669 , n322670 , n322671 , n322672 , n322673 , 
 n322674 , n322675 , n322676 , n322677 , n322678 , n32253 , n322680 , n322681 , n322682 , n322683 , 
 n322684 , n322685 , n322686 , n322687 , n32262 , n322689 , n322690 , n322691 , n322692 , n322693 , 
 n322694 , n32269 , n322696 , n322697 , n32272 , n322699 , n322700 , n32275 , n322702 , n322703 , 
 n322704 , n322705 , n322706 , n322707 , n322708 , n322709 , n322710 , n322711 , n322712 , n322713 , 
 n322714 , n322715 , n322716 , n322717 , n32292 , n322719 , n322720 , n322721 , n32296 , n322723 , 
 n32298 , n322725 , n322726 , n322727 , n322728 , n322729 , n322730 , n322731 , n322732 , n322733 , 
 n322734 , n322735 , n32310 , n322737 , n322738 , n32313 , n322740 , n322741 , n322742 , n322743 , 
 n32318 , n322745 , n322746 , n322747 , n322748 , n322749 , n322750 , n322751 , n322752 , n322753 , 
 n32328 , n322755 , n322756 , n32331 , n322758 , n322759 , n322760 , n322761 , n322762 , n322763 , 
 n322764 , n322765 , n322766 , n322767 , n32342 , n322769 , n322770 , n322771 , n322772 , n32347 , 
 n322774 , n322775 , n32350 , n322777 , n322778 , n322779 , n322780 , n322781 , n322782 , n322783 , 
 n322784 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n322792 , n32367 , 
 n322794 , n32369 , n32370 , n322797 , n322798 , n32373 , n322800 , n322801 , n32376 , n322803 , 
 n322804 , n32379 , n322806 , n322807 , n322808 , n322809 , n322810 , n322811 , n322812 , n32387 , 
 n322814 , n32389 , n322816 , n322817 , n322818 , n32393 , n322820 , n322821 , n322822 , n322823 , 
 n322824 , n322825 , n322826 , n322827 , n322828 , n322829 , n322830 , n322831 , n322832 , n322833 , 
 n322834 , n322835 , n322836 , n322837 , n32412 , n322839 , n322840 , n322841 , n322842 , n322843 , 
 n322844 , n322845 , n322846 , n32421 , n322848 , n322849 , n32424 , n322851 , n322852 , n32427 , 
 n322854 , n322855 , n32430 , n322857 , n322858 , n322859 , n322860 , n322861 , n322862 , n322863 , 
 n322864 , n322865 , n322866 , n322867 , n32442 , n322869 , n32444 , n322871 , n322872 , n32447 , 
 n322874 , n322875 , n322876 , n322877 , n322878 , n32453 , n32454 , n322881 , n32456 , n322883 , 
 n322884 , n32459 , n322886 , n32461 , n322888 , n322889 , n32464 , n322891 , n322892 , n322893 , 
 n32468 , n322895 , n322896 , n322897 , n322898 , n322899 , n322900 , n322901 , n32476 , n322903 , 
 n322904 , n322905 , n322906 , n322907 , n322908 , n322909 , n322910 , n322911 , n322912 , n322913 , 
 n32488 , n322915 , n32490 , n322917 , n322918 , n322919 , n32494 , n322921 , n32496 , n322923 , 
 n322924 , n32499 , n322926 , n322927 , n322928 , n322929 , n32504 , n322931 , n32506 , n322933 , 
 n322934 , n322935 , n32510 , n322937 , n32512 , n322939 , n322940 , n32515 , n322942 , n322943 , 
 n322944 , n32519 , n32520 , n322947 , n322948 , n32523 , n322950 , n32525 , n322952 , n322953 , 
 n322954 , n322955 , n322956 , n322957 , n32532 , n32533 , n322960 , n322961 , n322962 , n322963 , 
 n322964 , n32539 , n322966 , n322967 , n322968 , n32543 , n322970 , n322971 , n322972 , n32547 , 
 n322974 , n322975 , n322976 , n322977 , n322978 , n322979 , n322980 , n322981 , n322982 , n32557 , 
 n322984 , n322985 , n322986 , n322987 , n322988 , n322989 , n322990 , n322991 , n322992 , n322993 , 
 n322994 , n32569 , n322996 , n322997 , n322998 , n322999 , n32574 , n323001 , n323002 , n323003 , 
 n323004 , n32579 , n323006 , n323007 , n323008 , n323009 , n323010 , n323011 , n32586 , n323013 , 
 n323014 , n32589 , n32590 , n323017 , n323018 , n323019 , n323020 , n323021 , n323022 , n323023 , 
 n323024 , n323025 , n323026 , n323027 , n323028 , n323029 , n323030 , n323031 , n323032 , n323033 , 
 n32608 , n323035 , n323036 , n323037 , n323038 , n323039 , n323040 , n323041 , n32616 , n323043 , 
 n323044 , n323045 , n323046 , n323047 , n32622 , n323049 , n323050 , n323051 , n323052 , n323053 , 
 n32628 , n323055 , n323056 , n323057 , n32632 , n323059 , n323060 , n323061 , n32636 , n323063 , 
 n32638 , n32639 , n323066 , n323067 , n32642 , n323069 , n323070 , n323071 , n323072 , n323073 , 
 n32648 , n323075 , n323076 , n32651 , n323078 , n32653 , n323080 , n323081 , n323082 , n323083 , 
 n32658 , n323085 , n32660 , n32661 , n323088 , n323089 , n323090 , n323091 , n323092 , n32667 , 
 n32668 , n32669 , n32670 , n32671 , n323098 , n323099 , n32674 , n323101 , n323102 , n32677 , 
 n323104 , n323105 , n323106 , n32681 , n323108 , n32683 , n32684 , n323111 , n323112 , n323113 , 
 n323114 , n323115 , n323116 , n323117 , n323118 , n32693 , n323120 , n323121 , n323122 , n32697 , 
 n323124 , n323125 , n32700 , n323127 , n323128 , n32703 , n32704 , n323131 , n32706 , n32707 , 
 n323134 , n323135 , n32710 , n32711 , n32712 , n32713 , n32714 , n323141 , n323142 , n32717 , 
 n323144 , n323145 , n32720 , n32721 , n32722 , n32723 , n323150 , n323151 , n32726 , n32727 , 
 n32728 , n32729 , n323156 , n323157 , n32732 , n32733 , n32734 , n32735 , n32736 , n323163 , 
 n32738 , n32739 , n32740 , n323167 , n323168 , n32743 , n323170 , n323171 , n32746 , n32747 , 
 n32748 , n32749 , n32750 , n323177 , n323178 , n32753 , n323180 , n323181 , n32756 , n32757 , 
 n32758 , n32759 , n32760 , n323187 , n323188 , n323189 , n323190 , n32765 , n323192 , n32767 , 
 n32768 , n32769 , n323196 , n323197 , n323198 , n32773 , n323200 , n32775 , n32776 , n323203 , 
 n32778 , n323205 , n323206 , n323207 , n32782 , n32783 , n323210 , n323211 , n32786 , n32787 , 
 n32788 , n32789 , n323216 , n323217 , n32792 , n32793 , n32794 , n323221 , n323222 , n32797 , 
 n323224 , n323225 , n32800 , n32801 , n323228 , n32803 , n32804 , n323231 , n323232 , n32807 , 
 n32808 , n32809 , n32810 , n323237 , n323238 , n323239 , n323240 , n323241 , n323242 , n323243 , 
 n323244 , n323245 , n32820 , n32821 , n323248 , n32823 , n323250 , n323251 , n32826 , n323253 , 
 n323254 , n32829 , n32830 , n323257 , n32832 , n32833 , n32834 , n323261 , n323262 , n323263 , 
 n32838 , n323265 , n323266 , n32841 , n32842 , n323269 , n323270 , n32845 , n323272 , n323273 , 
 n32848 , n32849 , n32850 , n323277 , n32852 , n32853 , n323280 , n32855 , n323282 , n32857 , 
 n32858 , n323285 , n323286 , n32861 , n323288 , n323289 , n32864 , n323291 , n323292 , n323293 , 
 n32868 , n323295 , n32870 , n32871 , n323298 , n323299 , n32874 , n323301 , n323302 , n32877 , 
 n323304 , n323305 , n32880 , n323307 , n32882 , n323309 , n32884 , n32885 , n32886 , n323313 , 
 n323314 , n32889 , n323316 , n323317 , n32892 , n323319 , n323320 , n323321 , n32896 , n32897 , 
 n323324 , n323325 , n323326 , n323327 , n323328 , n32903 , n32904 , n323331 , n32906 , n323333 , 
 n323334 , n323335 , n32910 , n323337 , n32912 , n32913 , n323340 , n323341 , n32916 , n323343 , 
 n323344 , n32919 , n323346 , n323347 , n323348 , n323349 , n323350 , n32925 , n32926 , n323353 , 
 n323354 , n323355 , n323356 , n323357 , n323358 , n323359 , n323360 , n32935 , n323362 , n32937 , 
 n323364 , n32939 , n32940 , n323367 , n323368 , n32943 , n323370 , n323371 , n32946 , n323373 , 
 n323374 , n32949 , n323376 , n323377 , n32952 , n32953 , n32954 , n323381 , n323382 , n323383 , 
 n32958 , n323385 , n323386 , n32961 , n32962 , n32963 , n323390 , n323391 , n32966 , n32967 , 
 n32968 , n323395 , n323396 , n32971 , n32972 , n323399 , n323400 , n32975 , n323402 , n323403 , 
 n32978 , n323405 , n323406 , n32981 , n32982 , n32983 , n32984 , n323411 , n323412 , n32987 , 
 n32988 , n323415 , n323416 , n323417 , n323418 , n323419 , n323420 , n32995 , n323422 , n323423 , 
 n32998 , n323425 , n323426 , n33001 , n323428 , n323429 , n33004 , n33005 , n33006 , n33007 , 
 n33008 , n33009 , n33010 , n323437 , n33012 , n323439 , n323440 , n33015 , n33016 , n33017 , 
 n33018 , n33019 , n323446 , n323447 , n33022 , n323449 , n323450 , n33025 , n33026 , n33027 , 
 n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n323460 , n323461 , n323462 , n33037 , 
 n33038 , n323465 , n323466 , n323467 , n323468 , n323469 , n323470 , n323471 , n33046 , n323473 , 
 n323474 , n323475 , n33050 , n323477 , n323478 , n33053 , n323480 , n323481 , n33056 , n323483 , 
 n323484 , n33059 , n323486 , n323487 , n33062 , n323489 , n33064 , n323491 , n33066 , n33067 , 
 n323494 , n323495 , n33070 , n323497 , n323498 , n33073 , n323500 , n323501 , n33076 , n33077 , 
 n33078 , n323505 , n323506 , n33081 , n323508 , n33083 , n323510 , n323511 , n33086 , n323513 , 
 n323514 , n33089 , n323516 , n323517 , n323518 , n323519 , n323520 , n323521 , n33096 , n323523 , 
 n33098 , n33099 , n323526 , n323527 , n33102 , n323529 , n323530 , n33105 , n323532 , n323533 , 
 n33108 , n323535 , n33110 , n323537 , n323538 , n33113 , n323540 , n323541 , n33116 , n323543 , 
 n323544 , n323545 , n323546 , n323547 , n33122 , n33123 , n33124 , n323551 , n323552 , n33127 , 
 n323554 , n323555 , n33130 , n33131 , n33132 , n323559 , n323560 , n33135 , n33136 , n33137 , 
 n33138 , n323565 , n323566 , n33141 , n33142 , n33143 , n323570 , n323571 , n33146 , n33147 , 
 n33148 , n323575 , n323576 , n33151 , n323578 , n323579 , n33154 , n323581 , n33156 , n323583 , 
 n323584 , n33159 , n323586 , n323587 , n323588 , n33163 , n323590 , n323591 , n323592 , n33167 , 
 n33168 , n33169 , n33170 , n33171 , n323598 , n323599 , n33174 , n323601 , n323602 , n33177 , 
 n33178 , n33179 , n33180 , n33181 , n323608 , n323609 , n33184 , n33185 , n33186 , n323613 , 
 n323614 , n33189 , n33190 , n323617 , n323618 , n323619 , n323620 , n33195 , n33196 , n33197 , 
 n33198 , n33199 , n33200 , n323627 , n33202 , n323629 , n323630 , n323631 , n323632 , n33207 , 
 n323634 , n323635 , n323636 , n33211 , n323638 , n33213 , n323640 , n323641 , n33216 , n323643 , 
 n323644 , n33219 , n33220 , n33221 , n323648 , n323649 , n33224 , n323651 , n323652 , n33227 , 
 n323654 , n33229 , n33230 , n33231 , n33232 , n323659 , n33234 , n323661 , n33236 , n323663 , 
 n323664 , n33239 , n323666 , n323667 , n323668 , n323669 , n33244 , n323671 , n323672 , n33247 , 
 n323674 , n323675 , n33250 , n323677 , n323678 , n33253 , n323680 , n323681 , n33256 , n323683 , 
 n33258 , n323685 , n33260 , n323687 , n33262 , n33263 , n323690 , n323691 , n33266 , n323693 , 
 n323694 , n33269 , n323696 , n323697 , n323698 , n33273 , n33274 , n323701 , n33276 , n323703 , 
 n323704 , n33279 , n33280 , n323707 , n323708 , n33283 , n33284 , n323711 , n323712 , n33287 , 
 n33288 , n33289 , n33290 , n323717 , n323718 , n33293 , n33294 , n33295 , n33296 , n33297 , 
 n323724 , n33299 , n33300 , n33301 , n323728 , n323729 , n33304 , n33305 , n33306 , n323733 , 
 n323734 , n33309 , n33310 , n33311 , n323738 , n33313 , n33314 , n33315 , n33316 , n33317 , 
 n33318 , n323745 , n323746 , n33321 , n33322 , n33323 , n33324 , n323751 , n323752 , n33327 , 
 n33328 , n33329 , n323756 , n323757 , n33332 , n33333 , n33334 , n33335 , n323762 , n323763 , 
 n33338 , n33339 , n33340 , n323767 , n323768 , n33343 , n323770 , n323771 , n33346 , n323773 , 
 n323774 , n33349 , n323776 , n33351 , n323778 , n323779 , n33354 , n33355 , n33356 , n33357 , 
 n33358 , n33359 , n33360 , n323787 , n33362 , n323789 , n33364 , n323791 , n33366 , n33367 , 
 n323794 , n323795 , n33370 , n33371 , n323798 , n33373 , n33374 , n33375 , n33376 , n33377 , 
 n33378 , n33379 , n33380 , n323807 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , 
 n33388 , n33389 , n33390 , n323817 , n33392 , n33393 , n33394 , n33395 , n323822 , n33397 , 
 n323824 , n323825 , n33400 , n323827 , n323828 , n323829 , n323830 , n323831 , n33406 , n323833 , 
 n33408 , n323835 , n323836 , n33411 , n33412 , n33413 , n323840 , n323841 , n33416 , n323843 , 
 n323844 , n323845 , n323846 , n33421 , n323848 , n33423 , n33424 , n323851 , n33426 , n33427 , 
 n33428 , n33429 , n33430 , n33431 , n323858 , n323859 , n33434 , n33435 , n323862 , n323863 , 
 n33438 , n33439 , n33440 , n323867 , n33442 , n323869 , n33444 , n33445 , n323872 , n323873 , 
 n33448 , n33449 , n33450 , n33451 , n33452 , n323879 , n323880 , n33455 , n33456 , n33457 , 
 n323884 , n323885 , n33460 , n33461 , n323888 , n323889 , n33464 , n33465 , n33466 , n323893 , 
 n323894 , n33469 , n33470 , n33471 , n323898 , n323899 , n33474 , n323901 , n33476 , n33477 , 
 n33478 , n323905 , n323906 , n33481 , n33482 , n33483 , n33484 , n323911 , n33486 , n33487 , 
 n33488 , n323915 , n323916 , n33491 , n33492 , n33493 , n323920 , n323921 , n33496 , n33497 , 
 n33498 , n33499 , n323926 , n323927 , n33502 , n33503 , n323930 , n323931 , n33506 , n33507 , 
 n33508 , n323935 , n323936 , n33511 , n33512 , n33513 , n323940 , n323941 , n33516 , n33517 , 
 n33518 , n323945 , n323946 , n33521 , n33522 , n33523 , n323950 , n33525 , n33526 , n33527 , 
 n33528 , n33529 , n33530 , n33531 , n33532 , n323959 , n33534 , n33535 , n323962 , n33537 , 
 n33538 , n33539 , n33540 , n323967 , n323968 , n323969 , n33544 , n33545 , n33546 , n33547 , 
 n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , 
 n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , 
 n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n324001 , n324002 , n33577 , 
 n33578 , n33579 , n324006 , n324007 , n324008 , n324009 , n33584 , n33585 , n33586 , n33587 , 
 n324014 , n324015 , n324016 , n33591 , n33592 , n33593 , n324020 , n33595 , n33596 , n33597 , 
 n324024 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , 
 n33608 , n33609 , n33610 , n33611 , n33612 , n324039 , n33614 , n33615 , n33616 , n33617 , 
 n324044 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n324051 , n33626 , n33627 , 
 n324054 , n324055 , n33630 , n33631 , n324058 , n324059 , n33634 , n33635 , n33636 , n33637 , 
 n324064 , n324065 , n33640 , n33641 , n33642 , n324069 , n324070 , n324071 , n324072 , n324073 , 
 n33648 , n33649 , n324076 , n33651 , n324078 , n324079 , n324080 , n324081 , n324082 , n324083 , 
 n33658 , n33659 , n324086 , n324087 , n33662 , n33663 , n33664 , n324091 , n33666 , n33667 , 
 n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n324103 , 
 n324104 , n33679 , n324106 , n324107 , n33682 , n324109 , n33684 , n33685 , n324112 , n324113 , 
 n33688 , n324115 , n324116 , n33691 , n324118 , n33693 , n33694 , n33695 , n33696 , n33697 , 
 n33698 , n33699 , n33700 , n33701 , n324128 , n33703 , n324130 , n324131 , n33706 , n324133 , 
 n33708 , n33709 , n324136 , n324137 , n33712 , n324139 , n324140 , n33715 , n324142 , n33717 , 
 n324144 , n33719 , n324146 , n324147 , n324148 , n33723 , n324150 , n324151 , n33726 , n324153 , 
 n324154 , n324155 , n324156 , n324157 , n324158 , n324159 , n33734 , n33735 , n324162 , n324163 , 
 n33738 , n324165 , n324166 , n33741 , n324168 , n324169 , n33744 , n33745 , n33746 , n324173 , 
 n324174 , n33749 , n324176 , n33751 , n33752 , n324179 , n324180 , n33755 , n324182 , n324183 , 
 n33758 , n324185 , n33760 , n33761 , n324188 , n324189 , n33764 , n324191 , n324192 , n33767 , 
 n324194 , n324195 , n324196 , n33771 , n324198 , n324199 , n33774 , n324201 , n33776 , n33777 , 
 n324204 , n324205 , n33780 , n324207 , n324208 , n33783 , n324210 , n33785 , n324212 , n324213 , 
 n33788 , n324215 , n324216 , n33791 , n324218 , n33793 , n33794 , n324221 , n324222 , n33797 , 
 n324224 , n324225 , n33800 , n324227 , n33802 , n324229 , n324230 , n33805 , n324232 , n33807 , 
 n33808 , n33809 , n324236 , n33811 , n324238 , n33813 , n33814 , n324241 , n324242 , n33817 , 
 n324244 , n324245 , n33820 , n324247 , n324248 , n324249 , n324250 , n33825 , n324252 , n324253 , 
 n33828 , n324255 , n33830 , n324257 , n324258 , n324259 , n33834 , n324261 , n324262 , n33837 , 
 n324264 , n324265 , n33840 , n324267 , n324268 , n33843 , n324270 , n324271 , n33846 , n324273 , 
 n33848 , n33849 , n324276 , n324277 , n33852 , n324279 , n324280 , n33855 , n324282 , n324283 , 
 n33858 , n33859 , n33860 , n324287 , n33862 , n33863 , n33864 , n324291 , n324292 , n33867 , 
 n324294 , n324295 , n33870 , n324297 , n33872 , n33873 , n324300 , n324301 , n33876 , n324303 , 
 n324304 , n33879 , n324306 , n324307 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , 
 n324314 , n33889 , n324316 , n324317 , n324318 , n324319 , n324320 , n33895 , n33896 , n33897 , 
 n33898 , n324325 , n33900 , n33901 , n33902 , n324329 , n324330 , n33905 , n324332 , n33907 , 
 n33908 , n324335 , n33910 , n33911 , n324338 , n33913 , n324340 , n324341 , n33916 , n33917 , 
 n324344 , n324345 , n324346 , n33921 , n324348 , n324349 , n33924 , n324351 , n33926 , n33927 , 
 n324354 , n324355 , n33930 , n324357 , n324358 , n33933 , n324360 , n33935 , n324362 , n324363 , 
 n324364 , n33939 , n324366 , n33941 , n324368 , n324369 , n324370 , n33945 , n324372 , n33947 , 
 n324374 , n324375 , n324376 , n33951 , n324378 , n33953 , n33954 , n33955 , n324382 , n33957 , 
 n33958 , n324385 , n33960 , n33961 , n33962 , n324389 , n324390 , n33965 , n33966 , n33967 , 
 n324394 , n324395 , n33970 , n33971 , n33972 , n324399 , n324400 , n33975 , n33976 , n33977 , 
 n324404 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n324411 , n33986 , n33987 , 
 n33988 , n33989 , n324416 , n324417 , n33992 , n324419 , n33994 , n324421 , n33996 , n33997 , 
 n33998 , n33999 , n324426 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , 
 n324434 , n34009 , n34010 , n34011 , n34012 , n324439 , n34014 , n34015 , n34016 , n324443 , 
 n324444 , n34019 , n34020 , n34021 , n324448 , n34023 , n34024 , n34025 , n34026 , n324453 , 
 n34028 , n34029 , n34030 , n34031 , n34032 , n324459 , n34034 , n34035 , n34036 , n34037 , 
 n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , 
 n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , 
 n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , 
 n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , 
 n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , 
 n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n324522 , n324523 , 
 n34098 , n324525 , n324526 , n34101 , n324528 , n34103 , n34104 , n324531 , n324532 , n34107 , 
 n324534 , n324535 , n34110 , n324537 , n34112 , n324539 , n324540 , n34115 , n324542 , n324543 , 
 n34118 , n324545 , n34120 , n34121 , n324548 , n324549 , n34124 , n324551 , n324552 , n34127 , 
 n324554 , n34129 , n34130 , n34131 , n324558 , n324559 , n34134 , n324561 , n34136 , n324563 , 
 n324564 , n324565 , n324566 , n34141 , n324568 , n324569 , n324570 , n34145 , n324572 , n34147 , 
 n324574 , n324575 , n34150 , n324577 , n324578 , n34153 , n324580 , n34155 , n34156 , n324583 , 
 n324584 , n34159 , n324586 , n324587 , n34162 , n324589 , n34164 , n34165 , n34166 , n34167 , 
 n34168 , n34169 , n34170 , n324597 , n324598 , n34173 , n324600 , n34175 , n34176 , n34177 , 
 n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , 
 n324614 , n324615 , n34190 , n324617 , n324618 , n324619 , n34194 , n34195 , n34196 , n324623 , 
 n34198 , n324625 , n34200 , n34201 , n324628 , n34203 , n34204 , n34205 , n324632 , n34207 , 
 n34208 , n34209 , n324636 , n324637 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , 
 n324644 , n324645 , n34220 , n34221 , n34222 , n324649 , n34224 , n34225 , n324652 , n324653 , 
 n34228 , n34229 , n324656 , n324657 , n34232 , n34233 , n324660 , n324661 , n324662 , n34237 , 
 n324664 , n324665 , n34240 , n34241 , n324668 , n324669 , n324670 , n324671 , n34246 , n324673 , 
 n324674 , n34249 , n324676 , n34251 , n34252 , n324679 , n324680 , n324681 , n34256 , n324683 , 
 n324684 , n34259 , n324686 , n324687 , n34262 , n324689 , n324690 , n324691 , n34266 , n324693 , 
 n34268 , n34269 , n324696 , n324697 , n324698 , n34273 , n324700 , n324701 , n34276 , n324703 , 
 n324704 , n34279 , n324706 , n324707 , n34282 , n324709 , n324710 , n34285 , n324712 , n34287 , 
 n324714 , n324715 , n324716 , n324717 , n34292 , n324719 , n324720 , n324721 , n34296 , n324723 , 
 n324724 , n34299 , n324726 , n324727 , n34302 , n324729 , n34304 , n324731 , n34306 , n34307 , 
 n324734 , n324735 , n324736 , n34311 , n324738 , n324739 , n34314 , n324741 , n324742 , n34317 , 
 n324744 , n324745 , n324746 , n34321 , n324748 , n34323 , n34324 , n324751 , n324752 , n324753 , 
 n34328 , n324755 , n324756 , n34331 , n324758 , n324759 , n34334 , n324761 , n324762 , n34337 , 
 n34338 , n324765 , n324766 , n324767 , n324768 , n324769 , n324770 , n324771 , n34346 , n324773 , 
 n34348 , n34349 , n324776 , n34351 , n34352 , n34353 , n324780 , n324781 , n34356 , n34357 , 
 n34358 , n324785 , n324786 , n324787 , n324788 , n34363 , n324790 , n324791 , n34366 , n324793 , 
 n324794 , n34369 , n324796 , n324797 , n34372 , n324799 , n34374 , n34375 , n324802 , n324803 , 
 n324804 , n34379 , n324806 , n324807 , n34382 , n324809 , n324810 , n34385 , n324812 , n324813 , 
 n34388 , n34389 , n324816 , n324817 , n34392 , n324819 , n34394 , n324821 , n34396 , n34397 , 
 n324824 , n324825 , n34400 , n324827 , n324828 , n34403 , n324830 , n324831 , n34406 , n324833 , 
 n324834 , n34409 , n324836 , n324837 , n324838 , n324839 , n34414 , n324841 , n324842 , n34417 , 
 n324844 , n34419 , n34420 , n324847 , n324848 , n324849 , n34424 , n324851 , n324852 , n34427 , 
 n324854 , n324855 , n34430 , n324857 , n324858 , n34433 , n324860 , n324861 , n34436 , n324863 , 
 n324864 , n34439 , n324866 , n34441 , n34442 , n324869 , n324870 , n324871 , n34446 , n324873 , 
 n324874 , n34449 , n324876 , n324877 , n324878 , n324879 , n324880 , n34455 , n34456 , n324883 , 
 n324884 , n34459 , n324886 , n324887 , n34462 , n324889 , n324890 , n34465 , n324892 , n34467 , 
 n34468 , n324895 , n324896 , n324897 , n34472 , n324899 , n324900 , n34475 , n324902 , n324903 , 
 n34478 , n324905 , n324906 , n34481 , n324908 , n324909 , n34484 , n324911 , n324912 , n34487 , 
 n324914 , n34489 , n324916 , n34491 , n34492 , n324919 , n324920 , n34495 , n324922 , n324923 , 
 n34498 , n324925 , n324926 , n324927 , n324928 , n34503 , n324930 , n324931 , n34506 , n324933 , 
 n34508 , n34509 , n324936 , n324937 , n34512 , n324939 , n324940 , n34515 , n324942 , n324943 , 
 n34518 , n324945 , n34520 , n324947 , n34522 , n34523 , n324950 , n324951 , n34526 , n324953 , 
 n324954 , n34529 , n324956 , n324957 , n34532 , n324959 , n324960 , n34535 , n324962 , n324963 , 
 n34538 , n324965 , n324966 , n324967 , n34542 , n324969 , n324970 , n34545 , n34546 , n324973 , 
 n34548 , n324975 , n324976 , n34551 , n34552 , n324979 , n324980 , n324981 , n34556 , n34557 , 
 n324984 , n34559 , n324986 , n324987 , n34562 , n34563 , n324990 , n324991 , n34566 , n34567 , 
 n34568 , n34569 , n324996 , n324997 , n324998 , n34573 , n325000 , n325001 , n34576 , n325003 , 
 n34578 , n325005 , n325006 , n34581 , n325008 , n34583 , n34584 , n34585 , n325012 , n325013 , 
 n325014 , n34589 , n325016 , n325017 , n34592 , n325019 , n34594 , n34595 , n325022 , n325023 , 
 n34598 , n325025 , n34600 , n34601 , n34602 , n325029 , n325030 , n325031 , n34606 , n325033 , 
 n325034 , n34609 , n325036 , n34611 , n34612 , n325039 , n34614 , n34615 , n325042 , n325043 , 
 n34618 , n325045 , n325046 , n34621 , n325048 , n325049 , n34624 , n325051 , n34626 , n34627 , 
 n325054 , n325055 , n34630 , n325057 , n325058 , n325059 , n34634 , n325061 , n325062 , n34637 , 
 n325064 , n325065 , n325066 , n34641 , n325068 , n34643 , n34644 , n325071 , n325072 , n325073 , 
 n34648 , n325075 , n325076 , n34651 , n325078 , n325079 , n34654 , n325081 , n325082 , n34657 , 
 n325084 , n34659 , n325086 , n34661 , n34662 , n325089 , n34664 , n325091 , n34666 , n325093 , 
 n325094 , n34669 , n325096 , n325097 , n34672 , n325099 , n325100 , n34675 , n325102 , n325103 , 
 n34678 , n325105 , n325106 , n34681 , n34682 , n34683 , n325110 , n325111 , n34686 , n34687 , 
 n34688 , n325115 , n325116 , n34691 , n325118 , n34693 , n34694 , n34695 , n34696 , n325123 , 
 n325124 , n34699 , n325126 , n34701 , n34702 , n34703 , n34704 , n34705 , n325132 , n325133 , 
 n34708 , n325135 , n34710 , n34711 , n34712 , n34713 , n34714 , n325141 , n34716 , n34717 , 
 n325144 , n34719 , n34720 , n34721 , n34722 , n325149 , n325150 , n34725 , n325152 , n34727 , 
 n34728 , n34729 , n325156 , n34731 , n325158 , n34733 , n34734 , n325161 , n325162 , n34737 , 
 n325164 , n325165 , n34740 , n325167 , n34742 , n34743 , n34744 , n325171 , n34746 , n325173 , 
 n34748 , n34749 , n325176 , n325177 , n34752 , n325179 , n325180 , n34755 , n325182 , n34757 , 
 n34758 , n34759 , n325186 , n34761 , n34762 , n34763 , n325190 , n325191 , n34766 , n34767 , 
 n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , 
 n34778 , n34779 , n34780 , n34781 , n325208 , n34783 , n325210 , n34785 , n325212 , n325213 , 
 n34788 , n34789 , n325216 , n34791 , n325218 , n34793 , n325220 , n325221 , n34796 , n34797 , 
 n325224 , n34799 , n325226 , n34801 , n34802 , n325229 , n325230 , n34805 , n325232 , n325233 , 
 n34808 , n325235 , n325236 , n325237 , n34812 , n325239 , n34814 , n34815 , n325242 , n325243 , 
 n34818 , n325245 , n325246 , n34821 , n325248 , n325249 , n34824 , n325251 , n34826 , n325253 , 
 n34828 , n34829 , n325256 , n325257 , n34832 , n325259 , n325260 , n34835 , n325262 , n325263 , 
 n34838 , n325265 , n325266 , n325267 , n34842 , n325269 , n34844 , n34845 , n325272 , n325273 , 
 n34848 , n325275 , n325276 , n34851 , n325278 , n325279 , n34854 , n325281 , n34856 , n34857 , 
 n325284 , n325285 , n34860 , n325287 , n325288 , n34863 , n325290 , n34865 , n325292 , n325293 , 
 n325294 , n325295 , n34870 , n325297 , n325298 , n34873 , n325300 , n325301 , n325302 , n325303 , 
 n34878 , n325305 , n34880 , n325307 , n34882 , n325309 , n34884 , n34885 , n325312 , n325313 , 
 n34888 , n325315 , n325316 , n34891 , n325318 , n325319 , n34894 , n325321 , n34896 , n34897 , 
 n325324 , n325325 , n34900 , n325327 , n325328 , n34903 , n325330 , n34905 , n325332 , n325333 , 
 n34908 , n325335 , n325336 , n34911 , n34912 , n325339 , n34914 , n325341 , n34916 , n325343 , 
 n325344 , n325345 , n325346 , n325347 , n34922 , n325349 , n325350 , n325351 , n325352 , n34927 , 
 n325354 , n34929 , n325356 , n325357 , n34932 , n34933 , n325360 , n34935 , n325362 , n325363 , 
 n34938 , n34939 , n34940 , n34941 , n34942 , n325369 , n34944 , n325371 , n325372 , n34947 , 
 n34948 , n34949 , n34950 , n325377 , n325378 , n34953 , n34954 , n34955 , n34956 , n34957 , 
 n325384 , n325385 , n34960 , n325387 , n325388 , n34963 , n34964 , n325391 , n325392 , n325393 , 
 n325394 , n34969 , n34970 , n34971 , n34972 , n325399 , n325400 , n325401 , n34976 , n325403 , 
 n34978 , n34979 , n325406 , n325407 , n34982 , n325409 , n34984 , n325411 , n325412 , n34987 , 
 n325414 , n34989 , n34990 , n34991 , n34992 , n34993 , n325420 , n325421 , n34996 , n325423 , 
 n34998 , n34999 , n35000 , n35001 , n35002 , n325429 , n325430 , n35005 , n325432 , n35007 , 
 n35008 , n35009 , n35010 , n325437 , n325438 , n35013 , n325440 , n35015 , n325442 , n35017 , 
 n35018 , n325445 , n35020 , n35021 , n35022 , n35023 , n35024 , n325451 , n35026 , n35027 , 
 n35028 , n35029 , n325456 , n325457 , n35032 , n35033 , n325460 , n35035 , n35036 , n35037 , 
 n35038 , n35039 , n325466 , n325467 , n35042 , n325469 , n325470 , n325471 , n35046 , n325473 , 
 n35048 , n35049 , n325476 , n325477 , n35052 , n325479 , n325480 , n35055 , n35056 , n35057 , 
 n325484 , n325485 , n325486 , n35061 , n325488 , n35063 , n325490 , n325491 , n35066 , n35067 , 
 n325494 , n325495 , n35070 , n35071 , n325498 , n325499 , n325500 , n35075 , n35076 , n325503 , 
 n35078 , n35079 , n325506 , n325507 , n35082 , n325509 , n325510 , n35085 , n35086 , n35087 , 
 n325514 , n35089 , n325516 , n325517 , n325518 , n325519 , n35094 , n325521 , n325522 , n35097 , 
 n325524 , n325525 , n35100 , n325527 , n325528 , n35103 , n35104 , n35105 , n325532 , n35107 , 
 n35108 , n35109 , n35110 , n35111 , n325538 , n325539 , n35114 , n325541 , n35116 , n35117 , 
 n325544 , n325545 , n325546 , n35121 , n325548 , n325549 , n325550 , n35125 , n35126 , n35127 , 
 n325554 , n35129 , n35130 , n325557 , n325558 , n35133 , n35134 , n35135 , n35136 , n35137 , 
 n325564 , n325565 , n325566 , n325567 , n325568 , n35143 , n35144 , n35145 , n35146 , n325573 , 
 n325574 , n35149 , n35150 , n35151 , n325578 , n325579 , n35154 , n325581 , n35156 , n325583 , 
 n325584 , n35159 , n35160 , n35161 , n35162 , n325589 , n35164 , n325591 , n325592 , n325593 , 
 n35168 , n325595 , n325596 , n35171 , n325598 , n325599 , n35174 , n35175 , n35176 , n35177 , 
 n325604 , n325605 , n35180 , n325607 , n35182 , n325609 , n325610 , n35185 , n325612 , n35187 , 
 n325614 , n35189 , n325616 , n325617 , n35192 , n325619 , n35194 , n35195 , n35196 , n35197 , 
 n35198 , n35199 , n325626 , n325627 , n35202 , n35203 , n35204 , n35205 , n325632 , n325633 , 
 n35208 , n35209 , n35210 , n325637 , n325638 , n325639 , n35214 , n325641 , n35216 , n35217 , 
 n325644 , n325645 , n35220 , n35221 , n325648 , n325649 , n325650 , n35225 , n35226 , n325653 , 
 n35228 , n35229 , n325656 , n325657 , n35232 , n35233 , n35234 , n325661 , n325662 , n35237 , 
 n325664 , n325665 , n35240 , n325667 , n35242 , n35243 , n35244 , n35245 , n35246 , n325673 , 
 n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n325682 , n35257 , 
 n35258 , n325685 , n325686 , n35261 , n35262 , n325689 , n325690 , n35265 , n35266 , n35267 , 
 n35268 , n35269 , n325696 , n325697 , n35272 , n325699 , n35274 , n35275 , n35276 , n325703 , 
 n35278 , n35279 , n35280 , n35281 , n325708 , n35283 , n35284 , n35285 , n35286 , n35287 , 
 n35288 , n325715 , n35290 , n35291 , n325718 , n325719 , n35294 , n325721 , n325722 , n35297 , 
 n325724 , n325725 , n35300 , n325727 , n325728 , n325729 , n325730 , n325731 , n325732 , n35307 , 
 n325734 , n35309 , n35310 , n325737 , n325738 , n35313 , n325740 , n325741 , n35316 , n325743 , 
 n325744 , n325745 , n325746 , n35321 , n325748 , n325749 , n35324 , n325751 , n325752 , n35327 , 
 n35328 , n325755 , n325756 , n35331 , n35332 , n35333 , n325760 , n325761 , n35336 , n35337 , 
 n325764 , n325765 , n35340 , n35341 , n35342 , n35343 , n35344 , n325771 , n325772 , n35347 , 
 n35348 , n35349 , n35350 , n325777 , n325778 , n35353 , n35354 , n35355 , n35356 , n35357 , 
 n325784 , n325785 , n35360 , n35361 , n35362 , n325789 , n325790 , n35365 , n35366 , n35367 , 
 n325794 , n325795 , n35370 , n35371 , n325798 , n325799 , n35374 , n325801 , n325802 , n35377 , 
 n325804 , n35379 , n325806 , n325807 , n325808 , n325809 , n35384 , n325811 , n325812 , n35387 , 
 n325814 , n325815 , n35390 , n35391 , n325818 , n35393 , n35394 , n35395 , n325822 , n325823 , 
 n35398 , n35399 , n325826 , n325827 , n325828 , n35403 , n325830 , n325831 , n35406 , n35407 , 
 n35408 , n325835 , n325836 , n35411 , n325838 , n325839 , n325840 , n35415 , n35416 , n35417 , 
 n325844 , n325845 , n325846 , n325847 , n325848 , n325849 , n35424 , n325851 , n325852 , n325853 , 
 n325854 , n325855 , n35430 , n35431 , n35432 , n325859 , n35434 , n35435 , n325862 , n325863 , 
 n325864 , n325865 , n35440 , n325867 , n325868 , n325869 , n325870 , n325871 , n325872 , n325873 , 
 n35448 , n35449 , n325876 , n35451 , n35452 , n35453 , n325880 , n35455 , n35456 , n325883 , 
 n325884 , n35459 , n35460 , n325887 , n325888 , n35463 , n325890 , n325891 , n35466 , n35467 , 
 n325894 , n325895 , n325896 , n35471 , n325898 , n325899 , n325900 , n325901 , n325902 , n35477 , 
 n325904 , n325905 , n35480 , n325907 , n325908 , n35483 , n325910 , n325911 , n325912 , n325913 , 
 n35488 , n325915 , n325916 , n325917 , n325918 , n35493 , n325920 , n325921 , n325922 , n325923 , 
 n35498 , n325925 , n35500 , n35501 , n35502 , n325929 , n325930 , n35505 , n325932 , n325933 , 
 n35508 , n325935 , n35510 , n35511 , n325938 , n325939 , n35514 , n325941 , n35516 , n35517 , 
 n325944 , n325945 , n35520 , n325947 , n35522 , n35523 , n325950 , n325951 , n35526 , n325953 , 
 n35528 , n35529 , n325956 , n325957 , n35532 , n325959 , n325960 , n35535 , n325962 , n35537 , 
 n325964 , n325965 , n35540 , n325967 , n325968 , n325969 , n325970 , n35545 , n325972 , n325973 , 
 n35548 , n325975 , n35550 , n325977 , n325978 , n35553 , n325980 , n325981 , n35556 , n325983 , 
 n35558 , n35559 , n325986 , n325987 , n35562 , n325989 , n325990 , n35565 , n325992 , n35567 , 
 n35568 , n325995 , n325996 , n35571 , n325998 , n35573 , n35574 , n35575 , n326002 , n326003 , 
 n35578 , n326005 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , 
 n35588 , n326015 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , 
 n35598 , n35599 , n326026 , n326027 , n326028 , n326029 , n326030 , n326031 , n35606 , n326033 , 
 n35608 , n35609 , n326036 , n326037 , n35612 , n35613 , n326040 , n326041 , n35616 , n326043 , 
 n326044 , n35619 , n326046 , n326047 , n35622 , n326049 , n326050 , n35625 , n326052 , n326053 , 
 n326054 , n326055 , n35630 , n326057 , n35632 , n326059 , n35634 , n326061 , n326062 , n326063 , 
 n326064 , n35639 , n35640 , n35641 , n35642 , n326069 , n35644 , n326071 , n326072 , n326073 , 
 n35648 , n326075 , n326076 , n35651 , n326078 , n326079 , n326080 , n35655 , n326082 , n326083 , 
 n326084 , n35659 , n326086 , n326087 , n326088 , n326089 , n326090 , n35665 , n326092 , n326093 , 
 n326094 , n35669 , n326096 , n35671 , n326098 , n326099 , n326100 , n35675 , n326102 , n326103 , 
 n326104 , n35679 , n326106 , n326107 , n35682 , n326109 , n326110 , n35685 , n326112 , n35687 , 
 n35688 , n326115 , n35690 , n326117 , n326118 , n326119 , n35694 , n326121 , n35696 , n35697 , 
 n35698 , n35699 , n35700 , n35701 , n326128 , n326129 , n35704 , n326131 , n326132 , n35707 , 
 n326134 , n35709 , n35710 , n326137 , n326138 , n35713 , n326140 , n326141 , n35716 , n326143 , 
 n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , 
 n35728 , n326155 , n326156 , n35731 , n35732 , n35733 , n35734 , n326161 , n326162 , n35737 , 
 n35738 , n35739 , n326166 , n326167 , n35742 , n326169 , n35744 , n35745 , n35746 , n35747 , 
 n35748 , n326175 , n35750 , n35751 , n35752 , n35753 , n326180 , n326181 , n35756 , n326183 , 
 n35758 , n326185 , n326186 , n326187 , n35762 , n35763 , n35764 , n326191 , n326192 , n35767 , 
 n35768 , n35769 , n326196 , n35771 , n35772 , n326199 , n35774 , n326201 , n35776 , n35777 , 
 n326204 , n35779 , n35780 , n35781 , n35782 , n326209 , n35784 , n35785 , n35786 , n35787 , 
 n35788 , n35789 , n35790 , n35791 , n326218 , n35793 , n35794 , n35795 , n326222 , n326223 , 
 n35798 , n326225 , n326226 , n326227 , n35802 , n326229 , n35804 , n35805 , n326232 , n326233 , 
 n35808 , n326235 , n326236 , n326237 , n35812 , n326239 , n326240 , n35815 , n326242 , n326243 , 
 n35818 , n326245 , n326246 , n35821 , n326248 , n326249 , n35824 , n326251 , n35826 , n326253 , 
 n326254 , n326255 , n326256 , n35831 , n326258 , n326259 , n326260 , n326261 , n326262 , n326263 , 
 n326264 , n326265 , n326266 , n326267 , n35842 , n326269 , n326270 , n35845 , n326272 , n326273 , 
 n35848 , n326275 , n326276 , n35851 , n326278 , n326279 , n326280 , n35855 , n326282 , n326283 , 
 n35858 , n326285 , n35860 , n35861 , n35862 , n326289 , n326290 , n326291 , n326292 , n326293 , 
 n326294 , n326295 , n326296 , n35871 , n35872 , n326299 , n326300 , n35875 , n35876 , n35877 , 
 n326304 , n35879 , n326306 , n326307 , n35882 , n35883 , n326310 , n326311 , n326312 , n35887 , 
 n326314 , n326315 , n326316 , n326317 , n326318 , n326319 , n326320 , n326321 , n326322 , n326323 , 
 n326324 , n326325 , n35900 , n326327 , n35902 , n326329 , n326330 , n326331 , n35906 , n326333 , 
 n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n326340 , n35915 , n326342 , n35917 , 
 n35918 , n35919 , n35920 , n35921 , n326348 , n35923 , n35924 , n35925 , n35926 , n35927 , 
 n35928 , n35929 , n35930 , n326357 , n326358 , n35933 , n326360 , n326361 , n35936 , n326363 , 
 n35938 , n35939 , n326366 , n326367 , n35942 , n326369 , n326370 , n35945 , n326372 , n35947 , 
 n326374 , n35949 , n326376 , n35951 , n35952 , n326379 , n326380 , n35955 , n326382 , n326383 , 
 n35958 , n326385 , n326386 , n326387 , n35962 , n326389 , n35964 , n326391 , n326392 , n35967 , 
 n326394 , n326395 , n326396 , n35971 , n326398 , n35973 , n35974 , n35975 , n35976 , n35977 , 
 n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n326410 , n326411 , n35986 , n326413 , 
 n326414 , n35989 , n326416 , n326417 , n35992 , n326419 , n35994 , n326421 , n35996 , n35997 , 
 n326424 , n326425 , n36000 , n326427 , n326428 , n36003 , n326430 , n326431 , n36006 , n36007 , 
 n326434 , n36009 , n326436 , n326437 , n36012 , n326439 , n36014 , n36015 , n326442 , n36017 , 
 n326444 , n36019 , n36020 , n326447 , n326448 , n36023 , n326450 , n326451 , n36026 , n326453 , 
 n326454 , n36029 , n326456 , n326457 , n36032 , n326459 , n326460 , n36035 , n326462 , n326463 , 
 n36038 , n326465 , n326466 , n326467 , n36042 , n326469 , n326470 , n36045 , n36046 , n326473 , 
 n326474 , n36049 , n36050 , n326477 , n36052 , n36053 , n36054 , n36055 , n326482 , n36057 , 
 n326484 , n36059 , n36060 , n326487 , n326488 , n36063 , n326490 , n326491 , n36066 , n326493 , 
 n326494 , n36069 , n36070 , n36071 , n36072 , n326499 , n326500 , n326501 , n36076 , n326503 , 
 n36078 , n326505 , n326506 , n326507 , n326508 , n36083 , n326510 , n326511 , n326512 , n326513 , 
 n36088 , n326515 , n36090 , n36091 , n326518 , n326519 , n326520 , n326521 , n326522 , n326523 , 
 n36098 , n326525 , n36100 , n36101 , n326528 , n326529 , n36104 , n326531 , n326532 , n36107 , 
 n326534 , n36109 , n36110 , n36111 , n326538 , n36113 , n326540 , n36115 , n326542 , n36117 , 
 n36118 , n36119 , n36120 , n326547 , n326548 , n36123 , n326550 , n36125 , n326552 , n326553 , 
 n326554 , n326555 , n36130 , n36131 , n36132 , n326559 , n36134 , n36135 , n36136 , n36137 , 
 n36138 , n36139 , n36140 , n326567 , n36142 , n326569 , n326570 , n36145 , n326572 , n326573 , 
 n326574 , n326575 , n36150 , n36151 , n36152 , n326579 , n36154 , n36155 , n36156 , n36157 , 
 n36158 , n326585 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n326593 , 
 n36168 , n326595 , n36170 , n326597 , n326598 , n36173 , n326600 , n326601 , n36176 , n326603 , 
 n36178 , n326605 , n36180 , n326607 , n326608 , n36183 , n326610 , n36185 , n36186 , n36187 , 
 n36188 , n36189 , n36190 , n36191 , n326618 , n36193 , n36194 , n36195 , n326622 , n36197 , 
 n326624 , n36199 , n326626 , n326627 , n36202 , n326629 , n36204 , n36205 , n36206 , n36207 , 
 n326634 , n36209 , n326636 , n326637 , n36212 , n326639 , n326640 , n36215 , n36216 , n36217 , 
 n36218 , n326645 , n36220 , n36221 , n326648 , n326649 , n36224 , n326651 , n326652 , n36227 , 
 n326654 , n36229 , n326656 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , 
 n36238 , n36239 , n36240 , n36241 , n36242 , n326669 , n36244 , n326671 , n326672 , n36247 , 
 n36248 , n36249 , n36250 , n326677 , n36252 , n36253 , n326680 , n326681 , n36256 , n326683 , 
 n326684 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n326691 , n36266 , n36267 , 
 n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , 
 n36278 , n36279 , n36280 , n326707 , n326708 , n36283 , n326710 , n36285 , n36286 , n326713 , 
 n36288 , n326715 , n326716 , n36291 , n326718 , n326719 , n36294 , n326721 , n326722 , n36297 , 
 n36298 , n36299 , n36300 , n36301 , n36302 , n326729 , n36304 , n326731 , n326732 , n36307 , 
 n326734 , n326735 , n36310 , n36311 , n36312 , n36313 , n326740 , n326741 , n326742 , n36317 , 
 n326744 , n326745 , n326746 , n326747 , n36322 , n326749 , n326750 , n36325 , n326752 , n326753 , 
 n36328 , n326755 , n326756 , n326757 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , 
 n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , 
 n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , 
 n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , 
 n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , 
 n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , 
 n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n326820 , n36395 , n36396 , n36397 , 
 n36398 , n326825 , n326826 , n36401 , n36402 , n36403 , n36404 , n326831 , n326832 , n326833 , 
 n36408 , n326835 , n36410 , n36411 , n326838 , n36413 , n326840 , n36415 , n326842 , n326843 , 
 n36418 , n326845 , n326846 , n36421 , n326848 , n36423 , n326850 , n36425 , n36426 , n36427 , 
 n326854 , n36429 , n326856 , n36431 , n326858 , n36433 , n36434 , n326861 , n326862 , n326863 , 
 n36438 , n326865 , n326866 , n36441 , n326868 , n326869 , n36444 , n326871 , n326872 , n36447 , 
 n326874 , n326875 , n36450 , n326877 , n326878 , n326879 , n36454 , n326881 , n36456 , n326883 , 
 n326884 , n326885 , n326886 , n36461 , n326888 , n326889 , n36464 , n326891 , n326892 , n36467 , 
 n36468 , n326895 , n36470 , n326897 , n326898 , n326899 , n36474 , n36475 , n326902 , n326903 , 
 n326904 , n36479 , n326906 , n326907 , n36482 , n326909 , n326910 , n36485 , n326912 , n326913 , 
 n326914 , n326915 , n36490 , n326917 , n326918 , n36493 , n326920 , n326921 , n326922 , n326923 , 
 n326924 , n326925 , n326926 , n326927 , n326928 , n326929 , n326930 , n326931 , n326932 , n326933 , 
 n326934 , n326935 , n326936 , n326937 , n326938 , n326939 , n326940 , n326941 , n326942 , n36517 , 
 n36518 , n36519 , n326946 , n326947 , n36522 , n326949 , n36524 , n36525 , n36526 , n36527 , 
 n36528 , n36529 , n36530 , n326957 , n36532 , n36533 , n326960 , n36535 , n36536 , n36537 , 
 n36538 , n326965 , n36540 , n36541 , n36542 , n326969 , n36544 , n36545 , n326972 , n326973 , 
 n36548 , n326975 , n326976 , n36551 , n326978 , n36553 , n36554 , n36555 , n36556 , n36557 , 
 n36558 , n326985 , n326986 , n36561 , n326988 , n326989 , n326990 , n36565 , n326992 , n326993 , 
 n36568 , n326995 , n326996 , n36571 , n326998 , n36573 , n327000 , n36575 , n36576 , n327003 , 
 n327004 , n36579 , n327006 , n327007 , n36582 , n327009 , n36584 , n36585 , n327012 , n327013 , 
 n36588 , n327015 , n327016 , n36591 , n327018 , n327019 , n36594 , n327021 , n327022 , n36597 , 
 n327024 , n327025 , n36600 , n327027 , n36602 , n327029 , n327030 , n36605 , n36606 , n36607 , 
 n327034 , n36609 , n327036 , n327037 , n327038 , n36613 , n327040 , n327041 , n36616 , n327043 , 
 n327044 , n327045 , n327046 , n36621 , n327048 , n36623 , n327050 , n36625 , n36626 , n36627 , 
 n36628 , n327055 , n327056 , n327057 , n36632 , n327059 , n327060 , n36635 , n327062 , n327063 , 
 n327064 , n327065 , n327066 , n36641 , n327068 , n327069 , n36644 , n327071 , n36646 , n36647 , 
 n327074 , n36649 , n327076 , n36651 , n36652 , n327079 , n36654 , n327081 , n327082 , n36657 , 
 n327084 , n327085 , n36660 , n327087 , n36662 , n327089 , n36664 , n36665 , n327092 , n327093 , 
 n36668 , n327095 , n327096 , n327097 , n327098 , n36673 , n327100 , n36675 , n327102 , n36677 , 
 n36678 , n36679 , n36680 , n327107 , n36682 , n327109 , n327110 , n36685 , n327112 , n327113 , 
 n327114 , n36689 , n327116 , n36691 , n36692 , n327119 , n36694 , n327121 , n36696 , n327123 , 
 n327124 , n327125 , n327126 , n327127 , n36702 , n327129 , n327130 , n327131 , n327132 , n36707 , 
 n327134 , n327135 , n36710 , n327137 , n327138 , n36713 , n327140 , n36715 , n327142 , n327143 , 
 n327144 , n36719 , n36720 , n327147 , n327148 , n327149 , n327150 , n327151 , n327152 , n327153 , 
 n36728 , n327155 , n327156 , n327157 , n327158 , n327159 , n327160 , n327161 , n327162 , n36737 , 
 n327164 , n327165 , n36740 , n327167 , n327168 , n327169 , n36744 , n327171 , n327172 , n327173 , 
 n327174 , n327175 , n327176 , n327177 , n327178 , n36753 , n327180 , n327181 , n36756 , n327183 , 
 n327184 , n327185 , n327186 , n327187 , n327188 , n327189 , n327190 , n327191 , n327192 , n327193 , 
 n327194 , n327195 , n327196 , n327197 , n327198 , n327199 , n36774 , n327201 , n327202 , n327203 , 
 n327204 , n327205 , n327206 , n327207 , n327208 , n327209 , n327210 , n327211 , n36786 , n36787 , 
 n36788 , n327215 , n327216 , n327217 , n327218 , n36793 , n327220 , n327221 , n327222 , n327223 , 
 n327224 , n327225 , n327226 , n327227 , n327228 , n327229 , n36804 , n327231 , n36806 , n327233 , 
 n327234 , n327235 , n327236 , n327237 , n327238 , n36813 , n327240 , n36815 , n36816 , n327243 , 
 n327244 , n36819 , n327246 , n327247 , n36822 , n327249 , n327250 , n327251 , n327252 , n327253 , 
 n327254 , n327255 , n327256 , n327257 , n327258 , n327259 , n327260 , n327261 , n327262 , n327263 , 
 n327264 , n36839 , n327266 , n327267 , n327268 , n327269 , n327270 , n327271 , n327272 , n36847 , 
 n327274 , n327275 , n36850 , n327277 , n327278 , n327279 , n327280 , n327281 , n327282 , n327283 , 
 n327284 , n327285 , n327286 , n327287 , n36862 , n36863 , n327290 , n327291 , n36866 , n327293 , 
 n327294 , n327295 , n36870 , n327297 , n327298 , n327299 , n36874 , n327301 , n327302 , n327303 , 
 n327304 , n327305 , n36880 , n327307 , n327308 , n327309 , n36884 , n327311 , n327312 , n36887 , 
 n327314 , n327315 , n36890 , n327317 , n36892 , n327319 , n327320 , n36895 , n327322 , n327323 , 
 n327324 , n36899 , n327326 , n327327 , n36902 , n36903 , n36904 , n36905 , n36906 , n327333 , 
 n327334 , n36909 , n327336 , n327337 , n327338 , n327339 , n327340 , n36915 , n36916 , n36917 , 
 n327344 , n327345 , n327346 , n327347 , n36922 , n327349 , n327350 , n327351 , n36926 , n327353 , 
 n327354 , n327355 , n36930 , n327357 , n327358 , n327359 , n36934 , n327361 , n327362 , n327363 , 
 n36938 , n327365 , n327366 , n36941 , n327368 , n36943 , n36944 , n327371 , n327372 , n36947 , 
 n327374 , n327375 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n327383 , 
 n36958 , n327385 , n327386 , n36961 , n327388 , n327389 , n36964 , n36965 , n36966 , n36967 , 
 n327394 , n327395 , n36970 , n327397 , n36972 , n327399 , n327400 , n327401 , n36976 , n327403 , 
 n327404 , n327405 , n327406 , n36981 , n327408 , n327409 , n36984 , n327411 , n36986 , n327413 , 
 n327414 , n36989 , n327416 , n36991 , n36992 , n36993 , n36994 , n36995 , n327422 , n36997 , 
 n327424 , n36999 , n37000 , n327427 , n37002 , n327429 , n37004 , n327431 , n37006 , n327433 , 
 n327434 , n37009 , n37010 , n37011 , n37012 , n327439 , n327440 , n37015 , n327442 , n37017 , 
 n327444 , n327445 , n327446 , n37021 , n327448 , n327449 , n327450 , n37025 , n327452 , n327453 , 
 n37028 , n327455 , n37030 , n37031 , n327458 , n37033 , n327460 , n327461 , n37036 , n327463 , 
 n37038 , n37039 , n327466 , n37041 , n327468 , n327469 , n37044 , n327471 , n327472 , n37047 , 
 n327474 , n327475 , n37050 , n37051 , n37052 , n37053 , n327480 , n327481 , n37056 , n327483 , 
 n37058 , n327485 , n327486 , n37061 , n327488 , n327489 , n327490 , n37065 , n327492 , n37067 , 
 n37068 , n327495 , n37070 , n327497 , n327498 , n327499 , n327500 , n327501 , n37076 , n37077 , 
 n327504 , n327505 , n327506 , n37081 , n327508 , n327509 , n327510 , n327511 , n327512 , n37087 , 
 n327514 , n327515 , n327516 , n37091 , n327518 , n327519 , n327520 , n327521 , n327522 , n327523 , 
 n327524 , n327525 , n327526 , n37101 , n327528 , n37103 , n327530 , n327531 , n37106 , n327533 , 
 n327534 , n327535 , n327536 , n327537 , n327538 , n327539 , n327540 , n327541 , n327542 , n37117 , 
 n327544 , n327545 , n327546 , n37121 , n37122 , n37123 , n327550 , n327551 , n327552 , n327553 , 
 n327554 , n327555 , n327556 , n327557 , n327558 , n327559 , n37134 , n37135 , n37136 , n327563 , 
 n37138 , n327565 , n327566 , n37141 , n37142 , n327569 , n327570 , n327571 , n37146 , n327573 , 
 n327574 , n327575 , n327576 , n327577 , n327578 , n327579 , n327580 , n327581 , n37156 , n327583 , 
 n327584 , n37159 , n327586 , n327587 , n327588 , n37163 , n327590 , n37165 , n327592 , n327593 , 
 n327594 , n327595 , n327596 , n327597 , n327598 , n327599 , n37174 , n327601 , n327602 , n327603 , 
 n327604 , n327605 , n327606 , n37181 , n327608 , n327609 , n327610 , n37185 , n327612 , n327613 , 
 n327614 , n327615 , n327616 , n37191 , n327618 , n327619 , n327620 , n327621 , n327622 , n327623 , 
 n327624 , n37199 , n327626 , n327627 , n37202 , n327629 , n37204 , n327631 , n327632 , n327633 , 
 n327634 , n327635 , n327636 , n327637 , n327638 , n37213 , n37214 , n37215 , n37216 , n327643 , 
 n327644 , n327645 , n327646 , n37221 , n327648 , n327649 , n37224 , n37225 , n37226 , n327653 , 
 n37228 , n327655 , n327656 , n37231 , n37232 , n37233 , n37234 , n327661 , n37236 , n327663 , 
 n327664 , n327665 , n37240 , n327667 , n327668 , n327669 , n327670 , n327671 , n327672 , n37247 , 
 n327674 , n327675 , n327676 , n37251 , n327678 , n327679 , n327680 , n327681 , n327682 , n327683 , 
 n37258 , n327685 , n327686 , n37261 , n327688 , n327689 , n37264 , n327691 , n327692 , n37267 , 
 n327694 , n327695 , n327696 , n327697 , n37272 , n327699 , n37274 , n327701 , n327702 , n327703 , 
 n37278 , n37279 , n327706 , n327707 , n37282 , n327709 , n327710 , n327711 , n37286 , n327713 , 
 n327714 , n327715 , n327716 , n327717 , n327718 , n327719 , n37294 , n37295 , n37296 , n37297 , 
 n37298 , n327725 , n327726 , n37301 , n327728 , n327729 , n37304 , n37305 , n37306 , n327733 , 
 n327734 , n37309 , n37310 , n327737 , n327738 , n327739 , n327740 , n327741 , n327742 , n327743 , 
 n327744 , n327745 , n327746 , n327747 , n327748 , n37323 , n327750 , n327751 , n37326 , n327753 , 
 n327754 , n327755 , n37330 , n37331 , n37332 , n37333 , n327760 , n327761 , n327762 , n327763 , 
 n327764 , n327765 , n327766 , n327767 , n327768 , n327769 , n327770 , n327771 , n327772 , n327773 , 
 n327774 , n327775 , n37350 , n327777 , n327778 , n37353 , n327780 , n327781 , n327782 , n327783 , 
 n327784 , n327785 , n327786 , n327787 , n327788 , n327789 , n327790 , n327791 , n327792 , n327793 , 
 n327794 , n327795 , n37370 , n37371 , n327798 , n327799 , n327800 , n327801 , n327802 , n327803 , 
 n327804 , n37379 , n327806 , n327807 , n37382 , n37383 , n327810 , n327811 , n327812 , n37387 , 
 n327814 , n327815 , n327816 , n327817 , n37392 , n327819 , n37394 , n327821 , n327822 , n37397 , 
 n327824 , n327825 , n37400 , n37401 , n37402 , n37403 , n327830 , n37405 , n327832 , n327833 , 
 n37408 , n327835 , n327836 , n37411 , n327838 , n327839 , n37414 , n327841 , n37416 , n37417 , 
 n37418 , n37419 , n327846 , n37421 , n37422 , n37423 , n37424 , n327851 , n327852 , n37427 , 
 n327854 , n37429 , n327856 , n327857 , n327858 , n37433 , n327860 , n327861 , n37436 , n327863 , 
 n37438 , n327865 , n37440 , n37441 , n327868 , n37443 , n327870 , n37445 , n327872 , n37447 , 
 n37448 , n37449 , n37450 , n327877 , n327878 , n37453 , n327880 , n37455 , n327882 , n327883 , 
 n37458 , n327885 , n327886 , n37461 , n37462 , n37463 , n37464 , n327891 , n37466 , n327893 , 
 n327894 , n37469 , n327896 , n327897 , n37472 , n37473 , n37474 , n37475 , n327902 , n37477 , 
 n37478 , n37479 , n37480 , n327907 , n327908 , n327909 , n37484 , n327911 , n327912 , n37487 , 
 n327914 , n327915 , n327916 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , 
 n37498 , n37499 , n327926 , n37501 , n37502 , n37503 , n37504 , n327931 , n37506 , n327933 , 
 n327934 , n37509 , n327936 , n327937 , n327938 , n37513 , n37514 , n327941 , n37516 , n327943 , 
 n327944 , n37519 , n327946 , n37521 , n37522 , n327949 , n327950 , n37525 , n327952 , n327953 , 
 n37528 , n37529 , n327956 , n37531 , n327958 , n327959 , n37534 , n327961 , n327962 , n37537 , 
 n327964 , n327965 , n37540 , n37541 , n37542 , n37543 , n327970 , n327971 , n327972 , n37547 , 
 n327974 , n327975 , n327976 , n37551 , n327978 , n327979 , n327980 , n37555 , n327982 , n37557 , 
 n37558 , n327985 , n37560 , n327987 , n327988 , n37563 , n37564 , n37565 , n37566 , n327993 , 
 n327994 , n327995 , n37570 , n327997 , n327998 , n37573 , n328000 , n328001 , n328002 , n328003 , 
 n37578 , n328005 , n37580 , n37581 , n328008 , n37583 , n328010 , n328011 , n37586 , n37587 , 
 n37588 , n37589 , n328016 , n328017 , n328018 , n37593 , n328020 , n328021 , n37596 , n328023 , 
 n328024 , n328025 , n328026 , n328027 , n328028 , n328029 , n328030 , n37605 , n328032 , n328033 , 
 n328034 , n328035 , n328036 , n328037 , n328038 , n37613 , n328040 , n328041 , n328042 , n328043 , 
 n328044 , n328045 , n328046 , n37621 , n37622 , n328049 , n328050 , n328051 , n37626 , n37627 , 
 n328054 , n328055 , n37630 , n328057 , n328058 , n328059 , n37634 , n37635 , n328062 , n37637 , 
 n328064 , n37639 , n328066 , n37641 , n328068 , n37643 , n328070 , n37645 , n328072 , n328073 , 
 n37648 , n37649 , n37650 , n37651 , n328078 , n37653 , n328080 , n37655 , n328082 , n37657 , 
 n328084 , n328085 , n37660 , n328087 , n328088 , n37663 , n328090 , n328091 , n37666 , n328093 , 
 n328094 , n37669 , n37670 , n37671 , n37672 , n328099 , n328100 , n328101 , n37676 , n328103 , 
 n328104 , n328105 , n328106 , n328107 , n328108 , n328109 , n328110 , n328111 , n328112 , n37687 , 
 n328114 , n37689 , n328116 , n328117 , n37692 , n37693 , n328120 , n37695 , n37696 , n37697 , 
 n37698 , n328125 , n328126 , n328127 , n37702 , n328129 , n328130 , n328131 , n37706 , n328133 , 
 n37708 , n328135 , n328136 , n37711 , n328138 , n328139 , n328140 , n328141 , n328142 , n328143 , 
 n328144 , n328145 , n37720 , n328147 , n328148 , n328149 , n328150 , n37725 , n328152 , n328153 , 
 n328154 , n328155 , n328156 , n37731 , n328158 , n328159 , n328160 , n328161 , n328162 , n328163 , 
 n328164 , n328165 , n328166 , n37741 , n328168 , n328169 , n37744 , n328171 , n328172 , n328173 , 
 n37748 , n328175 , n328176 , n328177 , n328178 , n328179 , n328180 , n37755 , n328182 , n328183 , 
 n328184 , n328185 , n328186 , n37761 , n37762 , n328189 , n37764 , n328191 , n37766 , n328193 , 
 n328194 , n328195 , n328196 , n328197 , n328198 , n37773 , n37774 , n37775 , n328202 , n328203 , 
 n37778 , n328205 , n328206 , n328207 , n328208 , n328209 , n37784 , n328211 , n328212 , n328213 , 
 n328214 , n328215 , n328216 , n328217 , n328218 , n328219 , n328220 , n328221 , n328222 , n328223 , 
 n328224 , n328225 , n328226 , n328227 , n328228 , n37803 , n328230 , n328231 , n328232 , n328233 , 
 n37808 , n37809 , n37810 , n328237 , n328238 , n328239 , n328240 , n37815 , n328242 , n328243 , 
 n37818 , n328245 , n328246 , n328247 , n328248 , n328249 , n37824 , n328251 , n328252 , n37827 , 
 n328254 , n328255 , n328256 , n328257 , n37832 , n328259 , n328260 , n328261 , n328262 , n328263 , 
 n328264 , n328265 , n328266 , n328267 , n328268 , n328269 , n328270 , n37845 , n328272 , n328273 , 
 n328274 , n328275 , n328276 , n328277 , n37852 , n328279 , n328280 , n328281 , n328282 , n328283 , 
 n328284 , n37859 , n328286 , n328287 , n328288 , n328289 , n37864 , n328291 , n328292 , n328293 , 
 n328294 , n328295 , n37870 , n328297 , n328298 , n328299 , n328300 , n37875 , n328302 , n37877 , 
 n37878 , n328305 , n328306 , n328307 , n328308 , n328309 , n328310 , n328311 , n328312 , n37887 , 
 n328314 , n328315 , n37890 , n328317 , n328318 , n328319 , n328320 , n328321 , n328322 , n328323 , 
 n328324 , n328325 , n328326 , n328327 , n328328 , n328329 , n328330 , n328331 , n328332 , n328333 , 
 n328334 , n328335 , n37910 , n37911 , n328338 , n328339 , n37914 , n328341 , n328342 , n328343 , 
 n37918 , n328345 , n328346 , n328347 , n328348 , n37923 , n328350 , n37925 , n328352 , n328353 , 
 n328354 , n328355 , n328356 , n328357 , n328358 , n328359 , n328360 , n328361 , n37936 , n37937 , 
 n328364 , n37939 , n328366 , n328367 , n328368 , n328369 , n37944 , n328371 , n37946 , n328373 , 
 n328374 , n328375 , n328376 , n328377 , n328378 , n328379 , n328380 , n328381 , n328382 , n328383 , 
 n328384 , n328385 , n328386 , n328387 , n328388 , n328389 , n328390 , n328391 , n328392 , n328393 , 
 n37968 , n37969 , n328396 , n328397 , n328398 , n328399 , n328400 , n328401 , n37976 , n328403 , 
 n37978 , n37979 , n328406 , n328407 , n328408 , n328409 , n328410 , n328411 , n328412 , n328413 , 
 n37988 , n37989 , n328416 , n328417 , n328418 , n328419 , n328420 , n328421 , n328422 , n328423 , 
 n328424 , n328425 , n328426 , n328427 , n38002 , n38003 , n328430 , n328431 , n38006 , n328433 , 
 n328434 , n328435 , n38010 , n328437 , n328438 , n38013 , n328440 , n328441 , n38016 , n328443 , 
 n328444 , n38019 , n328446 , n38021 , n328448 , n328449 , n38024 , n328451 , n328452 , n328453 , 
 n328454 , n38029 , n328456 , n328457 , n38032 , n328459 , n328460 , n38035 , n328462 , n328463 , 
 n38038 , n38039 , n328466 , n328467 , n328468 , n328469 , n38044 , n328471 , n328472 , n328473 , 
 n328474 , n328475 , n328476 , n328477 , n328478 , n328479 , n328480 , n38055 , n328482 , n38057 , 
 n328484 , n328485 , n328486 , n38061 , n38062 , n38063 , n328490 , n328491 , n328492 , n328493 , 
 n328494 , n328495 , n328496 , n328497 , n38072 , n328499 , n328500 , n328501 , n328502 , n328503 , 
 n328504 , n328505 , n328506 , n328507 , n328508 , n328509 , n328510 , n38085 , n328512 , n328513 , 
 n328514 , n328515 , n328516 , n328517 , n38092 , n328519 , n328520 , n38095 , n328522 , n328523 , 
 n328524 , n328525 , n328526 , n328527 , n38102 , n38103 , n38104 , n38105 , n38106 , n328533 , 
 n328534 , n328535 , n328536 , n38111 , n328538 , n38113 , n38114 , n328541 , n328542 , n328543 , 
 n328544 , n38119 , n38120 , n328547 , n328548 , n328549 , n328550 , n328551 , n38126 , n328553 , 
 n38128 , n38129 , n38130 , n38131 , n328558 , n38133 , n328560 , n328561 , n328562 , n328563 , 
 n328564 , n38139 , n328566 , n38141 , n328568 , n328569 , n38144 , n328571 , n328572 , n328573 , 
 n328574 , n328575 , n328576 , n328577 , n38152 , n38153 , n328580 , n38155 , n38156 , n328583 , 
 n38158 , n328585 , n328586 , n328587 , n328588 , n328589 , n328590 , n328591 , n38166 , n328593 , 
 n328594 , n328595 , n328596 , n328597 , n328598 , n328599 , n328600 , n38175 , n328602 , n328603 , 
 n38178 , n328605 , n328606 , n38181 , n38182 , n328609 , n38184 , n328611 , n328612 , n328613 , 
 n38188 , n328615 , n38190 , n328617 , n328618 , n328619 , n328620 , n328621 , n328622 , n328623 , 
 n328624 , n328625 , n328626 , n328627 , n328628 , n328629 , n38204 , n328631 , n328632 , n38207 , 
 n328634 , n328635 , n328636 , n328637 , n328638 , n328639 , n38214 , n328641 , n328642 , n38217 , 
 n328644 , n328645 , n328646 , n328647 , n328648 , n328649 , n328650 , n328651 , n328652 , n328653 , 
 n328654 , n328655 , n328656 , n328657 , n38232 , n38233 , n328660 , n328661 , n328662 , n328663 , 
 n328664 , n38239 , n328666 , n328667 , n328668 , n328669 , n38244 , n38245 , n38246 , n38247 , 
 n38248 , n328675 , n38250 , n38251 , n328678 , n38253 , n328680 , n328681 , n38256 , n328683 , 
 n328684 , n328685 , n328686 , n328687 , n38262 , n328689 , n328690 , n328691 , n328692 , n38267 , 
 n38268 , n328695 , n38270 , n38271 , n38272 , n38273 , n328700 , n38275 , n328702 , n328703 , 
 n328704 , n38279 , n328706 , n328707 , n328708 , n38283 , n38284 , n328711 , n328712 , n328713 , 
 n328714 , n38289 , n328716 , n328717 , n328718 , n328719 , n38294 , n328721 , n328722 , n328723 , 
 n38298 , n328725 , n328726 , n38301 , n328728 , n328729 , n38304 , n328731 , n328732 , n38307 , 
 n328734 , n38309 , n328736 , n328737 , n328738 , n328739 , n328740 , n328741 , n328742 , n328743 , 
 n328744 , n328745 , n328746 , n328747 , n328748 , n38323 , n328750 , n328751 , n328752 , n328753 , 
 n38328 , n328755 , n328756 , n328757 , n328758 , n38333 , n328760 , n328761 , n328762 , n328763 , 
 n328764 , n328765 , n328766 , n328767 , n328768 , n328769 , n328770 , n328771 , n328772 , n328773 , 
 n328774 , n328775 , n328776 , n328777 , n38352 , n328779 , n328780 , n328781 , n38356 , n328783 , 
 n328784 , n38359 , n328786 , n328787 , n38362 , n38363 , n38364 , n328791 , n328792 , n328793 , 
 n328794 , n328795 , n328796 , n38371 , n328798 , n328799 , n328800 , n328801 , n328802 , n328803 , 
 n328804 , n38379 , n328806 , n328807 , n38382 , n38383 , n38384 , n328811 , n328812 , n328813 , 
 n328814 , n328815 , n328816 , n38391 , n328818 , n328819 , n328820 , n328821 , n328822 , n328823 , 
 n328824 , n38399 , n328826 , n328827 , n38402 , n328829 , n38404 , n328831 , n328832 , n328833 , 
 n328834 , n328835 , n328836 , n328837 , n328838 , n38413 , n328840 , n38415 , n38416 , n328843 , 
 n328844 , n328845 , n38420 , n328847 , n38422 , n328849 , n38424 , n38425 , n328852 , n328853 , 
 n38428 , n328855 , n328856 , n328857 , n328858 , n328859 , n328860 , n38435 , n38436 , n328863 , 
 n328864 , n38439 , n328866 , n328867 , n328868 , n328869 , n328870 , n328871 , n38446 , n328873 , 
 n328874 , n328875 , n328876 , n38451 , n38452 , n328879 , n328880 , n328881 , n38456 , n328883 , 
 n328884 , n328885 , n38460 , n328887 , n328888 , n328889 , n328890 , n328891 , n38466 , n328893 , 
 n38468 , n328895 , n328896 , n328897 , n328898 , n38473 , n328900 , n328901 , n38476 , n328903 , 
 n328904 , n38479 , n328906 , n38481 , n328908 , n328909 , n328910 , n328911 , n328912 , n38487 , 
 n328914 , n38489 , n328916 , n328917 , n38492 , n328919 , n38494 , n38495 , n38496 , n38497 , 
 n328924 , n328925 , n38500 , n328927 , n328928 , n328929 , n328930 , n328931 , n328932 , n38507 , 
 n328934 , n328935 , n38510 , n328937 , n328938 , n328939 , n328940 , n328941 , n38516 , n328943 , 
 n328944 , n38519 , n38520 , n328947 , n328948 , n328949 , n328950 , n328951 , n328952 , n328953 , 
 n328954 , n328955 , n328956 , n328957 , n328958 , n328959 , n38534 , n328961 , n328962 , n38537 , 
 n328964 , n328965 , n328966 , n328967 , n328968 , n328969 , n328970 , n38545 , n328972 , n328973 , 
 n328974 , n328975 , n328976 , n328977 , n38552 , n328979 , n328980 , n328981 , n328982 , n328983 , 
 n328984 , n328985 , n328986 , n38561 , n328988 , n328989 , n328990 , n328991 , n328992 , n38567 , 
 n328994 , n328995 , n328996 , n328997 , n328998 , n328999 , n329000 , n329001 , n38576 , n329003 , 
 n329004 , n329005 , n38580 , n329007 , n329008 , n38583 , n329010 , n329011 , n38586 , n329013 , 
 n329014 , n329015 , n329016 , n329017 , n329018 , n329019 , n329020 , n329021 , n329022 , n329023 , 
 n329024 , n329025 , n38600 , n329027 , n329028 , n329029 , n329030 , n329031 , n329032 , n329033 , 
 n329034 , n329035 , n38610 , n329037 , n329038 , n329039 , n329040 , n329041 , n329042 , n329043 , 
 n329044 , n329045 , n329046 , n38621 , n329048 , n329049 , n329050 , n38625 , n329052 , n329053 , 
 n38628 , n329055 , n329056 , n38631 , n38632 , n329059 , n329060 , n329061 , n329062 , n329063 , 
 n329064 , n329065 , n329066 , n38641 , n329068 , n329069 , n329070 , n329071 , n329072 , n38647 , 
 n329074 , n329075 , n38650 , n329077 , n329078 , n38653 , n38654 , n329081 , n329082 , n329083 , 
 n329084 , n329085 , n38660 , n329087 , n329088 , n38663 , n329090 , n329091 , n329092 , n329093 , 
 n329094 , n329095 , n38670 , n329097 , n329098 , n329099 , n329100 , n329101 , n329102 , n329103 , 
 n329104 , n38679 , n38680 , n329107 , n329108 , n329109 , n329110 , n329111 , n329112 , n329113 , 
 n329114 , n329115 , n329116 , n329117 , n329118 , n329119 , n38694 , n38695 , n329122 , n329123 , 
 n329124 , n38699 , n329126 , n329127 , n38702 , n329129 , n329130 , n329131 , n38706 , n329133 , 
 n329134 , n329135 , n38710 , n38711 , n329138 , n329139 , n329140 , n329141 , n329142 , n38717 , 
 n329144 , n329145 , n38720 , n329147 , n329148 , n329149 , n329150 , n329151 , n329152 , n329153 , 
 n329154 , n329155 , n38730 , n329157 , n329158 , n329159 , n329160 , n329161 , n329162 , n329163 , 
 n329164 , n38739 , n38740 , n329167 , n329168 , n329169 , n38744 , n329171 , n329172 , n38747 , 
 n329174 , n329175 , n329176 , n329177 , n329178 , n38753 , n329180 , n329181 , n329182 , n329183 , 
 n329184 , n329185 , n329186 , n329187 , n38762 , n329189 , n329190 , n38765 , n329192 , n329193 , 
 n329194 , n38769 , n329196 , n329197 , n329198 , n38773 , n329200 , n329201 , n329202 , n38777 , 
 n329204 , n329205 , n329206 , n329207 , n329208 , n329209 , n329210 , n329211 , n329212 , n38787 , 
 n329214 , n329215 , n329216 , n38791 , n329218 , n329219 , n38794 , n38795 , n38796 , n38797 , 
 n329224 , n329225 , n329226 , n38801 , n38802 , n38803 , n329230 , n329231 , n38806 , n38807 , 
 n329234 , n38809 , n38810 , n329237 , n38812 , n329239 , n329240 , n38815 , n329242 , n329243 , 
 n329244 , n38819 , n38820 , n38821 , n38822 , n329249 , n329250 , n329251 , n38826 , n329253 , 
 n38828 , n329255 , n329256 , n38831 , n329258 , n329259 , n38834 , n329261 , n329262 , n329263 , 
 n38838 , n329265 , n329266 , n38841 , n329268 , n329269 , n38844 , n329271 , n329272 , n38847 , 
 n329274 , n329275 , n38850 , n329277 , n329278 , n38853 , n329280 , n329281 , n38856 , n329283 , 
 n329284 , n38859 , n329286 , n329287 , n38862 , n329289 , n329290 , n329291 , n329292 , n329293 , 
 n38868 , n38869 , n38870 , n329297 , n329298 , n38873 , n329300 , n329301 , n38876 , n329303 , 
 n38878 , n329305 , n329306 , n329307 , n329308 , n329309 , n329310 , n38885 , n329312 , n329313 , 
 n38888 , n329315 , n329316 , n38891 , n329318 , n329319 , n329320 , n329321 , n329322 , n329323 , 
 n329324 , n329325 , n329326 , n329327 , n329328 , n329329 , n329330 , n329331 , n329332 , n329333 , 
 n38908 , n329335 , n38910 , n38911 , n329338 , n38913 , n329340 , n329341 , n38916 , n329343 , 
 n329344 , n38919 , n329346 , n329347 , n329348 , n329349 , n329350 , n329351 , n329352 , n38927 , 
 n329354 , n38929 , n38930 , n329357 , n329358 , n329359 , n329360 , n329361 , n329362 , n38937 , 
 n329364 , n329365 , n329366 , n329367 , n329368 , n38943 , n329370 , n329371 , n38946 , n329373 , 
 n329374 , n38949 , n329376 , n329377 , n329378 , n329379 , n329380 , n38955 , n329382 , n329383 , 
 n329384 , n38959 , n329386 , n329387 , n329388 , n329389 , n329390 , n38965 , n329392 , n329393 , 
 n329394 , n38969 , n329396 , n329397 , n38972 , n329399 , n38974 , n38975 , n38976 , n38977 , 
 n329404 , n38979 , n38980 , n38981 , n329408 , n329409 , n329410 , n329411 , n329412 , n329413 , 
 n38988 , n329415 , n38990 , n329417 , n329418 , n38993 , n329420 , n38995 , n329422 , n329423 , 
 n38998 , n329425 , n329426 , n39001 , n329428 , n39003 , n329430 , n329431 , n329432 , n329433 , 
 n39008 , n329435 , n329436 , n329437 , n329438 , n329439 , n39014 , n329441 , n329442 , n329443 , 
 n329444 , n329445 , n329446 , n329447 , n329448 , n329449 , n39024 , n329451 , n329452 , n329453 , 
 n39028 , n329455 , n329456 , n39031 , n329458 , n39033 , n39034 , n329461 , n39036 , n329463 , 
 n39038 , n39039 , n329466 , n39041 , n329468 , n329469 , n39044 , n329471 , n329472 , n39047 , 
 n329474 , n39049 , n39050 , n39051 , n39052 , n329479 , n39054 , n39055 , n39056 , n329483 , 
 n329484 , n329485 , n329486 , n329487 , n329488 , n329489 , n329490 , n329491 , n329492 , n39067 , 
 n329494 , n329495 , n329496 , n39071 , n329498 , n39073 , n329500 , n329501 , n329502 , n39077 , 
 n329504 , n39079 , n329506 , n329507 , n39082 , n329509 , n329510 , n39085 , n329512 , n329513 , 
 n329514 , n329515 , n329516 , n329517 , n329518 , n329519 , n39094 , n329521 , n329522 , n39097 , 
 n329524 , n329525 , n39100 , n329527 , n329528 , n39103 , n329530 , n39105 , n329532 , n329533 , 
 n329534 , n39109 , n39110 , n329537 , n329538 , n39113 , n329540 , n39115 , n329542 , n329543 , 
 n329544 , n329545 , n329546 , n329547 , n329548 , n39123 , n329550 , n329551 , n329552 , n329553 , 
 n329554 , n39129 , n329556 , n329557 , n329558 , n329559 , n39134 , n329561 , n329562 , n39137 , 
 n39138 , n329565 , n39140 , n39141 , n329568 , n329569 , n329570 , n329571 , n329572 , n329573 , 
 n329574 , n329575 , n39150 , n39151 , n329578 , n39153 , n329580 , n329581 , n39156 , n329583 , 
 n329584 , n329585 , n39160 , n329587 , n329588 , n329589 , n329590 , n39165 , n329592 , n329593 , 
 n39168 , n329595 , n329596 , n329597 , n329598 , n329599 , n329600 , n329601 , n39176 , n329603 , 
 n329604 , n39179 , n329606 , n39181 , n329608 , n329609 , n39184 , n329611 , n329612 , n39187 , 
 n329614 , n329615 , n39190 , n329617 , n39192 , n39193 , n329620 , n329621 , n39196 , n39197 , 
 n329624 , n329625 , n329626 , n329627 , n329628 , n329629 , n329630 , n329631 , n329632 , n329633 , 
 n329634 , n39209 , n329636 , n329637 , n39212 , n329639 , n329640 , n329641 , n39216 , n39217 , 
 n329644 , n39219 , n39220 , n39221 , n39222 , n39223 , n329650 , n329651 , n329652 , n329653 , 
 n39228 , n329655 , n39230 , n329657 , n39232 , n329659 , n329660 , n329661 , n329662 , n39237 , 
 n329664 , n329665 , n39240 , n329667 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , 
 n39248 , n329675 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n329682 , n329683 , 
 n329684 , n329685 , n39260 , n329687 , n329688 , n39263 , n329690 , n39265 , n39266 , n39267 , 
 n329694 , n329695 , n329696 , n39271 , n329698 , n329699 , n39274 , n329701 , n39276 , n39277 , 
 n329704 , n329705 , n329706 , n39281 , n329708 , n39283 , n329710 , n329711 , n329712 , n39287 , 
 n329714 , n329715 , n39290 , n329717 , n39292 , n329719 , n329720 , n39295 , n329722 , n329723 , 
 n39298 , n329725 , n39300 , n39301 , n39302 , n329729 , n329730 , n39305 , n329732 , n329733 , 
 n329734 , n329735 , n39310 , n39311 , n329738 , n329739 , n329740 , n329741 , n329742 , n329743 , 
 n329744 , n329745 , n329746 , n329747 , n39322 , n329749 , n329750 , n39325 , n39326 , n329753 , 
 n329754 , n329755 , n329756 , n39331 , n329758 , n39333 , n39334 , n39335 , n329762 , n329763 , 
 n329764 , n329765 , n329766 , n329767 , n39342 , n39343 , n329770 , n329771 , n329772 , n329773 , 
 n329774 , n329775 , n329776 , n329777 , n329778 , n329779 , n329780 , n329781 , n329782 , n39357 , 
 n39358 , n39359 , n329786 , n39361 , n329788 , n329789 , n329790 , n329791 , n329792 , n329793 , 
 n329794 , n39369 , n39370 , n329797 , n329798 , n329799 , n39374 , n39375 , n39376 , n39377 , 
 n39378 , n329805 , n39380 , n39381 , n329808 , n329809 , n329810 , n39385 , n329812 , n39387 , 
 n39388 , n329815 , n329816 , n39391 , n329818 , n329819 , n39394 , n39395 , n39396 , n329823 , 
 n39398 , n329825 , n329826 , n329827 , n329828 , n329829 , n329830 , n329831 , n329832 , n329833 , 
 n329834 , n329835 , n329836 , n329837 , n39412 , n329839 , n329840 , n39415 , n329842 , n329843 , 
 n39418 , n329845 , n329846 , n329847 , n329848 , n329849 , n329850 , n329851 , n39426 , n329853 , 
 n329854 , n39429 , n329856 , n329857 , n39432 , n329859 , n329860 , n39435 , n329862 , n329863 , 
 n329864 , n39439 , n329866 , n329867 , n39442 , n329869 , n329870 , n329871 , n39446 , n329873 , 
 n329874 , n329875 , n39450 , n329877 , n329878 , n329879 , n329880 , n39455 , n329882 , n329883 , 
 n329884 , n329885 , n329886 , n39461 , n329888 , n39463 , n329890 , n329891 , n329892 , n39467 , 
 n329894 , n329895 , n329896 , n329897 , n329898 , n329899 , n329900 , n329901 , n329902 , n329903 , 
 n39478 , n329905 , n39480 , n329907 , n329908 , n39483 , n329910 , n329911 , n329912 , n329913 , 
 n329914 , n329915 , n329916 , n39491 , n329918 , n39493 , n329920 , n329921 , n329922 , n39497 , 
 n329924 , n39499 , n329926 , n329927 , n39502 , n329929 , n329930 , n39505 , n329932 , n329933 , 
 n39508 , n329935 , n329936 , n329937 , n329938 , n329939 , n329940 , n329941 , n329942 , n329943 , 
 n329944 , n329945 , n39520 , n329947 , n329948 , n329949 , n329950 , n329951 , n329952 , n329953 , 
 n329954 , n329955 , n39530 , n39531 , n329958 , n39533 , n329960 , n329961 , n39536 , n329963 , 
 n329964 , n329965 , n329966 , n329967 , n329968 , n329969 , n329970 , n329971 , n329972 , n329973 , 
 n329974 , n329975 , n329976 , n329977 , n329978 , n329979 , n329980 , n39555 , n329982 , n39557 , 
 n39558 , n39559 , n39560 , n329987 , n39562 , n329989 , n329990 , n329991 , n329992 , n329993 , 
 n39568 , n329995 , n329996 , n39571 , n329998 , n329999 , n39574 , n330001 , n330002 , n39577 , 
 n330004 , n39579 , n330006 , n330007 , n330008 , n330009 , n330010 , n330011 , n330012 , n330013 , 
 n330014 , n39589 , n39590 , n39591 , n330018 , n39593 , n330020 , n330021 , n39596 , n330023 , 
 n39598 , n330025 , n39600 , n39601 , n330028 , n39603 , n330030 , n330031 , n39606 , n330033 , 
 n330034 , n330035 , n330036 , n39611 , n330038 , n39613 , n330040 , n39615 , n330042 , n330043 , 
 n330044 , n330045 , n330046 , n39621 , n330048 , n330049 , n330050 , n330051 , n330052 , n330053 , 
 n330054 , n330055 , n330056 , n330057 , n39632 , n39633 , n330060 , n39635 , n39636 , n330063 , 
 n330064 , n330065 , n39640 , n330067 , n330068 , n39643 , n330070 , n330071 , n330072 , n330073 , 
 n330074 , n330075 , n330076 , n330077 , n39652 , n330079 , n330080 , n39655 , n330082 , n330083 , 
 n330084 , n39659 , n330086 , n330087 , n330088 , n330089 , n330090 , n39665 , n39666 , n39667 , 
 n39668 , n39669 , n330096 , n39671 , n39672 , n330099 , n39674 , n330101 , n330102 , n330103 , 
 n39678 , n330105 , n330106 , n330107 , n330108 , n39683 , n330110 , n330111 , n330112 , n330113 , 
 n330114 , n330115 , n330116 , n330117 , n330118 , n330119 , n39694 , n39695 , n39696 , n330123 , 
 n39698 , n330125 , n330126 , n330127 , n39702 , n330129 , n330130 , n39705 , n330132 , n39707 , 
 n330134 , n330135 , n39710 , n39711 , n330138 , n330139 , n39714 , n330141 , n330142 , n39717 , 
 n330144 , n39719 , n330146 , n330147 , n330148 , n39723 , n39724 , n39725 , n39726 , n330153 , 
 n39728 , n330155 , n330156 , n330157 , n330158 , n330159 , n330160 , n330161 , n330162 , n330163 , 
 n330164 , n39739 , n330166 , n330167 , n330168 , n330169 , n39744 , n39745 , n39746 , n39747 , 
 n330174 , n330175 , n39750 , n330177 , n330178 , n330179 , n330180 , n39755 , n330182 , n330183 , 
 n39758 , n39759 , n330186 , n39761 , n330188 , n330189 , n330190 , n39765 , n330192 , n330193 , 
 n39768 , n330195 , n330196 , n39771 , n39772 , n39773 , n330200 , n39775 , n39776 , n330203 , 
 n39778 , n39779 , n330206 , n330207 , n39782 , n330209 , n330210 , n39785 , n330212 , n330213 , 
 n330214 , n330215 , n39790 , n330217 , n330218 , n39793 , n330220 , n330221 , n39796 , n330223 , 
 n330224 , n39799 , n39800 , n330227 , n39802 , n39803 , n330230 , n330231 , n330232 , n39807 , 
 n330234 , n330235 , n330236 , n330237 , n330238 , n330239 , n39814 , n330241 , n39816 , n39817 , 
 n39818 , n39819 , n330246 , n330247 , n330248 , n330249 , n330250 , n39825 , n330252 , n330253 , 
 n39828 , n330255 , n330256 , n330257 , n330258 , n39833 , n330260 , n330261 , n39836 , n330263 , 
 n330264 , n39839 , n39840 , n330267 , n39842 , n330269 , n330270 , n39845 , n39846 , n39847 , 
 n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n330280 , n330281 , n39856 , n330283 , 
 n330284 , n39859 , n330286 , n330287 , n330288 , n330289 , n330290 , n330291 , n330292 , n330293 , 
 n39868 , n330295 , n330296 , n330297 , n330298 , n39873 , n39874 , n39875 , n39876 , n330303 , 
 n330304 , n330305 , n330306 , n330307 , n330308 , n330309 , n330310 , n330311 , n330312 , n330313 , 
 n330314 , n330315 , n330316 , n39891 , n330318 , n330319 , n330320 , n39895 , n330322 , n330323 , 
 n39898 , n330325 , n330326 , n39901 , n330328 , n330329 , n330330 , n330331 , n330332 , n330333 , 
 n39908 , n330335 , n330336 , n39911 , n330338 , n330339 , n330340 , n330341 , n330342 , n330343 , 
 n330344 , n330345 , n330346 , n330347 , n330348 , n330349 , n330350 , n330351 , n330352 , n330353 , 
 n330354 , n39929 , n39930 , n39931 , n330358 , n39933 , n330360 , n330361 , n330362 , n330363 , 
 n330364 , n330365 , n330366 , n330367 , n330368 , n39943 , n330370 , n330371 , n330372 , n330373 , 
 n330374 , n330375 , n330376 , n330377 , n330378 , n330379 , n330380 , n330381 , n39956 , n330383 , 
 n330384 , n330385 , n330386 , n39961 , n330388 , n330389 , n330390 , n330391 , n39966 , n330393 , 
 n330394 , n330395 , n330396 , n330397 , n330398 , n330399 , n330400 , n39975 , n330402 , n330403 , 
 n39978 , n330405 , n330406 , n39981 , n330408 , n330409 , n330410 , n330411 , n330412 , n330413 , 
 n330414 , n330415 , n330416 , n39991 , n330418 , n39993 , n39994 , n39995 , n330422 , n330423 , 
 n330424 , n330425 , n330426 , n330427 , n330428 , n330429 , n330430 , n330431 , n40006 , n330433 , 
 n40008 , n330435 , n330436 , n330437 , n330438 , n40013 , n330440 , n330441 , n330442 , n330443 , 
 n40018 , n330445 , n330446 , n40021 , n330448 , n40023 , n330450 , n330451 , n330452 , n330453 , 
 n40028 , n330455 , n330456 , n40031 , n330458 , n330459 , n330460 , n330461 , n330462 , n40037 , 
 n330464 , n330465 , n40040 , n330467 , n330468 , n330469 , n330470 , n330471 , n330472 , n330473 , 
 n330474 , n330475 , n330476 , n40051 , n330478 , n330479 , n330480 , n330481 , n40056 , n40057 , 
 n330484 , n40059 , n40060 , n330487 , n330488 , n330489 , n330490 , n330491 , n330492 , n40067 , 
 n330494 , n330495 , n330496 , n330497 , n330498 , n40073 , n40074 , n40075 , n40076 , n330503 , 
 n40078 , n330505 , n330506 , n330507 , n330508 , n330509 , n40084 , n330511 , n330512 , n330513 , 
 n330514 , n40089 , n330516 , n40091 , n40092 , n330519 , n330520 , n330521 , n330522 , n330523 , 
 n330524 , n330525 , n330526 , n330527 , n330528 , n330529 , n330530 , n330531 , n40106 , n40107 , 
 n330534 , n330535 , n40110 , n330537 , n330538 , n40113 , n330540 , n40115 , n330542 , n330543 , 
 n330544 , n330545 , n330546 , n40121 , n330548 , n330549 , n330550 , n330551 , n40126 , n40127 , 
 n40128 , n330555 , n330556 , n330557 , n40132 , n330559 , n330560 , n330561 , n330562 , n40137 , 
 n330564 , n40139 , n330566 , n330567 , n40142 , n330569 , n40144 , n40145 , n40146 , n330573 , 
 n330574 , n40149 , n330576 , n330577 , n330578 , n330579 , n330580 , n330581 , n330582 , n330583 , 
 n330584 , n40159 , n330586 , n330587 , n40162 , n330589 , n330590 , n40165 , n330592 , n330593 , 
 n330594 , n330595 , n330596 , n330597 , n330598 , n330599 , n330600 , n330601 , n330602 , n330603 , 
 n330604 , n330605 , n330606 , n330607 , n330608 , n330609 , n40184 , n40185 , n40186 , n330613 , 
 n330614 , n330615 , n330616 , n330617 , n330618 , n330619 , n330620 , n330621 , n330622 , n330623 , 
 n40198 , n330625 , n330626 , n330627 , n330628 , n330629 , n330630 , n330631 , n330632 , n330633 , 
 n330634 , n330635 , n330636 , n330637 , n330638 , n330639 , n330640 , n330641 , n40216 , n330643 , 
 n330644 , n40219 , n330646 , n330647 , n40222 , n330649 , n330650 , n40225 , n330652 , n330653 , 
 n40228 , n330655 , n330656 , n40231 , n330658 , n330659 , n330660 , n330661 , n330662 , n330663 , 
 n330664 , n330665 , n330666 , n330667 , n330668 , n330669 , n330670 , n330671 , n330672 , n330673 , 
 n330674 , n330675 , n330676 , n330677 , n330678 , n330679 , n330680 , n40255 , n40256 , n330683 , 
 n40258 , n330685 , n40260 , n330687 , n330688 , n330689 , n330690 , n330691 , n330692 , n330693 , 
 n330694 , n330695 , n330696 , n330697 , n330698 , n330699 , n330700 , n330701 , n330702 , n330703 , 
 n330704 , n330705 , n330706 , n330707 , n40282 , n330709 , n330710 , n330711 , n330712 , n40287 , 
 n330714 , n330715 , n330716 , n330717 , n330718 , n330719 , n330720 , n330721 , n330722 , n330723 , 
 n330724 , n40299 , n330726 , n330727 , n330728 , n330729 , n330730 , n330731 , n330732 , n330733 , 
 n40308 , n330735 , n40310 , n330737 , n330738 , n330739 , n330740 , n40315 , n330742 , n330743 , 
 n40318 , n330745 , n330746 , n330747 , n330748 , n330749 , n330750 , n330751 , n330752 , n40327 , 
 n330754 , n330755 , n40330 , n330757 , n40332 , n40333 , n330760 , n330761 , n330762 , n330763 , 
 n330764 , n330765 , n330766 , n330767 , n330768 , n330769 , n330770 , n330771 , n330772 , n330773 , 
 n330774 , n330775 , n330776 , n330777 , n330778 , n330779 , n330780 , n40355 , n40356 , n330783 , 
 n40358 , n330785 , n330786 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , 
 n330794 , n40369 , n330796 , n330797 , n40372 , n40373 , n40374 , n40375 , n330802 , n330803 , 
 n40378 , n330805 , n330806 , n330807 , n40382 , n330809 , n330810 , n40385 , n40386 , n40387 , 
 n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , 
 n40398 , n40399 , n330826 , n40401 , n330828 , n330829 , n330830 , n330831 , n330832 , n330833 , 
 n330834 , n330835 , n330836 , n40411 , n330838 , n40413 , n330840 , n40415 , n40416 , n40417 , 
 n40418 , n330845 , n40420 , n330847 , n40422 , n330849 , n330850 , n330851 , n330852 , n40427 , 
 n330854 , n330855 , n330856 , n330857 , n330858 , n40433 , n40434 , n40435 , n330862 , n40437 , 
 n330864 , n330865 , n40440 , n40441 , n330868 , n40443 , n330870 , n330871 , n40446 , n40447 , 
 n330874 , n330875 , n330876 , n40451 , n40452 , n40453 , n40454 , n330881 , n330882 , n330883 , 
 n330884 , n330885 , n330886 , n330887 , n330888 , n330889 , n330890 , n40465 , n330892 , n40467 , 
 n40468 , n330895 , n330896 , n330897 , n40472 , n330899 , n40474 , n330901 , n40476 , n330903 , 
 n40478 , n330905 , n330906 , n40481 , n330908 , n330909 , n330910 , n40485 , n330912 , n330913 , 
 n40488 , n330915 , n330916 , n40491 , n330918 , n330919 , n330920 , n330921 , n330922 , n330923 , 
 n330924 , n330925 , n330926 , n330927 , n330928 , n330929 , n40504 , n330931 , n330932 , n40507 , 
 n330934 , n330935 , n40510 , n330937 , n330938 , n40513 , n330940 , n330941 , n40516 , n330943 , 
 n330944 , n40519 , n40520 , n330947 , n330948 , n330949 , n40524 , n330951 , n330952 , n40527 , 
 n330954 , n330955 , n40530 , n330957 , n330958 , n40533 , n330960 , n330961 , n40536 , n330963 , 
 n330964 , n330965 , n330966 , n330967 , n40542 , n330969 , n330970 , n40545 , n330972 , n330973 , 
 n40548 , n330975 , n330976 , n40551 , n40552 , n330979 , n40554 , n330981 , n40556 , n40557 , 
 n330984 , n330985 , n40560 , n330987 , n330988 , n330989 , n330990 , n330991 , n330992 , n330993 , 
 n330994 , n330995 , n330996 , n40571 , n330998 , n40573 , n40574 , n331001 , n331002 , n331003 , 
 n331004 , n331005 , n331006 , n331007 , n331008 , n331009 , n40584 , n331011 , n40586 , n331013 , 
 n331014 , n40589 , n331016 , n331017 , n40592 , n331019 , n331020 , n40595 , n40596 , n331023 , 
 n40598 , n331025 , n331026 , n331027 , n331028 , n40603 , n331030 , n331031 , n331032 , n40607 , 
 n331034 , n331035 , n331036 , n331037 , n331038 , n331039 , n40614 , n331041 , n331042 , n331043 , 
 n331044 , n331045 , n40620 , n331047 , n331048 , n40623 , n331050 , n331051 , n40626 , n40627 , 
 n40628 , n40629 , n331056 , n331057 , n40632 , n331059 , n40634 , n331061 , n331062 , n331063 , 
 n40638 , n331065 , n331066 , n331067 , n331068 , n331069 , n331070 , n331071 , n40646 , n331073 , 
 n40648 , n331075 , n331076 , n331077 , n331078 , n331079 , n331080 , n331081 , n331082 , n331083 , 
 n331084 , n40659 , n331086 , n331087 , n331088 , n331089 , n40664 , n331091 , n331092 , n331093 , 
 n331094 , n331095 , n40670 , n331097 , n331098 , n40673 , n331100 , n40675 , n331102 , n331103 , 
 n40678 , n331105 , n331106 , n40681 , n331108 , n331109 , n331110 , n331111 , n331112 , n40687 , 
 n331114 , n331115 , n40690 , n40691 , n40692 , n40693 , n331120 , n331121 , n331122 , n40697 , 
 n331124 , n331125 , n331126 , n40701 , n331128 , n331129 , n331130 , n331131 , n40706 , n331133 , 
 n331134 , n331135 , n331136 , n40711 , n40712 , n331139 , n331140 , n331141 , n40716 , n331143 , 
 n331144 , n40719 , n331146 , n40721 , n331148 , n331149 , n40724 , n40725 , n331152 , n40727 , 
 n331154 , n331155 , n40730 , n331157 , n331158 , n40733 , n40734 , n40735 , n40736 , n331163 , 
 n331164 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n331171 , n40746 , n331173 , 
 n331174 , n40749 , n40750 , n40751 , n331178 , n331179 , n331180 , n331181 , n40756 , n331183 , 
 n331184 , n331185 , n331186 , n331187 , n40762 , n331189 , n331190 , n331191 , n40766 , n331193 , 
 n331194 , n40769 , n331196 , n331197 , n40772 , n331199 , n331200 , n331201 , n331202 , n40777 , 
 n331204 , n331205 , n40780 , n331207 , n331208 , n331209 , n331210 , n331211 , n331212 , n331213 , 
 n331214 , n331215 , n331216 , n331217 , n331218 , n40793 , n331220 , n331221 , n331222 , n40797 , 
 n331224 , n331225 , n331226 , n331227 , n331228 , n331229 , n331230 , n331231 , n331232 , n331233 , 
 n331234 , n40809 , n40810 , n331237 , n40812 , n40813 , n331240 , n40815 , n331242 , n40817 , 
 n40818 , n331245 , n331246 , n331247 , n331248 , n331249 , n331250 , n331251 , n40826 , n331253 , 
 n331254 , n331255 , n331256 , n40831 , n331258 , n331259 , n331260 , n40835 , n331262 , n331263 , 
 n40838 , n40839 , n331266 , n331267 , n331268 , n331269 , n331270 , n331271 , n331272 , n331273 , 
 n40848 , n331275 , n331276 , n40851 , n331278 , n331279 , n40854 , n331281 , n331282 , n331283 , 
 n40858 , n40859 , n40860 , n40861 , n40862 , n331289 , n331290 , n331291 , n331292 , n331293 , 
 n331294 , n331295 , n331296 , n331297 , n331298 , n331299 , n331300 , n331301 , n331302 , n331303 , 
 n40878 , n331305 , n331306 , n40881 , n331308 , n331309 , n331310 , n331311 , n331312 , n331313 , 
 n331314 , n331315 , n331316 , n331317 , n331318 , n40893 , n40894 , n331321 , n40896 , n40897 , 
 n40898 , n40899 , n331326 , n331327 , n331328 , n331329 , n331330 , n331331 , n40906 , n331333 , 
 n331334 , n331335 , n40910 , n331337 , n331338 , n40913 , n40914 , n40915 , n331342 , n331343 , 
 n331344 , n331345 , n331346 , n331347 , n331348 , n331349 , n331350 , n331351 , n331352 , n40927 , 
 n331354 , n331355 , n40930 , n331357 , n331358 , n40933 , n331360 , n331361 , n331362 , n331363 , 
 n331364 , n331365 , n331366 , n40941 , n40942 , n331369 , n40944 , n331371 , n331372 , n40947 , 
 n40948 , n40949 , n40950 , n331377 , n331378 , n40953 , n331380 , n331381 , n40956 , n331383 , 
 n40958 , n331385 , n331386 , n331387 , n331388 , n331389 , n331390 , n331391 , n40966 , n331393 , 
 n331394 , n40969 , n331396 , n331397 , n331398 , n331399 , n331400 , n331401 , n331402 , n331403 , 
 n331404 , n331405 , n331406 , n40981 , n331408 , n331409 , n40984 , n331411 , n331412 , n40987 , 
 n331414 , n40989 , n40990 , n331417 , n331418 , n331419 , n331420 , n331421 , n331422 , n40997 , 
 n331424 , n331425 , n331426 , n331427 , n331428 , n331429 , n41004 , n331431 , n331432 , n331433 , 
 n331434 , n331435 , n331436 , n41011 , n331438 , n331439 , n41014 , n41015 , n331442 , n41017 , 
 n41018 , n331445 , n331446 , n41021 , n331448 , n331449 , n331450 , n331451 , n41026 , n331453 , 
 n331454 , n331455 , n331456 , n331457 , n41032 , n331459 , n331460 , n331461 , n331462 , n331463 , 
 n41038 , n331465 , n331466 , n41041 , n331468 , n331469 , n331470 , n331471 , n331472 , n331473 , 
 n331474 , n41049 , n331476 , n331477 , n41052 , n331479 , n331480 , n331481 , n331482 , n331483 , 
 n331484 , n331485 , n41060 , n331487 , n331488 , n331489 , n331490 , n331491 , n41066 , n331493 , 
 n331494 , n331495 , n331496 , n331497 , n331498 , n331499 , n331500 , n331501 , n331502 , n331503 , 
 n331504 , n331505 , n331506 , n331507 , n331508 , n41083 , n331510 , n331511 , n41086 , n41087 , 
 n41088 , n41089 , n331516 , n41091 , n41092 , n41093 , n41094 , n331521 , n331522 , n331523 , 
 n331524 , n331525 , n331526 , n331527 , n41102 , n331529 , n331530 , n331531 , n331532 , n41107 , 
 n41108 , n331535 , n331536 , n331537 , n41112 , n331539 , n331540 , n331541 , n331542 , n41117 , 
 n331544 , n331545 , n41120 , n331547 , n331548 , n41123 , n41124 , n331551 , n41126 , n41127 , 
 n331554 , n41129 , n331556 , n331557 , n41132 , n331559 , n41134 , n331561 , n331562 , n41137 , 
 n41138 , n41139 , n331566 , n331567 , n331568 , n331569 , n41144 , n331571 , n331572 , n331573 , 
 n331574 , n331575 , n331576 , n331577 , n331578 , n41153 , n331580 , n331581 , n331582 , n41157 , 
 n331584 , n41159 , n331586 , n331587 , n331588 , n331589 , n331590 , n331591 , n331592 , n331593 , 
 n331594 , n41169 , n41170 , n41171 , n41172 , n331599 , n331600 , n41175 , n331602 , n331603 , 
 n331604 , n331605 , n331606 , n331607 , n331608 , n331609 , n41184 , n331611 , n331612 , n41187 , 
 n41188 , n41189 , n41190 , n331617 , n331618 , n331619 , n41194 , n331621 , n331622 , n331623 , 
 n331624 , n331625 , n331626 , n331627 , n331628 , n41203 , n331630 , n331631 , n41206 , n331633 , 
 n41208 , n41209 , n331636 , n331637 , n331638 , n41213 , n331640 , n331641 , n41216 , n331643 , 
 n41218 , n331645 , n331646 , n331647 , n331648 , n331649 , n41224 , n331651 , n331652 , n331653 , 
 n41228 , n331655 , n331656 , n331657 , n331658 , n41233 , n331660 , n331661 , n331662 , n41237 , 
 n331664 , n331665 , n331666 , n331667 , n331668 , n331669 , n331670 , n331671 , n331672 , n331673 , 
 n331674 , n331675 , n331676 , n41251 , n331678 , n41253 , n41254 , n331681 , n331682 , n331683 , 
 n331684 , n331685 , n331686 , n331687 , n331688 , n331689 , n331690 , n331691 , n331692 , n331693 , 
 n331694 , n331695 , n331696 , n331697 , n331698 , n331699 , n331700 , n331701 , n331702 , n331703 , 
 n41278 , n41279 , n41280 , n41281 , n331708 , n331709 , n41284 , n331711 , n41286 , n331713 , 
 n331714 , n331715 , n41290 , n331717 , n331718 , n331719 , n331720 , n331721 , n331722 , n331723 , 
 n41298 , n41299 , n331726 , n331727 , n331728 , n331729 , n331730 , n331731 , n331732 , n331733 , 
 n331734 , n331735 , n331736 , n41311 , n331738 , n41313 , n331740 , n331741 , n331742 , n41317 , 
 n331744 , n331745 , n331746 , n331747 , n331748 , n331749 , n41324 , n331751 , n331752 , n331753 , 
 n331754 , n331755 , n331756 , n331757 , n331758 , n331759 , n331760 , n331761 , n331762 , n331763 , 
 n331764 , n331765 , n331766 , n331767 , n331768 , n331769 , n331770 , n41345 , n331772 , n41347 , 
 n331774 , n331775 , n331776 , n331777 , n331778 , n41353 , n331780 , n331781 , n331782 , n331783 , 
 n41358 , n41359 , n41360 , n331787 , n41362 , n331789 , n41364 , n331791 , n331792 , n331793 , 
 n41368 , n331795 , n331796 , n331797 , n41372 , n331799 , n41374 , n331801 , n331802 , n331803 , 
 n331804 , n331805 , n331806 , n331807 , n41382 , n331809 , n331810 , n331811 , n41386 , n331813 , 
 n41388 , n331815 , n331816 , n331817 , n41392 , n331819 , n331820 , n331821 , n331822 , n331823 , 
 n331824 , n41399 , n331826 , n331827 , n331828 , n331829 , n331830 , n331831 , n41406 , n331833 , 
 n331834 , n41409 , n331836 , n41411 , n41412 , n331839 , n41414 , n331841 , n331842 , n331843 , 
 n41418 , n41419 , n41420 , n331847 , n331848 , n41423 , n331850 , n331851 , n331852 , n331853 , 
 n331854 , n331855 , n41430 , n331857 , n331858 , n41433 , n331860 , n331861 , n41436 , n331863 , 
 n331864 , n41439 , n331866 , n331867 , n331868 , n331869 , n331870 , n331871 , n331872 , n331873 , 
 n331874 , n41449 , n331876 , n331877 , n331878 , n331879 , n331880 , n41455 , n41456 , n331883 , 
 n41458 , n41459 , n331886 , n331887 , n331888 , n41463 , n41464 , n41465 , n41466 , n41467 , 
 n331894 , n41469 , n331896 , n41471 , n331898 , n331899 , n331900 , n331901 , n331902 , n331903 , 
 n41478 , n331905 , n331906 , n331907 , n41482 , n331909 , n331910 , n41485 , n331912 , n331913 , 
 n331914 , n331915 , n41490 , n331917 , n331918 , n41493 , n41494 , n331921 , n331922 , n41497 , 
 n331924 , n41499 , n331926 , n331927 , n331928 , n41503 , n331930 , n331931 , n331932 , n331933 , 
 n331934 , n331935 , n331936 , n41511 , n331938 , n331939 , n331940 , n331941 , n331942 , n331943 , 
 n331944 , n331945 , n331946 , n41521 , n331948 , n41523 , n331950 , n41525 , n331952 , n331953 , 
 n41528 , n331955 , n331956 , n41531 , n331958 , n331959 , n41534 , n41535 , n331962 , n331963 , 
 n331964 , n331965 , n331966 , n331967 , n331968 , n331969 , n331970 , n331971 , n331972 , n331973 , 
 n331974 , n331975 , n331976 , n41551 , n41552 , n41553 , n331980 , n331981 , n331982 , n331983 , 
 n331984 , n331985 , n331986 , n331987 , n331988 , n41563 , n41564 , n331991 , n331992 , n41567 , 
 n331994 , n331995 , n331996 , n331997 , n331998 , n331999 , n41574 , n332001 , n332002 , n41577 , 
 n41578 , n332005 , n332006 , n41581 , n332008 , n332009 , n332010 , n332011 , n332012 , n41587 , 
 n332014 , n41589 , n41590 , n332017 , n332018 , n41593 , n332020 , n41595 , n41596 , n332023 , 
 n41598 , n41599 , n41600 , n332027 , n332028 , n332029 , n332030 , n41605 , n332032 , n332033 , 
 n332034 , n332035 , n332036 , n332037 , n332038 , n332039 , n332040 , n332041 , n332042 , n41617 , 
 n332044 , n332045 , n332046 , n332047 , n332048 , n332049 , n332050 , n332051 , n41626 , n332053 , 
 n332054 , n41629 , n332056 , n41631 , n332058 , n332059 , n41634 , n332061 , n332062 , n41637 , 
 n332064 , n332065 , n332066 , n332067 , n41642 , n332069 , n332070 , n332071 , n332072 , n332073 , 
 n332074 , n332075 , n332076 , n332077 , n332078 , n332079 , n332080 , n332081 , n41656 , n332083 , 
 n332084 , n41659 , n332086 , n332087 , n41662 , n332089 , n332090 , n332091 , n332092 , n41667 , 
 n332094 , n332095 , n41670 , n41671 , n41672 , n41673 , n332100 , n332101 , n41676 , n332103 , 
 n332104 , n332105 , n41680 , n332107 , n332108 , n332109 , n41684 , n332111 , n332112 , n332113 , 
 n332114 , n41689 , n332116 , n332117 , n41692 , n332119 , n332120 , n41695 , n332122 , n41697 , 
 n41698 , n332125 , n332126 , n41701 , n332128 , n332129 , n41704 , n332131 , n332132 , n41707 , 
 n41708 , n41709 , n332136 , n332137 , n332138 , n332139 , n332140 , n332141 , n332142 , n41717 , 
 n332144 , n332145 , n332146 , n332147 , n332148 , n332149 , n332150 , n41725 , n332152 , n332153 , 
 n332154 , n332155 , n332156 , n41731 , n41732 , n332159 , n332160 , n332161 , n332162 , n41737 , 
 n41738 , n41739 , n41740 , n41741 , n332168 , n332169 , n332170 , n332171 , n41746 , n332173 , 
 n332174 , n332175 , n332176 , n332177 , n332178 , n41753 , n332180 , n41755 , n41756 , n332183 , 
 n41758 , n332185 , n332186 , n332187 , n332188 , n41763 , n332190 , n332191 , n332192 , n332193 , 
 n41768 , n332195 , n332196 , n41771 , n332198 , n332199 , n41774 , n41775 , n332202 , n332203 , 
 n332204 , n332205 , n332206 , n332207 , n332208 , n332209 , n332210 , n332211 , n41786 , n41787 , 
 n41788 , n332215 , n332216 , n332217 , n332218 , n332219 , n332220 , n332221 , n332222 , n332223 , 
 n332224 , n41799 , n332226 , n41801 , n41802 , n332229 , n41804 , n332231 , n332232 , n332233 , 
 n332234 , n332235 , n332236 , n332237 , n332238 , n332239 , n332240 , n332241 , n332242 , n332243 , 
 n332244 , n332245 , n332246 , n332247 , n332248 , n332249 , n332250 , n41825 , n332252 , n332253 , 
 n332254 , n332255 , n41830 , n41831 , n332258 , n41833 , n332260 , n41835 , n41836 , n332263 , 
 n332264 , n332265 , n332266 , n41841 , n332268 , n332269 , n41844 , n41845 , n332272 , n332273 , 
 n332274 , n41849 , n332276 , n332277 , n332278 , n332279 , n41854 , n332281 , n332282 , n41857 , 
 n332284 , n332285 , n332286 , n332287 , n332288 , n41863 , n332290 , n332291 , n41866 , n332293 , 
 n332294 , n332295 , n332296 , n332297 , n332298 , n332299 , n332300 , n332301 , n332302 , n332303 , 
 n332304 , n332305 , n41880 , n41881 , n41882 , n332309 , n41884 , n332311 , n41886 , n41887 , 
 n41888 , n332315 , n332316 , n332317 , n332318 , n41893 , n332320 , n332321 , n332322 , n332323 , 
 n41898 , n332325 , n332326 , n41901 , n332328 , n41903 , n41904 , n332331 , n332332 , n332333 , 
 n332334 , n41909 , n332336 , n332337 , n332338 , n332339 , n332340 , n332341 , n332342 , n41917 , 
 n332344 , n332345 , n332346 , n332347 , n332348 , n332349 , n332350 , n41925 , n332352 , n332353 , 
 n41928 , n332355 , n332356 , n41931 , n332358 , n41933 , n332360 , n332361 , n41936 , n41937 , 
 n41938 , n41939 , n332366 , n332367 , n332368 , n41943 , n332370 , n332371 , n332372 , n41947 , 
 n332374 , n332375 , n332376 , n41951 , n332378 , n41953 , n332380 , n332381 , n332382 , n332383 , 
 n41958 , n332385 , n332386 , n41961 , n332388 , n332389 , n332390 , n332391 , n41966 , n41967 , 
 n41968 , n41969 , n41970 , n332397 , n41972 , n332399 , n332400 , n41975 , n41976 , n332403 , 
 n41978 , n332405 , n332406 , n41981 , n332408 , n332409 , n332410 , n332411 , n332412 , n332413 , 
 n332414 , n332415 , n332416 , n332417 , n41992 , n41993 , n41994 , n41995 , n332422 , n332423 , 
 n332424 , n332425 , n332426 , n332427 , n42002 , n332429 , n332430 , n42005 , n332432 , n332433 , 
 n332434 , n42009 , n332436 , n332437 , n42012 , n332439 , n42014 , n42015 , n332442 , n332443 , 
 n332444 , n332445 , n332446 , n332447 , n332448 , n332449 , n332450 , n332451 , n42026 , n332453 , 
 n332454 , n332455 , n42030 , n332457 , n332458 , n332459 , n332460 , n332461 , n42036 , n42037 , 
 n42038 , n332465 , n42040 , n42041 , n332468 , n332469 , n332470 , n332471 , n332472 , n42047 , 
 n332474 , n332475 , n332476 , n42051 , n332478 , n332479 , n332480 , n42055 , n332482 , n332483 , 
 n332484 , n42059 , n332486 , n332487 , n332488 , n42063 , n332490 , n332491 , n332492 , n332493 , 
 n42068 , n332495 , n332496 , n332497 , n42072 , n332499 , n332500 , n332501 , n42076 , n332503 , 
 n332504 , n42079 , n332506 , n332507 , n332508 , n42083 , n332510 , n332511 , n42086 , n332513 , 
 n332514 , n42089 , n42090 , n42091 , n42092 , n332519 , n332520 , n42095 , n332522 , n332523 , 
 n332524 , n42099 , n332526 , n332527 , n332528 , n42103 , n332530 , n332531 , n332532 , n332533 , 
 n42108 , n332535 , n332536 , n332537 , n42112 , n332539 , n332540 , n332541 , n332542 , n42117 , 
 n332544 , n332545 , n332546 , n332547 , n42122 , n332549 , n42124 , n332551 , n332552 , n42127 , 
 n332554 , n332555 , n42130 , n42131 , n42132 , n42133 , n332560 , n332561 , n332562 , n42137 , 
 n332564 , n332565 , n42140 , n332567 , n332568 , n332569 , n332570 , n42145 , n332572 , n332573 , 
 n42148 , n332575 , n332576 , n42151 , n332578 , n332579 , n332580 , n42155 , n332582 , n332583 , 
 n42158 , n332585 , n332586 , n332587 , n332588 , n42163 , n332590 , n332591 , n42166 , n42167 , 
 n42168 , n332595 , n42170 , n332597 , n42172 , n42173 , n332600 , n42175 , n332602 , n42177 , 
 n332604 , n42179 , n332606 , n332607 , n42182 , n42183 , n42184 , n42185 , n332612 , n332613 , 
 n332614 , n42189 , n332616 , n332617 , n332618 , n332619 , n332620 , n42195 , n42196 , n42197 , 
 n42198 , n42199 , n332626 , n332627 , n332628 , n42203 , n332630 , n332631 , n332632 , n42207 , 
 n332634 , n332635 , n332636 , n332637 , n42212 , n332639 , n332640 , n332641 , n332642 , n332643 , 
 n42218 , n332645 , n332646 , n42221 , n332648 , n332649 , n332650 , n42225 , n332652 , n332653 , 
 n42228 , n42229 , n42230 , n42231 , n332658 , n332659 , n332660 , n42235 , n332662 , n332663 , 
 n42238 , n332665 , n332666 , n332667 , n332668 , n332669 , n332670 , n42245 , n332672 , n332673 , 
 n42248 , n332675 , n332676 , n332677 , n332678 , n332679 , n42254 , n332681 , n332682 , n42257 , 
 n332684 , n42259 , n332686 , n42261 , n42262 , n332689 , n42264 , n332691 , n332692 , n42267 , 
 n332694 , n332695 , n42270 , n42271 , n42272 , n42273 , n332700 , n332701 , n42276 , n332703 , 
 n42278 , n332705 , n332706 , n332707 , n42282 , n332709 , n332710 , n332711 , n332712 , n332713 , 
 n332714 , n332715 , n332716 , n332717 , n42292 , n332719 , n332720 , n332721 , n332722 , n42297 , 
 n42298 , n42299 , n332726 , n42301 , n332728 , n42303 , n42304 , n42305 , n42306 , n332733 , 
 n42308 , n42309 , n42310 , n332737 , n332738 , n332739 , n332740 , n332741 , n332742 , n332743 , 
 n42318 , n332745 , n42320 , n332747 , n332748 , n332749 , n42324 , n332751 , n332752 , n332753 , 
 n332754 , n332755 , n332756 , n332757 , n332758 , n42333 , n42334 , n332761 , n332762 , n42337 , 
 n332764 , n42339 , n332766 , n332767 , n332768 , n332769 , n332770 , n42345 , n42346 , n42347 , 
 n332774 , n332775 , n332776 , n332777 , n42352 , n332779 , n332780 , n332781 , n332782 , n332783 , 
 n332784 , n332785 , n42360 , n42361 , n332788 , n332789 , n42364 , n42365 , n42366 , n332793 , 
 n332794 , n332795 , n332796 , n332797 , n42372 , n332799 , n332800 , n332801 , n332802 , n332803 , 
 n42378 , n332805 , n42380 , n332807 , n42382 , n332809 , n332810 , n42385 , n332812 , n332813 , 
 n42388 , n332815 , n332816 , n332817 , n42392 , n332819 , n42394 , n332821 , n332822 , n332823 , 
 n42398 , n332825 , n42400 , n332827 , n332828 , n332829 , n332830 , n42405 , n332832 , n42407 , 
 n42408 , n42409 , n332836 , n42411 , n42412 , n332839 , n332840 , n332841 , n332842 , n332843 , 
 n332844 , n332845 , n332846 , n332847 , n332848 , n332849 , n332850 , n42425 , n332852 , n332853 , 
 n42428 , n42429 , n332856 , n332857 , n332858 , n332859 , n332860 , n332861 , n332862 , n42437 , 
 n42438 , n42439 , n332866 , n332867 , n332868 , n332869 , n42444 , n42445 , n42446 , n42447 , 
 n332874 , n332875 , n332876 , n42451 , n332878 , n332879 , n332880 , n332881 , n42456 , n332883 , 
 n332884 , n332885 , n332886 , n42461 , n42462 , n42463 , n42464 , n42465 , n332892 , n332893 , 
 n332894 , n42469 , n332896 , n332897 , n332898 , n332899 , n332900 , n332901 , n332902 , n332903 , 
 n332904 , n332905 , n332906 , n332907 , n332908 , n42483 , n332910 , n332911 , n332912 , n332913 , 
 n332914 , n332915 , n42490 , n332917 , n332918 , n332919 , n332920 , n42495 , n332922 , n42497 , 
 n332924 , n332925 , n332926 , n332927 , n332928 , n42503 , n332930 , n332931 , n332932 , n332933 , 
 n42508 , n42509 , n332936 , n332937 , n332938 , n332939 , n42514 , n332941 , n332942 , n42517 , 
 n42518 , n332945 , n332946 , n332947 , n332948 , n42523 , n332950 , n332951 , n332952 , n332953 , 
 n42528 , n332955 , n332956 , n42531 , n332958 , n332959 , n332960 , n332961 , n332962 , n332963 , 
 n332964 , n332965 , n42540 , n42541 , n332968 , n332969 , n42544 , n332971 , n332972 , n332973 , 
 n332974 , n42549 , n42550 , n332977 , n42552 , n42553 , n332980 , n332981 , n42556 , n332983 , 
 n42558 , n332985 , n332986 , n332987 , n332988 , n42563 , n332990 , n332991 , n332992 , n332993 , 
 n332994 , n332995 , n42570 , n332997 , n332998 , n332999 , n333000 , n42575 , n42576 , n42577 , 
 n333004 , n333005 , n333006 , n333007 , n333008 , n42583 , n333010 , n333011 , n42586 , n333013 , 
 n333014 , n42589 , n333016 , n42591 , n333018 , n333019 , n333020 , n333021 , n42596 , n42597 , 
 n333024 , n333025 , n333026 , n42601 , n42602 , n333029 , n333030 , n42605 , n333032 , n333033 , 
 n333034 , n333035 , n333036 , n333037 , n333038 , n333039 , n333040 , n333041 , n42616 , n333043 , 
 n333044 , n42619 , n42620 , n333047 , n42622 , n333049 , n333050 , n333051 , n333052 , n333053 , 
 n333054 , n42629 , n333056 , n333057 , n333058 , n42633 , n333060 , n333061 , n333062 , n333063 , 
 n42638 , n42639 , n333066 , n42641 , n42642 , n333069 , n42644 , n333071 , n42646 , n333073 , 
 n42648 , n42649 , n333076 , n42651 , n333078 , n333079 , n333080 , n42655 , n42656 , n333083 , 
 n333084 , n333085 , n42660 , n42661 , n333088 , n333089 , n42664 , n333091 , n333092 , n333093 , 
 n42668 , n333095 , n333096 , n333097 , n42672 , n333099 , n333100 , n333101 , n42676 , n333103 , 
 n42678 , n333105 , n333106 , n42681 , n333108 , n333109 , n333110 , n42685 , n333112 , n333113 , 
 n333114 , n42689 , n42690 , n333117 , n333118 , n333119 , n42694 , n333121 , n42696 , n333123 , 
 n333124 , n42699 , n333126 , n333127 , n333128 , n42703 , n42704 , n42705 , n42706 , n42707 , 
 n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n333140 , n42715 , n42716 , n333143 , 
 n42718 , n42719 , n42720 , n42721 , n333148 , n333149 , n333150 , n42725 , n333152 , n42727 , 
 n42728 , n333155 , n42730 , n42731 , n42732 , n42733 , n333160 , n333161 , n333162 , n42737 , 
 n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , 
 n333174 , n42749 , n42750 , n333177 , n42752 , n42753 , n42754 , n42755 , n333182 , n333183 , 
 n333184 , n333185 , n42760 , n42761 , n333188 , n42763 , n42764 , n42765 , n42766 , n333193 , 
 n333194 , n333195 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , 
 n333204 , n42779 , n42780 , n333207 , n42782 , n42783 , n42784 , n42785 , n333212 , n333213 , 
 n333214 , n333215 , n42790 , n42791 , n333218 , n42793 , n42794 , n42795 , n42796 , n333223 , 
 n333224 , n333225 , n333226 , n42801 , n42802 , n333229 , n42804 , n42805 , n42806 , n42807 , 
 n333234 , n333235 , n333236 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , 
 n42818 , n42819 , n42820 , n42821 , n42822 , n333249 , n42824 , n42825 , n333252 , n42827 , 
 n42828 , n42829 , n42830 , n333257 , n333258 , n333259 , n42834 , n333261 , n42836 , n42837 , 
 n333264 , n42839 , n42840 , n42841 , n42842 , n333269 , n333270 , n333271 , n333272 , n42847 , 
 n42848 , n333275 , n42850 , n42851 , n42852 , n42853 , n333280 , n333281 , n333282 , n333283 , 
 n42858 , n42859 , n333286 , n42861 , n42862 , n42863 , n42864 , n333291 , n333292 , n42867 , 
 n333294 , n42869 , n333296 , n42871 , n333298 , n333299 , n333300 , n42875 , n333302 , n42877 , 
 n333304 , n333305 , n333306 , n42881 , n333308 , n42883 , n333310 , n333311 , n333312 , n42887 , 
 n333314 , n42889 , n333316 , n333317 , n333318 , n42893 , n333320 , n42895 , n333322 , n333323 , 
 n333324 , n42899 , n333326 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , 
 n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , 
 n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , 
 n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , 
 n42938 , n333365 , n42940 , n333367 , n42942 , n333369 , n333370 , n333371 , n42946 , n333373 , 
 n333374 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , 
 n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , 
 n42968 , n333395 , n42970 , n333397 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , 
 n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , 
 n42988 , n42989 , n42990 , n42991 , n333418 , n42993 , n333420 , n42995 , n42996 , n42997 , 
 n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , 
 n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , 
 n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , 
 n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , 
 n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , 
 n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , 
 n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , 
 n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , 
 n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n333510 , n333511 , n333512 , n43087 , 
 n43088 , n333515 , n43090 , n43091 , n43092 , n43093 , n333520 , n333521 , n333522 , n333523 , 
 n43098 , n43099 , n333526 , n43101 , n43102 , n43103 , n43104 , n333531 , n333532 , n333533 , 
 n333534 , n333535 , n43110 , n333537 , n43112 , n43113 , n43114 , n43115 , n333542 , n333543 , 
 n333544 , n43119 , n333546 , n43121 , n43122 , n333549 , n43124 , n43125 , n43126 , n43127 , 
 n333554 , n333555 , n333556 , n333557 , n43132 , n43133 , n333560 , n43135 , n43136 , n43137 , 
 n43138 , n333565 , n333566 , n333567 , n333568 , n43143 , n43144 , n333571 , n43146 , n333573 , 
 n43148 , n43149 , n333576 , n333577 , n333578 , n333579 , n43154 , n43155 , n333582 , n43157 , 
 n43158 , n43159 , n43160 , n333587 , n333588 , n333589 , n333590 , n43165 , n43166 , n333593 , 
 n43168 , n43169 , n43170 , n43171 , n333598 , n333599 , n333600 , n333601 , n43176 , n43177 , 
 n333604 , n43179 , n43180 , n43181 , n43182 , n333609 , n333610 , n333611 , n333612 , n43187 , 
 n43188 , n333615 , n43190 , n43191 , n43192 , n43193 , n333620 , n333621 , n333622 , n333623 , 
 n43198 , n43199 , n333626 , n43201 , n43202 , n43203 , n43204 , n333631 , n333632 , n333633 , 
 n333634 , n43209 , n43210 , n333637 , n43212 , n43213 , n43214 , n43215 , n333642 , n333643 , 
 n333644 , n333645 , n43220 , n43221 , n333648 , n43223 , n43224 , n43225 , n43226 , n333653 , 
 n333654 , n333655 , n333656 , n43231 , n43232 , n333659 , n43234 , n43235 , n43236 , n43237 , 
 n333664 , n333665 , n333666 , n333667 , n43242 , n43243 , n333670 , n43245 , n43246 , n43247 , 
 n43248 , n333675 , n333676 , n43251 , n333678 , n333679 , n43254 , n43255 , n333682 , n43257 , 
 n43258 , n43259 , n43260 , n333687 , n333688 , n333689 , n333690 , n43265 , n43266 , n333693 , 
 n43268 , n43269 , n43270 , n43271 , n333698 , n333699 , n43274 , n333701 , n333702 , n43277 , 
 n43278 , n333705 , n43280 , n43281 , n43282 , n43283 , n333710 , n333711 , n43286 , n333713 , 
 n333714 , n43289 , n43290 , n333717 , n43292 , n43293 , n43294 , n43295 , n333722 , n333723 , 
 n43298 , n43299 , n333726 , n333727 , n43302 , n43303 , n333730 , n43305 , n43306 , n43307 , 
 n43308 , n333735 , n43310 , n333737 , n43312 , n333739 , n333740 , n43315 , n43316 , n333743 , 
 n43318 , n43319 , n43320 , n43321 , n333748 , n43323 , n333750 , n333751 , n333752 , n43327 , 
 n43328 , n333755 , n43330 , n43331 , n43332 , n43333 , n333760 , n333761 , n43336 , n333763 , 
 n333764 , n43339 , n43340 , n333767 , n43342 , n43343 , n43344 , n43345 , n333772 , n333773 , 
 n333774 , n333775 , n43350 , n43351 , n333778 , n43353 , n333780 , n43355 , n43356 , n333783 , 
 n333784 , n43359 , n333786 , n333787 , n333788 , n43363 , n333790 , n333791 , n43366 , n333793 , 
 n43368 , n333795 , n333796 , n333797 , n333798 , n43373 , n43374 , n333801 , n43376 , n43377 , 
 n43378 , n43379 , n333806 , n333807 , n333808 , n333809 , n43384 , n43385 , n333812 , n43387 , 
 n43388 , n333815 , n43390 , n333817 , n43392 , n43393 , n333820 , n333821 , n43396 , n43397 , 
 n333824 , n43399 , n43400 , n43401 , n43402 , n333829 , n333830 , n333831 , n333832 , n43407 , 
 n43408 , n333835 , n43410 , n43411 , n43412 , n43413 , n333840 , n333841 , n43416 , n333843 , 
 n333844 , n333845 , n333846 , n43421 , n43422 , n43423 , n43424 , n333851 , n333852 , n333853 , 
 n333854 , n43429 , n43430 , n333857 , n43432 , n43433 , n43434 , n43435 , n333862 , n333863 , 
 n333864 , n43439 , n333866 , n333867 , n333868 , n333869 , n333870 , n43445 , n333872 , n43447 , 
 n333874 , n333875 , n333876 , n333877 , n333878 , n333879 , n333880 , n333881 , n333882 , n333883 , 
 n333884 , n43459 , n333886 , n333887 , n333888 , n43463 , n333890 , n333891 , n333892 , n333893 , 
 n333894 , n43469 , n333896 , n333897 , n43472 , n333899 , n333900 , n333901 , n333902 , n333903 , 
 n43478 , n333905 , n333906 , n43481 , n333908 , n333909 , n43484 , n333911 , n43486 , n333913 , 
 n333914 , n333915 , n43490 , n333917 , n43492 , n333919 , n333920 , n43495 , n43496 , n43497 , 
 n43498 , n333925 , n333926 , n333927 , n333928 , n333929 , n333930 , n43505 , n333932 , n333933 , 
 n333934 , n333935 , n333936 , n333937 , n333938 , n43513 , n333940 , n333941 , n43516 , n43517 , 
 n333944 , n43519 , n333946 , n333947 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , 
 n333954 , n43529 , n333956 , n43531 , n43532 , n43533 , n333960 , n43535 , n333962 , n333963 , 
 n333964 , n43539 , n333966 , n43541 , n333968 , n43543 , n333970 , n43545 , n333972 , n333973 , 
 n43548 , n333975 , n333976 , n333977 , n43552 , n43553 , n43554 , n43555 , n333982 , n333983 , 
 n43558 , n333985 , n333986 , n43561 , n333988 , n333989 , n333990 , n333991 , n333992 , n333993 , 
 n333994 , n333995 , n333996 , n333997 , n333998 , n333999 , n334000 , n334001 , n334002 , n43577 , 
 n334004 , n334005 , n43580 , n334007 , n334008 , n334009 , n334010 , n334011 , n334012 , n334013 , 
 n334014 , n334015 , n334016 , n43591 , n43592 , n334019 , n43594 , n43595 , n334022 , n334023 , 
 n334024 , n334025 , n43600 , n334027 , n43602 , n43603 , n43604 , n334031 , n334032 , n43607 , 
 n43608 , n43609 , n334036 , n43611 , n334038 , n43613 , n334040 , n334041 , n334042 , n43617 , 
 n334044 , n334045 , n43620 , n334047 , n334048 , n43623 , n334050 , n334051 , n334052 , n334053 , 
 n43628 , n334055 , n334056 , n334057 , n334058 , n334059 , n334060 , n334061 , n334062 , n334063 , 
 n334064 , n334065 , n334066 , n43641 , n334068 , n334069 , n43644 , n334071 , n334072 , n43647 , 
 n334074 , n334075 , n334076 , n334077 , n334078 , n334079 , n43654 , n334081 , n43656 , n43657 , 
 n43658 , n334085 , n334086 , n43661 , n334088 , n334089 , n43664 , n334091 , n43666 , n334093 , 
 n334094 , n334095 , n334096 , n334097 , n334098 , n43673 , n334100 , n334101 , n43676 , n334103 , 
 n334104 , n43679 , n334106 , n334107 , n43682 , n334109 , n334110 , n334111 , n334112 , n43687 , 
 n334114 , n334115 , n43690 , n334117 , n334118 , n334119 , n334120 , n334121 , n334122 , n43697 , 
 n334124 , n334125 , n43700 , n334127 , n334128 , n43703 , n43704 , n334131 , n43706 , n334133 , 
 n334134 , n43709 , n334136 , n334137 , n334138 , n334139 , n43714 , n43715 , n334142 , n334143 , 
 n334144 , n334145 , n334146 , n334147 , n334148 , n334149 , n334150 , n334151 , n334152 , n334153 , 
 n43728 , n334155 , n334156 , n334157 , n334158 , n334159 , n334160 , n334161 , n334162 , n334163 , 
 n334164 , n334165 , n334166 , n43741 , n334168 , n334169 , n334170 , n43745 , n334172 , n334173 , 
 n334174 , n334175 , n334176 , n334177 , n334178 , n334179 , n334180 , n43755 , n334182 , n334183 , 
 n43758 , n334185 , n334186 , n334187 , n43762 , n334189 , n334190 , n43765 , n334192 , n334193 , 
 n43768 , n334195 , n334196 , n334197 , n43772 , n334199 , n334200 , n334201 , n334202 , n334203 , 
 n334204 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n334213 , 
 n43788 , n334215 , n334216 , n334217 , n334218 , n334219 , n334220 , n43795 , n43796 , n43797 , 
 n334224 , n43799 , n334226 , n43801 , n334228 , n43803 , n334230 , n334231 , n334232 , n334233 , 
 n43808 , n334235 , n334236 , n334237 , n43812 , n334239 , n334240 , n334241 , n334242 , n334243 , 
 n334244 , n334245 , n334246 , n334247 , n334248 , n334249 , n334250 , n334251 , n334252 , n334253 , 
 n334254 , n43829 , n334256 , n334257 , n334258 , n334259 , n334260 , n334261 , n334262 , n334263 , 
 n334264 , n334265 , n334266 , n334267 , n334268 , n334269 , n334270 , n334271 , n334272 , n334273 , 
 n334274 , n43849 , n334276 , n43851 , n43852 , n43853 , n43854 , n334281 , n43856 , n43857 , 
 n334284 , n43859 , n334286 , n334287 , n43862 , n334289 , n334290 , n334291 , n334292 , n334293 , 
 n334294 , n334295 , n43870 , n334297 , n334298 , n334299 , n334300 , n43875 , n334302 , n334303 , 
 n334304 , n334305 , n334306 , n43881 , n334308 , n334309 , n43884 , n334311 , n334312 , n334313 , 
 n334314 , n334315 , n334316 , n43891 , n43892 , n334319 , n334320 , n334321 , n334322 , n334323 , 
 n334324 , n334325 , n334326 , n334327 , n334328 , n43903 , n334330 , n43905 , n334332 , n334333 , 
 n334334 , n334335 , n334336 , n334337 , n334338 , n334339 , n334340 , n334341 , n334342 , n334343 , 
 n334344 , n334345 , n43920 , n43921 , n334348 , n43923 , n334350 , n334351 , n334352 , n334353 , 
 n334354 , n334355 , n334356 , n334357 , n334358 , n334359 , n334360 , n334361 , n334362 , n334363 , 
 n334364 , n334365 , n334366 , n334367 , n334368 , n334369 , n334370 , n43945 , n334372 , n334373 , 
 n43948 , n43949 , n334376 , n334377 , n43952 , n334379 , n334380 , n43955 , n334382 , n334383 , 
 n43958 , n334385 , n334386 , n43961 , n334388 , n334389 , n334390 , n43965 , n334392 , n43967 , 
 n43968 , n43969 , n334396 , n334397 , n43972 , n334399 , n43974 , n334401 , n334402 , n334403 , 
 n43978 , n334405 , n334406 , n43981 , n43982 , n43983 , n43984 , n43985 , n334412 , n334413 , 
 n334414 , n43989 , n334416 , n334417 , n334418 , n334419 , n43994 , n334421 , n334422 , n334423 , 
 n43998 , n334425 , n334426 , n44001 , n334428 , n44003 , n44004 , n334431 , n44006 , n334433 , 
 n334434 , n44009 , n334436 , n334437 , n334438 , n334439 , n44014 , n334441 , n334442 , n44017 , 
 n334444 , n334445 , n44020 , n44021 , n334448 , n44023 , n334450 , n334451 , n44026 , n334453 , 
 n334454 , n334455 , n334456 , n334457 , n44032 , n334459 , n334460 , n44035 , n334462 , n334463 , 
 n44038 , n44039 , n44040 , n334467 , n334468 , n44043 , n44044 , n44045 , n334472 , n334473 , 
 n44048 , n334475 , n44050 , n334477 , n334478 , n44053 , n44054 , n44055 , n334482 , n334483 , 
 n44058 , n44059 , n44060 , n334487 , n334488 , n334489 , n334490 , n334491 , n334492 , n44067 , 
 n334494 , n334495 , n44070 , n334497 , n334498 , n334499 , n44074 , n334501 , n334502 , n44077 , 
 n334504 , n334505 , n44080 , n334507 , n334508 , n334509 , n334510 , n44085 , n334512 , n334513 , 
 n44088 , n334515 , n334516 , n334517 , n44092 , n334519 , n334520 , n334521 , n334522 , n44097 , 
 n334524 , n334525 , n44100 , n334527 , n334528 , n44103 , n334530 , n334531 , n334532 , n44107 , 
 n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n334542 , n44117 , 
 n334544 , n334545 , n44120 , n44121 , n44122 , n334549 , n44124 , n334551 , n334552 , n334553 , 
 n334554 , n44129 , n334556 , n44131 , n334558 , n334559 , n44134 , n334561 , n334562 , n44137 , 
 n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , 
 n44148 , n44149 , n334576 , n44151 , n44152 , n44153 , n44154 , n334581 , n334582 , n334583 , 
 n334584 , n334585 , n44160 , n334587 , n334588 , n44163 , n44164 , n334591 , n44166 , n44167 , 
 n334594 , n44169 , n334596 , n334597 , n44172 , n334599 , n334600 , n334601 , n334602 , n44177 , 
 n44178 , n334605 , n334606 , n44181 , n334608 , n334609 , n44184 , n334611 , n334612 , n44187 , 
 n334614 , n44189 , n334616 , n334617 , n44192 , n44193 , n334620 , n334621 , n44196 , n334623 , 
 n334624 , n44199 , n334626 , n334627 , n44202 , n44203 , n334630 , n334631 , n44206 , n334633 , 
 n334634 , n44209 , n334636 , n334637 , n44212 , n334639 , n334640 , n44215 , n334642 , n334643 , 
 n334644 , n44219 , n334646 , n334647 , n44222 , n334649 , n334650 , n44225 , n334652 , n334653 , 
 n44228 , n334655 , n334656 , n44231 , n44232 , n44233 , n334660 , n44235 , n334662 , n334663 , 
 n334664 , n44239 , n334666 , n334667 , n334668 , n44243 , n334670 , n44245 , n334672 , n44247 , 
 n334674 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n334682 , n44257 , 
 n334684 , n334685 , n44260 , n44261 , n44262 , n334689 , n334690 , n44265 , n334692 , n334693 , 
 n44268 , n334695 , n334696 , n44271 , n334698 , n334699 , n44274 , n334701 , n334702 , n334703 , 
 n44278 , n44279 , n44280 , n44281 , n334708 , n334709 , n44284 , n334711 , n334712 , n44287 , 
 n334714 , n334715 , n44290 , n334717 , n334718 , n44293 , n334720 , n334721 , n44296 , n334723 , 
 n334724 , n44299 , n334726 , n44301 , n334728 , n334729 , n334730 , n44305 , n334732 , n334733 , 
 n44308 , n334735 , n334736 , n44311 , n334738 , n334739 , n44314 , n334741 , n334742 , n44317 , 
 n44318 , n334745 , n334746 , n44321 , n334748 , n334749 , n44324 , n334751 , n334752 , n44327 , 
 n334754 , n44329 , n44330 , n334757 , n44332 , n334759 , n44334 , n334761 , n334762 , n44337 , 
 n334764 , n334765 , n44340 , n334767 , n334768 , n44343 , n44344 , n334771 , n44346 , n334773 , 
 n44348 , n334775 , n334776 , n44351 , n334778 , n334779 , n334780 , n44355 , n44356 , n334783 , 
 n44358 , n334785 , n44360 , n334787 , n44362 , n44363 , n44364 , n334791 , n334792 , n44367 , 
 n334794 , n334795 , n44370 , n334797 , n334798 , n334799 , n44374 , n44375 , n334802 , n334803 , 
 n44378 , n334805 , n334806 , n44381 , n334808 , n334809 , n44384 , n334811 , n44386 , n334813 , 
 n334814 , n334815 , n334816 , n334817 , n334818 , n334819 , n334820 , n334821 , n334822 , n44397 , 
 n334824 , n334825 , n334826 , n334827 , n334828 , n44403 , n334830 , n334831 , n44406 , n334833 , 
 n334834 , n44409 , n334836 , n334837 , n44412 , n334839 , n334840 , n44415 , n44416 , n44417 , 
 n44418 , n44419 , n334846 , n44421 , n334848 , n334849 , n334850 , n334851 , n334852 , n334853 , 
 n44428 , n334855 , n334856 , n44431 , n334858 , n334859 , n44434 , n334861 , n334862 , n44437 , 
 n334864 , n334865 , n334866 , n44441 , n44442 , n334869 , n334870 , n334871 , n334872 , n44447 , 
 n44448 , n334875 , n334876 , n44451 , n44452 , n334879 , n334880 , n44455 , n44456 , n334883 , 
 n334884 , n334885 , n334886 , n334887 , n334888 , n334889 , n334890 , n44465 , n44466 , n44467 , 
 n44468 , n44469 , n334896 , n334897 , n334898 , n334899 , n334900 , n44475 , n334902 , n44477 , 
 n44478 , n44479 , n44480 , n334907 , n44482 , n334909 , n334910 , n44485 , n334912 , n334913 , 
 n334914 , n334915 , n44490 , n334917 , n44492 , n44493 , n44494 , n334921 , n334922 , n44497 , 
 n334924 , n334925 , n334926 , n334927 , n334928 , n334929 , n334930 , n334931 , n334932 , n334933 , 
 n334934 , n334935 , n334936 , n334937 , n44512 , n334939 , n334940 , n334941 , n334942 , n44517 , 
 n334944 , n44519 , n334946 , n334947 , n334948 , n44523 , n334950 , n334951 , n44526 , n44527 , 
 n334954 , n44529 , n334956 , n334957 , n334958 , n44533 , n334960 , n334961 , n44536 , n44537 , 
 n334964 , n44539 , n44540 , n334967 , n44542 , n334969 , n334970 , n44545 , n334972 , n334973 , 
 n334974 , n334975 , n44550 , n334977 , n334978 , n334979 , n334980 , n334981 , n334982 , n334983 , 
 n334984 , n44559 , n44560 , n44561 , n334988 , n44563 , n334990 , n334991 , n44566 , n334993 , 
 n334994 , n334995 , n334996 , n334997 , n334998 , n334999 , n335000 , n335001 , n335002 , n335003 , 
 n335004 , n44579 , n335006 , n335007 , n44582 , n335009 , n335010 , n44585 , n335012 , n335013 , 
 n44588 , n335015 , n335016 , n335017 , n44592 , n335019 , n335020 , n335021 , n44596 , n335023 , 
 n335024 , n335025 , n44600 , n335027 , n335028 , n44603 , n335030 , n335031 , n44606 , n335033 , 
 n335034 , n44609 , n335036 , n335037 , n44612 , n335039 , n335040 , n335041 , n335042 , n44617 , 
 n335044 , n335045 , n44620 , n335047 , n44622 , n335049 , n335050 , n335051 , n335052 , n335053 , 
 n335054 , n44629 , n335056 , n335057 , n44632 , n335059 , n335060 , n44635 , n335062 , n335063 , 
 n44638 , n335065 , n335066 , n44641 , n44642 , n335069 , n44644 , n335071 , n44646 , n335073 , 
 n335074 , n44649 , n335076 , n335077 , n335078 , n44653 , n335080 , n335081 , n44656 , n335083 , 
 n335084 , n44659 , n335086 , n335087 , n44662 , n44663 , n335090 , n44665 , n335092 , n44667 , 
 n335094 , n335095 , n44670 , n335097 , n335098 , n44673 , n44674 , n335101 , n335102 , n44677 , 
 n335104 , n335105 , n44680 , n335107 , n335108 , n44683 , n335110 , n44685 , n335112 , n44687 , 
 n335114 , n335115 , n44690 , n335117 , n335118 , n335119 , n44694 , n335121 , n335122 , n44697 , 
 n335124 , n335125 , n44700 , n335127 , n335128 , n44703 , n335130 , n335131 , n44706 , n44707 , 
 n335134 , n335135 , n44710 , n335137 , n335138 , n44713 , n335140 , n335141 , n44716 , n335143 , 
 n44718 , n335145 , n335146 , n44721 , n335148 , n44723 , n335150 , n44725 , n335152 , n335153 , 
 n335154 , n335155 , n44730 , n335157 , n335158 , n335159 , n335160 , n335161 , n335162 , n44737 , 
 n335164 , n335165 , n335166 , n335167 , n44742 , n335169 , n335170 , n335171 , n335172 , n335173 , 
 n44748 , n335175 , n335176 , n335177 , n335178 , n335179 , n44754 , n335181 , n44756 , n335183 , 
 n335184 , n335185 , n335186 , n335187 , n335188 , n44763 , n335190 , n335191 , n335192 , n44767 , 
 n335194 , n335195 , n335196 , n335197 , n335198 , n335199 , n335200 , n335201 , n335202 , n44777 , 
 n335204 , n335205 , n335206 , n44781 , n335208 , n44783 , n44784 , n44785 , n335212 , n44787 , 
 n335214 , n44789 , n335216 , n335217 , n335218 , n335219 , n335220 , n335221 , n44796 , n335223 , 
 n335224 , n335225 , n335226 , n335227 , n44802 , n335229 , n335230 , n335231 , n44806 , n44807 , 
 n44808 , n335235 , n335236 , n44811 , n335238 , n44813 , n44814 , n335241 , n335242 , n335243 , 
 n335244 , n335245 , n335246 , n335247 , n44822 , n335249 , n335250 , n335251 , n44826 , n44827 , 
 n335254 , n335255 , n335256 , n335257 , n335258 , n44833 , n335260 , n335261 , n335262 , n335263 , 
 n335264 , n335265 , n335266 , n335267 , n335268 , n335269 , n335270 , n335271 , n335272 , n335273 , 
 n335274 , n44849 , n335276 , n44851 , n335278 , n335279 , n44854 , n44855 , n335282 , n44857 , 
 n335284 , n335285 , n44860 , n44861 , n44862 , n44863 , n44864 , n335291 , n44866 , n44867 , 
 n335294 , n44869 , n44870 , n335297 , n335298 , n335299 , n335300 , n335301 , n335302 , n44877 , 
 n335304 , n335305 , n335306 , n335307 , n44882 , n44883 , n44884 , n44885 , n335312 , n44887 , 
 n335314 , n44889 , n335316 , n335317 , n335318 , n44893 , n335320 , n44895 , n44896 , n44897 , 
 n335324 , n335325 , n335326 , n335327 , n44902 , n335329 , n335330 , n335331 , n335332 , n335333 , 
 n335334 , n335335 , n335336 , n335337 , n335338 , n335339 , n335340 , n335341 , n335342 , n335343 , 
 n44918 , n335345 , n335346 , n335347 , n335348 , n335349 , n335350 , n335351 , n335352 , n335353 , 
 n335354 , n335355 , n335356 , n335357 , n335358 , n44933 , n335360 , n335361 , n335362 , n335363 , 
 n335364 , n44939 , n44940 , n335367 , n44942 , n335369 , n44944 , n335371 , n335372 , n335373 , 
 n335374 , n335375 , n335376 , n335377 , n44952 , n335379 , n335380 , n335381 , n335382 , n44957 , 
 n335384 , n335385 , n335386 , n335387 , n44962 , n335389 , n44964 , n44965 , n335392 , n335393 , 
 n335394 , n335395 , n44970 , n335397 , n335398 , n335399 , n335400 , n44975 , n44976 , n335403 , 
 n44978 , n335405 , n335406 , n335407 , n335408 , n335409 , n335410 , n44985 , n335412 , n335413 , 
 n44988 , n335415 , n335416 , n335417 , n335418 , n335419 , n335420 , n335421 , n335422 , n335423 , 
 n44998 , n335425 , n335426 , n335427 , n45002 , n335429 , n335430 , n335431 , n45006 , n45007 , 
 n335434 , n335435 , n45010 , n335437 , n335438 , n335439 , n335440 , n335441 , n45016 , n335443 , 
 n45018 , n335445 , n335446 , n335447 , n335448 , n335449 , n335450 , n335451 , n45026 , n335453 , 
 n45028 , n335455 , n335456 , n335457 , n335458 , n45033 , n335460 , n335461 , n45036 , n335463 , 
 n335464 , n335465 , n335466 , n335467 , n335468 , n335469 , n45044 , n335471 , n335472 , n335473 , 
 n335474 , n335475 , n335476 , n335477 , n335478 , n45053 , n335480 , n335481 , n45056 , n335483 , 
 n335484 , n45059 , n335486 , n335487 , n335488 , n45063 , n45064 , n45065 , n335492 , n335493 , 
 n45068 , n45069 , n45070 , n335497 , n335498 , n335499 , n335500 , n335501 , n335502 , n335503 , 
 n335504 , n45079 , n335506 , n335507 , n335508 , n335509 , n45084 , n45085 , n335512 , n335513 , 
 n335514 , n335515 , n335516 , n335517 , n45092 , n335519 , n335520 , n45095 , n45096 , n335523 , 
 n335524 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n335532 , n335533 , 
 n335534 , n335535 , n335536 , n335537 , n335538 , n335539 , n335540 , n45115 , n45116 , n335543 , 
 n335544 , n335545 , n335546 , n335547 , n335548 , n45123 , n335550 , n335551 , n335552 , n335553 , 
 n335554 , n45129 , n45130 , n335557 , n335558 , n335559 , n335560 , n45135 , n335562 , n335563 , 
 n45138 , n335565 , n335566 , n335567 , n45142 , n335569 , n335570 , n335571 , n335572 , n335573 , 
 n335574 , n45149 , n335576 , n335577 , n335578 , n335579 , n45154 , n335581 , n335582 , n335583 , 
 n335584 , n335585 , n335586 , n45161 , n335588 , n335589 , n45164 , n335591 , n335592 , n335593 , 
 n335594 , n335595 , n335596 , n335597 , n335598 , n45173 , n335600 , n335601 , n335602 , n45177 , 
 n45178 , n335605 , n45180 , n45181 , n335608 , n335609 , n335610 , n335611 , n335612 , n335613 , 
 n45188 , n335615 , n335616 , n335617 , n45192 , n45193 , n45194 , n335621 , n335622 , n335623 , 
 n45198 , n45199 , n45200 , n335627 , n335628 , n45203 , n335630 , n335631 , n335632 , n335633 , 
 n335634 , n335635 , n335636 , n335637 , n45212 , n335639 , n45214 , n335641 , n335642 , n335643 , 
 n45218 , n335645 , n335646 , n335647 , n335648 , n45223 , n45224 , n335651 , n45226 , n335653 , 
 n335654 , n45229 , n335656 , n45231 , n335658 , n335659 , n335660 , n335661 , n335662 , n335663 , 
 n335664 , n45239 , n335666 , n335667 , n335668 , n335669 , n45244 , n45245 , n45246 , n335673 , 
 n335674 , n335675 , n335676 , n45251 , n45252 , n45253 , n45254 , n335681 , n335682 , n335683 , 
 n335684 , n335685 , n335686 , n335687 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , 
 n45268 , n45269 , n45270 , n335697 , n335698 , n335699 , n335700 , n335701 , n335702 , n335703 , 
 n335704 , n45279 , n45280 , n335707 , n335708 , n335709 , n45284 , n335711 , n335712 , n45287 , 
 n335714 , n335715 , n335716 , n45291 , n45292 , n45293 , n45294 , n335721 , n335722 , n45297 , 
 n335724 , n335725 , n335726 , n335727 , n335728 , n45303 , n335730 , n335731 , n335732 , n335733 , 
 n45308 , n335735 , n335736 , n335737 , n335738 , n45313 , n335740 , n45315 , n335742 , n45317 , 
 n45318 , n335745 , n335746 , n45321 , n335748 , n335749 , n335750 , n335751 , n335752 , n45327 , 
 n335754 , n335755 , n335756 , n45331 , n45332 , n335759 , n45334 , n45335 , n45336 , n45337 , 
 n335764 , n335765 , n335766 , n45341 , n45342 , n45343 , n45344 , n335771 , n335772 , n335773 , 
 n335774 , n335775 , n45350 , n335777 , n335778 , n335779 , n45354 , n335781 , n335782 , n335783 , 
 n335784 , n335785 , n335786 , n335787 , n335788 , n335789 , n335790 , n335791 , n335792 , n335793 , 
 n45368 , n45369 , n45370 , n45371 , n335798 , n335799 , n335800 , n335801 , n335802 , n335803 , 
 n335804 , n335805 , n335806 , n335807 , n45382 , n45383 , n335810 , n335811 , n335812 , n335813 , 
 n335814 , n335815 , n45390 , n335817 , n335818 , n45393 , n45394 , n335821 , n45396 , n335823 , 
 n335824 , n45399 , n45400 , n335827 , n335828 , n335829 , n335830 , n45405 , n335832 , n335833 , 
 n335834 , n335835 , n335836 , n45411 , n45412 , n45413 , n335840 , n45415 , n335842 , n335843 , 
 n45418 , n335845 , n335846 , n335847 , n335848 , n335849 , n335850 , n335851 , n335852 , n45427 , 
 n45428 , n45429 , n335856 , n335857 , n335858 , n335859 , n45434 , n45435 , n45436 , n45437 , 
 n45438 , n335865 , n335866 , n335867 , n335868 , n335869 , n335870 , n335871 , n335872 , n335873 , 
 n335874 , n335875 , n335876 , n335877 , n45452 , n335879 , n335880 , n335881 , n335882 , n335883 , 
 n335884 , n335885 , n45460 , n335887 , n335888 , n335889 , n335890 , n335891 , n335892 , n335893 , 
 n45468 , n45469 , n335896 , n335897 , n335898 , n335899 , n335900 , n335901 , n335902 , n335903 , 
 n335904 , n335905 , n335906 , n335907 , n335908 , n335909 , n335910 , n335911 , n335912 , n45487 , 
 n335914 , n335915 , n335916 , n335917 , n45492 , n335919 , n335920 , n335921 , n335922 , n335923 , 
 n335924 , n335925 , n335926 , n335927 , n335928 , n335929 , n335930 , n45505 , n45506 , n335933 , 
 n335934 , n335935 , n335936 , n335937 , n335938 , n45513 , n45514 , n45515 , n45516 , n45517 , 
 n45518 , n45519 , n45520 , n335947 , n45522 , n45523 , n335950 , n335951 , n45526 , n335953 , 
 n335954 , n335955 , n45530 , n335957 , n335958 , n335959 , n45534 , n335961 , n335962 , n335963 , 
 n335964 , n335965 , n335966 , n335967 , n335968 , n335969 , n335970 , n45545 , n335972 , n45547 , 
 n45548 , n335975 , n335976 , n45551 , n335978 , n335979 , n335980 , n45555 , n335982 , n335983 , 
 n335984 , n45559 , n335986 , n45561 , n335988 , n45563 , n45564 , n335991 , n335992 , n45567 , 
 n45568 , n335995 , n335996 , n335997 , n335998 , n335999 , n336000 , n336001 , n336002 , n336003 , 
 n336004 , n336005 , n336006 , n336007 , n336008 , n45583 , n336010 , n336011 , n336012 , n336013 , 
 n336014 , n336015 , n336016 , n336017 , n336018 , n336019 , n336020 , n336021 , n336022 , n336023 , 
 n336024 , n336025 , n336026 , n336027 , n336028 , n336029 , n336030 , n336031 , n45606 , n336033 , 
 n336034 , n336035 , n45610 , n45611 , n45612 , n336039 , n336040 , n45615 , n336042 , n336043 , 
 n336044 , n336045 , n336046 , n336047 , n336048 , n336049 , n336050 , n336051 , n336052 , n336053 , 
 n336054 , n45629 , n336056 , n45631 , n45632 , n336059 , n336060 , n336061 , n336062 , n45637 , 
 n336064 , n45639 , n45640 , n336067 , n336068 , n45643 , n336070 , n336071 , n336072 , n336073 , 
 n336074 , n336075 , n336076 , n45651 , n336078 , n336079 , n336080 , n336081 , n336082 , n336083 , 
 n336084 , n336085 , n336086 , n336087 , n336088 , n336089 , n336090 , n336091 , n336092 , n336093 , 
 n336094 , n336095 , n336096 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , 
 n336104 , n45679 , n45680 , n336107 , n336108 , n336109 , n336110 , n336111 , n336112 , n45687 , 
 n336114 , n336115 , n336116 , n45691 , n45692 , n336119 , n45694 , n45695 , n336122 , n336123 , 
 n336124 , n336125 , n336126 , n336127 , n336128 , n45703 , n45704 , n336131 , n336132 , n336133 , 
 n336134 , n336135 , n336136 , n45711 , n336138 , n336139 , n336140 , n336141 , n336142 , n336143 , 
 n336144 , n336145 , n336146 , n336147 , n45722 , n45723 , n336150 , n45725 , n45726 , n336153 , 
 n45728 , n45729 , n45730 , n45731 , n336158 , n336159 , n45734 , n336161 , n45736 , n336163 , 
 n336164 , n336165 , n45740 , n336167 , n336168 , n45743 , n45744 , n45745 , n45746 , n45747 , 
 n336174 , n45749 , n45750 , n45751 , n45752 , n336179 , n336180 , n336181 , n45756 , n336183 , 
 n336184 , n336185 , n45760 , n336187 , n336188 , n336189 , n336190 , n45765 , n336192 , n336193 , 
 n45768 , n336195 , n45770 , n45771 , n336198 , n336199 , n45774 , n336201 , n336202 , n45777 , 
 n336204 , n45779 , n336206 , n336207 , n45782 , n336209 , n336210 , n45785 , n45786 , n45787 , 
 n45788 , n336215 , n45790 , n336217 , n336218 , n45793 , n336220 , n336221 , n336222 , n45797 , 
 n336224 , n336225 , n336226 , n336227 , n45802 , n336229 , n336230 , n336231 , n336232 , n45807 , 
 n336234 , n336235 , n336236 , n45811 , n336238 , n336239 , n45814 , n336241 , n336242 , n45817 , 
 n336244 , n336245 , n45820 , n336247 , n336248 , n45823 , n336250 , n336251 , n336252 , n45827 , 
 n336254 , n336255 , n336256 , n45831 , n336258 , n336259 , n336260 , n45835 , n336262 , n45837 , 
 n336264 , n336265 , n45840 , n45841 , n336268 , n45843 , n336270 , n336271 , n45846 , n336273 , 
 n336274 , n45849 , n45850 , n45851 , n45852 , n336279 , n336280 , n336281 , n45856 , n336283 , 
 n336284 , n336285 , n45860 , n336287 , n336288 , n336289 , n45864 , n336291 , n45866 , n45867 , 
 n336294 , n45869 , n336296 , n336297 , n45872 , n45873 , n45874 , n45875 , n336302 , n336303 , 
 n336304 , n45879 , n336306 , n336307 , n336308 , n45883 , n336310 , n336311 , n336312 , n45887 , 
 n45888 , n45889 , n45890 , n336317 , n336318 , n45893 , n336320 , n336321 , n336322 , n45897 , 
 n336324 , n336325 , n336326 , n45901 , n336328 , n336329 , n336330 , n336331 , n45906 , n336333 , 
 n45908 , n336335 , n336336 , n45911 , n336338 , n336339 , n336340 , n336341 , n336342 , n45917 , 
 n336344 , n336345 , n336346 , n45921 , n336348 , n336349 , n336350 , n336351 , n45926 , n336353 , 
 n336354 , n336355 , n336356 , n45931 , n45932 , n45933 , n45934 , n45935 , n336362 , n336363 , 
 n336364 , n45939 , n336366 , n336367 , n336368 , n336369 , n45944 , n336371 , n336372 , n336373 , 
 n336374 , n45949 , n45950 , n45951 , n45952 , n45953 , n336380 , n336381 , n45956 , n336383 , 
 n336384 , n336385 , n45960 , n336387 , n336388 , n336389 , n336390 , n336391 , n45966 , n45967 , 
 n45968 , n45969 , n45970 , n336397 , n336398 , n336399 , n336400 , n45975 , n336402 , n336403 , 
 n45978 , n336405 , n336406 , n336407 , n45982 , n336409 , n45984 , n45985 , n336412 , n45987 , 
 n336414 , n336415 , n45990 , n336417 , n336418 , n45993 , n45994 , n336421 , n336422 , n336423 , 
 n45998 , n336425 , n336426 , n336427 , n336428 , n336429 , n46004 , n46005 , n46006 , n46007 , 
 n46008 , n336435 , n46010 , n46011 , n336438 , n336439 , n336440 , n46015 , n336442 , n336443 , 
 n336444 , n46019 , n336446 , n336447 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , 
 n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , 
 n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , 
 n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , 
 n46058 , n336485 , n46060 , n336487 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , 
 n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , 
 n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , 
 n46088 , n46089 , n46090 , n46091 , n46092 , n336519 , n46094 , n336521 , n336522 , n46097 , 
 n336524 , n46099 , n46100 , n46101 , n46102 , n336529 , n336530 , n336531 , n46106 , n336533 , 
 n46108 , n46109 , n46110 , n336537 , n336538 , n336539 , n46114 , n336541 , n336542 , n46117 , 
 n336544 , n336545 , n46120 , n336547 , n336548 , n46123 , n336550 , n336551 , n336552 , n336553 , 
 n46128 , n336555 , n336556 , n46131 , n336558 , n336559 , n46134 , n336561 , n46136 , n336563 , 
 n46138 , n336565 , n46140 , n46141 , n336568 , n46143 , n336570 , n46145 , n336572 , n46147 , 
 n46148 , n336575 , n336576 , n46151 , n336578 , n46153 , n336580 , n46155 , n46156 , n336583 , 
 n336584 , n46159 , n46160 , n336587 , n336588 , n46163 , n336590 , n336591 , n46166 , n336593 , 
 n336594 , n46169 , n336596 , n336597 , n46172 , n46173 , n336600 , n336601 , n46176 , n336603 , 
 n46178 , n336605 , n336606 , n336607 , n46182 , n336609 , n336610 , n46185 , n46186 , n46187 , 
 n46188 , n336615 , n336616 , n46191 , n336618 , n336619 , n46194 , n336621 , n336622 , n46197 , 
 n336624 , n336625 , n336626 , n46201 , n336628 , n336629 , n336630 , n46205 , n336632 , n336633 , 
 n46208 , n336635 , n336636 , n336637 , n46212 , n336639 , n336640 , n46215 , n336642 , n336643 , 
 n336644 , n46219 , n336646 , n336647 , n336648 , n46223 , n336650 , n336651 , n336652 , n336653 , 
 n46228 , n46229 , n46230 , n46231 , n336658 , n336659 , n336660 , n46235 , n336662 , n336663 , 
 n336664 , n46239 , n336666 , n336667 , n46242 , n336669 , n336670 , n336671 , n46246 , n336673 , 
 n336674 , n336675 , n46250 , n336677 , n46252 , n46253 , n46254 , n336681 , n46256 , n336683 , 
 n46258 , n336685 , n46260 , n46261 , n336688 , n336689 , n46264 , n336691 , n336692 , n336693 , 
 n46268 , n336695 , n336696 , n46272 , n336698 , n46274 , n336700 , n336701 , n336702 , n336703 , 
 n46279 , n46280 , n336706 , n336707 , n336708 , n336709 , n46285 , n336711 , n336712 , n336713 , 
 n336714 , n46290 , n336716 , n336717 , n336718 , n336719 , n336720 , n46296 , n46297 , n46298 , 
 n46299 , n46300 , n336726 , n336727 , n336728 , n336729 , n46305 , n336731 , n336732 , n336733 , 
 n336734 , n46310 , n336736 , n336737 , n336738 , n336739 , n46315 , n46316 , n46317 , n46318 , 
 n336744 , n336745 , n336746 , n336747 , n46323 , n336749 , n336750 , n336751 , n46327 , n46328 , 
 n336754 , n336755 , n46331 , n336757 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , 
 n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n336773 , 
 n46349 , n336775 , n336776 , n46352 , n46353 , n336779 , n336780 , n336781 , n336782 , n336783 , 
 n46359 , n46360 , n46361 , n46362 , n46363 , n336789 , n46365 , n46366 , n46367 , n46368 , 
 n46369 , n46370 , n46371 , n46372 , n336798 , n46374 , n336800 , n336801 , n46377 , n46378 , 
 n336804 , n336805 , n336806 , n336807 , n336808 , n46384 , n336810 , n46386 , n46387 , n46388 , 
 n46389 , n336815 , n46391 , n336817 , n336818 , n46394 , n46395 , n336821 , n336822 , n336823 , 
 n46399 , n46400 , n46401 , n336827 , n46403 , n46404 , n46405 , n46406 , n46407 , n336833 , 
 n46409 , n46410 , n336836 , n336837 , n336838 , n46414 , n46415 , n336841 , n46417 , n46418 , 
 n46419 , n46420 , n336846 , n46422 , n46423 , n336849 , n336850 , n336851 , n336852 , n46428 , 
 n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n336860 , n46436 , n46437 , n336863 , 
 n336864 , n336865 , n46441 , n46442 , n336868 , n46444 , n336870 , n46446 , n336872 , n46448 , 
 n46449 , n336875 , n46451 , n336877 , n336878 , n46454 , n46455 , n336881 , n336882 , n336883 , 
 n46459 , n336885 , n46461 , n46462 , n46463 , n46464 , n46465 , n336891 , n336892 , n46468 , 
 n336894 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , 
 n336904 , n46480 , n336906 , n46482 , n46483 , n336909 , n46485 , n336911 , n46487 , n46488 , 
 n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , 
 n336924 , n46500 , n336926 , n46502 , n46503 , n336929 , n46505 , n336931 , n46507 , n46508 , 
 n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n336941 , n46517 , n336943 , 
 n46519 , n46520 , n336946 , n46522 , n336948 , n46524 , n46525 , n46526 , n46527 , n46528 , 
 n46529 , n46530 , n46531 , n336957 , n46533 , n336959 , n46535 , n46536 , n336962 , n46538 , 
 n336964 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , 
 n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , 
 n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , 
 n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , 
 n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , 
 n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , 
 n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , 
 n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , 
 n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , 
 n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , 
 n46639 , n46640 , n337066 , n337067 , n46643 , n337069 , n46645 , n46646 , n46647 , n46648 , 
 n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n337082 , n46658 , 
 n337084 , n46660 , n337086 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , 
 n46669 , n337095 , n337096 , n46672 , n337098 , n337099 , n337100 , n46676 , n337102 , n337103 , 
 n337104 , n46680 , n337106 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , 
 n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , 
 n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n337131 , n337132 , n46708 , 
 n337134 , n337135 , n46711 , n337137 , n46713 , n337139 , n46715 , n46716 , n46717 , n46718 , 
 n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , 
 n46729 , n46730 , n46731 , n337157 , n337158 , n46734 , n337160 , n337161 , n337162 , n337163 , 
 n46739 , n337165 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , 
 n46749 , n337175 , n337176 , n46752 , n337178 , n46754 , n46755 , n46756 , n46757 , n46758 , 
 n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , 
 n46769 , n46770 , n46771 , n46772 , n337198 , n337199 , n337200 , n46776 , n337202 , n46778 , 
 n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , 
 n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , 
 n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , 
 n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , 
 n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , 
 n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , 
 n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , 
 n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , 
 n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , 
 n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , 
 n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , 
 n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , 
 n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , 
 n46909 , n46910 , n46911 , n337337 , n337338 , n46914 , n46915 , n337341 , n46917 , n46918 , 
 n46919 , n46920 , n337346 , n46922 , n46923 , n337349 , n337350 , n337351 , n46927 , n337353 , 
 n337354 , n337355 , n46931 , n337357 , n337358 , n337359 , n337360 , n46936 , n337362 , n337363 , 
 n337364 , n337365 , n46941 , n337367 , n337368 , n337369 , n46945 , n337371 , n337372 , n337373 , 
 n337374 , n46950 , n46951 , n46952 , n46953 , n46954 , n337380 , n46956 , n46957 , n46958 , 
 n46959 , n46960 , n337386 , n337387 , n46963 , n337389 , n46965 , n337391 , n337392 , n46968 , 
 n337394 , n46970 , n46971 , n46972 , n46973 , n46974 , C0n , C0 ;
buf ( n768 , n0 );
buf ( n769 , n1 );
buf ( n770 , n2 );
buf ( n771 , n3 );
buf ( n772 , n4 );
buf ( n773 , n5 );
buf ( n774 , n6 );
buf ( n775 , n7 );
buf ( n776 , n8 );
buf ( n777 , n9 );
buf ( n778 , n10 );
buf ( n779 , n11 );
buf ( n780 , n12 );
buf ( n781 , n13 );
buf ( n782 , n14 );
buf ( n783 , n15 );
buf ( n784 , n16 );
buf ( n785 , n17 );
buf ( n786 , n18 );
buf ( n787 , n19 );
buf ( n788 , n20 );
buf ( n789 , n21 );
buf ( n790 , n22 );
buf ( n791 , n23 );
buf ( n792 , n24 );
buf ( n793 , n25 );
buf ( n794 , n26 );
buf ( n795 , n27 );
buf ( n796 , n28 );
buf ( n797 , n29 );
buf ( n798 , n30 );
buf ( n799 , n31 );
buf ( n800 , n32 );
buf ( n801 , n33 );
buf ( n802 , n34 );
buf ( n803 , n35 );
buf ( n804 , n36 );
buf ( n805 , n37 );
buf ( n806 , n38 );
buf ( n807 , n39 );
buf ( n808 , n40 );
buf ( n809 , n41 );
buf ( n810 , n42 );
buf ( n811 , n43 );
buf ( n812 , n44 );
buf ( n813 , n45 );
buf ( n814 , n46 );
buf ( n815 , n47 );
buf ( n816 , n48 );
buf ( n817 , n49 );
buf ( n818 , n50 );
buf ( n819 , n51 );
buf ( n820 , n52 );
buf ( n821 , n53 );
buf ( n822 , n54 );
buf ( n823 , n55 );
buf ( n824 , n56 );
buf ( n825 , n57 );
buf ( n826 , n58 );
buf ( n827 , n59 );
buf ( n828 , n60 );
buf ( n829 , n61 );
buf ( n830 , n62 );
buf ( n831 , n63 );
buf ( n832 , n64 );
buf ( n833 , n65 );
buf ( n834 , n66 );
buf ( n835 , n67 );
buf ( n836 , n68 );
buf ( n837 , n69 );
buf ( n838 , n70 );
buf ( n839 , n71 );
buf ( n840 , n72 );
buf ( n841 , n73 );
buf ( n842 , n74 );
buf ( n843 , n75 );
buf ( n844 , n76 );
buf ( n845 , n77 );
buf ( n846 , n78 );
buf ( n847 , n79 );
buf ( n848 , n80 );
buf ( n849 , n81 );
buf ( n850 , n82 );
buf ( n851 , n83 );
buf ( n852 , n84 );
buf ( n853 , n85 );
buf ( n854 , n86 );
buf ( n855 , n87 );
buf ( n856 , n88 );
buf ( n857 , n89 );
buf ( n858 , n90 );
buf ( n859 , n91 );
buf ( n860 , n92 );
buf ( n861 , n93 );
buf ( n862 , n94 );
buf ( n863 , n95 );
buf ( n864 , n96 );
buf ( n865 , n97 );
buf ( n866 , n98 );
buf ( n867 , n99 );
buf ( n868 , n100 );
buf ( n869 , n101 );
buf ( n870 , n102 );
buf ( n871 , n103 );
buf ( n872 , n104 );
buf ( n873 , n105 );
buf ( n874 , n106 );
buf ( n875 , n107 );
buf ( n876 , n108 );
buf ( n877 , n109 );
buf ( n878 , n110 );
buf ( n879 , n111 );
buf ( n880 , n112 );
buf ( n881 , n113 );
buf ( n882 , n114 );
buf ( n883 , n115 );
buf ( n884 , n116 );
buf ( n885 , n117 );
buf ( n886 , n118 );
buf ( n887 , n119 );
buf ( n888 , n120 );
buf ( n889 , n121 );
buf ( n890 , n122 );
buf ( n891 , n123 );
buf ( n892 , n124 );
buf ( n893 , n125 );
buf ( n894 , n126 );
buf ( n895 , n127 );
buf ( n128 , n896 );
buf ( n129 , n897 );
buf ( n130 , n898 );
buf ( n131 , n899 );
buf ( n132 , n900 );
buf ( n133 , n901 );
buf ( n134 , n902 );
buf ( n135 , n903 );
buf ( n136 , n904 );
buf ( n137 , n905 );
buf ( n138 , n906 );
buf ( n139 , n907 );
buf ( n140 , n908 );
buf ( n141 , n909 );
buf ( n142 , n910 );
buf ( n143 , n911 );
buf ( n144 , n912 );
buf ( n145 , n913 );
buf ( n146 , n914 );
buf ( n147 , n915 );
buf ( n148 , n916 );
buf ( n149 , n917 );
buf ( n150 , n918 );
buf ( n151 , n919 );
buf ( n152 , n920 );
buf ( n153 , n921 );
buf ( n154 , n922 );
buf ( n155 , n923 );
buf ( n156 , n924 );
buf ( n157 , n925 );
buf ( n158 , n926 );
buf ( n159 , n927 );
buf ( n160 , n928 );
buf ( n161 , n929 );
buf ( n162 , n930 );
buf ( n163 , n931 );
buf ( n164 , n932 );
buf ( n165 , n933 );
buf ( n166 , n934 );
buf ( n167 , n935 );
buf ( n168 , n936 );
buf ( n169 , n937 );
buf ( n170 , n938 );
buf ( n171 , n939 );
buf ( n172 , n940 );
buf ( n173 , n941 );
buf ( n174 , n942 );
buf ( n175 , n943 );
buf ( n176 , n944 );
buf ( n177 , n945 );
buf ( n178 , n946 );
buf ( n179 , n947 );
buf ( n180 , n948 );
buf ( n181 , n949 );
buf ( n182 , n950 );
buf ( n183 , n951 );
buf ( n184 , n952 );
buf ( n185 , n953 );
buf ( n186 , n954 );
buf ( n187 , n955 );
buf ( n188 , n956 );
buf ( n189 , n957 );
buf ( n190 , n958 );
buf ( n191 , n959 );
buf ( n192 , n960 );
buf ( n193 , n961 );
buf ( n194 , n962 );
buf ( n195 , n963 );
buf ( n196 , n964 );
buf ( n197 , n965 );
buf ( n198 , n966 );
buf ( n199 , n967 );
buf ( n200 , n968 );
buf ( n201 , n969 );
buf ( n202 , n970 );
buf ( n203 , n971 );
buf ( n204 , n972 );
buf ( n205 , n973 );
buf ( n206 , n974 );
buf ( n207 , n975 );
buf ( n208 , n976 );
buf ( n209 , n977 );
buf ( n210 , n978 );
buf ( n211 , n979 );
buf ( n212 , n980 );
buf ( n213 , n981 );
buf ( n214 , n982 );
buf ( n215 , n983 );
buf ( n216 , n984 );
buf ( n217 , n985 );
buf ( n218 , n986 );
buf ( n219 , n987 );
buf ( n220 , n988 );
buf ( n221 , n989 );
buf ( n222 , n990 );
buf ( n223 , n991 );
buf ( n224 , n992 );
buf ( n225 , n993 );
buf ( n226 , n994 );
buf ( n227 , n995 );
buf ( n228 , n996 );
buf ( n229 , n997 );
buf ( n230 , n998 );
buf ( n231 , n999 );
buf ( n232 , n1000 );
buf ( n233 , n1001 );
buf ( n234 , n1002 );
buf ( n235 , n1003 );
buf ( n236 , n1004 );
buf ( n237 , n1005 );
buf ( n238 , n1006 );
buf ( n239 , n1007 );
buf ( n240 , n1008 );
buf ( n241 , n1009 );
buf ( n242 , n1010 );
buf ( n243 , n1011 );
buf ( n244 , n1012 );
buf ( n245 , n1013 );
buf ( n246 , n1014 );
buf ( n247 , n1015 );
buf ( n248 , n1016 );
buf ( n249 , n1017 );
buf ( n250 , n1018 );
buf ( n251 , n1019 );
buf ( n252 , n1020 );
buf ( n253 , n1021 );
buf ( n254 , n1022 );
buf ( n255 , n1023 );
buf ( n256 , n1024 );
buf ( n257 , n1025 );
buf ( n258 , n1026 );
buf ( n259 , n1027 );
buf ( n260 , n1028 );
buf ( n261 , n1029 );
buf ( n262 , n1030 );
buf ( n263 , n1031 );
buf ( n264 , n1032 );
buf ( n265 , n1033 );
buf ( n266 , n1034 );
buf ( n267 , n1035 );
buf ( n268 , n1036 );
buf ( n269 , n1037 );
buf ( n270 , n1038 );
buf ( n271 , n1039 );
buf ( n272 , n1040 );
buf ( n273 , n1041 );
buf ( n274 , n1042 );
buf ( n275 , n1043 );
buf ( n276 , n1044 );
buf ( n277 , n1045 );
buf ( n278 , n1046 );
buf ( n279 , n1047 );
buf ( n280 , n1048 );
buf ( n281 , n1049 );
buf ( n282 , n1050 );
buf ( n283 , n1051 );
buf ( n284 , n1052 );
buf ( n285 , n1053 );
buf ( n286 , n1054 );
buf ( n287 , n1055 );
buf ( n288 , n1056 );
buf ( n289 , n1057 );
buf ( n290 , n1058 );
buf ( n291 , n1059 );
buf ( n292 , n1060 );
buf ( n293 , n1061 );
buf ( n294 , n1062 );
buf ( n295 , n1063 );
buf ( n296 , n1064 );
buf ( n297 , n1065 );
buf ( n298 , n1066 );
buf ( n299 , n1067 );
buf ( n300 , n1068 );
buf ( n301 , n1069 );
buf ( n302 , n1070 );
buf ( n303 , n1071 );
buf ( n304 , n1072 );
buf ( n305 , n1073 );
buf ( n306 , n1074 );
buf ( n307 , n1075 );
buf ( n308 , n1076 );
buf ( n309 , n1077 );
buf ( n310 , n1078 );
buf ( n311 , n1079 );
buf ( n312 , n1080 );
buf ( n313 , n1081 );
buf ( n314 , n1082 );
buf ( n315 , n1083 );
buf ( n316 , n1084 );
buf ( n317 , n1085 );
buf ( n318 , n1086 );
buf ( n319 , n1087 );
buf ( n320 , n1088 );
buf ( n321 , n1089 );
buf ( n322 , n1090 );
buf ( n323 , n1091 );
buf ( n324 , n1092 );
buf ( n325 , n1093 );
buf ( n326 , n1094 );
buf ( n327 , n1095 );
buf ( n328 , n1096 );
buf ( n329 , n1097 );
buf ( n330 , n1098 );
buf ( n331 , n1099 );
buf ( n332 , n1100 );
buf ( n333 , n1101 );
buf ( n334 , n1102 );
buf ( n335 , n1103 );
buf ( n336 , n1104 );
buf ( n337 , n1105 );
buf ( n338 , n1106 );
buf ( n339 , n1107 );
buf ( n340 , n1108 );
buf ( n341 , n1109 );
buf ( n342 , n1110 );
buf ( n343 , n1111 );
buf ( n344 , n1112 );
buf ( n345 , n1113 );
buf ( n346 , n1114 );
buf ( n347 , n1115 );
buf ( n348 , n1116 );
buf ( n349 , n1117 );
buf ( n350 , n1118 );
buf ( n351 , n1119 );
buf ( n352 , n1120 );
buf ( n353 , n1121 );
buf ( n354 , n1122 );
buf ( n355 , n1123 );
buf ( n356 , n1124 );
buf ( n357 , n1125 );
buf ( n358 , n1126 );
buf ( n359 , n1127 );
buf ( n360 , n1128 );
buf ( n361 , n1129 );
buf ( n362 , n1130 );
buf ( n363 , n1131 );
buf ( n364 , n1132 );
buf ( n365 , n1133 );
buf ( n366 , n1134 );
buf ( n367 , n1135 );
buf ( n368 , n1136 );
buf ( n369 , n1137 );
buf ( n370 , n1138 );
buf ( n371 , n1139 );
buf ( n372 , n1140 );
buf ( n373 , n1141 );
buf ( n374 , n1142 );
buf ( n375 , n1143 );
buf ( n376 , n1144 );
buf ( n377 , n1145 );
buf ( n378 , n1146 );
buf ( n379 , n1147 );
buf ( n380 , n1148 );
buf ( n381 , n1149 );
buf ( n382 , n1150 );
buf ( n383 , n1151 );
buf ( n896 , n46607 );
buf ( n897 , n46617 );
buf ( n898 , n46628 );
buf ( n899 , n46566 );
buf ( n900 , n46597 );
buf ( n901 , n46586 );
buf ( n902 , n46576 );
buf ( n903 , n335196 );
buf ( n904 , n335255 );
buf ( n905 , n44870 );
buf ( n906 , n334974 );
buf ( n907 , n335317 );
buf ( n908 , n44940 );
buf ( n909 , n335403 );
buf ( n910 , n335007 );
buf ( n911 , n335504 );
buf ( n912 , n335571 );
buf ( n913 , n46875 );
buf ( n914 , n335622 );
buf ( n915 , n335656 );
buf ( n916 , n335483 );
buf ( n917 , n335440 );
buf ( n918 , n46865 );
buf ( n919 , n45270 );
buf ( n920 , n335750 );
buf ( n921 , n335779 );
buf ( n922 , n335807 );
buf ( n923 , n335829 );
buf ( n924 , n45438 );
buf ( n925 , n335888 );
buf ( n926 , n335681 );
buf ( n927 , n46911 );
buf ( n928 , n45515 );
buf ( n929 , n46721 );
buf ( n930 , n336695 );
buf ( n931 , n46760 );
buf ( n932 , n46770 );
buf ( n933 , n335984 );
buf ( n934 , n335962 );
buf ( n935 , n335997 );
buf ( n936 , n336044 );
buf ( n937 , n336215 );
buf ( n938 , n336081 );
buf ( n939 , n45672 );
buf ( n940 , n336139 );
buf ( n941 , n336158 );
buf ( n942 , n336179 );
buf ( n943 , n46923 );
buf ( n944 , n336691 );
buf ( n945 , n46792 );
buf ( n946 , n46814 );
buf ( n947 , n336677 );
buf ( n948 , n46905 );
buf ( n949 , n336279 );
buf ( n950 , n336302 );
buf ( n951 , n336317 );
buf ( n952 , n336362 );
buf ( n953 , n336380 );
buf ( n954 , n46833 );
buf ( n955 , n336397 );
buf ( n956 , n46822 );
buf ( n957 , n336435 );
buf ( n958 , n336438 );
buf ( n959 , n336658 );
buf ( n960 , n46498 );
buf ( n961 , n327055 );
buf ( n962 , n327107 );
buf ( n963 , n46515 );
buf ( n964 , n46705 );
buf ( n965 , n46531 );
buf ( n966 , n46547 );
buf ( n967 , n46556 );
buf ( n968 , n326645 );
buf ( n969 , n326677 );
buf ( n970 , n46669 );
buf ( n971 , n46478 );
buf ( n972 , n326740 );
buf ( n973 , n46636 );
buf ( n974 , n46652 );
buf ( n975 , n327243 );
buf ( n976 , n327295 );
buf ( n977 , n327345 );
buf ( n978 , n327394 );
buf ( n979 , n327603 );
buf ( n980 , n327439 );
buf ( n981 , n327215 );
buf ( n982 , n327643 );
buf ( n983 , n46688 );
buf ( n984 , n327157 );
buf ( n985 , n327676 );
buf ( n986 , n46887 );
buf ( n987 , n327506 );
buf ( n988 , n327545 );
buf ( n989 , n327480 );
buf ( n990 , n327571 );
buf ( n991 , n336726 );
buf ( n992 , n327798 );
buf ( n993 , n327830 );
buf ( n994 , n327851 );
buf ( n995 , n46748 );
buf ( n996 , n46731 );
buf ( n997 , n327733 );
buf ( n998 , n327707 );
buf ( n999 , n327907 );
buf ( n1000 , n327891 );
buf ( n1001 , n328049 );
buf ( n1002 , n327931 );
buf ( n1003 , n337346 );
buf ( n1004 , n327970 );
buf ( n1005 , n327993 );
buf ( n1006 , n328016 );
buf ( n1007 , n46959 );
buf ( n1008 , n328099 );
buf ( n1009 , n46897 );
buf ( n1010 , n328158 );
buf ( n1011 , n328507 );
buf ( n1012 , n46782 );
buf ( n1013 , n328184 );
buf ( n1014 , n328125 );
buf ( n1015 , n337106 );
buf ( n1016 , n328214 );
buf ( n1017 , n328232 );
buf ( n1018 , n328254 );
buf ( n1019 , n46850 );
buf ( n1020 , n328318 );
buf ( n1021 , n328433 );
buf ( n1022 , n328462 );
buf ( n1023 , n328471 );
buf ( n1024 , C0 );
buf ( n1025 , C0 );
buf ( n1026 , C0 );
buf ( n1027 , C0 );
buf ( n1028 , C0 );
buf ( n1029 , C0 );
buf ( n1030 , C0 );
buf ( n1031 , C0 );
buf ( n1032 , C0 );
buf ( n1033 , C0 );
buf ( n1034 , C0 );
buf ( n1035 , C0 );
buf ( n1036 , C0 );
buf ( n1037 , C0 );
buf ( n1038 , C0 );
buf ( n1039 , C0 );
buf ( n1040 , C0 );
buf ( n1041 , C0 );
buf ( n1042 , C0 );
buf ( n1043 , C0 );
buf ( n1044 , C0 );
buf ( n1045 , C0 );
buf ( n1046 , C0 );
buf ( n1047 , C0 );
buf ( n1048 , C0 );
buf ( n1049 , C0 );
buf ( n1050 , C0 );
buf ( n1051 , C0 );
buf ( n1052 , C0 );
buf ( n1053 , C0 );
buf ( n1054 , C0 );
buf ( n1055 , C0 );
buf ( n1056 , C0 );
buf ( n1057 , C0 );
buf ( n1058 , C0 );
buf ( n1059 , C0 );
buf ( n1060 , C0 );
buf ( n1061 , C0 );
buf ( n1062 , C0 );
buf ( n1063 , C0 );
buf ( n1064 , C0 );
buf ( n1065 , C0 );
buf ( n1066 , C0 );
buf ( n1067 , C0 );
buf ( n1068 , C0 );
buf ( n1069 , C0 );
buf ( n1070 , C0 );
buf ( n1071 , C0 );
buf ( n1072 , C0 );
buf ( n1073 , C0 );
buf ( n1074 , C0 );
buf ( n1075 , C0 );
buf ( n1076 , C0 );
buf ( n1077 , C0 );
buf ( n1078 , C0 );
buf ( n1079 , C0 );
buf ( n1080 , C0 );
buf ( n1081 , C0 );
buf ( n1082 , C0 );
buf ( n1083 , C0 );
buf ( n1084 , C0 );
buf ( n1085 , C0 );
buf ( n1086 , C0 );
buf ( n1087 , n331326 );
buf ( n1088 , n331516 );
buf ( n1089 , n331377 );
buf ( n1090 , n331617 );
buf ( n1091 , n331657 );
buf ( n1092 , n331708 );
buf ( n1093 , n40552 );
buf ( n1094 , n331025 );
buf ( n1095 , n331056 );
buf ( n1096 , n331120 );
buf ( n1097 , n331163 );
buf ( n1098 , n331986 );
buf ( n1099 , n330760 );
buf ( n1100 , n331556 );
buf ( n1101 , n331417 );
buf ( n1102 , n331450 );
buf ( n1103 , n331810 );
buf ( n1104 , n331878 );
buf ( n1105 , n331926 );
buf ( n1106 , n41360 );
buf ( n1107 , n332017 );
buf ( n1108 , n332070 );
buf ( n1109 , n332100 );
buf ( n1110 , n332405 );
buf ( n1111 , n332160 );
buf ( n1112 , n332210 );
buf ( n1113 , n332137 );
buf ( n1114 , n332254 );
buf ( n1115 , n332277 );
buf ( n1116 , n41887 );
buf ( n1117 , n332339 );
buf ( n1118 , n332366 );
buf ( n1119 , n332626 );
buf ( n1120 , n332612 );
buf ( n1121 , n332560 );
buf ( n1122 , n332519 );
buf ( n1123 , n332658 );
buf ( n1124 , n332700 );
buf ( n1125 , n332470 );
buf ( n1126 , n332442 );
buf ( n1127 , n332721 );
buf ( n1128 , n46807 );
buf ( n1129 , n46974 );
buf ( n1130 , n46799 );
buf ( n1131 , n333099 );
buf ( n1132 , n333126 );
buf ( n1133 , n333108 );
buf ( n1134 , n333112 );
buf ( n1135 , n332764 );
buf ( n1136 , n337380 );
buf ( n1137 , n332781 );
buf ( n1138 , n332874 );
buf ( n1139 , n332892 );
buf ( n1140 , n332924 );
buf ( n1141 , n42518 );
buf ( n1142 , n332836 );
buf ( n1143 , n332959 );
buf ( n1144 , n46844 );
buf ( n1145 , n332980 );
buf ( n1146 , n332999 );
buf ( n1147 , n333013 );
buf ( n1148 , n333032 );
buf ( n1149 , n42620 );
buf ( n1150 , n333049 );
buf ( n1151 , n333071 );
not ( n291647 , n831 );
buf ( n291648 , n849 );
xor ( n1221 , n830 , n787 );
buf ( n291650 , n1221 );
not ( n291651 , n291650 );
not ( n291652 , n831 );
nand ( n291653 , n291652 , n830 );
buf ( n291654 , n291653 );
not ( n291655 , n291654 );
buf ( n291656 , n291655 );
buf ( n291657 , n291656 );
not ( n291658 , n291657 );
or ( n291659 , n291651 , n291658 );
buf ( n291660 , n786 );
buf ( n291661 , n830 );
xor ( n291662 , n291660 , n291661 );
buf ( n291663 , n291662 );
buf ( n291664 , n291663 );
buf ( n291665 , n831 );
nand ( n1238 , n291664 , n291665 );
buf ( n291667 , n1238 );
buf ( n291668 , n291667 );
nand ( n1241 , n291659 , n291668 );
buf ( n291670 , n1241 );
buf ( n1243 , n291670 );
buf ( n291672 , n799 );
buf ( n291673 , n819 );
or ( n291674 , n291672 , n291673 );
buf ( n291675 , n820 );
nand ( n1248 , n291674 , n291675 );
buf ( n1249 , n1248 );
buf ( n1250 , n1249 );
buf ( n1251 , n799 );
buf ( n1252 , n819 );
nand ( n1253 , n1251 , n1252 );
buf ( n1254 , n1253 );
buf ( n1255 , n1254 );
buf ( n291684 , n818 );
and ( n291685 , n1250 , n1255 , n291684 );
buf ( n291686 , n291685 );
buf ( n291687 , n291686 );
xor ( n291688 , n1243 , n291687 );
buf ( n291689 , n291688 );
buf ( n291690 , n291689 );
buf ( n1263 , n788 );
buf ( n1264 , n830 );
xor ( n1265 , n1263 , n1264 );
buf ( n1266 , n1265 );
buf ( n1267 , n1266 );
not ( n1268 , n1267 );
not ( n291697 , n831 );
nand ( n1270 , n291697 , n830 );
not ( n1271 , n1270 );
buf ( n291700 , n1271 );
not ( n291701 , n291700 );
or ( n1274 , n1268 , n291701 );
buf ( n291703 , n1221 );
buf ( n291704 , n831 );
nand ( n291705 , n291703 , n291704 );
buf ( n291706 , n291705 );
buf ( n291707 , n291706 );
nand ( n291708 , n1274 , n291707 );
buf ( n291709 , n291708 );
buf ( n291710 , n291709 );
xor ( n291711 , n820 , n798 );
buf ( n291712 , n291711 );
not ( n291713 , n291712 );
xor ( n291714 , n821 , n822 );
and ( n291715 , n821 , n820 );
not ( n291716 , n821 );
not ( n1289 , n820 );
and ( n291718 , n291716 , n1289 );
nor ( n291719 , n291715 , n291718 );
not ( n1292 , n291719 );
nor ( n291721 , n291714 , n1292 );
buf ( n291722 , n291721 );
buf ( n291723 , n291722 );
not ( n291724 , n291723 );
or ( n1297 , n291713 , n291724 );
not ( n291726 , n821 );
not ( n1299 , n822 );
not ( n291728 , n1299 );
or ( n1301 , n291726 , n291728 );
buf ( n291730 , n821 );
not ( n291731 , n291730 );
buf ( n291732 , n291731 );
nand ( n291733 , n291732 , n822 );
nand ( n291734 , n1301 , n291733 );
buf ( n291735 , n291734 );
buf ( n291736 , n797 );
buf ( n291737 , n820 );
xor ( n291738 , n291736 , n291737 );
buf ( n291739 , n291738 );
buf ( n1312 , n291739 );
nand ( n1313 , n291735 , n1312 );
buf ( n1314 , n1313 );
buf ( n291743 , n1314 );
nand ( n1316 , n1297 , n291743 );
buf ( n1317 , n1316 );
buf ( n291746 , n1317 );
xor ( n1319 , n291710 , n291746 );
xor ( n291748 , n822 , n796 );
buf ( n291749 , n291748 );
not ( n1322 , n291749 );
and ( n1323 , n824 , n823 );
not ( n1324 , n824 );
not ( n1325 , n823 );
and ( n1326 , n1324 , n1325 );
nor ( n291755 , n1323 , n1326 );
not ( n1328 , n291755 );
xor ( n291757 , n823 , n822 );
nand ( n1330 , n1328 , n291757 );
buf ( n291759 , n1330 );
not ( n1332 , n291759 );
buf ( n291761 , n1332 );
buf ( n291762 , n291761 );
not ( n291763 , n291762 );
or ( n1336 , n1322 , n291763 );
xor ( n291765 , n823 , n824 );
not ( n1338 , n291765 );
not ( n1339 , n1338 );
buf ( n291768 , n1339 );
xor ( n291769 , n822 , n795 );
buf ( n1342 , n291769 );
nand ( n1343 , n291768 , n1342 );
buf ( n1344 , n1343 );
buf ( n291773 , n1344 );
nand ( n1346 , n1336 , n291773 );
buf ( n291775 , n1346 );
buf ( n291776 , n291775 );
and ( n1349 , n1319 , n291776 );
and ( n1350 , n291710 , n291746 );
or ( n1351 , n1349 , n1350 );
buf ( n291780 , n1351 );
buf ( n291781 , n291780 );
xor ( n1354 , n291690 , n291781 );
xor ( n1355 , n819 , n820 );
not ( n1356 , n1355 );
not ( n1357 , n1356 );
buf ( n291786 , n1357 );
buf ( n291787 , n291786 );
buf ( n291788 , n291787 );
buf ( n291789 , n291788 );
buf ( n291790 , n799 );
and ( n291791 , n291789 , n291790 );
buf ( n291792 , n291791 );
buf ( n291793 , n291792 );
xor ( n291794 , n828 , n790 );
buf ( n291795 , n291794 );
not ( n291796 , n291795 );
xor ( n291797 , n829 , n830 );
buf ( n291798 , n291797 );
not ( n291799 , n291798 );
buf ( n291800 , n291799 );
xor ( n1373 , n829 , n828 );
nand ( n291802 , n291800 , n1373 );
buf ( n1375 , n291802 );
not ( n1376 , n1375 );
buf ( n291805 , n1376 );
buf ( n291806 , n291805 );
buf ( n291807 , n291806 );
buf ( n291808 , n291807 );
buf ( n291809 , n291808 );
not ( n291810 , n291809 );
or ( n1383 , n291796 , n291810 );
buf ( n291812 , n291797 );
buf ( n291813 , n291812 );
buf ( n1386 , n789 );
buf ( n1387 , n828 );
xor ( n1388 , n1386 , n1387 );
buf ( n1389 , n1388 );
buf ( n291818 , n1389 );
nand ( n1391 , n291813 , n291818 );
buf ( n291820 , n1391 );
buf ( n291821 , n291820 );
nand ( n291822 , n1383 , n291821 );
buf ( n291823 , n291822 );
buf ( n291824 , n291823 );
xor ( n1397 , n291793 , n291824 );
xor ( n291826 , n824 , n794 );
buf ( n291827 , n291826 );
not ( n291828 , n291827 );
not ( n291829 , n825 );
nand ( n1402 , n291829 , n826 );
not ( n291831 , n826 );
nand ( n291832 , n291831 , n825 );
xor ( n1405 , n824 , n825 );
nand ( n1406 , n1402 , n291832 , n1405 );
not ( n291835 , n1406 );
buf ( n291836 , n291835 );
buf ( n291837 , n291836 );
buf ( n291838 , n291837 );
buf ( n291839 , n291838 );
not ( n291840 , n291839 );
or ( n1413 , n291828 , n291840 );
xor ( n291842 , n825 , n826 );
buf ( n291843 , n291842 );
buf ( n291844 , n291843 );
xor ( n291845 , n824 , n793 );
buf ( n291846 , n291845 );
nand ( n1419 , n291844 , n291846 );
buf ( n1420 , n1419 );
buf ( n291849 , n1420 );
nand ( n1422 , n1413 , n291849 );
buf ( n291851 , n1422 );
buf ( n291852 , n291851 );
and ( n1425 , n1397 , n291852 );
and ( n291854 , n291793 , n291824 );
or ( n291855 , n1425 , n291854 );
buf ( n291856 , n291855 );
buf ( n291857 , n291856 );
xor ( n291858 , n1354 , n291857 );
buf ( n291859 , n291858 );
buf ( n291860 , n291859 );
xor ( n291861 , n291710 , n291746 );
xor ( n1434 , n291861 , n291776 );
buf ( n291863 , n1434 );
buf ( n291864 , n291863 );
xor ( n291865 , n291793 , n291824 );
xor ( n291866 , n291865 , n291852 );
buf ( n291867 , n291866 );
buf ( n291868 , n291867 );
xor ( n291869 , n291864 , n291868 );
xor ( n1442 , n826 , n793 );
buf ( n291871 , n1442 );
not ( n291872 , n291871 );
xor ( n1445 , n828 , n827 );
not ( n291874 , n827 );
and ( n291875 , n826 , n291874 );
not ( n1448 , n826 );
and ( n291877 , n1448 , n827 );
nor ( n291878 , n291875 , n291877 );
nor ( n291879 , n1445 , n291878 );
buf ( n291880 , n291879 );
buf ( n1453 , n291880 );
buf ( n291882 , n1453 );
not ( n291883 , n291882 );
or ( n1456 , n291872 , n291883 );
xor ( n291885 , n828 , n827 );
buf ( n291886 , n291885 );
buf ( n291887 , n291886 );
buf ( n291888 , n792 );
buf ( n291889 , n826 );
xor ( n1462 , n291888 , n291889 );
buf ( n291891 , n1462 );
buf ( n291892 , n291891 );
nand ( n1465 , n291887 , n291892 );
buf ( n291894 , n1465 );
buf ( n291895 , n291894 );
nand ( n1468 , n1456 , n291895 );
buf ( n1469 , n1468 );
buf ( n291898 , n820 );
buf ( n291899 , n799 );
xor ( n1472 , n291898 , n291899 );
buf ( n291901 , n1472 );
not ( n1474 , n291901 );
buf ( n291903 , n291722 );
not ( n291904 , n291903 );
or ( n1477 , n1474 , n291904 );
buf ( n291906 , n291734 );
buf ( n291907 , n291906 );
buf ( n291908 , n291711 );
nand ( n291909 , n291907 , n291908 );
buf ( n291910 , n291909 );
nand ( n291911 , n1477 , n291910 );
xor ( n291912 , n1469 , n291911 );
buf ( n291913 , n799 );
buf ( n291914 , n821 );
or ( n291915 , n291913 , n291914 );
buf ( n291916 , n822 );
nand ( n1489 , n291915 , n291916 );
buf ( n291918 , n1489 );
buf ( n291919 , n291918 );
buf ( n291920 , n799 );
buf ( n291921 , n821 );
nand ( n291922 , n291920 , n291921 );
buf ( n291923 , n291922 );
buf ( n291924 , n291923 );
buf ( n291925 , n820 );
nand ( n1498 , n291919 , n291924 , n291925 );
buf ( n291927 , n1498 );
buf ( n291928 , n291927 );
not ( n291929 , n291928 );
xor ( n291930 , n828 , n791 );
buf ( n291931 , n291930 );
not ( n291932 , n291931 );
buf ( n291933 , n291808 );
not ( n1506 , n291933 );
or ( n1507 , n291932 , n1506 );
xor ( n1508 , n829 , n830 );
buf ( n291937 , n1508 );
buf ( n291938 , n291937 );
buf ( n291939 , n291938 );
buf ( n291940 , n291939 );
buf ( n291941 , n291794 );
nand ( n291942 , n291940 , n291941 );
buf ( n291943 , n291942 );
buf ( n291944 , n291943 );
nand ( n291945 , n1507 , n291944 );
buf ( n291946 , n291945 );
buf ( n291947 , n291946 );
not ( n291948 , n291947 );
or ( n1521 , n291929 , n291948 );
buf ( n291950 , n291946 );
buf ( n291951 , n291927 );
or ( n1524 , n291950 , n291951 );
nand ( n1525 , n1521 , n1524 );
buf ( n291954 , n1525 );
and ( n1527 , n291912 , n291954 );
and ( n291956 , n1469 , n291911 );
or ( n291957 , n1527 , n291956 );
buf ( n291958 , n291957 );
and ( n1531 , n291869 , n291958 );
and ( n291960 , n291864 , n291868 );
or ( n291961 , n1531 , n291960 );
buf ( n291962 , n291961 );
buf ( n291963 , n291962 );
xor ( n291964 , n291860 , n291963 );
not ( n291965 , n291739 );
not ( n291966 , n291722 );
or ( n1539 , n291965 , n291966 );
xor ( n291968 , n821 , n822 );
buf ( n291969 , n291968 );
buf ( n291970 , n291969 );
xor ( n1543 , n820 , n796 );
buf ( n291972 , n1543 );
nand ( n291973 , n291970 , n291972 );
buf ( n291974 , n291973 );
nand ( n291975 , n1539 , n291974 );
xor ( n1548 , n818 , n799 );
buf ( n291977 , n1548 );
not ( n1550 , n291977 );
xor ( n291979 , n818 , n819 );
nand ( n291980 , n1356 , n291979 );
not ( n1553 , n291980 );
buf ( n291982 , n1553 );
buf ( n291983 , n291982 );
buf ( n291984 , n291983 );
buf ( n291985 , n291984 );
not ( n291986 , n291985 );
or ( n1559 , n1550 , n291986 );
xor ( n291988 , n819 , n820 );
buf ( n291989 , n291988 );
buf ( n1562 , n291989 );
xor ( n291991 , n818 , n798 );
buf ( n291992 , n291991 );
nand ( n291993 , n1562 , n291992 );
buf ( n291994 , n291993 );
buf ( n291995 , n291994 );
nand ( n291996 , n1559 , n291995 );
buf ( n291997 , n291996 );
xor ( n1570 , n291975 , n291997 );
buf ( n291999 , n791 );
buf ( n1572 , n826 );
xor ( n1573 , n291999 , n1572 );
buf ( n292002 , n1573 );
not ( n292003 , n292002 );
not ( n1576 , n1453 );
or ( n292005 , n292003 , n1576 );
not ( n292006 , n1445 );
not ( n1579 , n292006 );
buf ( n1580 , n1579 );
buf ( n292009 , n1580 );
buf ( n1582 , n790 );
buf ( n292011 , n826 );
xor ( n292012 , n1582 , n292011 );
buf ( n292013 , n292012 );
buf ( n292014 , n292013 );
nand ( n1587 , n292009 , n292014 );
buf ( n292016 , n1587 );
nand ( n1589 , n292005 , n292016 );
xor ( n292018 , n1570 , n1589 );
buf ( n292019 , n292018 );
buf ( n292020 , n291769 );
not ( n292021 , n292020 );
buf ( n292022 , n291761 );
not ( n292023 , n292022 );
or ( n292024 , n292021 , n292023 );
xnor ( n1597 , n823 , n824 );
buf ( n292026 , n1597 );
not ( n1599 , n292026 );
buf ( n1600 , n1599 );
buf ( n1601 , n1600 );
xor ( n292030 , n822 , n794 );
buf ( n1603 , n292030 );
nand ( n1604 , n1601 , n1603 );
buf ( n1605 , n1604 );
buf ( n292034 , n1605 );
nand ( n292035 , n292024 , n292034 );
buf ( n292036 , n292035 );
buf ( n292037 , n292036 );
not ( n292038 , n291845 );
not ( n1611 , n291835 );
or ( n292040 , n292038 , n1611 );
xor ( n1613 , n825 , n826 );
buf ( n292042 , n1613 );
xor ( n1615 , n824 , n792 );
buf ( n292044 , n1615 );
nand ( n1617 , n292042 , n292044 );
buf ( n292046 , n1617 );
nand ( n1619 , n292040 , n292046 );
buf ( n292048 , n1619 );
xor ( n292049 , n292037 , n292048 );
buf ( n292050 , n291808 );
buf ( n292051 , n1389 );
nand ( n292052 , n292050 , n292051 );
buf ( n292053 , n292052 );
buf ( n292054 , n292053 );
buf ( n292055 , n291812 );
buf ( n292056 , n788 );
buf ( n292057 , n828 );
xor ( n1630 , n292056 , n292057 );
buf ( n292059 , n1630 );
buf ( n292060 , n292059 );
nand ( n1633 , n292055 , n292060 );
buf ( n292062 , n1633 );
buf ( n1635 , n292062 );
nand ( n1636 , n292054 , n1635 );
buf ( n1637 , n1636 );
buf ( n292066 , n1637 );
xor ( n1639 , n292049 , n292066 );
buf ( n292068 , n1639 );
buf ( n292069 , n292068 );
xor ( n292070 , n292019 , n292069 );
buf ( n292071 , n291891 );
not ( n292072 , n292071 );
buf ( n292073 , n1453 );
not ( n1646 , n292073 );
or ( n1647 , n292072 , n1646 );
buf ( n292076 , n291886 );
buf ( n292077 , n292002 );
nand ( n292078 , n292076 , n292077 );
buf ( n292079 , n292078 );
buf ( n292080 , n292079 );
nand ( n1653 , n1647 , n292080 );
buf ( n1654 , n1653 );
buf ( n292083 , n1654 );
buf ( n292084 , n291946 );
not ( n292085 , n292084 );
buf ( n1658 , n291927 );
nor ( n1659 , n292085 , n1658 );
buf ( n292088 , n1659 );
buf ( n292089 , n292088 );
xor ( n1662 , n292083 , n292089 );
not ( n292091 , n1271 );
buf ( n292092 , n789 );
buf ( n292093 , n830 );
xor ( n1666 , n292092 , n292093 );
buf ( n1667 , n1666 );
not ( n292096 , n1667 );
or ( n1669 , n292091 , n292096 );
buf ( n292098 , n1266 );
buf ( n292099 , n831 );
nand ( n1672 , n292098 , n292099 );
buf ( n292101 , n1672 );
nand ( n292102 , n1669 , n292101 );
not ( n1675 , n291748 );
buf ( n292104 , n291765 );
buf ( n292105 , n292104 );
not ( n1678 , n292105 );
or ( n292107 , n1675 , n1678 );
xor ( n292108 , n822 , n797 );
nand ( n292109 , n292108 , n291761 );
nand ( n292110 , n292107 , n292109 );
xor ( n1683 , n292102 , n292110 );
xor ( n292112 , n824 , n795 );
not ( n292113 , n292112 );
not ( n1686 , n291838 );
or ( n292115 , n292113 , n1686 );
buf ( n292116 , n291843 );
buf ( n292117 , n291826 );
nand ( n292118 , n292116 , n292117 );
buf ( n292119 , n292118 );
nand ( n1692 , n292115 , n292119 );
and ( n1693 , n1683 , n1692 );
and ( n1694 , n292102 , n292110 );
or ( n1695 , n1693 , n1694 );
buf ( n292124 , n1695 );
and ( n292125 , n1662 , n292124 );
and ( n1698 , n292083 , n292089 );
or ( n292127 , n292125 , n1698 );
buf ( n292128 , n292127 );
buf ( n292129 , n292128 );
xor ( n292130 , n292070 , n292129 );
buf ( n292131 , n292130 );
buf ( n292132 , n292131 );
and ( n1705 , n291964 , n292132 );
and ( n1706 , n291860 , n291963 );
or ( n1707 , n1705 , n1706 );
buf ( n292136 , n1707 );
buf ( n292137 , n292136 );
xor ( n1710 , n291648 , n292137 );
xor ( n1711 , n817 , n818 );
buf ( n1712 , n1711 );
buf ( n292141 , n1712 );
buf ( n292142 , n799 );
and ( n292143 , n292141 , n292142 );
buf ( n292144 , n292143 );
buf ( n292145 , n292144 );
buf ( n292146 , n291663 );
not ( n1719 , n292146 );
buf ( n292148 , n1271 );
not ( n1721 , n292148 );
or ( n292150 , n1719 , n1721 );
buf ( n292151 , n785 );
buf ( n292152 , n830 );
xor ( n292153 , n292151 , n292152 );
buf ( n292154 , n292153 );
buf ( n292155 , n292154 );
buf ( n292156 , n831 );
nand ( n1729 , n292155 , n292156 );
buf ( n292158 , n1729 );
buf ( n292159 , n292158 );
nand ( n1732 , n292150 , n292159 );
buf ( n292161 , n1732 );
buf ( n292162 , n292161 );
xor ( n1735 , n292145 , n292162 );
buf ( n292164 , n292059 );
not ( n1737 , n292164 );
buf ( n292166 , n291802 );
not ( n1739 , n292166 );
buf ( n292168 , n1739 );
buf ( n292169 , n292168 );
not ( n292170 , n292169 );
or ( n1743 , n1737 , n292170 );
buf ( n292172 , n291812 );
buf ( n292173 , n787 );
buf ( n292174 , n828 );
xor ( n292175 , n292173 , n292174 );
buf ( n292176 , n292175 );
buf ( n1749 , n292176 );
nand ( n1750 , n292172 , n1749 );
buf ( n1751 , n1750 );
buf ( n292180 , n1751 );
nand ( n1753 , n1743 , n292180 );
buf ( n292182 , n1753 );
buf ( n292183 , n292182 );
xor ( n1756 , n1735 , n292183 );
buf ( n292185 , n1756 );
buf ( n1758 , n292185 );
buf ( n292187 , n1589 );
not ( n1760 , n292187 );
buf ( n292189 , n291739 );
not ( n292190 , n292189 );
buf ( n292191 , n291722 );
not ( n292192 , n292191 );
or ( n292193 , n292190 , n292192 );
buf ( n292194 , n291974 );
nand ( n292195 , n292193 , n292194 );
buf ( n292196 , n292195 );
buf ( n292197 , n292196 );
not ( n1770 , n292197 );
or ( n292199 , n1760 , n1770 );
or ( n1772 , n1589 , n292196 );
nand ( n1773 , n1772 , n291997 );
buf ( n292202 , n1773 );
nand ( n1775 , n292199 , n292202 );
buf ( n292204 , n1775 );
buf ( n292205 , n292204 );
xor ( n1778 , n1758 , n292205 );
xor ( n1779 , n292037 , n292048 );
and ( n1780 , n1779 , n292066 );
and ( n292209 , n292037 , n292048 );
or ( n1782 , n1780 , n292209 );
buf ( n292211 , n1782 );
buf ( n292212 , n292211 );
xor ( n292213 , n1778 , n292212 );
buf ( n292214 , n292213 );
buf ( n292215 , n292214 );
xor ( n1788 , n292019 , n292069 );
and ( n1789 , n1788 , n292129 );
and ( n1790 , n292019 , n292069 );
or ( n292219 , n1789 , n1790 );
buf ( n292220 , n292219 );
buf ( n292221 , n292220 );
xor ( n1794 , n292215 , n292221 );
buf ( n292223 , n291670 );
buf ( n292224 , n291686 );
and ( n1797 , n292223 , n292224 );
buf ( n292226 , n1797 );
buf ( n1799 , n292226 );
buf ( n292228 , n291991 );
not ( n1801 , n292228 );
buf ( n292230 , n291984 );
not ( n292231 , n292230 );
or ( n292232 , n1801 , n292231 );
buf ( n292233 , n291989 );
buf ( n292234 , n797 );
buf ( n292235 , n818 );
xor ( n292236 , n292234 , n292235 );
buf ( n292237 , n292236 );
buf ( n292238 , n292237 );
nand ( n292239 , n292233 , n292238 );
buf ( n292240 , n292239 );
buf ( n292241 , n292240 );
nand ( n292242 , n292232 , n292241 );
buf ( n292243 , n292242 );
buf ( n292244 , n292243 );
xor ( n1817 , n1799 , n292244 );
buf ( n292246 , n1543 );
not ( n1819 , n292246 );
buf ( n292248 , n291903 );
not ( n292249 , n292248 );
or ( n292250 , n1819 , n292249 );
buf ( n292251 , n291969 );
buf ( n292252 , n795 );
buf ( n292253 , n820 );
xor ( n1826 , n292252 , n292253 );
buf ( n292255 , n1826 );
buf ( n292256 , n292255 );
nand ( n1829 , n292251 , n292256 );
buf ( n292258 , n1829 );
buf ( n292259 , n292258 );
nand ( n1832 , n292250 , n292259 );
buf ( n292261 , n1832 );
buf ( n292262 , n292261 );
xor ( n1835 , n1817 , n292262 );
buf ( n292264 , n1835 );
buf ( n292265 , n292264 );
not ( n1838 , n292013 );
not ( n292267 , n291880 );
or ( n1840 , n1838 , n292267 );
buf ( n292269 , n291886 );
buf ( n1842 , n789 );
buf ( n292271 , n826 );
xor ( n292272 , n1842 , n292271 );
buf ( n292273 , n292272 );
buf ( n292274 , n292273 );
nand ( n1847 , n292269 , n292274 );
buf ( n292276 , n1847 );
nand ( n292277 , n1840 , n292276 );
not ( n1850 , n292277 );
buf ( n292279 , n1613 );
buf ( n1852 , n791 );
buf ( n292281 , n824 );
xor ( n292282 , n1852 , n292281 );
buf ( n292283 , n292282 );
buf ( n292284 , n292283 );
nand ( n292285 , n292279 , n292284 );
buf ( n292286 , n292285 );
nand ( n292287 , n1615 , n291835 );
and ( n292288 , n292286 , n292287 );
not ( n1861 , n292288 );
and ( n292290 , n1850 , n1861 );
and ( n292291 , n292288 , n292277 );
nor ( n1864 , n292290 , n292291 );
not ( n292293 , n1864 );
not ( n1866 , n292030 );
not ( n1867 , n291761 );
or ( n1868 , n1866 , n1867 );
buf ( n292297 , n292105 );
buf ( n292298 , n793 );
buf ( n292299 , n822 );
xor ( n292300 , n292298 , n292299 );
buf ( n292301 , n292300 );
buf ( n292302 , n292301 );
nand ( n292303 , n292297 , n292302 );
buf ( n292304 , n292303 );
nand ( n1877 , n1868 , n292304 );
not ( n292306 , n1877 );
nand ( n292307 , n292293 , n292306 );
nand ( n1880 , n1877 , n1864 );
nand ( n292309 , n292307 , n1880 );
buf ( n292310 , n292309 );
xor ( n292311 , n292265 , n292310 );
xor ( n292312 , n291690 , n291781 );
and ( n292313 , n292312 , n291857 );
and ( n292314 , n291690 , n291781 );
or ( n1887 , n292313 , n292314 );
buf ( n292316 , n1887 );
buf ( n292317 , n292316 );
xor ( n292318 , n292311 , n292317 );
buf ( n292319 , n292318 );
buf ( n292320 , n292319 );
xor ( n292321 , n1794 , n292320 );
buf ( n292322 , n292321 );
buf ( n292323 , n292322 );
and ( n1896 , n1710 , n292323 );
and ( n292325 , n291648 , n292137 );
or ( n292326 , n1896 , n292325 );
buf ( n292327 , n292326 );
not ( n1900 , n292327 );
or ( n1901 , n291647 , n1900 );
buf ( n292330 , n831 );
not ( n1903 , n292330 );
buf ( n292332 , n881 );
buf ( n292333 , n292136 );
xor ( n292334 , n292332 , n292333 );
buf ( n292335 , n292322 );
and ( n292336 , n292334 , n292335 );
and ( n292337 , n292332 , n292333 );
or ( n1910 , n292336 , n292337 );
buf ( n292339 , n1910 );
buf ( n1912 , n292339 );
nand ( n1913 , n1903 , n1912 );
buf ( n1914 , n1913 );
nand ( n292343 , n1901 , n1914 );
buf ( n1916 , n292343 );
buf ( n292345 , n831 );
not ( n292346 , n292345 );
buf ( n292347 , n841 );
or ( n292348 , n799 , n813 );
nand ( n292349 , n292348 , n814 );
buf ( n292350 , n292349 );
buf ( n292351 , n799 );
buf ( n292352 , n813 );
nand ( n1925 , n292351 , n292352 );
buf ( n292354 , n1925 );
buf ( n292355 , n292354 );
buf ( n292356 , n812 );
nand ( n292357 , n292350 , n292355 , n292356 );
buf ( n292358 , n292357 );
buf ( n292359 , n292358 );
not ( n292360 , n292359 );
and ( n1933 , n291697 , n830 );
not ( n1934 , n1933 );
and ( n292363 , n781 , n830 );
not ( n1936 , n781 );
buf ( n292365 , n830 );
not ( n292366 , n292365 );
buf ( n292367 , n292366 );
and ( n292368 , n1936 , n292367 );
nor ( n292369 , n292363 , n292368 );
not ( n292370 , n292369 );
or ( n292371 , n1934 , n292370 );
buf ( n292372 , n780 );
buf ( n292373 , n830 );
xor ( n292374 , n292372 , n292373 );
buf ( n292375 , n292374 );
buf ( n292376 , n292375 );
buf ( n292377 , n831 );
nand ( n1950 , n292376 , n292377 );
buf ( n1951 , n1950 );
nand ( n292380 , n292371 , n1951 );
buf ( n292381 , n292380 );
nand ( n292382 , n292360 , n292381 );
buf ( n292383 , n292382 );
buf ( n292384 , n292383 );
xor ( n292385 , n818 , n792 );
buf ( n1958 , n292385 );
not ( n1959 , n1958 );
not ( n1960 , n291979 );
xor ( n1961 , n819 , n820 );
nor ( n1962 , n1960 , n1961 );
buf ( n292391 , n1962 );
buf ( n1964 , n292391 );
buf ( n292393 , n1964 );
buf ( n1966 , n292393 );
not ( n1967 , n1966 );
or ( n1968 , n1959 , n1967 );
buf ( n1969 , n291788 );
buf ( n292398 , n791 );
buf ( n292399 , n818 );
xor ( n292400 , n292398 , n292399 );
buf ( n292401 , n292400 );
buf ( n292402 , n292401 );
nand ( n292403 , n1969 , n292402 );
buf ( n292404 , n292403 );
buf ( n292405 , n292404 );
nand ( n1978 , n1968 , n292405 );
buf ( n292407 , n1978 );
buf ( n292408 , n292407 );
not ( n292409 , n292408 );
buf ( n292410 , n292409 );
buf ( n292411 , n292410 );
xor ( n292412 , n292384 , n292411 );
buf ( n292413 , n790 );
buf ( n292414 , n820 );
xor ( n292415 , n292413 , n292414 );
buf ( n292416 , n292415 );
buf ( n292417 , n292416 );
not ( n292418 , n292417 );
buf ( n292419 , n291722 );
not ( n1992 , n292419 );
or ( n292421 , n292418 , n1992 );
not ( n292422 , n291968 );
not ( n1995 , n292422 );
buf ( n292424 , n1995 );
buf ( n1997 , n789 );
buf ( n1998 , n820 );
xor ( n1999 , n1997 , n1998 );
buf ( n292428 , n1999 );
buf ( n292429 , n292428 );
nand ( n292430 , n292424 , n292429 );
buf ( n292431 , n292430 );
buf ( n292432 , n292431 );
nand ( n292433 , n292421 , n292432 );
buf ( n292434 , n292433 );
buf ( n292435 , n292434 );
xor ( n292436 , n292412 , n292435 );
buf ( n292437 , n292436 );
buf ( n292438 , n292437 );
not ( n292439 , n292358 );
and ( n292440 , n292380 , n292439 );
not ( n292441 , n292380 );
and ( n2014 , n292441 , n292358 );
nor ( n292443 , n292440 , n2014 );
not ( n292444 , n292443 );
not ( n2017 , n292444 );
not ( n292446 , n2017 );
not ( n292447 , n292369 );
not ( n2020 , n831 );
or ( n292449 , n292447 , n2020 );
xor ( n292450 , n830 , n782 );
nand ( n2023 , n292450 , n1271 );
nand ( n292452 , n292449 , n2023 );
not ( n292453 , n292452 );
xor ( n2026 , n814 , n813 );
nand ( n292455 , n2026 , n799 );
nand ( n292456 , n292453 , n292455 );
not ( n2029 , n292456 );
buf ( n292458 , n788 );
buf ( n292459 , n824 );
xor ( n2032 , n292458 , n292459 );
buf ( n292461 , n2032 );
not ( n2034 , n292461 );
not ( n292463 , n826 );
nand ( n292464 , n292463 , n825 );
not ( n2037 , n824 );
not ( n2038 , n825 );
not ( n292467 , n2038 );
or ( n292468 , n2037 , n292467 );
not ( n2041 , n824 );
nand ( n292470 , n2041 , n825 );
nand ( n292471 , n292468 , n292470 );
nand ( n2044 , n292464 , n1402 , n292471 );
not ( n292473 , n2044 );
not ( n2046 , n292473 );
or ( n2047 , n2034 , n2046 );
buf ( n2048 , n291843 );
buf ( n292477 , n787 );
buf ( n292478 , n824 );
xor ( n292479 , n292477 , n292478 );
buf ( n292480 , n292479 );
buf ( n292481 , n292480 );
nand ( n292482 , n2048 , n292481 );
buf ( n292483 , n292482 );
nand ( n292484 , n2047 , n292483 );
not ( n292485 , n292484 );
or ( n2058 , n2029 , n292485 );
not ( n292487 , n292455 );
not ( n292488 , n292453 );
nand ( n2061 , n292487 , n292488 );
nand ( n2062 , n2058 , n2061 );
not ( n2063 , n2062 );
or ( n2064 , n292446 , n2063 );
not ( n2065 , n292444 );
not ( n2066 , n2062 );
not ( n292495 , n2066 );
or ( n2068 , n2065 , n292495 );
buf ( n292497 , n798 );
buf ( n292498 , n814 );
xor ( n292499 , n292497 , n292498 );
buf ( n292500 , n292499 );
not ( n292501 , n292500 );
xor ( n292502 , n815 , n816 );
not ( n2075 , n292502 );
xor ( n292504 , n814 , n815 );
nand ( n292505 , n2075 , n292504 );
not ( n2078 , n292505 );
buf ( n2079 , n2078 );
buf ( n292508 , n2079 );
buf ( n292509 , n292508 );
not ( n292510 , n292509 );
or ( n292511 , n292501 , n292510 );
and ( n2084 , n816 , n815 );
not ( n2085 , n816 );
not ( n2086 , n815 );
and ( n2087 , n2085 , n2086 );
nor ( n2088 , n2084 , n2087 );
buf ( n2089 , n2088 );
buf ( n292518 , n2089 );
buf ( n292519 , n292518 );
buf ( n292520 , n797 );
buf ( n292521 , n814 );
xor ( n292522 , n292520 , n292521 );
buf ( n292523 , n292522 );
buf ( n292524 , n292523 );
nand ( n2097 , n292519 , n292524 );
buf ( n292526 , n2097 );
nand ( n292527 , n292511 , n292526 );
not ( n2100 , n292527 );
xor ( n292529 , n816 , n796 );
not ( n292530 , n292529 );
not ( n2103 , n817 );
nand ( n2104 , n2103 , n816 );
not ( n292533 , n2104 );
not ( n2106 , n816 );
nand ( n292535 , n2106 , n817 );
not ( n292536 , n292535 );
or ( n2109 , n292533 , n292536 );
not ( n292538 , n818 );
and ( n292539 , n817 , n292538 );
not ( n2112 , n817 );
and ( n292541 , n2112 , n818 );
nor ( n292542 , n292539 , n292541 );
nand ( n292543 , n2109 , n292542 );
buf ( n292544 , n292543 );
not ( n2117 , n292544 );
buf ( n2118 , n2117 );
not ( n292547 , n2118 );
or ( n2120 , n292530 , n292547 );
buf ( n292549 , n1712 );
buf ( n292550 , n795 );
buf ( n292551 , n816 );
xor ( n292552 , n292550 , n292551 );
buf ( n292553 , n292552 );
buf ( n292554 , n292553 );
nand ( n2127 , n292549 , n292554 );
buf ( n292556 , n2127 );
nand ( n292557 , n2120 , n292556 );
buf ( n292558 , n784 );
buf ( n292559 , n828 );
xor ( n292560 , n292558 , n292559 );
buf ( n292561 , n292560 );
not ( n2134 , n292561 );
not ( n292563 , n292168 );
or ( n292564 , n2134 , n292563 );
buf ( n292565 , n291812 );
buf ( n292566 , n783 );
buf ( n292567 , n828 );
xor ( n2140 , n292566 , n292567 );
buf ( n2141 , n2140 );
buf ( n2142 , n2141 );
nand ( n2143 , n292565 , n2142 );
buf ( n292572 , n2143 );
nand ( n2145 , n292564 , n292572 );
or ( n2146 , n292557 , n2145 );
not ( n2147 , n2146 );
or ( n292576 , n2100 , n2147 );
nand ( n292577 , n2145 , n292557 );
nand ( n2150 , n292576 , n292577 );
nand ( n292579 , n2068 , n2150 );
nand ( n2152 , n2064 , n292579 );
buf ( n292581 , n2152 );
xor ( n2154 , n292438 , n292581 );
xor ( n2155 , n820 , n792 );
buf ( n292584 , n2155 );
not ( n2157 , n292584 );
buf ( n292586 , n291722 );
not ( n2159 , n292586 );
or ( n2160 , n2157 , n2159 );
buf ( n292589 , n1995 );
buf ( n2162 , n791 );
buf ( n292591 , n820 );
xor ( n292592 , n2162 , n292591 );
buf ( n292593 , n292592 );
buf ( n292594 , n292593 );
nand ( n292595 , n292589 , n292594 );
buf ( n292596 , n292595 );
buf ( n292597 , n292596 );
nand ( n2170 , n2160 , n292597 );
buf ( n292599 , n2170 );
buf ( n292600 , n786 );
buf ( n292601 , n826 );
xor ( n292602 , n292600 , n292601 );
buf ( n292603 , n292602 );
not ( n292604 , n292603 );
not ( n2177 , n291880 );
or ( n292606 , n292604 , n2177 );
buf ( n292607 , n1579 );
buf ( n292608 , n785 );
buf ( n292609 , n826 );
xor ( n2182 , n292608 , n292609 );
buf ( n292611 , n2182 );
buf ( n292612 , n292611 );
nand ( n2185 , n292607 , n292612 );
buf ( n292614 , n2185 );
nand ( n2187 , n292606 , n292614 );
nand ( n292616 , n292599 , n2187 );
buf ( n292617 , n2155 );
not ( n2190 , n292617 );
buf ( n292619 , n291722 );
not ( n292620 , n292619 );
or ( n292621 , n2190 , n292620 );
buf ( n292622 , n292596 );
nand ( n292623 , n292621 , n292622 );
buf ( n292624 , n292623 );
or ( n2197 , n292624 , n2187 );
xor ( n292626 , n822 , n790 );
buf ( n292627 , n292626 );
not ( n2200 , n292627 );
buf ( n292629 , n1330 );
not ( n2202 , n292629 );
buf ( n292631 , n2202 );
buf ( n292632 , n292631 );
not ( n292633 , n292632 );
or ( n2206 , n2200 , n292633 );
buf ( n292635 , n292105 );
buf ( n292636 , n789 );
buf ( n292637 , n822 );
xor ( n292638 , n292636 , n292637 );
buf ( n292639 , n292638 );
buf ( n292640 , n292639 );
nand ( n2213 , n292635 , n292640 );
buf ( n292642 , n2213 );
buf ( n292643 , n292642 );
nand ( n292644 , n2206 , n292643 );
buf ( n292645 , n292644 );
nand ( n292646 , n2197 , n292645 );
nand ( n2219 , n292616 , n292646 );
not ( n2220 , n2219 );
xor ( n292649 , n818 , n793 );
not ( n2222 , n292649 );
not ( n292651 , n1553 );
or ( n292652 , n2222 , n292651 );
buf ( n292653 , n291988 );
buf ( n292654 , n292385 );
nand ( n292655 , n292653 , n292654 );
buf ( n292656 , n292655 );
nand ( n292657 , n292652 , n292656 );
buf ( n292658 , n292593 );
not ( n2231 , n292658 );
and ( n292660 , n821 , n822 );
not ( n292661 , n821 );
not ( n2234 , n822 );
and ( n292663 , n292661 , n2234 );
nor ( n292664 , n292660 , n292663 );
not ( n2237 , n292664 );
xor ( n2238 , n820 , n821 );
nand ( n292667 , n2237 , n2238 );
not ( n292668 , n292667 );
buf ( n292669 , n292668 );
not ( n292670 , n292669 );
or ( n292671 , n2231 , n292670 );
nand ( n292672 , n292416 , n291714 );
buf ( n292673 , n292672 );
nand ( n292674 , n292671 , n292673 );
buf ( n292675 , n292674 );
xor ( n2248 , n292657 , n292675 );
not ( n292677 , n292611 );
not ( n2250 , n291880 );
or ( n292679 , n292677 , n2250 );
buf ( n292680 , n1579 );
buf ( n292681 , n784 );
buf ( n292682 , n826 );
xor ( n292683 , n292681 , n292682 );
buf ( n292684 , n292683 );
buf ( n292685 , n292684 );
nand ( n292686 , n292680 , n292685 );
buf ( n292687 , n292686 );
nand ( n2260 , n292679 , n292687 );
xor ( n2261 , n2248 , n2260 );
not ( n2262 , n2261 );
nand ( n2263 , n2220 , n2262 );
not ( n2264 , n2263 );
buf ( n292693 , n292553 );
not ( n2266 , n292693 );
buf ( n292695 , n2118 );
not ( n292696 , n292695 );
or ( n2269 , n2266 , n292696 );
buf ( n292698 , n1711 );
not ( n292699 , n292698 );
buf ( n292700 , n292699 );
not ( n292701 , n292700 );
xor ( n2274 , n816 , n794 );
nand ( n292703 , n292701 , n2274 );
buf ( n292704 , n292703 );
nand ( n2277 , n2269 , n292704 );
buf ( n2278 , n2277 );
nand ( n292707 , n291835 , n292480 );
xor ( n2280 , n824 , n786 );
buf ( n292709 , n2280 );
buf ( n292710 , n1613 );
nand ( n2283 , n292709 , n292710 );
buf ( n2284 , n2283 );
and ( n292713 , n292707 , n2284 );
xor ( n292714 , n2278 , n292713 );
buf ( n292715 , n292523 );
not ( n292716 , n292715 );
not ( n2289 , n292502 );
xor ( n292718 , n814 , n815 );
and ( n292719 , n2289 , n292718 );
buf ( n292720 , n292719 );
not ( n292721 , n292720 );
or ( n292722 , n292716 , n292721 );
buf ( n2295 , n2089 );
buf ( n292724 , n2295 );
buf ( n292725 , n292724 );
buf ( n292726 , n292725 );
buf ( n292727 , n796 );
buf ( n292728 , n814 );
xor ( n292729 , n292727 , n292728 );
buf ( n292730 , n292729 );
buf ( n292731 , n292730 );
nand ( n292732 , n292726 , n292731 );
buf ( n292733 , n292732 );
buf ( n292734 , n292733 );
nand ( n292735 , n292722 , n292734 );
buf ( n292736 , n292735 );
and ( n2309 , n292714 , n292736 );
not ( n292738 , n292714 );
buf ( n292739 , n292736 );
not ( n2312 , n292739 );
buf ( n292741 , n2312 );
and ( n292742 , n292738 , n292741 );
nor ( n2315 , n2309 , n292742 );
not ( n292744 , n2315 );
not ( n292745 , n292744 );
or ( n2318 , n2264 , n292745 );
nand ( n292747 , n2219 , n2261 );
nand ( n292748 , n2318 , n292747 );
buf ( n292749 , n292748 );
and ( n292750 , n2154 , n292749 );
and ( n292751 , n292438 , n292581 );
or ( n2324 , n292750 , n292751 );
buf ( n292753 , n2324 );
buf ( n292754 , n292753 );
buf ( n292755 , n292639 );
not ( n2328 , n292755 );
buf ( n292757 , n292631 );
not ( n2330 , n292757 );
or ( n292759 , n2328 , n2330 );
buf ( n2332 , n292104 );
buf ( n2333 , n788 );
buf ( n2334 , n822 );
xor ( n2335 , n2333 , n2334 );
buf ( n292764 , n2335 );
buf ( n2337 , n292764 );
nand ( n2338 , n2332 , n2337 );
buf ( n2339 , n2338 );
buf ( n2340 , n2339 );
nand ( n2341 , n292759 , n2340 );
buf ( n2342 , n2341 );
not ( n292771 , n2342 );
buf ( n292772 , n2141 );
not ( n2345 , n292772 );
buf ( n292774 , n292168 );
not ( n2347 , n292774 );
or ( n292776 , n2345 , n2347 );
buf ( n292777 , n291939 );
buf ( n292778 , n782 );
buf ( n292779 , n828 );
xor ( n2352 , n292778 , n292779 );
buf ( n2353 , n2352 );
buf ( n292782 , n2353 );
nand ( n2355 , n292777 , n292782 );
buf ( n292784 , n2355 );
buf ( n292785 , n292784 );
nand ( n2358 , n292776 , n292785 );
buf ( n292787 , n2358 );
not ( n2360 , n292787 );
or ( n2361 , n292771 , n2360 );
buf ( n2362 , n2342 );
buf ( n292791 , n292787 );
nor ( n292792 , n2362 , n292791 );
buf ( n292793 , n292792 );
xor ( n2366 , n814 , n813 );
not ( n2367 , n812 );
and ( n2368 , n813 , n2367 );
not ( n292797 , n813 );
and ( n2370 , n292797 , n812 );
nor ( n292799 , n2368 , n2370 );
nor ( n2372 , n2366 , n292799 );
buf ( n2373 , n2372 );
buf ( n292802 , n2373 );
buf ( n2375 , n292802 );
buf ( n2376 , n2375 );
buf ( n292805 , n2376 );
xor ( n2378 , n812 , n799 );
buf ( n292807 , n2378 );
and ( n292808 , n292805 , n292807 );
not ( n2381 , n2366 );
not ( n292810 , n2381 );
buf ( n2383 , n292810 );
buf ( n292812 , n2383 );
xor ( n292813 , n812 , n798 );
buf ( n292814 , n292813 );
and ( n292815 , n292812 , n292814 );
nor ( n2388 , n292808 , n292815 );
buf ( n292817 , n2388 );
or ( n292818 , n292793 , n292817 );
nand ( n292819 , n2361 , n292818 );
buf ( n292820 , n292819 );
xor ( n2393 , n292657 , n292675 );
and ( n292822 , n2393 , n2260 );
and ( n292823 , n292657 , n292675 );
or ( n2396 , n292822 , n292823 );
buf ( n292825 , n2396 );
xor ( n292826 , n292820 , n292825 );
not ( n292827 , n2278 );
not ( n2400 , n292713 );
not ( n2401 , n2400 );
or ( n292830 , n292827 , n2401 );
nor ( n292831 , n2278 , n2400 );
or ( n2404 , n292831 , n292741 );
nand ( n2405 , n292830 , n2404 );
buf ( n292834 , n2405 );
xor ( n292835 , n292826 , n292834 );
buf ( n292836 , n292835 );
buf ( n292837 , n292836 );
xor ( n2410 , n811 , n812 );
buf ( n292839 , n2410 );
buf ( n2412 , n292839 );
buf ( n292841 , n2412 );
buf ( n2414 , n292841 );
buf ( n292843 , n799 );
and ( n292844 , n2414 , n292843 );
buf ( n292845 , n292844 );
buf ( n292846 , n292845 );
buf ( n292847 , n292375 );
not ( n2420 , n292847 );
buf ( n292849 , n291656 );
not ( n2422 , n292849 );
or ( n292851 , n2420 , n2422 );
buf ( n292852 , n779 );
buf ( n292853 , n830 );
xor ( n292854 , n292852 , n292853 );
buf ( n292855 , n292854 );
buf ( n292856 , n292855 );
buf ( n292857 , n831 );
nand ( n292858 , n292856 , n292857 );
buf ( n292859 , n292858 );
buf ( n292860 , n292859 );
nand ( n292861 , n292851 , n292860 );
buf ( n292862 , n292861 );
buf ( n292863 , n292862 );
xor ( n292864 , n292846 , n292863 );
buf ( n292865 , n2280 );
not ( n2438 , n292865 );
buf ( n292867 , n291838 );
not ( n292868 , n292867 );
or ( n2441 , n2438 , n292868 );
buf ( n292870 , n1613 );
buf ( n292871 , n292870 );
xor ( n292872 , n824 , n785 );
buf ( n292873 , n292872 );
nand ( n2446 , n292871 , n292873 );
buf ( n292875 , n2446 );
buf ( n292876 , n292875 );
nand ( n292877 , n2441 , n292876 );
buf ( n292878 , n292877 );
buf ( n292879 , n292878 );
xor ( n292880 , n292864 , n292879 );
buf ( n292881 , n292880 );
buf ( n292882 , n292881 );
buf ( n292883 , n2274 );
not ( n2456 , n292883 );
not ( n292885 , n816 );
nand ( n292886 , n292885 , n817 );
not ( n2459 , n292886 );
not ( n292888 , n2104 );
or ( n292889 , n2459 , n292888 );
xnor ( n2462 , n817 , n818 );
nand ( n292891 , n292889 , n2462 );
not ( n292892 , n292891 );
buf ( n292893 , n292892 );
not ( n292894 , n292893 );
or ( n2467 , n2456 , n292894 );
buf ( n292896 , n1712 );
buf ( n292897 , n793 );
buf ( n292898 , n816 );
xor ( n292899 , n292897 , n292898 );
buf ( n292900 , n292899 );
buf ( n292901 , n292900 );
nand ( n2474 , n292896 , n292901 );
buf ( n292903 , n2474 );
buf ( n292904 , n292903 );
nand ( n292905 , n2467 , n292904 );
buf ( n292906 , n292905 );
not ( n292907 , n292906 );
not ( n2480 , n292907 );
not ( n292909 , n292730 );
not ( n2482 , n2078 );
or ( n292911 , n292909 , n2482 );
buf ( n292912 , n292725 );
buf ( n292913 , n795 );
buf ( n292914 , n814 );
xor ( n292915 , n292913 , n292914 );
buf ( n292916 , n292915 );
buf ( n292917 , n292916 );
nand ( n292918 , n292912 , n292917 );
buf ( n292919 , n292918 );
nand ( n292920 , n292911 , n292919 );
not ( n292921 , n292920 );
not ( n292922 , n292921 );
or ( n292923 , n2480 , n292922 );
nand ( n2496 , n292920 , n292906 );
nand ( n292925 , n292923 , n2496 );
buf ( n292926 , n2353 );
not ( n2499 , n292926 );
buf ( n292928 , n291805 );
not ( n292929 , n292928 );
or ( n2502 , n2499 , n292929 );
buf ( n292931 , n291812 );
buf ( n2504 , n781 );
buf ( n292933 , n828 );
xor ( n2506 , n2504 , n292933 );
buf ( n292935 , n2506 );
buf ( n292936 , n292935 );
nand ( n2509 , n292931 , n292936 );
buf ( n292938 , n2509 );
buf ( n292939 , n292938 );
nand ( n2512 , n2502 , n292939 );
buf ( n2513 , n2512 );
buf ( n292942 , n2513 );
not ( n2515 , n292942 );
buf ( n2516 , n2515 );
and ( n292945 , n292925 , n2516 );
not ( n2518 , n292925 );
and ( n292947 , n2518 , n2513 );
nor ( n2520 , n292945 , n292947 );
buf ( n292949 , n2520 );
xor ( n2522 , n292882 , n292949 );
buf ( n292951 , n292764 );
not ( n292952 , n292951 );
buf ( n292953 , n291761 );
not ( n292954 , n292953 );
or ( n292955 , n292952 , n292954 );
buf ( n292956 , n1600 );
xor ( n2529 , n822 , n787 );
buf ( n292958 , n2529 );
nand ( n2531 , n292956 , n292958 );
buf ( n2532 , n2531 );
buf ( n292961 , n2532 );
nand ( n2534 , n292955 , n292961 );
buf ( n2535 , n2534 );
buf ( n292964 , n292813 );
not ( n292965 , n292964 );
buf ( n292966 , n2376 );
not ( n2539 , n292966 );
or ( n292968 , n292965 , n2539 );
buf ( n292969 , n2383 );
buf ( n292970 , n797 );
buf ( n292971 , n812 );
xor ( n292972 , n292970 , n292971 );
buf ( n292973 , n292972 );
buf ( n292974 , n292973 );
nand ( n292975 , n292969 , n292974 );
buf ( n292976 , n292975 );
buf ( n292977 , n292976 );
nand ( n292978 , n292968 , n292977 );
buf ( n292979 , n292978 );
xor ( n292980 , n2535 , n292979 );
buf ( n292981 , n783 );
buf ( n292982 , n826 );
xor ( n2555 , n292981 , n292982 );
buf ( n292984 , n2555 );
buf ( n292985 , n292984 );
not ( n292986 , n292985 );
buf ( n292987 , n291886 );
not ( n292988 , n292987 );
or ( n292989 , n292986 , n292988 );
buf ( n292990 , n1453 );
buf ( n292991 , n292684 );
nand ( n292992 , n292990 , n292991 );
buf ( n292993 , n292992 );
buf ( n292994 , n292993 );
nand ( n2567 , n292989 , n292994 );
buf ( n292996 , n2567 );
xor ( n292997 , n292980 , n292996 );
buf ( n292998 , n292997 );
xor ( n292999 , n2522 , n292998 );
buf ( n293000 , n292999 );
buf ( n293001 , n293000 );
xor ( n293002 , n292837 , n293001 );
xor ( n2575 , n292438 , n292581 );
xor ( n2576 , n2575 , n292749 );
buf ( n293005 , n2576 );
buf ( n293006 , n293005 );
and ( n2579 , n293002 , n293006 );
and ( n2580 , n292837 , n293001 );
or ( n293009 , n2579 , n2580 );
buf ( n293010 , n293009 );
buf ( n2583 , n293010 );
xor ( n2584 , n292754 , n2583 );
xor ( n293013 , n292882 , n292949 );
and ( n293014 , n293013 , n292998 );
and ( n2587 , n292882 , n292949 );
or ( n293016 , n293014 , n2587 );
buf ( n293017 , n293016 );
buf ( n293018 , n293017 );
buf ( n293019 , n292383 );
not ( n293020 , n293019 );
buf ( n293021 , n292410 );
not ( n2594 , n293021 );
or ( n293023 , n293020 , n2594 );
buf ( n293024 , n292434 );
nand ( n2597 , n293023 , n293024 );
buf ( n293026 , n2597 );
buf ( n293027 , n293026 );
buf ( n293028 , n292383 );
not ( n2601 , n293028 );
buf ( n293030 , n292407 );
nand ( n293031 , n2601 , n293030 );
buf ( n293032 , n293031 );
buf ( n293033 , n293032 );
nand ( n293034 , n293027 , n293033 );
buf ( n293035 , n293034 );
buf ( n293036 , n293035 );
not ( n2609 , n2529 );
not ( n293038 , n292631 );
or ( n2611 , n2609 , n293038 );
buf ( n293040 , n292105 );
buf ( n293041 , n786 );
buf ( n293042 , n822 );
xor ( n2615 , n293041 , n293042 );
buf ( n293044 , n2615 );
buf ( n293045 , n293044 );
nand ( n293046 , n293040 , n293045 );
buf ( n293047 , n293046 );
nand ( n2620 , n2611 , n293047 );
xor ( n293049 , n810 , n799 );
not ( n293050 , n293049 );
xnor ( n293051 , n810 , n811 );
buf ( n293052 , n293051 );
buf ( n293053 , n2410 );
nor ( n293054 , n293052 , n293053 );
buf ( n293055 , n293054 );
buf ( n293056 , n293055 );
buf ( n293057 , n293056 );
buf ( n293058 , n293057 );
not ( n2631 , n293058 );
or ( n293060 , n293050 , n2631 );
buf ( n293061 , n292841 );
xor ( n2634 , n810 , n798 );
buf ( n293063 , n2634 );
nand ( n293064 , n293061 , n293063 );
buf ( n293065 , n293064 );
nand ( n2638 , n293060 , n293065 );
xor ( n293067 , n2620 , n2638 );
buf ( n293068 , n292973 );
not ( n293069 , n293068 );
buf ( n2642 , n2376 );
not ( n2643 , n2642 );
or ( n2644 , n293069 , n2643 );
buf ( n2645 , n2383 );
xor ( n2646 , n812 , n796 );
buf ( n293075 , n2646 );
nand ( n293076 , n2645 , n293075 );
buf ( n293077 , n293076 );
buf ( n293078 , n293077 );
nand ( n2651 , n2644 , n293078 );
buf ( n2652 , n2651 );
xor ( n293081 , n293067 , n2652 );
buf ( n293082 , n293081 );
xor ( n293083 , n293036 , n293082 );
xor ( n293084 , n824 , n784 );
and ( n293085 , n292870 , n293084 );
and ( n2658 , n291838 , n292872 );
nor ( n293087 , n293085 , n2658 );
not ( n2660 , n293087 );
not ( n2661 , n292900 );
not ( n293090 , n2118 );
or ( n293091 , n2661 , n293090 );
buf ( n293092 , n1712 );
xor ( n293093 , n816 , n792 );
buf ( n293094 , n293093 );
nand ( n2667 , n293092 , n293094 );
buf ( n2668 , n2667 );
nand ( n293097 , n293091 , n2668 );
not ( n2670 , n293097 );
xor ( n2671 , n2660 , n2670 );
buf ( n293100 , n292916 );
not ( n2673 , n293100 );
buf ( n293102 , n292719 );
not ( n2675 , n293102 );
or ( n293104 , n2673 , n2675 );
buf ( n293105 , n292725 );
buf ( n293106 , n794 );
buf ( n293107 , n814 );
xor ( n2680 , n293106 , n293107 );
buf ( n2681 , n2680 );
buf ( n293110 , n2681 );
nand ( n2683 , n293105 , n293110 );
buf ( n2684 , n2683 );
buf ( n293113 , n2684 );
nand ( n2686 , n293104 , n293113 );
buf ( n293115 , n2686 );
not ( n2688 , n293115 );
xor ( n293117 , n2671 , n2688 );
buf ( n293118 , n293117 );
xor ( n2691 , n293083 , n293118 );
buf ( n293120 , n2691 );
buf ( n293121 , n293120 );
xor ( n293122 , n293018 , n293121 );
buf ( n293123 , n292401 );
not ( n2696 , n293123 );
buf ( n293125 , n292393 );
not ( n293126 , n293125 );
or ( n2699 , n2696 , n293126 );
buf ( n293128 , n291788 );
xor ( n293129 , n818 , n790 );
buf ( n293130 , n293129 );
nand ( n293131 , n293128 , n293130 );
buf ( n293132 , n293131 );
buf ( n293133 , n293132 );
nand ( n2706 , n2699 , n293133 );
buf ( n293135 , n2706 );
buf ( n293136 , n293135 );
buf ( n293137 , n799 );
buf ( n293138 , n811 );
or ( n2711 , n293137 , n293138 );
buf ( n293140 , n812 );
nand ( n2713 , n2711 , n293140 );
buf ( n293142 , n2713 );
buf ( n293143 , n293142 );
buf ( n293144 , n799 );
buf ( n293145 , n811 );
nand ( n293146 , n293144 , n293145 );
buf ( n293147 , n293146 );
buf ( n293148 , n293147 );
buf ( n293149 , n810 );
and ( n2722 , n293143 , n293148 , n293149 );
buf ( n293151 , n2722 );
buf ( n293152 , n292935 );
not ( n2725 , n293152 );
buf ( n2726 , n291805 );
not ( n2727 , n2726 );
or ( n2728 , n2725 , n2727 );
buf ( n2729 , n291939 );
buf ( n293158 , n780 );
buf ( n293159 , n828 );
xor ( n293160 , n293158 , n293159 );
buf ( n293161 , n293160 );
buf ( n293162 , n293161 );
nand ( n293163 , n2729 , n293162 );
buf ( n293164 , n293163 );
buf ( n293165 , n293164 );
nand ( n293166 , n2728 , n293165 );
buf ( n293167 , n293166 );
xor ( n2740 , n293151 , n293167 );
buf ( n293169 , n2740 );
xor ( n2742 , n293136 , n293169 );
not ( n2743 , n2513 );
not ( n293172 , n292906 );
or ( n293173 , n2743 , n293172 );
buf ( n293174 , n2513 );
buf ( n293175 , n292906 );
nor ( n293176 , n293174 , n293175 );
buf ( n293177 , n293176 );
or ( n2750 , n292921 , n293177 );
nand ( n293179 , n293173 , n2750 );
buf ( n293180 , n293179 );
xor ( n2753 , n2742 , n293180 );
buf ( n293182 , n2753 );
buf ( n293183 , n293182 );
xor ( n2756 , n292820 , n292825 );
and ( n293185 , n2756 , n292834 );
and ( n293186 , n292820 , n292825 );
or ( n2759 , n293185 , n293186 );
buf ( n293188 , n2759 );
buf ( n293189 , n293188 );
xor ( n2762 , n293183 , n293189 );
xor ( n293191 , n292846 , n292863 );
and ( n2764 , n293191 , n292879 );
and ( n293193 , n292846 , n292863 );
or ( n293194 , n2764 , n293193 );
buf ( n293195 , n293194 );
buf ( n293196 , n293195 );
buf ( n293197 , n292855 );
not ( n293198 , n293197 );
buf ( n293199 , n1271 );
not ( n2772 , n293199 );
or ( n293201 , n293198 , n2772 );
xor ( n293202 , n830 , n778 );
buf ( n293203 , n293202 );
buf ( n293204 , n831 );
nand ( n2777 , n293203 , n293204 );
buf ( n293206 , n2777 );
buf ( n293207 , n293206 );
nand ( n293208 , n293201 , n293207 );
buf ( n293209 , n293208 );
buf ( n293210 , n292428 );
not ( n293211 , n293210 );
not ( n2784 , n820 );
nand ( n293213 , n2784 , n291732 );
nand ( n293214 , n820 , n821 );
and ( n2787 , n2237 , n293213 , n293214 );
buf ( n293216 , n2787 );
not ( n2789 , n293216 );
or ( n293218 , n293211 , n2789 );
xor ( n293219 , n788 , n820 );
nand ( n2792 , n291969 , n293219 );
buf ( n293221 , n2792 );
nand ( n293222 , n293218 , n293221 );
buf ( n293223 , n293222 );
buf ( n293224 , n293223 );
xor ( n2797 , n293209 , n293224 );
buf ( n293226 , n292984 );
not ( n293227 , n293226 );
buf ( n293228 , n291880 );
not ( n293229 , n293228 );
or ( n293230 , n293227 , n293229 );
buf ( n293231 , n291886 );
buf ( n293232 , n782 );
buf ( n293233 , n826 );
xor ( n2806 , n293232 , n293233 );
buf ( n2807 , n2806 );
buf ( n293236 , n2807 );
nand ( n2809 , n293231 , n293236 );
buf ( n293238 , n2809 );
buf ( n293239 , n293238 );
nand ( n293240 , n293230 , n293239 );
buf ( n293241 , n293240 );
xor ( n2814 , n2797 , n293241 );
buf ( n293243 , n2814 );
xor ( n293244 , n293196 , n293243 );
buf ( n293245 , n2535 );
buf ( n293246 , n292996 );
or ( n2819 , n293245 , n293246 );
buf ( n293248 , n292979 );
nand ( n293249 , n2819 , n293248 );
buf ( n293250 , n293249 );
nand ( n2823 , n292996 , n2535 );
nand ( n293252 , n293250 , n2823 );
buf ( n293253 , n293252 );
xor ( n2826 , n293244 , n293253 );
buf ( n293255 , n2826 );
buf ( n293256 , n293255 );
xor ( n2829 , n2762 , n293256 );
buf ( n293258 , n2829 );
buf ( n293259 , n293258 );
xor ( n2832 , n293122 , n293259 );
buf ( n293261 , n2832 );
buf ( n293262 , n293261 );
and ( n2835 , n2584 , n293262 );
and ( n293264 , n292754 , n2583 );
or ( n293265 , n2835 , n293264 );
buf ( n293266 , n293265 );
buf ( n293267 , n293266 );
xor ( n293268 , n292347 , n293267 );
nand ( n293269 , n293167 , n293151 );
not ( n2842 , n293209 );
not ( n293271 , n293224 );
or ( n293272 , n2842 , n293271 );
or ( n2845 , n293209 , n293223 );
nand ( n293274 , n2845 , n293241 );
nand ( n2847 , n293272 , n293274 );
xor ( n2848 , n293269 , n2847 );
xor ( n293277 , n2620 , n2638 );
and ( n293278 , n293277 , n2652 );
and ( n2851 , n2620 , n2638 );
or ( n293280 , n293278 , n2851 );
xnor ( n293281 , n2848 , n293280 );
buf ( n293282 , n293281 );
xor ( n293283 , n293196 , n293243 );
and ( n2856 , n293283 , n293253 );
and ( n293285 , n293196 , n293243 );
or ( n293286 , n2856 , n293285 );
buf ( n293287 , n293286 );
buf ( n293288 , n293287 );
xor ( n293289 , n293282 , n293288 );
xor ( n2862 , n293036 , n293082 );
and ( n293291 , n2862 , n293118 );
and ( n2864 , n293036 , n293082 );
or ( n2865 , n293291 , n2864 );
buf ( n293294 , n2865 );
buf ( n293295 , n293294 );
xor ( n2868 , n293289 , n293295 );
buf ( n293297 , n2868 );
buf ( n293298 , n293297 );
xor ( n2871 , n293018 , n293121 );
and ( n293300 , n2871 , n293259 );
and ( n2873 , n293018 , n293121 );
or ( n2874 , n293300 , n2873 );
buf ( n293303 , n2874 );
buf ( n293304 , n293303 );
xor ( n2877 , n293298 , n293304 );
not ( n293306 , n293093 );
not ( n293307 , n292892 );
or ( n2880 , n293306 , n293307 );
buf ( n293309 , n1712 );
buf ( n293310 , n791 );
buf ( n293311 , n816 );
xor ( n293312 , n293310 , n293311 );
buf ( n293313 , n293312 );
buf ( n293314 , n293313 );
nand ( n293315 , n293309 , n293314 );
buf ( n293316 , n293315 );
nand ( n293317 , n2880 , n293316 );
buf ( n293318 , n2681 );
not ( n293319 , n293318 );
nand ( n2892 , n2289 , n292718 );
not ( n2893 , n2892 );
buf ( n293322 , n2893 );
not ( n2895 , n293322 );
or ( n2896 , n293319 , n2895 );
buf ( n293325 , n2089 );
buf ( n293326 , n793 );
buf ( n293327 , n814 );
xor ( n293328 , n293326 , n293327 );
buf ( n293329 , n293328 );
buf ( n293330 , n293329 );
nand ( n293331 , n293325 , n293330 );
buf ( n293332 , n293331 );
buf ( n293333 , n293332 );
nand ( n293334 , n2896 , n293333 );
buf ( n293335 , n293334 );
xor ( n2908 , n293317 , n293335 );
buf ( n293337 , n293044 );
not ( n293338 , n293337 );
buf ( n293339 , n292631 );
not ( n293340 , n293339 );
or ( n293341 , n293338 , n293340 );
buf ( n293342 , n292105 );
buf ( n293343 , n785 );
buf ( n293344 , n822 );
xor ( n293345 , n293343 , n293344 );
buf ( n293346 , n293345 );
buf ( n293347 , n293346 );
nand ( n293348 , n293342 , n293347 );
buf ( n293349 , n293348 );
buf ( n293350 , n293349 );
nand ( n293351 , n293341 , n293350 );
buf ( n293352 , n293351 );
buf ( n293353 , n293352 );
not ( n293354 , n293353 );
buf ( n293355 , n293354 );
and ( n2928 , n2908 , n293355 );
not ( n2929 , n2908 );
and ( n2930 , n2929 , n293352 );
nor ( n293359 , n2928 , n2930 );
buf ( n293360 , n293359 );
not ( n293361 , n293360 );
buf ( n293362 , n293361 );
buf ( n293363 , n293362 );
not ( n293364 , n293363 );
not ( n293365 , n293097 );
not ( n2938 , n2660 );
or ( n293367 , n293365 , n2938 );
not ( n2940 , n2670 );
not ( n2941 , n293087 );
or ( n293370 , n2940 , n2941 );
nand ( n293371 , n293370 , n293115 );
nand ( n2944 , n293367 , n293371 );
buf ( n293373 , n293219 );
not ( n293374 , n293373 );
buf ( n293375 , n292668 );
not ( n293376 , n293375 );
or ( n293377 , n293374 , n293376 );
not ( n2950 , n820 );
not ( n293379 , n787 );
not ( n293380 , n293379 );
or ( n2953 , n2950 , n293380 );
nand ( n293382 , n2784 , n787 );
nand ( n293383 , n2953 , n293382 );
nand ( n2956 , n291969 , n293383 );
buf ( n293385 , n2956 );
nand ( n2958 , n293377 , n293385 );
buf ( n293387 , n2958 );
buf ( n293388 , n293387 );
not ( n293389 , n293388 );
buf ( n293390 , n2807 );
not ( n293391 , n293390 );
not ( n293392 , n291885 );
xor ( n2965 , n826 , n827 );
and ( n293394 , n293392 , n2965 );
buf ( n2967 , n293394 );
not ( n2968 , n2967 );
or ( n2969 , n293391 , n2968 );
buf ( n293398 , n781 );
buf ( n293399 , n826 );
xor ( n2972 , n293398 , n293399 );
buf ( n293401 , n2972 );
not ( n293402 , n292006 );
nand ( n2975 , n293401 , n293402 );
buf ( n293404 , n2975 );
nand ( n293405 , n2969 , n293404 );
buf ( n293406 , n293405 );
buf ( n293407 , n293406 );
not ( n2980 , n293407 );
buf ( n293409 , n2980 );
buf ( n293410 , n293409 );
not ( n293411 , n293410 );
and ( n293412 , n293389 , n293411 );
buf ( n293413 , n293387 );
buf ( n293414 , n293409 );
and ( n293415 , n293413 , n293414 );
nor ( n2988 , n293412 , n293415 );
buf ( n2989 , n2988 );
buf ( n293418 , n2989 );
not ( n2991 , n291788 );
xor ( n293420 , n818 , n789 );
not ( n293421 , n293420 );
or ( n2994 , n2991 , n293421 );
not ( n293423 , n1961 );
not ( n2996 , n291979 );
not ( n2997 , n2996 );
nand ( n2998 , n293423 , n2997 , n293129 );
nand ( n2999 , n2994 , n2998 );
buf ( n293428 , n2999 );
and ( n3001 , n293418 , n293428 );
not ( n3002 , n293418 );
buf ( n293431 , n2999 );
not ( n3004 , n293431 );
buf ( n293433 , n3004 );
buf ( n293434 , n293433 );
and ( n293435 , n3002 , n293434 );
nor ( n3008 , n3001 , n293435 );
buf ( n293437 , n3008 );
xor ( n3010 , n2944 , n293437 );
buf ( n293439 , n3010 );
not ( n293440 , n293439 );
or ( n3013 , n293364 , n293440 );
buf ( n293442 , n3010 );
buf ( n293443 , n293362 );
or ( n3016 , n293442 , n293443 );
nand ( n3017 , n3013 , n3016 );
buf ( n293446 , n3017 );
buf ( n3019 , n293446 );
buf ( n293448 , n293202 );
not ( n293449 , n293448 );
buf ( n293450 , n830 );
not ( n3023 , n293450 );
buf ( n293452 , n831 );
nor ( n3025 , n3023 , n293452 );
buf ( n293454 , n3025 );
buf ( n293455 , n293454 );
not ( n3028 , n293455 );
or ( n293457 , n293449 , n3028 );
xor ( n3030 , n830 , n777 );
buf ( n293459 , n3030 );
buf ( n293460 , n831 );
nand ( n3033 , n293459 , n293460 );
buf ( n293462 , n3033 );
buf ( n293463 , n293462 );
nand ( n3036 , n293457 , n293463 );
buf ( n293465 , n3036 );
buf ( n293466 , n293465 );
not ( n293467 , n2634 );
xnor ( n293468 , n810 , n811 );
nor ( n3041 , n293468 , n2410 );
not ( n3042 , n3041 );
or ( n293471 , n293467 , n3042 );
xor ( n3044 , n810 , n797 );
nand ( n3045 , n3044 , n2410 );
nand ( n293474 , n293471 , n3045 );
buf ( n293475 , n293474 );
xor ( n3048 , n293466 , n293475 );
buf ( n293477 , n2646 );
not ( n293478 , n293477 );
buf ( n293479 , n2373 );
not ( n3052 , n293479 );
or ( n3053 , n293478 , n3052 );
buf ( n293482 , n292810 );
xor ( n3055 , n812 , n795 );
buf ( n293484 , n3055 );
nand ( n293485 , n293482 , n293484 );
buf ( n293486 , n293485 );
buf ( n293487 , n293486 );
nand ( n3060 , n3053 , n293487 );
buf ( n293489 , n3060 );
buf ( n293490 , n293489 );
xor ( n3063 , n3048 , n293490 );
buf ( n293492 , n3063 );
xor ( n293493 , n293136 , n293169 );
and ( n3066 , n293493 , n293180 );
and ( n293495 , n293136 , n293169 );
or ( n3068 , n3066 , n293495 );
buf ( n293497 , n3068 );
xor ( n3070 , n293492 , n293497 );
buf ( n293499 , n293084 );
not ( n3072 , n293499 );
buf ( n293501 , n291835 );
not ( n3074 , n293501 );
or ( n293503 , n3072 , n3074 );
buf ( n293504 , n291843 );
buf ( n293505 , n783 );
buf ( n293506 , n824 );
xor ( n3079 , n293505 , n293506 );
buf ( n3080 , n3079 );
buf ( n293509 , n3080 );
nand ( n293510 , n293504 , n293509 );
buf ( n293511 , n293510 );
buf ( n293512 , n293511 );
nand ( n293513 , n293503 , n293512 );
buf ( n293514 , n293513 );
not ( n3087 , n293514 );
buf ( n293516 , n293161 );
not ( n3089 , n293516 );
buf ( n3090 , n291805 );
not ( n3091 , n3090 );
or ( n3092 , n3089 , n3091 );
and ( n3093 , n829 , n830 );
not ( n3094 , n829 );
and ( n293523 , n3094 , n292367 );
nor ( n3096 , n3093 , n293523 );
not ( n293525 , n3096 );
not ( n293526 , n293525 );
buf ( n293527 , n779 );
buf ( n293528 , n828 );
xor ( n293529 , n293527 , n293528 );
buf ( n293530 , n293529 );
nand ( n293531 , n293526 , n293530 );
buf ( n293532 , n293531 );
nand ( n293533 , n3092 , n293532 );
buf ( n293534 , n293533 );
not ( n293535 , n293534 );
not ( n3108 , n809 );
not ( n293537 , n810 );
not ( n293538 , n293537 );
or ( n3111 , n3108 , n293538 );
not ( n3112 , n809 );
nand ( n293541 , n3112 , n810 );
nand ( n3114 , n3111 , n293541 );
buf ( n293543 , n3114 );
buf ( n293544 , n799 );
and ( n293545 , n293543 , n293544 );
buf ( n293546 , n293545 );
not ( n3119 , n293546 );
nand ( n293548 , n293535 , n3119 );
not ( n293549 , n293548 );
not ( n3122 , n293549 );
or ( n3123 , n3087 , n3122 );
nand ( n3124 , n293534 , n293546 );
not ( n3125 , n3124 );
nand ( n3126 , n3125 , n293514 );
nand ( n293555 , n3123 , n3126 );
not ( n293556 , n293534 );
buf ( n3129 , n293546 );
nor ( n293558 , n293556 , n293514 , n3129 );
nand ( n293559 , n293535 , n293546 );
nor ( n3132 , n293514 , n293559 );
or ( n3133 , n293555 , n293558 , n3132 );
xor ( n3134 , n3070 , n3133 );
buf ( n293563 , n3134 );
xor ( n293564 , n3019 , n293563 );
xor ( n3137 , n293183 , n293189 );
and ( n3138 , n3137 , n293256 );
and ( n3139 , n293183 , n293189 );
or ( n3140 , n3138 , n3139 );
buf ( n293569 , n3140 );
buf ( n293570 , n293569 );
xor ( n293571 , n293564 , n293570 );
buf ( n293572 , n293571 );
buf ( n293573 , n293572 );
xor ( n293574 , n2877 , n293573 );
buf ( n293575 , n293574 );
buf ( n293576 , n293575 );
and ( n3149 , n293268 , n293576 );
and ( n3150 , n292347 , n293267 );
or ( n293579 , n3149 , n3150 );
buf ( n293580 , n293579 );
buf ( n293581 , n293580 );
not ( n3154 , n293581 );
or ( n3155 , n292346 , n3154 );
buf ( n293584 , n831 );
not ( n293585 , n293584 );
buf ( n3158 , n873 );
buf ( n293587 , n293266 );
xor ( n3160 , n3158 , n293587 );
buf ( n293589 , n293575 );
and ( n3162 , n3160 , n293589 );
and ( n293591 , n3158 , n293587 );
or ( n293592 , n3162 , n293591 );
buf ( n293593 , n293592 );
buf ( n293594 , n293593 );
nand ( n3167 , n293585 , n293594 );
buf ( n293596 , n3167 );
buf ( n293597 , n293596 );
nand ( n293598 , n3155 , n293597 );
buf ( n293599 , n293598 );
buf ( n3172 , n293599 );
buf ( n293601 , n3172 );
buf ( n293602 , n831 );
not ( n3175 , n293602 );
buf ( n293604 , n3030 );
not ( n3177 , n293604 );
buf ( n293606 , n830 );
not ( n293607 , n293606 );
buf ( n3180 , n831 );
nor ( n3181 , n293607 , n3180 );
buf ( n3182 , n3181 );
buf ( n293611 , n3182 );
not ( n3184 , n293611 );
or ( n293613 , n3177 , n3184 );
buf ( n293614 , n776 );
buf ( n293615 , n830 );
xor ( n293616 , n293614 , n293615 );
buf ( n293617 , n293616 );
buf ( n293618 , n293617 );
buf ( n293619 , n831 );
nand ( n3192 , n293618 , n293619 );
buf ( n293621 , n3192 );
buf ( n293622 , n293621 );
nand ( n293623 , n293613 , n293622 );
buf ( n293624 , n293623 );
not ( n3197 , n293624 );
buf ( n293626 , n293401 );
not ( n293627 , n293626 );
buf ( n293628 , n291880 );
not ( n293629 , n293628 );
or ( n3202 , n293627 , n293629 );
buf ( n293631 , n291886 );
buf ( n293632 , n780 );
buf ( n293633 , n826 );
xor ( n293634 , n293632 , n293633 );
buf ( n293635 , n293634 );
buf ( n3208 , n293635 );
nand ( n3209 , n293631 , n3208 );
buf ( n3210 , n3209 );
buf ( n3211 , n3210 );
nand ( n3212 , n3202 , n3211 );
buf ( n3213 , n3212 );
xor ( n293642 , n3197 , n3213 );
buf ( n293643 , n799 );
buf ( n293644 , n808 );
xor ( n293645 , n293643 , n293644 );
buf ( n293646 , n293645 );
buf ( n293647 , n293646 );
not ( n293648 , n293647 );
xor ( n293649 , n809 , n810 );
not ( n3222 , n293649 );
xor ( n3223 , n808 , n809 );
nand ( n293652 , n3222 , n3223 );
buf ( n3225 , n293652 );
not ( n293654 , n3225 );
buf ( n293655 , n293654 );
buf ( n3228 , n293655 );
not ( n3229 , n3228 );
or ( n3230 , n293648 , n3229 );
not ( n293659 , n3222 );
buf ( n293660 , n798 );
buf ( n3233 , n808 );
xor ( n3234 , n293660 , n3233 );
buf ( n3235 , n3234 );
nand ( n293664 , n293659 , n3235 );
buf ( n293665 , n293664 );
nand ( n293666 , n3230 , n293665 );
buf ( n293667 , n293666 );
xor ( n3240 , n293642 , n293667 );
not ( n293669 , n3240 );
buf ( n293670 , n293669 );
not ( n3243 , n293670 );
buf ( n3244 , n293346 );
not ( n3245 , n3244 );
buf ( n3246 , n292631 );
not ( n3247 , n3246 );
or ( n3248 , n3245 , n3247 );
buf ( n3249 , n1600 );
buf ( n293678 , n784 );
buf ( n293679 , n822 );
xor ( n293680 , n293678 , n293679 );
buf ( n293681 , n293680 );
buf ( n293682 , n293681 );
nand ( n293683 , n3249 , n293682 );
buf ( n293684 , n293683 );
buf ( n293685 , n293684 );
nand ( n293686 , n3248 , n293685 );
buf ( n293687 , n293686 );
buf ( n293688 , n3055 );
not ( n293689 , n293688 );
buf ( n293690 , n2373 );
not ( n293691 , n293690 );
or ( n293692 , n293689 , n293691 );
buf ( n293693 , n2026 );
buf ( n293694 , n794 );
buf ( n293695 , n812 );
xor ( n3268 , n293694 , n293695 );
buf ( n293697 , n3268 );
buf ( n293698 , n293697 );
nand ( n3271 , n293693 , n293698 );
buf ( n293700 , n3271 );
buf ( n293701 , n293700 );
nand ( n293702 , n293692 , n293701 );
buf ( n293703 , n293702 );
xnor ( n293704 , n293687 , n293703 );
buf ( n293705 , n293704 );
buf ( n293706 , n3044 );
not ( n293707 , n293706 );
buf ( n293708 , n293058 );
not ( n3281 , n293708 );
or ( n293710 , n293707 , n3281 );
buf ( n293711 , n292841 );
buf ( n293712 , n796 );
buf ( n293713 , n810 );
xor ( n293714 , n293712 , n293713 );
buf ( n293715 , n293714 );
buf ( n293716 , n293715 );
nand ( n293717 , n293711 , n293716 );
buf ( n293718 , n293717 );
buf ( n293719 , n293718 );
nand ( n3292 , n293710 , n293719 );
buf ( n3293 , n3292 );
buf ( n3294 , n3293 );
and ( n3295 , n293705 , n3294 );
not ( n293724 , n293705 );
buf ( n293725 , n3293 );
not ( n3298 , n293725 );
buf ( n3299 , n3298 );
buf ( n293728 , n3299 );
and ( n293729 , n293724 , n293728 );
nor ( n3302 , n3295 , n293729 );
buf ( n293731 , n3302 );
buf ( n293732 , n293731 );
not ( n3305 , n293732 );
buf ( n293734 , n3305 );
buf ( n293735 , n293734 );
not ( n3308 , n293735 );
or ( n3309 , n3243 , n3308 );
not ( n3310 , n3240 );
not ( n3311 , n293731 );
or ( n3312 , n3310 , n3311 );
not ( n293741 , n293317 );
not ( n3314 , n293352 );
or ( n293743 , n293741 , n3314 );
buf ( n293744 , n293317 );
not ( n3317 , n293744 );
buf ( n293746 , n3317 );
buf ( n293747 , n293746 );
not ( n293748 , n293747 );
buf ( n293749 , n293355 );
not ( n3322 , n293749 );
or ( n293751 , n293748 , n3322 );
buf ( n293752 , n293335 );
nand ( n293753 , n293751 , n293752 );
buf ( n293754 , n293753 );
nand ( n3327 , n293743 , n293754 );
nand ( n293756 , n3312 , n3327 );
buf ( n293757 , n293756 );
nand ( n3330 , n3309 , n293757 );
buf ( n3331 , n3330 );
not ( n293760 , n3331 );
buf ( n293761 , n293624 );
not ( n3334 , n293761 );
buf ( n293763 , n3213 );
not ( n293764 , n293763 );
or ( n3337 , n3334 , n293764 );
buf ( n293766 , n3197 );
not ( n293767 , n293766 );
buf ( n293768 , n3213 );
not ( n3341 , n293768 );
buf ( n293770 , n3341 );
buf ( n293771 , n293770 );
not ( n3344 , n293771 );
or ( n293773 , n293767 , n3344 );
buf ( n293774 , n293667 );
nand ( n293775 , n293773 , n293774 );
buf ( n293776 , n293775 );
buf ( n293777 , n293776 );
nand ( n293778 , n3337 , n293777 );
buf ( n293779 , n293778 );
not ( n293780 , n293779 );
not ( n293781 , n293313 );
not ( n3354 , n292892 );
or ( n293783 , n293781 , n3354 );
buf ( n293784 , n1712 );
buf ( n293785 , n790 );
buf ( n293786 , n816 );
xor ( n293787 , n293785 , n293786 );
buf ( n293788 , n293787 );
buf ( n293789 , n293788 );
nand ( n293790 , n293784 , n293789 );
buf ( n293791 , n293790 );
nand ( n3364 , n293783 , n293791 );
not ( n293793 , n3080 );
not ( n3366 , n292473 );
or ( n293795 , n293793 , n3366 );
buf ( n293796 , n1613 );
xor ( n3369 , n824 , n782 );
buf ( n293798 , n3369 );
nand ( n3371 , n293796 , n293798 );
buf ( n293800 , n3371 );
nand ( n293801 , n293795 , n293800 );
or ( n293802 , n3364 , n293801 );
buf ( n293803 , n293329 );
not ( n293804 , n293803 );
buf ( n293805 , n292509 );
not ( n3378 , n293805 );
or ( n3379 , n293804 , n3378 );
buf ( n3380 , n292725 );
buf ( n3381 , n792 );
buf ( n3382 , n814 );
xor ( n3383 , n3381 , n3382 );
buf ( n3384 , n3383 );
buf ( n3385 , n3384 );
nand ( n3386 , n3380 , n3385 );
buf ( n3387 , n3386 );
buf ( n3388 , n3387 );
nand ( n3389 , n3379 , n3388 );
buf ( n3390 , n3389 );
nand ( n293819 , n293802 , n3390 );
nand ( n3392 , n293801 , n3364 );
nand ( n293821 , n293819 , n3392 );
not ( n3394 , n293821 );
or ( n3395 , n293780 , n3394 );
not ( n293824 , n293779 );
buf ( n293825 , n293821 );
not ( n293826 , n293825 );
buf ( n293827 , n293826 );
nand ( n293828 , n293824 , n293827 );
nand ( n293829 , n3395 , n293828 );
buf ( n293830 , n3235 );
not ( n293831 , n293830 );
buf ( n293832 , n3222 );
buf ( n293833 , n3223 );
nand ( n293834 , n293832 , n293833 );
buf ( n293835 , n293834 );
not ( n3408 , n293835 );
buf ( n293837 , n3408 );
not ( n3410 , n293837 );
or ( n293839 , n293831 , n3410 );
buf ( n293840 , n797 );
buf ( n293841 , n808 );
xor ( n3414 , n293840 , n293841 );
buf ( n293843 , n3414 );
buf ( n3416 , n293843 );
buf ( n293845 , n3114 );
nand ( n293846 , n3416 , n293845 );
buf ( n293847 , n293846 );
buf ( n293848 , n293847 );
nand ( n293849 , n293839 , n293848 );
buf ( n293850 , n293849 );
buf ( n293851 , n293850 );
buf ( n293852 , n293635 );
not ( n3425 , n293852 );
buf ( n293854 , n291880 );
not ( n3427 , n293854 );
or ( n293856 , n3425 , n3427 );
buf ( n293857 , n1579 );
buf ( n293858 , n779 );
buf ( n293859 , n826 );
xor ( n3432 , n293858 , n293859 );
buf ( n293861 , n3432 );
buf ( n293862 , n293861 );
nand ( n293863 , n293857 , n293862 );
buf ( n293864 , n293863 );
buf ( n293865 , n293864 );
nand ( n293866 , n293856 , n293865 );
buf ( n293867 , n293866 );
buf ( n293868 , n293867 );
xor ( n3441 , n293851 , n293868 );
xor ( n3442 , n820 , n786 );
buf ( n293871 , n3442 );
not ( n293872 , n293871 );
buf ( n293873 , n291722 );
not ( n3446 , n293873 );
or ( n3447 , n293872 , n3446 );
buf ( n293876 , n291906 );
buf ( n293877 , n785 );
buf ( n293878 , n820 );
xor ( n293879 , n293877 , n293878 );
buf ( n293880 , n293879 );
buf ( n293881 , n293880 );
nand ( n293882 , n293876 , n293881 );
buf ( n293883 , n293882 );
buf ( n293884 , n293883 );
nand ( n3457 , n3447 , n293884 );
buf ( n3458 , n3457 );
buf ( n293887 , n3458 );
xor ( n293888 , n3441 , n293887 );
buf ( n293889 , n293888 );
and ( n293890 , n293829 , n293889 );
not ( n3463 , n293829 );
buf ( n293892 , n293889 );
not ( n3465 , n293892 );
buf ( n293894 , n3465 );
and ( n3467 , n3463 , n293894 );
nor ( n293896 , n293890 , n3467 );
not ( n3469 , n293896 );
not ( n293898 , n3469 );
or ( n3471 , n293760 , n293898 );
or ( n3472 , n3331 , n3469 );
nand ( n293901 , n3471 , n3472 );
xor ( n293902 , n807 , n808 );
buf ( n293903 , n293902 );
buf ( n293904 , n799 );
and ( n293905 , n293903 , n293904 );
buf ( n293906 , n293905 );
buf ( n293907 , n293906 );
buf ( n293908 , n778 );
buf ( n293909 , n828 );
xor ( n3482 , n293908 , n293909 );
buf ( n3483 , n3482 );
buf ( n293912 , n3483 );
not ( n3485 , n293912 );
buf ( n293914 , n291805 );
not ( n293915 , n293914 );
or ( n293916 , n3485 , n293915 );
buf ( n293917 , n777 );
buf ( n293918 , n828 );
xor ( n293919 , n293917 , n293918 );
buf ( n293920 , n293919 );
nand ( n3493 , n293920 , n3096 );
buf ( n293922 , n3493 );
nand ( n3495 , n293916 , n293922 );
buf ( n293924 , n3495 );
buf ( n293925 , n293924 );
xor ( n293926 , n293907 , n293925 );
buf ( n293927 , n3369 );
not ( n3500 , n293927 );
buf ( n293929 , n292473 );
not ( n3502 , n293929 );
or ( n293931 , n3500 , n3502 );
buf ( n293932 , n1613 );
buf ( n293933 , n781 );
buf ( n293934 , n824 );
xor ( n293935 , n293933 , n293934 );
buf ( n293936 , n293935 );
buf ( n293937 , n293936 );
nand ( n3510 , n293932 , n293937 );
buf ( n293939 , n3510 );
buf ( n293940 , n293939 );
nand ( n3513 , n293931 , n293940 );
buf ( n293942 , n3513 );
buf ( n293943 , n293942 );
xor ( n3516 , n293926 , n293943 );
buf ( n293945 , n3516 );
buf ( n293946 , n293945 );
buf ( n293947 , n3182 );
not ( n3520 , n293947 );
buf ( n293949 , n293617 );
not ( n3522 , n293949 );
or ( n293951 , n3520 , n3522 );
buf ( n293952 , n775 );
buf ( n293953 , n830 );
xor ( n3526 , n293952 , n293953 );
buf ( n293955 , n3526 );
buf ( n293956 , n293955 );
buf ( n293957 , n831 );
nand ( n3530 , n293956 , n293957 );
buf ( n293959 , n3530 );
buf ( n293960 , n293959 );
nand ( n3533 , n293951 , n293960 );
buf ( n293962 , n3533 );
buf ( n293963 , n293962 );
buf ( n293964 , n293697 );
not ( n3537 , n293964 );
xnor ( n3538 , n812 , n813 );
nor ( n3539 , n3538 , n2366 );
buf ( n293968 , n3539 );
not ( n3541 , n293968 );
or ( n3542 , n3537 , n3541 );
buf ( n293971 , n793 );
buf ( n293972 , n812 );
xor ( n3545 , n293971 , n293972 );
buf ( n293974 , n3545 );
buf ( n293975 , n293974 );
buf ( n293976 , n2366 );
nand ( n3549 , n293975 , n293976 );
buf ( n293978 , n3549 );
buf ( n293979 , n293978 );
nand ( n3552 , n3542 , n293979 );
buf ( n293981 , n3552 );
buf ( n293982 , n293981 );
xor ( n3555 , n293963 , n293982 );
buf ( n293984 , n293715 );
not ( n3557 , n293984 );
buf ( n293986 , n293058 );
not ( n293987 , n293986 );
or ( n3560 , n3557 , n293987 );
buf ( n293989 , n292841 );
buf ( n293990 , n795 );
buf ( n293991 , n810 );
xor ( n3564 , n293990 , n293991 );
buf ( n293993 , n3564 );
buf ( n293994 , n293993 );
nand ( n3567 , n293989 , n293994 );
buf ( n293996 , n3567 );
buf ( n293997 , n293996 );
nand ( n3570 , n3560 , n293997 );
buf ( n293999 , n3570 );
buf ( n294000 , n293999 );
xnor ( n3573 , n3555 , n294000 );
buf ( n294002 , n3573 );
buf ( n294003 , n294002 );
not ( n3576 , n294003 );
buf ( n294005 , n3576 );
buf ( n3578 , n294005 );
xor ( n3579 , n293946 , n3578 );
not ( n294008 , n1712 );
buf ( n294009 , n789 );
buf ( n294010 , n816 );
xor ( n3583 , n294009 , n294010 );
buf ( n294012 , n3583 );
not ( n294013 , n294012 );
or ( n294014 , n294008 , n294013 );
not ( n294015 , n292885 );
not ( n3588 , n817 );
or ( n294017 , n294015 , n3588 );
nand ( n294018 , n2103 , n816 );
nand ( n3591 , n294017 , n294018 );
nand ( n294020 , n293788 , n3591 , n292700 );
nand ( n294021 , n294014 , n294020 );
not ( n3594 , n294021 );
buf ( n294023 , n3594 );
not ( n294024 , n294023 );
buf ( n294025 , n3384 );
not ( n294026 , n294025 );
buf ( n294027 , n2078 );
not ( n3600 , n294027 );
or ( n294029 , n294026 , n3600 );
buf ( n3602 , n2089 );
buf ( n294031 , n791 );
buf ( n294032 , n814 );
xor ( n294033 , n294031 , n294032 );
buf ( n294034 , n294033 );
buf ( n294035 , n294034 );
nand ( n294036 , n3602 , n294035 );
buf ( n294037 , n294036 );
buf ( n294038 , n294037 );
nand ( n294039 , n294029 , n294038 );
buf ( n294040 , n294039 );
buf ( n294041 , n294040 );
not ( n3614 , n294041 );
and ( n294043 , n294024 , n3614 );
buf ( n294044 , n294040 );
buf ( n294045 , n3594 );
and ( n294046 , n294044 , n294045 );
nor ( n3619 , n294043 , n294046 );
buf ( n294048 , n3619 );
buf ( n294049 , n294048 );
buf ( n294050 , n293681 );
not ( n294051 , n294050 );
buf ( n294052 , n292631 );
not ( n294053 , n294052 );
or ( n3626 , n294051 , n294053 );
buf ( n3627 , n1600 );
buf ( n294056 , n783 );
buf ( n294057 , n822 );
xor ( n294058 , n294056 , n294057 );
buf ( n294059 , n294058 );
buf ( n294060 , n294059 );
nand ( n294061 , n3627 , n294060 );
buf ( n294062 , n294061 );
buf ( n294063 , n294062 );
nand ( n3636 , n3626 , n294063 );
buf ( n3637 , n3636 );
buf ( n3638 , n3637 );
xor ( n3639 , n294049 , n3638 );
buf ( n294068 , n3639 );
buf ( n294069 , n294068 );
not ( n3642 , n294069 );
buf ( n3643 , n3642 );
buf ( n294072 , n3643 );
xor ( n294073 , n3579 , n294072 );
buf ( n294074 , n294073 );
buf ( n3647 , n294074 );
not ( n294076 , n3647 );
and ( n294077 , n293901 , n294076 );
not ( n3650 , n293901 );
and ( n294079 , n3650 , n3647 );
nor ( n294080 , n294077 , n294079 );
not ( n3653 , n293383 );
not ( n294082 , n291722 );
or ( n3655 , n3653 , n294082 );
nand ( n3656 , n291969 , n3442 );
nand ( n294085 , n3655 , n3656 );
not ( n3658 , n294085 );
buf ( n294087 , n291984 );
buf ( n294088 , n293420 );
and ( n3661 , n294087 , n294088 );
buf ( n294090 , n291788 );
buf ( n3663 , n788 );
buf ( n294092 , n818 );
xor ( n294093 , n3663 , n294092 );
buf ( n294094 , n294093 );
buf ( n294095 , n294094 );
and ( n294096 , n294090 , n294095 );
nor ( n3669 , n3661 , n294096 );
buf ( n3670 , n3669 );
xor ( n294099 , n3658 , n3670 );
buf ( n294100 , n799 );
buf ( n294101 , n809 );
or ( n294102 , n294100 , n294101 );
buf ( n294103 , n810 );
nand ( n294104 , n294102 , n294103 );
buf ( n294105 , n294104 );
buf ( n3678 , n799 );
buf ( n294107 , n809 );
nand ( n294108 , n3678 , n294107 );
buf ( n294109 , n294108 );
and ( n3682 , n294105 , n294109 , n808 );
not ( n3683 , n293530 );
not ( n294112 , n291805 );
or ( n294113 , n3683 , n294112 );
nand ( n294114 , n3483 , n291939 );
nand ( n3687 , n294113 , n294114 );
or ( n294116 , n3682 , n3687 );
nand ( n294117 , n3687 , n3682 );
nand ( n3690 , n294116 , n294117 );
and ( n294119 , n294099 , n3690 );
not ( n294120 , n294099 );
not ( n3693 , n3690 );
and ( n294122 , n294120 , n3693 );
or ( n294123 , n294119 , n294122 );
buf ( n294124 , n294123 );
not ( n294125 , n294124 );
not ( n294126 , n293280 );
not ( n3699 , n2847 );
nand ( n3700 , n3699 , n293269 );
not ( n294129 , n3700 );
or ( n3702 , n294126 , n294129 );
not ( n294131 , n293269 );
nand ( n3704 , n294131 , n2847 );
nand ( n3705 , n3702 , n3704 );
buf ( n294134 , n3705 );
not ( n294135 , n294134 );
or ( n294136 , n294125 , n294135 );
buf ( n294137 , n3705 );
buf ( n294138 , n294123 );
or ( n294139 , n294137 , n294138 );
xor ( n3712 , n293801 , n3390 );
xor ( n294141 , n3712 , n3364 );
buf ( n294142 , n294141 );
nand ( n294143 , n294139 , n294142 );
buf ( n294144 , n294143 );
buf ( n294145 , n294144 );
nand ( n3718 , n294136 , n294145 );
buf ( n3719 , n3718 );
buf ( n294148 , n3719 );
and ( n3721 , n3658 , n3670 );
buf ( n294150 , n3721 );
buf ( n294151 , n3690 );
or ( n294152 , n294150 , n294151 );
buf ( n294153 , n3670 );
not ( n3726 , n294153 );
buf ( n294155 , n294085 );
nand ( n294156 , n3726 , n294155 );
buf ( n294157 , n294156 );
buf ( n294158 , n294157 );
nand ( n294159 , n294152 , n294158 );
buf ( n294160 , n294159 );
buf ( n294161 , n294160 );
xor ( n3734 , n293466 , n293475 );
and ( n294163 , n3734 , n293490 );
and ( n3736 , n293466 , n293475 );
or ( n294165 , n294163 , n3736 );
buf ( n294166 , n294165 );
buf ( n294167 , n293409 );
not ( n294168 , n294167 );
buf ( n294169 , n294168 );
buf ( n294170 , n294169 );
buf ( n294171 , n2999 );
or ( n3744 , n294170 , n294171 );
buf ( n294173 , n293387 );
nand ( n294174 , n3744 , n294173 );
buf ( n294175 , n294174 );
buf ( n294176 , n294175 );
buf ( n294177 , n2999 );
buf ( n294178 , n294169 );
nand ( n294179 , n294177 , n294178 );
buf ( n294180 , n294179 );
buf ( n294181 , n294180 );
nand ( n294182 , n294176 , n294181 );
buf ( n294183 , n294182 );
xor ( n294184 , n294166 , n294183 );
not ( n3757 , n293514 );
not ( n294186 , n293548 );
or ( n3759 , n3757 , n294186 );
nand ( n294188 , n3759 , n3124 );
and ( n294189 , n294184 , n294188 );
and ( n3762 , n294166 , n294183 );
or ( n294191 , n294189 , n3762 );
buf ( n3764 , n294191 );
xor ( n3765 , n294161 , n3764 );
buf ( n294194 , n294094 );
not ( n3767 , n294194 );
buf ( n294196 , n291984 );
not ( n3769 , n294196 );
or ( n294198 , n3767 , n3769 );
buf ( n294199 , n291989 );
buf ( n294200 , n787 );
buf ( n294201 , n818 );
xor ( n294202 , n294200 , n294201 );
buf ( n294203 , n294202 );
buf ( n294204 , n294203 );
nand ( n3777 , n294199 , n294204 );
buf ( n294206 , n3777 );
buf ( n294207 , n294206 );
nand ( n294208 , n294198 , n294207 );
buf ( n294209 , n294208 );
buf ( n294210 , n294209 );
not ( n294211 , n294117 );
buf ( n294212 , n294211 );
xor ( n3785 , n294210 , n294212 );
buf ( n294214 , n293703 );
buf ( n294215 , n293687 );
nor ( n294216 , n294214 , n294215 );
buf ( n294217 , n294216 );
buf ( n294218 , n294217 );
buf ( n294219 , n3299 );
or ( n3792 , n294218 , n294219 );
buf ( n294221 , n293703 );
buf ( n294222 , n293687 );
nand ( n294223 , n294221 , n294222 );
buf ( n294224 , n294223 );
buf ( n294225 , n294224 );
nand ( n3798 , n3792 , n294225 );
buf ( n294227 , n3798 );
buf ( n294228 , n294227 );
xor ( n294229 , n3785 , n294228 );
buf ( n294230 , n294229 );
buf ( n294231 , n294230 );
xor ( n3804 , n3765 , n294231 );
buf ( n294233 , n3804 );
buf ( n294234 , n294233 );
xor ( n294235 , n294148 , n294234 );
xor ( n294236 , n294166 , n294183 );
xor ( n3809 , n294236 , n294188 );
buf ( n294238 , n3809 );
buf ( n294239 , n293437 );
not ( n3812 , n294239 );
buf ( n294241 , n293359 );
not ( n294242 , n294241 );
or ( n294243 , n3812 , n294242 );
buf ( n294244 , n2944 );
nand ( n294245 , n294243 , n294244 );
buf ( n294246 , n294245 );
buf ( n3819 , n294246 );
buf ( n294248 , n293437 );
not ( n3821 , n294248 );
buf ( n294250 , n293362 );
nand ( n294251 , n3821 , n294250 );
buf ( n294252 , n294251 );
buf ( n294253 , n294252 );
nand ( n294254 , n3819 , n294253 );
buf ( n294255 , n294254 );
buf ( n294256 , n294255 );
xor ( n294257 , n294238 , n294256 );
not ( n294258 , n3327 );
and ( n3831 , n3240 , n294258 );
not ( n294260 , n3240 );
and ( n294261 , n294260 , n3327 );
nor ( n3834 , n3831 , n294261 );
and ( n294263 , n3834 , n293734 );
not ( n294264 , n3834 );
buf ( n294265 , n293734 );
not ( n294266 , n294265 );
buf ( n294267 , n294266 );
and ( n3840 , n294264 , n294267 );
nor ( n3841 , n294263 , n3840 );
buf ( n294270 , n3841 );
and ( n294271 , n294257 , n294270 );
and ( n3844 , n294238 , n294256 );
or ( n3845 , n294271 , n3844 );
buf ( n294274 , n3845 );
buf ( n294275 , n294274 );
xor ( n294276 , n294235 , n294275 );
buf ( n294277 , n294276 );
xor ( n294278 , n294080 , n294277 );
xor ( n294279 , n293492 , n293497 );
and ( n3852 , n294279 , n3133 );
and ( n294281 , n293492 , n293497 );
or ( n294282 , n3852 , n294281 );
buf ( n294283 , n294282 );
and ( n294284 , n3693 , n294099 );
not ( n294285 , n3693 );
not ( n3858 , n294099 );
and ( n294287 , n294285 , n3858 );
nor ( n294288 , n294284 , n294287 );
and ( n294289 , n294288 , n294141 );
not ( n3862 , n294288 );
not ( n294291 , n294141 );
and ( n3864 , n3862 , n294291 );
nor ( n3865 , n294289 , n3864 );
not ( n294294 , n3865 );
not ( n294295 , n294294 );
not ( n3868 , n3705 );
or ( n294297 , n294295 , n3868 );
not ( n3870 , n3705 );
nand ( n294299 , n3870 , n3865 );
nand ( n294300 , n294297 , n294299 );
buf ( n294301 , n294300 );
xor ( n294302 , n294283 , n294301 );
xor ( n294303 , n294238 , n294256 );
xor ( n3876 , n294303 , n294270 );
buf ( n294305 , n3876 );
buf ( n294306 , n294305 );
and ( n3879 , n294302 , n294306 );
and ( n3880 , n294283 , n294301 );
or ( n294309 , n3879 , n3880 );
buf ( n294310 , n294309 );
and ( n3883 , n294278 , n294310 );
and ( n294312 , n294080 , n294277 );
or ( n294313 , n3883 , n294312 );
xor ( n3886 , n838 , n294313 );
not ( n294315 , n293889 );
not ( n294316 , n293779 );
or ( n3889 , n294315 , n294316 );
buf ( n294318 , n293889 );
buf ( n294319 , n293779 );
or ( n3892 , n294318 , n294319 );
buf ( n294321 , n293821 );
nand ( n294322 , n3892 , n294321 );
buf ( n294323 , n294322 );
nand ( n3896 , n3889 , n294323 );
buf ( n294325 , n293920 );
not ( n294326 , n294325 );
xnor ( n294327 , n829 , n830 );
nand ( n3900 , n294327 , n1373 );
not ( n294329 , n3900 );
buf ( n294330 , n294329 );
not ( n3903 , n294330 );
or ( n294332 , n294326 , n3903 );
buf ( n3905 , n1508 );
buf ( n294334 , n776 );
buf ( n294335 , n828 );
xor ( n294336 , n294334 , n294335 );
buf ( n294337 , n294336 );
buf ( n294338 , n294337 );
nand ( n294339 , n3905 , n294338 );
buf ( n294340 , n294339 );
buf ( n294341 , n294340 );
nand ( n294342 , n294332 , n294341 );
buf ( n294343 , n294342 );
buf ( n294344 , n294343 );
or ( n3917 , n799 , n807 );
nand ( n3918 , n3917 , n808 );
buf ( n294347 , n3918 );
buf ( n294348 , n799 );
buf ( n294349 , n807 );
nand ( n3922 , n294348 , n294349 );
buf ( n294351 , n3922 );
buf ( n294352 , n294351 );
buf ( n294353 , n806 );
nand ( n3926 , n294347 , n294352 , n294353 );
buf ( n294355 , n3926 );
buf ( n294356 , n294355 );
and ( n294357 , n294344 , n294356 );
not ( n3930 , n294344 );
buf ( n294359 , n294355 );
not ( n294360 , n294359 );
buf ( n294361 , n294360 );
buf ( n294362 , n294361 );
and ( n294363 , n3930 , n294362 );
nor ( n3936 , n294357 , n294363 );
buf ( n3937 , n3936 );
not ( n294366 , n3937 );
buf ( n294367 , n293981 );
buf ( n294368 , n293962 );
or ( n294369 , n294367 , n294368 );
buf ( n294370 , n293999 );
nand ( n3943 , n294369 , n294370 );
buf ( n294372 , n3943 );
buf ( n294373 , n294372 );
buf ( n294374 , n293962 );
buf ( n294375 , n293981 );
nand ( n294376 , n294374 , n294375 );
buf ( n294377 , n294376 );
buf ( n294378 , n294377 );
nand ( n294379 , n294373 , n294378 );
buf ( n294380 , n294379 );
not ( n3953 , n294380 );
or ( n294382 , n294366 , n3953 );
buf ( n3955 , n294380 );
not ( n294384 , n3955 );
buf ( n294385 , n294384 );
buf ( n294386 , n3937 );
not ( n294387 , n294386 );
buf ( n294388 , n294387 );
nand ( n294389 , n294385 , n294388 );
nand ( n294390 , n294382 , n294389 );
or ( n3963 , n3637 , n294021 );
nand ( n294392 , n3963 , n294040 );
nand ( n294393 , n3637 , n294021 );
nand ( n3966 , n294392 , n294393 );
and ( n3967 , n294390 , n3966 );
not ( n294396 , n294390 );
not ( n3969 , n3966 );
and ( n294398 , n294396 , n3969 );
nor ( n294399 , n3967 , n294398 );
not ( n3972 , n294399 );
xor ( n3973 , n3896 , n3972 );
buf ( n294402 , n294012 );
not ( n3975 , n294402 );
nand ( n3976 , n292700 , n3591 );
not ( n3977 , n3976 );
buf ( n294406 , n3977 );
not ( n294407 , n294406 );
or ( n3980 , n3975 , n294407 );
buf ( n294409 , n1712 );
buf ( n3982 , n788 );
buf ( n294411 , n816 );
xor ( n294412 , n3982 , n294411 );
buf ( n294413 , n294412 );
buf ( n294414 , n294413 );
nand ( n294415 , n294409 , n294414 );
buf ( n294416 , n294415 );
buf ( n294417 , n294416 );
nand ( n3990 , n3980 , n294417 );
buf ( n294419 , n3990 );
buf ( n294420 , n294419 );
buf ( n294421 , n294034 );
not ( n3994 , n294421 );
buf ( n294423 , n2893 );
not ( n294424 , n294423 );
or ( n294425 , n3994 , n294424 );
buf ( n294426 , n2089 );
buf ( n294427 , n790 );
buf ( n4000 , n814 );
xor ( n4001 , n294427 , n4000 );
buf ( n4002 , n4001 );
buf ( n294431 , n4002 );
nand ( n4004 , n294426 , n294431 );
buf ( n294433 , n4004 );
buf ( n294434 , n294433 );
nand ( n4007 , n294425 , n294434 );
buf ( n294436 , n4007 );
buf ( n294437 , n294436 );
xor ( n4010 , n294420 , n294437 );
buf ( n294439 , n293936 );
not ( n294440 , n294439 );
buf ( n294441 , n291838 );
not ( n4014 , n294441 );
or ( n294443 , n294440 , n4014 );
buf ( n294444 , n292870 );
buf ( n294445 , n780 );
buf ( n294446 , n824 );
xor ( n4019 , n294445 , n294446 );
buf ( n4020 , n4019 );
buf ( n294449 , n4020 );
nand ( n294450 , n294444 , n294449 );
buf ( n294451 , n294450 );
buf ( n294452 , n294451 );
nand ( n294453 , n294443 , n294452 );
buf ( n294454 , n294453 );
buf ( n294455 , n294454 );
xor ( n294456 , n4010 , n294455 );
buf ( n294457 , n294456 );
not ( n4030 , n294059 );
and ( n4031 , n1338 , n291757 );
not ( n294460 , n4031 );
or ( n4033 , n4030 , n294460 );
buf ( n294462 , n292104 );
buf ( n4035 , n782 );
buf ( n294464 , n822 );
xor ( n294465 , n4035 , n294464 );
buf ( n294466 , n294465 );
buf ( n294467 , n294466 );
nand ( n4040 , n294462 , n294467 );
buf ( n294469 , n4040 );
nand ( n4042 , n4033 , n294469 );
not ( n4043 , n4042 );
buf ( n294472 , n293974 );
not ( n294473 , n294472 );
buf ( n294474 , n2373 );
not ( n4047 , n294474 );
or ( n294476 , n294473 , n4047 );
xor ( n4049 , n812 , n792 );
buf ( n294478 , n4049 );
not ( n294479 , n2381 );
buf ( n294480 , n294479 );
nand ( n294481 , n294478 , n294480 );
buf ( n294482 , n294481 );
buf ( n294483 , n294482 );
nand ( n294484 , n294476 , n294483 );
buf ( n294485 , n294484 );
not ( n294486 , n294485 );
or ( n294487 , n4043 , n294486 );
not ( n4060 , n294485 );
buf ( n294489 , n4042 );
not ( n294490 , n294489 );
buf ( n294491 , n294490 );
nand ( n4064 , n4060 , n294491 );
nand ( n294493 , n294487 , n4064 );
buf ( n294494 , n293993 );
not ( n4067 , n294494 );
buf ( n294496 , n293058 );
not ( n294497 , n294496 );
or ( n294498 , n4067 , n294497 );
buf ( n294499 , n292841 );
buf ( n294500 , n794 );
buf ( n4073 , n810 );
xor ( n4074 , n294500 , n4073 );
buf ( n4075 , n4074 );
buf ( n294504 , n4075 );
nand ( n4077 , n294499 , n294504 );
buf ( n4078 , n4077 );
buf ( n294507 , n4078 );
nand ( n4080 , n294498 , n294507 );
buf ( n294509 , n4080 );
not ( n4082 , n294509 );
and ( n294511 , n294493 , n4082 );
not ( n4084 , n294493 );
and ( n4085 , n4084 , n294509 );
nor ( n294514 , n294511 , n4085 );
not ( n294515 , n294514 );
xor ( n294516 , n294457 , n294515 );
buf ( n294517 , n293955 );
not ( n294518 , n294517 );
buf ( n294519 , n1933 );
not ( n4092 , n294519 );
or ( n294521 , n294518 , n4092 );
buf ( n294522 , n774 );
buf ( n294523 , n830 );
xor ( n294524 , n294522 , n294523 );
buf ( n294525 , n294524 );
buf ( n294526 , n294525 );
buf ( n294527 , n831 );
nand ( n294528 , n294526 , n294527 );
buf ( n294529 , n294528 );
buf ( n294530 , n294529 );
nand ( n294531 , n294521 , n294530 );
buf ( n294532 , n294531 );
buf ( n294533 , n294532 );
buf ( n294534 , n293880 );
not ( n4107 , n294534 );
buf ( n294536 , n292668 );
not ( n294537 , n294536 );
or ( n294538 , n4107 , n294537 );
buf ( n294539 , n291734 );
buf ( n294540 , n784 );
buf ( n294541 , n820 );
xor ( n4114 , n294540 , n294541 );
buf ( n294543 , n4114 );
buf ( n294544 , n294543 );
nand ( n4117 , n294539 , n294544 );
buf ( n294546 , n4117 );
buf ( n294547 , n294546 );
nand ( n294548 , n294538 , n294547 );
buf ( n294549 , n294548 );
buf ( n294550 , n294549 );
xor ( n4123 , n294533 , n294550 );
buf ( n294552 , n293843 );
not ( n294553 , n294552 );
buf ( n294554 , n293655 );
not ( n294555 , n294554 );
or ( n4128 , n294553 , n294555 );
buf ( n294557 , n293649 );
buf ( n294558 , n294557 );
buf ( n294559 , n796 );
buf ( n294560 , n808 );
xor ( n294561 , n294559 , n294560 );
buf ( n294562 , n294561 );
buf ( n294563 , n294562 );
nand ( n4136 , n294558 , n294563 );
buf ( n294565 , n4136 );
buf ( n294566 , n294565 );
nand ( n294567 , n4128 , n294566 );
buf ( n294568 , n294567 );
buf ( n294569 , n294568 );
not ( n4142 , n294569 );
xor ( n294571 , n4123 , n4142 );
buf ( n294572 , n294571 );
xor ( n4145 , n294516 , n294572 );
xnor ( n294574 , n3973 , n4145 );
buf ( n4147 , n294574 );
xor ( n4148 , n294148 , n294234 );
and ( n294577 , n4148 , n294275 );
and ( n4150 , n294148 , n294234 );
or ( n4151 , n294577 , n4150 );
buf ( n294580 , n4151 );
buf ( n294581 , n294580 );
xor ( n4154 , n4147 , n294581 );
xor ( n294583 , n294161 , n3764 );
and ( n4156 , n294583 , n294231 );
and ( n294585 , n294161 , n3764 );
or ( n4158 , n4156 , n294585 );
buf ( n294587 , n4158 );
xor ( n4160 , n294210 , n294212 );
and ( n4161 , n4160 , n294228 );
and ( n4162 , n294210 , n294212 );
or ( n294591 , n4161 , n4162 );
buf ( n294592 , n294591 );
buf ( n294593 , n294005 );
not ( n294594 , n294593 );
buf ( n294595 , n3643 );
not ( n4168 , n294595 );
or ( n294597 , n294594 , n4168 );
buf ( n294598 , n294002 );
not ( n294599 , n294598 );
buf ( n294600 , n294068 );
not ( n4173 , n294600 );
or ( n4174 , n294599 , n4173 );
buf ( n294603 , n293945 );
nand ( n294604 , n4174 , n294603 );
buf ( n294605 , n294604 );
buf ( n294606 , n294605 );
nand ( n294607 , n294597 , n294606 );
buf ( n294608 , n294607 );
xor ( n294609 , n294592 , n294608 );
xor ( n4182 , n293851 , n293868 );
and ( n294611 , n4182 , n293887 );
and ( n4184 , n293851 , n293868 );
or ( n4185 , n294611 , n4184 );
buf ( n294614 , n4185 );
xor ( n294615 , n293907 , n293925 );
and ( n294616 , n294615 , n293943 );
and ( n4189 , n293907 , n293925 );
or ( n294618 , n294616 , n4189 );
buf ( n294619 , n294618 );
and ( n4192 , n294614 , n294619 );
not ( n294621 , n294614 );
buf ( n294622 , n294619 );
not ( n4195 , n294622 );
buf ( n4196 , n4195 );
and ( n294625 , n294621 , n4196 );
nor ( n4198 , n4192 , n294625 );
buf ( n294627 , n799 );
buf ( n294628 , n806 );
xor ( n4201 , n294627 , n294628 );
buf ( n294630 , n4201 );
not ( n294631 , n294630 );
not ( n294632 , n807 );
nand ( n4205 , n294632 , n808 );
xor ( n294634 , n806 , n807 );
not ( n294635 , n808 );
nand ( n4208 , n294635 , n807 );
and ( n294637 , n4205 , n294634 , n4208 );
not ( n294638 , n294637 );
or ( n4211 , n294631 , n294638 );
buf ( n294640 , n293902 );
buf ( n294641 , n798 );
buf ( n294642 , n806 );
xor ( n4215 , n294641 , n294642 );
buf ( n294644 , n4215 );
buf ( n294645 , n294644 );
nand ( n294646 , n294640 , n294645 );
buf ( n294647 , n294646 );
nand ( n4220 , n4211 , n294647 );
not ( n294649 , n4220 );
buf ( n294650 , n293861 );
not ( n294651 , n294650 );
buf ( n294652 , n293394 );
not ( n4225 , n294652 );
or ( n294654 , n294651 , n4225 );
not ( n4227 , n292006 );
and ( n294656 , n778 , n826 );
not ( n4229 , n778 );
and ( n294658 , n4229 , n292463 );
nor ( n294659 , n294656 , n294658 );
nand ( n4232 , n4227 , n294659 );
buf ( n294661 , n4232 );
nand ( n294662 , n294654 , n294661 );
buf ( n294663 , n294662 );
and ( n4236 , n294649 , n294663 );
not ( n294665 , n294649 );
not ( n294666 , n294663 );
and ( n294667 , n294665 , n294666 );
nor ( n4240 , n4236 , n294667 );
buf ( n294669 , n786 );
buf ( n4242 , n818 );
xor ( n4243 , n294669 , n4242 );
buf ( n4244 , n4243 );
not ( n294673 , n4244 );
not ( n4246 , n291788 );
or ( n294675 , n294673 , n4246 );
nand ( n294676 , n291984 , n294203 );
nand ( n294677 , n294675 , n294676 );
and ( n4250 , n4240 , n294677 );
not ( n294679 , n4240 );
buf ( n294680 , n294677 );
not ( n4253 , n294680 );
buf ( n294682 , n4253 );
and ( n294683 , n294679 , n294682 );
or ( n294684 , n4250 , n294683 );
and ( n4257 , n4198 , n294684 );
not ( n294686 , n4198 );
and ( n294687 , n4240 , n294677 );
not ( n4260 , n4240 );
and ( n294689 , n4260 , n294682 );
nor ( n294690 , n294687 , n294689 );
buf ( n4263 , n294690 );
and ( n294692 , n294686 , n4263 );
nor ( n294693 , n4257 , n294692 );
xor ( n4266 , n294609 , n294693 );
xor ( n294695 , n294587 , n4266 );
buf ( n294696 , n3331 );
buf ( n294697 , n3469 );
or ( n4270 , n294696 , n294697 );
buf ( n294699 , n294074 );
nand ( n294700 , n4270 , n294699 );
buf ( n294701 , n294700 );
buf ( n294702 , n294701 );
buf ( n294703 , n3469 );
buf ( n294704 , n3331 );
nand ( n294705 , n294703 , n294704 );
buf ( n294706 , n294705 );
buf ( n294707 , n294706 );
nand ( n294708 , n294702 , n294707 );
buf ( n294709 , n294708 );
xor ( n294710 , n294695 , n294709 );
buf ( n294711 , n294710 );
xor ( n4284 , n4154 , n294711 );
buf ( n294713 , n4284 );
and ( n294714 , n3886 , n294713 );
and ( n294715 , n838 , n294313 );
or ( n4288 , n294714 , n294715 );
buf ( n294717 , n4288 );
not ( n294718 , n294717 );
or ( n294719 , n3175 , n294718 );
buf ( n294720 , n831 );
not ( n4293 , n294720 );
buf ( n294722 , n870 );
buf ( n294723 , n294713 );
xor ( n4296 , n294722 , n294723 );
buf ( n294725 , n294313 );
and ( n294726 , n4296 , n294725 );
and ( n294727 , n294722 , n294723 );
or ( n4300 , n294726 , n294727 );
buf ( n294729 , n4300 );
buf ( n294730 , n294729 );
nand ( n294731 , n4293 , n294730 );
buf ( n294732 , n294731 );
buf ( n294733 , n294732 );
nand ( n294734 , n294719 , n294733 );
buf ( n294735 , n294734 );
buf ( n294736 , n294735 );
buf ( n4309 , n294736 );
buf ( n294738 , n853 );
xor ( n4311 , n830 , n791 );
buf ( n294740 , n4311 );
not ( n4313 , n294740 );
buf ( n294742 , n1271 );
not ( n4315 , n294742 );
or ( n294744 , n4313 , n4315 );
buf ( n294745 , n790 );
buf ( n294746 , n830 );
xor ( n294747 , n294745 , n294746 );
buf ( n294748 , n294747 );
buf ( n294749 , n294748 );
buf ( n294750 , n831 );
nand ( n294751 , n294749 , n294750 );
buf ( n294752 , n294751 );
buf ( n294753 , n294752 );
nand ( n294754 , n294744 , n294753 );
buf ( n294755 , n294754 );
buf ( n294756 , n294755 );
xor ( n294757 , n822 , n799 );
buf ( n294758 , n294757 );
not ( n4331 , n294758 );
buf ( n294760 , n291761 );
not ( n294761 , n294760 );
or ( n4334 , n4331 , n294761 );
buf ( n294763 , n292105 );
xor ( n294764 , n822 , n798 );
buf ( n294765 , n294764 );
nand ( n294766 , n294763 , n294765 );
buf ( n294767 , n294766 );
buf ( n294768 , n294767 );
nand ( n294769 , n4334 , n294768 );
buf ( n294770 , n294769 );
buf ( n294771 , n294770 );
xor ( n294772 , n294756 , n294771 );
buf ( n4345 , n797 );
buf ( n294774 , n824 );
xor ( n294775 , n4345 , n294774 );
buf ( n294776 , n294775 );
buf ( n294777 , n294776 );
not ( n294778 , n294777 );
buf ( n294779 , n291838 );
not ( n294780 , n294779 );
or ( n294781 , n294778 , n294780 );
buf ( n294782 , n291842 );
xor ( n294783 , n824 , n796 );
buf ( n294784 , n294783 );
nand ( n4357 , n294782 , n294784 );
buf ( n294786 , n4357 );
buf ( n294787 , n294786 );
nand ( n294788 , n294781 , n294787 );
buf ( n294789 , n294788 );
buf ( n294790 , n294789 );
xor ( n4363 , n294772 , n294790 );
buf ( n294792 , n4363 );
not ( n294793 , n294792 );
buf ( n294794 , n793 );
buf ( n294795 , n830 );
xor ( n4368 , n294794 , n294795 );
buf ( n294797 , n4368 );
buf ( n294798 , n294797 );
not ( n4371 , n294798 );
buf ( n294800 , n291656 );
not ( n4373 , n294800 );
or ( n4374 , n4371 , n4373 );
buf ( n294803 , n831 );
xor ( n4376 , n830 , n792 );
buf ( n294805 , n4376 );
nand ( n4378 , n294803 , n294805 );
buf ( n294807 , n4378 );
buf ( n294808 , n294807 );
nand ( n4381 , n4374 , n294808 );
buf ( n294810 , n4381 );
buf ( n294811 , n799 );
buf ( n294812 , n825 );
or ( n4385 , n294811 , n294812 );
buf ( n294814 , n826 );
nand ( n294815 , n4385 , n294814 );
buf ( n294816 , n294815 );
buf ( n4389 , n294816 );
buf ( n294818 , n799 );
buf ( n294819 , n825 );
nand ( n294820 , n294818 , n294819 );
buf ( n294821 , n294820 );
buf ( n4394 , n294821 );
buf ( n294823 , n824 );
and ( n294824 , n4389 , n4394 , n294823 );
buf ( n294825 , n294824 );
and ( n4398 , n294810 , n294825 );
not ( n4399 , n291808 );
xor ( n294828 , n828 , n794 );
not ( n294829 , n294828 );
or ( n4402 , n4399 , n294829 );
buf ( n294831 , n291812 );
buf ( n294832 , n793 );
buf ( n294833 , n828 );
xor ( n294834 , n294832 , n294833 );
buf ( n294835 , n294834 );
buf ( n294836 , n294835 );
nand ( n294837 , n294831 , n294836 );
buf ( n294838 , n294837 );
nand ( n294839 , n4402 , n294838 );
xor ( n294840 , n4398 , n294839 );
buf ( n294841 , n796 );
buf ( n294842 , n826 );
xor ( n4415 , n294841 , n294842 );
buf ( n294844 , n4415 );
not ( n294845 , n294844 );
not ( n294846 , n1453 );
or ( n4419 , n294845 , n294846 );
buf ( n294848 , n291886 );
buf ( n294849 , n795 );
buf ( n294850 , n826 );
xor ( n294851 , n294849 , n294850 );
buf ( n294852 , n294851 );
buf ( n294853 , n294852 );
nand ( n4426 , n294848 , n294853 );
buf ( n294855 , n4426 );
nand ( n4428 , n4419 , n294855 );
and ( n4429 , n294840 , n4428 );
and ( n4430 , n4398 , n294839 );
or ( n4431 , n4429 , n4430 );
not ( n4432 , n4431 );
nand ( n294861 , n294793 , n4432 );
not ( n294862 , n294861 );
buf ( n294863 , n294852 );
not ( n4436 , n294863 );
buf ( n294865 , n1453 );
not ( n4438 , n294865 );
or ( n294867 , n4436 , n4438 );
buf ( n4440 , n1580 );
xor ( n294869 , n826 , n794 );
buf ( n294870 , n294869 );
nand ( n294871 , n4440 , n294870 );
buf ( n294872 , n294871 );
buf ( n294873 , n294872 );
nand ( n4446 , n294867 , n294873 );
buf ( n4447 , n4446 );
not ( n294876 , n291808 );
not ( n4449 , n294835 );
or ( n4450 , n294876 , n4449 );
buf ( n294879 , n291812 );
buf ( n294880 , n792 );
buf ( n294881 , n828 );
xor ( n4454 , n294880 , n294881 );
buf ( n294883 , n4454 );
buf ( n294884 , n294883 );
nand ( n294885 , n294879 , n294884 );
buf ( n294886 , n294885 );
nand ( n4459 , n4450 , n294886 );
buf ( n294888 , n799 );
buf ( n294889 , n823 );
or ( n294890 , n294888 , n294889 );
buf ( n294891 , n824 );
nand ( n4464 , n294890 , n294891 );
buf ( n294893 , n4464 );
buf ( n294894 , n294893 );
buf ( n294895 , n799 );
buf ( n294896 , n823 );
nand ( n4469 , n294895 , n294896 );
buf ( n294898 , n4469 );
buf ( n294899 , n294898 );
buf ( n294900 , n822 );
and ( n294901 , n294894 , n294899 , n294900 );
buf ( n294902 , n294901 );
not ( n4475 , n294902 );
and ( n294904 , n4459 , n4475 );
not ( n294905 , n4459 );
and ( n4478 , n294905 , n294902 );
nor ( n294907 , n294904 , n4478 );
xor ( n4480 , n4447 , n294907 );
buf ( n294909 , n292105 );
buf ( n294910 , n799 );
and ( n294911 , n294909 , n294910 );
buf ( n294912 , n294911 );
buf ( n294913 , n294912 );
buf ( n294914 , n291656 );
not ( n4487 , n294914 );
buf ( n294916 , n4376 );
not ( n294917 , n294916 );
or ( n294918 , n4487 , n294917 );
buf ( n294919 , n4311 );
buf ( n294920 , n831 );
nand ( n294921 , n294919 , n294920 );
buf ( n294922 , n294921 );
buf ( n294923 , n294922 );
nand ( n4496 , n294918 , n294923 );
buf ( n294925 , n4496 );
buf ( n294926 , n294925 );
xor ( n4499 , n294913 , n294926 );
buf ( n4500 , n798 );
buf ( n4501 , n824 );
xor ( n4502 , n4500 , n4501 );
buf ( n4503 , n4502 );
buf ( n294932 , n4503 );
not ( n4505 , n294932 );
buf ( n294934 , n291838 );
not ( n294935 , n294934 );
or ( n4508 , n4505 , n294935 );
buf ( n4509 , n292870 );
buf ( n4510 , n294776 );
nand ( n4511 , n4509 , n4510 );
buf ( n4512 , n4511 );
buf ( n294941 , n4512 );
nand ( n4514 , n4508 , n294941 );
buf ( n294943 , n4514 );
buf ( n294944 , n294943 );
and ( n4517 , n4499 , n294944 );
and ( n294946 , n294913 , n294926 );
or ( n294947 , n4517 , n294946 );
buf ( n294948 , n294947 );
xnor ( n294949 , n4480 , n294948 );
not ( n294950 , n294949 );
or ( n4523 , n294862 , n294950 );
nand ( n294952 , n294792 , n4431 );
nand ( n294953 , n4523 , n294952 );
buf ( n294954 , n294953 );
xor ( n4527 , n294738 , n294954 );
buf ( n294956 , n294748 );
not ( n294957 , n294956 );
buf ( n294958 , n1271 );
not ( n4531 , n294958 );
or ( n4532 , n294957 , n4531 );
buf ( n294961 , n1667 );
buf ( n294962 , n831 );
nand ( n294963 , n294961 , n294962 );
buf ( n294964 , n294963 );
buf ( n294965 , n294964 );
nand ( n4538 , n4532 , n294965 );
buf ( n294967 , n4538 );
buf ( n294968 , n294967 );
buf ( n294969 , n294764 );
not ( n4542 , n294969 );
buf ( n294971 , n291761 );
not ( n4544 , n294971 );
or ( n4545 , n4542 , n4544 );
buf ( n294974 , n292108 );
buf ( n294975 , n292105 );
nand ( n4548 , n294974 , n294975 );
buf ( n294977 , n4548 );
buf ( n294978 , n294977 );
nand ( n4551 , n4545 , n294978 );
buf ( n294980 , n4551 );
buf ( n294981 , n294980 );
xor ( n4554 , n294968 , n294981 );
buf ( n294983 , n1453 );
buf ( n294984 , n294869 );
nand ( n4557 , n294983 , n294984 );
buf ( n294986 , n4557 );
buf ( n4559 , n294986 );
buf ( n294988 , n1580 );
buf ( n294989 , n1442 );
nand ( n294990 , n294988 , n294989 );
buf ( n294991 , n294990 );
buf ( n294992 , n294991 );
nand ( n4565 , n4559 , n294992 );
buf ( n294994 , n4565 );
buf ( n294995 , n294994 );
xor ( n294996 , n4554 , n294995 );
buf ( n294997 , n294996 );
not ( n294998 , n294907 );
not ( n294999 , n294998 );
not ( n4572 , n4447 );
or ( n4573 , n294999 , n4572 );
not ( n295002 , n294907 );
not ( n295003 , n4447 );
not ( n4576 , n295003 );
or ( n295005 , n295002 , n4576 );
nand ( n295006 , n295005 , n294948 );
nand ( n4579 , n4573 , n295006 );
xor ( n295008 , n294997 , n4579 );
and ( n4581 , n4459 , n294902 );
xor ( n4582 , n294756 , n294771 );
and ( n295011 , n4582 , n294790 );
and ( n295012 , n294756 , n294771 );
or ( n4585 , n295011 , n295012 );
buf ( n295014 , n4585 );
xor ( n4587 , n4581 , n295014 );
buf ( n295016 , n291906 );
buf ( n295017 , n799 );
and ( n295018 , n295016 , n295017 );
buf ( n295019 , n295018 );
buf ( n295020 , n295019 );
buf ( n295021 , n294883 );
not ( n295022 , n295021 );
buf ( n295023 , n291808 );
not ( n295024 , n295023 );
or ( n295025 , n295022 , n295024 );
buf ( n295026 , n291939 );
buf ( n295027 , n291930 );
nand ( n295028 , n295026 , n295027 );
buf ( n295029 , n295028 );
buf ( n295030 , n295029 );
nand ( n4603 , n295025 , n295030 );
buf ( n295032 , n4603 );
buf ( n295033 , n295032 );
xor ( n295034 , n295020 , n295033 );
buf ( n295035 , n294783 );
not ( n295036 , n295035 );
buf ( n295037 , n291838 );
not ( n4610 , n295037 );
or ( n295039 , n295036 , n4610 );
buf ( n295040 , n291843 );
buf ( n295041 , n292112 );
nand ( n295042 , n295040 , n295041 );
buf ( n295043 , n295042 );
buf ( n295044 , n295043 );
nand ( n295045 , n295039 , n295044 );
buf ( n295046 , n295045 );
buf ( n295047 , n295046 );
xor ( n295048 , n295034 , n295047 );
buf ( n295049 , n295048 );
xor ( n4622 , n4587 , n295049 );
xor ( n295051 , n295008 , n4622 );
buf ( n295052 , n295051 );
and ( n4625 , n4527 , n295052 );
and ( n295054 , n294738 , n294954 );
or ( n295055 , n4625 , n295054 );
buf ( n295056 , n295055 );
and ( n295057 , n831 , n295056 );
not ( n4630 , n831 );
buf ( n295059 , n885 );
buf ( n295060 , n294953 );
xor ( n295061 , n295059 , n295060 );
buf ( n295062 , n295051 );
and ( n295063 , n295061 , n295062 );
and ( n295064 , n295059 , n295060 );
or ( n4637 , n295063 , n295064 );
buf ( n295066 , n4637 );
and ( n295067 , n4630 , n295066 );
or ( n4640 , n295057 , n295067 );
buf ( n4641 , n4640 );
buf ( n295070 , n854 );
buf ( n295071 , n797 );
buf ( n295072 , n826 );
xor ( n295073 , n295071 , n295072 );
buf ( n295074 , n295073 );
not ( n4647 , n295074 );
not ( n295076 , n291880 );
or ( n295077 , n4647 , n295076 );
buf ( n295078 , n1579 );
buf ( n295079 , n294844 );
nand ( n4652 , n295078 , n295079 );
buf ( n295081 , n4652 );
nand ( n295082 , n295077 , n295081 );
xor ( n295083 , n824 , n799 );
buf ( n295084 , n295083 );
not ( n295085 , n295084 );
buf ( n295086 , n291838 );
not ( n4659 , n295086 );
or ( n295088 , n295085 , n4659 );
buf ( n295089 , n292870 );
buf ( n295090 , n4503 );
nand ( n295091 , n295089 , n295090 );
buf ( n295092 , n295091 );
buf ( n295093 , n295092 );
nand ( n295094 , n295088 , n295093 );
buf ( n295095 , n295094 );
xor ( n295096 , n295082 , n295095 );
buf ( n295097 , n795 );
buf ( n295098 , n828 );
xor ( n295099 , n295097 , n295098 );
buf ( n295100 , n295099 );
buf ( n295101 , n295100 );
not ( n295102 , n295101 );
buf ( n295103 , n291808 );
not ( n4676 , n295103 );
or ( n295105 , n295102 , n4676 );
buf ( n295106 , n291939 );
buf ( n295107 , n294828 );
nand ( n295108 , n295106 , n295107 );
buf ( n295109 , n295108 );
buf ( n295110 , n295109 );
nand ( n295111 , n295105 , n295110 );
buf ( n295112 , n295111 );
and ( n295113 , n295096 , n295112 );
and ( n295114 , n295082 , n295095 );
or ( n4687 , n295113 , n295114 );
xor ( n295116 , n294913 , n294926 );
xor ( n295117 , n295116 , n294944 );
buf ( n295118 , n295117 );
or ( n295119 , n4687 , n295118 );
xor ( n4692 , n4398 , n294839 );
xor ( n4693 , n4692 , n4428 );
nand ( n295122 , n295119 , n4693 );
nand ( n295123 , n295118 , n4687 );
nand ( n4696 , n295122 , n295123 );
buf ( n295125 , n4696 );
xor ( n295126 , n295070 , n295125 );
and ( n4699 , n294792 , n4432 );
not ( n295128 , n294792 );
and ( n295129 , n295128 , n4431 );
or ( n4702 , n4699 , n295129 );
xor ( n4703 , n4702 , n294949 );
buf ( n295132 , n4703 );
and ( n4705 , n295126 , n295132 );
and ( n295134 , n295070 , n295125 );
or ( n295135 , n4705 , n295134 );
buf ( n295136 , n295135 );
and ( n295137 , n831 , n295136 );
not ( n4710 , n831 );
buf ( n295139 , n886 );
buf ( n295140 , n4696 );
xor ( n4713 , n295139 , n295140 );
buf ( n295142 , n4703 );
and ( n4715 , n4713 , n295142 );
and ( n295144 , n295139 , n295140 );
or ( n4717 , n4715 , n295144 );
buf ( n295146 , n4717 );
and ( n4719 , n4710 , n295146 );
or ( n295148 , n295137 , n4719 );
buf ( n4721 , n295148 );
buf ( n295150 , n4721 );
buf ( n295151 , n831 );
not ( n295152 , n295151 );
buf ( n295153 , n835 );
not ( n4726 , n3937 );
not ( n295155 , n294385 );
or ( n295156 , n4726 , n295155 );
nand ( n4729 , n295156 , n3966 );
buf ( n295158 , n4729 );
buf ( n295159 , n294380 );
buf ( n295160 , n294388 );
nand ( n4733 , n295159 , n295160 );
buf ( n295162 , n4733 );
buf ( n295163 , n295162 );
nand ( n295164 , n295158 , n295163 );
buf ( n295165 , n295164 );
buf ( n295166 , n295165 );
not ( n4739 , n294619 );
not ( n4740 , n294684 );
or ( n295169 , n4739 , n4740 );
not ( n4742 , n4196 );
not ( n295171 , n294690 );
or ( n4744 , n4742 , n295171 );
nand ( n295173 , n4744 , n294614 );
nand ( n4746 , n295169 , n295173 );
buf ( n295175 , n4746 );
xor ( n295176 , n295166 , n295175 );
not ( n295177 , n294572 );
not ( n4750 , n294515 );
or ( n4751 , n295177 , n4750 );
nand ( n295180 , n4751 , n294457 );
buf ( n295181 , n295180 );
not ( n295182 , n294572 );
nand ( n4755 , n295182 , n294514 );
buf ( n295184 , n4755 );
nand ( n4757 , n295181 , n295184 );
buf ( n295186 , n4757 );
buf ( n295187 , n295186 );
xor ( n4760 , n295176 , n295187 );
buf ( n295189 , n4760 );
not ( n4762 , n295189 );
xor ( n295191 , n294592 , n294608 );
and ( n4764 , n295191 , n294693 );
and ( n295193 , n294592 , n294608 );
or ( n4766 , n4764 , n295193 );
not ( n4767 , n4766 );
or ( n4768 , n4762 , n4767 );
or ( n295197 , n295189 , n4766 );
not ( n4770 , n294399 );
not ( n4771 , n3896 );
nand ( n4772 , n4770 , n4771 );
not ( n4773 , n4772 );
not ( n4774 , n4145 );
or ( n295203 , n4773 , n4774 );
nand ( n4776 , n294399 , n3896 );
nand ( n295205 , n295203 , n4776 );
nand ( n295206 , n295197 , n295205 );
nand ( n4779 , n4768 , n295206 );
not ( n295208 , n4779 );
not ( n4781 , n294659 );
nand ( n295210 , n826 , n827 );
not ( n4783 , n826 );
not ( n295212 , n827 );
nand ( n4785 , n4783 , n295212 );
nand ( n4786 , n295210 , n4785 );
nor ( n4787 , n4786 , n1445 );
not ( n4788 , n4787 );
or ( n4789 , n4781 , n4788 );
buf ( n295218 , n777 );
buf ( n295219 , n826 );
xor ( n4792 , n295218 , n295219 );
buf ( n295221 , n4792 );
nand ( n295222 , n295221 , n1579 );
nand ( n4795 , n4789 , n295222 );
buf ( n295224 , n4244 );
not ( n4797 , n295224 );
not ( n4798 , n291980 );
buf ( n295227 , n4798 );
not ( n295228 , n295227 );
or ( n4801 , n4797 , n295228 );
buf ( n295230 , n291988 );
buf ( n4803 , n295230 );
buf ( n295232 , n785 );
buf ( n295233 , n818 );
xor ( n295234 , n295232 , n295233 );
buf ( n295235 , n295234 );
buf ( n295236 , n295235 );
nand ( n295237 , n4803 , n295236 );
buf ( n295238 , n295237 );
buf ( n295239 , n295238 );
nand ( n295240 , n4801 , n295239 );
buf ( n295241 , n295240 );
xor ( n4814 , n4795 , n295241 );
buf ( n295243 , n294343 );
buf ( n4816 , n294361 );
and ( n4817 , n295243 , n4816 );
buf ( n295246 , n4817 );
and ( n4819 , n4814 , n295246 );
and ( n295248 , n4795 , n295241 );
or ( n4821 , n4819 , n295248 );
buf ( n295250 , n793 );
buf ( n295251 , n810 );
xor ( n295252 , n295250 , n295251 );
buf ( n295253 , n295252 );
buf ( n295254 , n295253 );
not ( n295255 , n295254 );
buf ( n295256 , n293058 );
not ( n295257 , n295256 );
or ( n4830 , n295255 , n295257 );
xor ( n295259 , n811 , n812 );
buf ( n295260 , n295259 );
buf ( n295261 , n792 );
buf ( n295262 , n810 );
xor ( n4835 , n295261 , n295262 );
buf ( n295264 , n4835 );
buf ( n295265 , n295264 );
nand ( n4838 , n295260 , n295265 );
buf ( n295267 , n4838 );
buf ( n295268 , n295267 );
nand ( n4841 , n4830 , n295268 );
buf ( n4842 , n4841 );
buf ( n295271 , n4842 );
buf ( n295272 , n295271 );
and ( n4845 , n781 , n822 );
not ( n4846 , n781 );
and ( n295275 , n4846 , n1299 );
nor ( n4848 , n4845 , n295275 );
not ( n4849 , n4848 );
not ( n4850 , n292631 );
or ( n4851 , n4849 , n4850 );
buf ( n295280 , n292104 );
buf ( n4853 , n780 );
buf ( n295282 , n822 );
xor ( n4855 , n4853 , n295282 );
buf ( n295284 , n4855 );
buf ( n295285 , n295284 );
nand ( n295286 , n295280 , n295285 );
buf ( n295287 , n295286 );
nand ( n4860 , n4851 , n295287 );
buf ( n295289 , n791 );
buf ( n295290 , n812 );
xor ( n4863 , n295289 , n295290 );
buf ( n295292 , n4863 );
buf ( n295293 , n295292 );
not ( n4866 , n295293 );
buf ( n295295 , n2373 );
not ( n4868 , n295295 );
or ( n295297 , n4866 , n4868 );
buf ( n295298 , n294479 );
buf ( n295299 , n790 );
buf ( n295300 , n812 );
xor ( n295301 , n295299 , n295300 );
buf ( n295302 , n295301 );
buf ( n295303 , n295302 );
nand ( n4876 , n295298 , n295303 );
buf ( n295305 , n4876 );
buf ( n295306 , n295305 );
nand ( n295307 , n295297 , n295306 );
buf ( n295308 , n295307 );
xor ( n4881 , n4860 , n295308 );
buf ( n295310 , n4881 );
xor ( n4883 , n295272 , n295310 );
buf ( n295312 , n4883 );
xor ( n4885 , n4821 , n295312 );
not ( n4886 , n291788 );
buf ( n295315 , n784 );
buf ( n295316 , n818 );
xor ( n4889 , n295315 , n295316 );
buf ( n4890 , n4889 );
not ( n295319 , n4890 );
or ( n295320 , n4886 , n295319 );
nand ( n4893 , n4798 , n295235 );
nand ( n295322 , n295320 , n4893 );
not ( n4895 , n295322 );
buf ( n295324 , n799 );
buf ( n295325 , n805 );
or ( n4898 , n295324 , n295325 );
buf ( n295327 , n806 );
nand ( n4900 , n4898 , n295327 );
buf ( n295329 , n4900 );
buf ( n295330 , n295329 );
buf ( n295331 , n799 );
buf ( n295332 , n805 );
nand ( n295333 , n295331 , n295332 );
buf ( n295334 , n295333 );
buf ( n295335 , n295334 );
buf ( n295336 , n804 );
and ( n4909 , n295330 , n295335 , n295336 );
buf ( n295338 , n4909 );
xor ( n4911 , n828 , n775 );
buf ( n295340 , n4911 );
not ( n295341 , n295340 );
buf ( n295342 , n291805 );
not ( n4915 , n295342 );
or ( n295344 , n295341 , n4915 );
buf ( n295345 , n1508 );
xor ( n4918 , n828 , n774 );
buf ( n295347 , n4918 );
nand ( n4920 , n295345 , n295347 );
buf ( n295349 , n4920 );
buf ( n295350 , n295349 );
nand ( n295351 , n295344 , n295350 );
buf ( n295352 , n295351 );
xor ( n295353 , n295338 , n295352 );
and ( n295354 , n4895 , n295353 );
not ( n4927 , n4895 );
not ( n295356 , n295353 );
and ( n295357 , n4927 , n295356 );
nor ( n295358 , n295354 , n295357 );
not ( n295359 , n295358 );
xor ( n4932 , n805 , n806 );
buf ( n295361 , n4932 );
buf ( n295362 , n295361 );
buf ( n295363 , n799 );
and ( n295364 , n295362 , n295363 );
buf ( n295365 , n295364 );
buf ( n295366 , n294337 );
not ( n295367 , n295366 );
buf ( n295368 , n292168 );
not ( n4941 , n295368 );
or ( n295370 , n295367 , n4941 );
buf ( n295371 , n1508 );
buf ( n295372 , n4911 );
nand ( n295373 , n295371 , n295372 );
buf ( n295374 , n295373 );
buf ( n295375 , n295374 );
nand ( n4948 , n295370 , n295375 );
buf ( n295377 , n4948 );
xor ( n4950 , n295365 , n295377 );
buf ( n295379 , n4020 );
not ( n4952 , n295379 );
buf ( n295381 , n292473 );
not ( n4954 , n295381 );
or ( n295383 , n4952 , n4954 );
buf ( n295384 , n291843 );
and ( n295385 , n779 , n824 );
not ( n295386 , n779 );
not ( n4959 , n824 );
and ( n4960 , n295386 , n4959 );
nor ( n4961 , n295385 , n4960 );
buf ( n295390 , n4961 );
nand ( n295391 , n295384 , n295390 );
buf ( n295392 , n295391 );
buf ( n295393 , n295392 );
nand ( n295394 , n295383 , n295393 );
buf ( n295395 , n295394 );
and ( n295396 , n4950 , n295395 );
and ( n4969 , n295365 , n295377 );
or ( n295398 , n295396 , n4969 );
not ( n4971 , n295398 );
or ( n4972 , n295359 , n4971 );
or ( n295401 , n295358 , n295398 );
nand ( n295402 , n4972 , n295401 );
xor ( n4975 , n4885 , n295402 );
not ( n295404 , n4975 );
not ( n295405 , n295404 );
xor ( n4978 , n4795 , n295241 );
xor ( n295407 , n4978 , n295246 );
not ( n295408 , n294562 );
xor ( n4981 , n810 , n809 );
not ( n295410 , n3223 );
nor ( n4983 , n4981 , n295410 );
not ( n295412 , n4983 );
or ( n4985 , n295408 , n295412 );
buf ( n295414 , n3114 );
buf ( n4987 , n795 );
buf ( n4988 , n808 );
xor ( n4989 , n4987 , n4988 );
buf ( n4990 , n4989 );
buf ( n295419 , n4990 );
nand ( n4992 , n295414 , n295419 );
buf ( n4993 , n4992 );
nand ( n295422 , n4985 , n4993 );
buf ( n295423 , n294644 );
not ( n295424 , n295423 );
and ( n295425 , n808 , n807 );
not ( n4998 , n808 );
not ( n295427 , n807 );
and ( n295428 , n4998 , n295427 );
nor ( n5001 , n295425 , n295428 );
not ( n295430 , n5001 );
xor ( n5003 , n806 , n807 );
nand ( n5004 , n295430 , n5003 );
not ( n295433 , n5004 );
buf ( n295434 , n295433 );
not ( n5007 , n295434 );
or ( n295436 , n295424 , n5007 );
buf ( n295437 , n293902 );
buf ( n295438 , n295437 );
xor ( n295439 , n806 , n797 );
buf ( n295440 , n295439 );
nand ( n5013 , n295438 , n295440 );
buf ( n295442 , n5013 );
buf ( n295443 , n295442 );
nand ( n295444 , n295436 , n295443 );
buf ( n295445 , n295444 );
xor ( n5018 , n295422 , n295445 );
buf ( n295447 , n294543 );
not ( n5020 , n295447 );
buf ( n295449 , n291722 );
not ( n295450 , n295449 );
or ( n5023 , n5020 , n295450 );
buf ( n295452 , n291906 );
buf ( n295453 , n783 );
buf ( n295454 , n820 );
xor ( n295455 , n295453 , n295454 );
buf ( n295456 , n295455 );
buf ( n295457 , n295456 );
nand ( n295458 , n295452 , n295457 );
buf ( n295459 , n295458 );
buf ( n295460 , n295459 );
nand ( n5033 , n5023 , n295460 );
buf ( n5034 , n5033 );
xor ( n295463 , n5018 , n5034 );
xor ( n5036 , n295407 , n295463 );
buf ( n295465 , n4002 );
not ( n5038 , n295465 );
buf ( n295467 , n2893 );
not ( n295468 , n295467 );
or ( n295469 , n5038 , n295468 );
buf ( n295470 , n789 );
buf ( n295471 , n814 );
xor ( n295472 , n295470 , n295471 );
buf ( n295473 , n295472 );
buf ( n295474 , n295473 );
and ( n295475 , n816 , n815 );
not ( n5048 , n816 );
and ( n5049 , n5048 , n2086 );
nor ( n295478 , n295475 , n5049 );
buf ( n5051 , n295478 );
buf ( n295480 , n5051 );
nand ( n5053 , n295474 , n295480 );
buf ( n295482 , n5053 );
buf ( n295483 , n295482 );
nand ( n295484 , n295469 , n295483 );
buf ( n295485 , n295484 );
buf ( n295486 , n295485 );
not ( n295487 , n295486 );
buf ( n295488 , n294413 );
not ( n295489 , n295488 );
buf ( n295490 , n3977 );
not ( n5063 , n295490 );
or ( n5064 , n295489 , n5063 );
and ( n5065 , n816 , n787 );
not ( n295494 , n816 );
and ( n295495 , n295494 , n293379 );
nor ( n295496 , n5065 , n295495 );
nand ( n295497 , n295496 , n1712 );
buf ( n295498 , n295497 );
nand ( n295499 , n5064 , n295498 );
buf ( n295500 , n295499 );
buf ( n295501 , n295500 );
not ( n295502 , n295501 );
buf ( n295503 , n295502 );
buf ( n295504 , n295503 );
not ( n295505 , n295504 );
and ( n295506 , n295487 , n295505 );
buf ( n295507 , n295485 );
buf ( n295508 , n295503 );
and ( n295509 , n295507 , n295508 );
nor ( n5082 , n295506 , n295509 );
buf ( n5083 , n5082 );
not ( n295512 , n294466 );
not ( n295513 , n4031 );
or ( n295514 , n295512 , n295513 );
nand ( n5087 , n1339 , n4848 );
nand ( n295516 , n295514 , n5087 );
not ( n5089 , n295516 );
and ( n5090 , n5083 , n5089 );
not ( n5091 , n5083 );
and ( n5092 , n5091 , n295516 );
nor ( n5093 , n5090 , n5092 );
and ( n5094 , n5036 , n5093 );
and ( n295523 , n295407 , n295463 );
or ( n5096 , n5094 , n295523 );
not ( n5097 , n5096 );
not ( n5098 , n295496 );
not ( n5099 , n292892 );
or ( n5100 , n5098 , n5099 );
not ( n5101 , n292700 );
xor ( n5102 , n816 , n786 );
nand ( n5103 , n5101 , n5102 );
nand ( n5104 , n5100 , n5103 );
buf ( n295533 , n295473 );
not ( n5106 , n295533 );
buf ( n295535 , n2078 );
not ( n5108 , n295535 );
or ( n295537 , n5106 , n5108 );
buf ( n295538 , n5051 );
buf ( n295539 , n788 );
buf ( n295540 , n814 );
xor ( n5113 , n295539 , n295540 );
buf ( n295542 , n5113 );
buf ( n295543 , n295542 );
nand ( n5116 , n295538 , n295543 );
buf ( n295545 , n5116 );
buf ( n295546 , n295545 );
nand ( n295547 , n295537 , n295546 );
buf ( n295548 , n295547 );
not ( n5121 , n295548 );
xor ( n5122 , n5104 , n5121 );
not ( n5123 , n291842 );
buf ( n295552 , n778 );
buf ( n295553 , n824 );
xor ( n5126 , n295552 , n295553 );
buf ( n295555 , n5126 );
not ( n5128 , n295555 );
or ( n5129 , n5123 , n5128 );
not ( n295558 , n824 );
not ( n5131 , n2038 );
or ( n5132 , n295558 , n5131 );
nand ( n5133 , n5132 , n292470 );
not ( n295562 , n291842 );
nand ( n295563 , n4961 , n5133 , n295562 );
nand ( n5136 , n5129 , n295563 );
not ( n5137 , n5136 );
xor ( n5138 , n5122 , n5137 );
buf ( n295567 , n773 );
buf ( n5140 , n830 );
xor ( n5141 , n295567 , n5140 );
buf ( n295570 , n5141 );
buf ( n5143 , n295570 );
not ( n5144 , n5143 );
buf ( n295573 , n293454 );
not ( n5146 , n295573 );
or ( n295575 , n5144 , n5146 );
buf ( n295576 , n772 );
buf ( n295577 , n830 );
xor ( n295578 , n295576 , n295577 );
buf ( n295579 , n295578 );
buf ( n295580 , n295579 );
buf ( n295581 , n831 );
nand ( n295582 , n295580 , n295581 );
buf ( n295583 , n295582 );
buf ( n295584 , n295583 );
nand ( n5157 , n295575 , n295584 );
buf ( n295586 , n5157 );
buf ( n295587 , n295586 );
buf ( n295588 , n4990 );
not ( n295589 , n295588 );
buf ( n295590 , n3408 );
not ( n295591 , n295590 );
or ( n5164 , n295589 , n295591 );
buf ( n295593 , n3114 );
buf ( n295594 , n794 );
buf ( n295595 , n808 );
xor ( n295596 , n295594 , n295595 );
buf ( n295597 , n295596 );
buf ( n295598 , n295597 );
nand ( n5171 , n295593 , n295598 );
buf ( n295600 , n5171 );
buf ( n295601 , n295600 );
nand ( n295602 , n5164 , n295601 );
buf ( n295603 , n295602 );
buf ( n295604 , n295603 );
xor ( n5177 , n295587 , n295604 );
buf ( n295606 , n295456 );
not ( n5179 , n295606 );
buf ( n295608 , n2787 );
not ( n295609 , n295608 );
or ( n295610 , n5179 , n295609 );
buf ( n295611 , n291969 );
buf ( n295612 , n782 );
buf ( n295613 , n820 );
xor ( n295614 , n295612 , n295613 );
buf ( n295615 , n295614 );
buf ( n295616 , n295615 );
nand ( n295617 , n295611 , n295616 );
buf ( n295618 , n295617 );
buf ( n295619 , n295618 );
nand ( n295620 , n295610 , n295619 );
buf ( n295621 , n295620 );
buf ( n295622 , n295621 );
xnor ( n5195 , n5177 , n295622 );
buf ( n5196 , n5195 );
and ( n295625 , n5138 , n5196 );
not ( n5198 , n5138 );
buf ( n295627 , n5196 );
not ( n5200 , n295627 );
buf ( n295629 , n5200 );
and ( n295630 , n5198 , n295629 );
nor ( n295631 , n295625 , n295630 );
buf ( n295632 , n295631 );
not ( n295633 , n295439 );
not ( n295634 , n294637 );
or ( n5207 , n295633 , n295634 );
buf ( n295636 , n293902 );
xor ( n295637 , n806 , n796 );
buf ( n295638 , n295637 );
nand ( n295639 , n295636 , n295638 );
buf ( n295640 , n295639 );
nand ( n295641 , n5207 , n295640 );
not ( n5214 , n295221 );
and ( n295643 , n293392 , n2965 );
not ( n295644 , n295643 );
or ( n295645 , n5214 , n295644 );
not ( n295646 , n292006 );
buf ( n295647 , n776 );
buf ( n295648 , n826 );
xor ( n295649 , n295647 , n295648 );
buf ( n295650 , n295649 );
nand ( n5223 , n295646 , n295650 );
nand ( n295652 , n295645 , n5223 );
xor ( n295653 , n295641 , n295652 );
buf ( n5226 , n295653 );
xor ( n295655 , n799 , n804 );
not ( n5228 , n295655 );
xor ( n295657 , n804 , n805 );
not ( n295658 , n4932 );
nand ( n5231 , n295657 , n295658 );
not ( n295660 , n5231 );
not ( n5233 , n295660 );
or ( n5234 , n5228 , n5233 );
buf ( n5235 , n798 );
buf ( n5236 , n804 );
xor ( n5237 , n5235 , n5236 );
buf ( n5238 , n5237 );
nand ( n295667 , n5238 , n295361 );
nand ( n5240 , n5234 , n295667 );
buf ( n295669 , n5240 );
xnor ( n295670 , n5226 , n295669 );
buf ( n295671 , n295670 );
buf ( n295672 , n295671 );
buf ( n295673 , n295672 );
buf ( n295674 , n295673 );
buf ( n5247 , n295674 );
not ( n295676 , n5247 );
buf ( n295677 , n295676 );
buf ( n295678 , n295677 );
and ( n295679 , n295632 , n295678 );
not ( n5252 , n295632 );
buf ( n295681 , n295674 );
and ( n5254 , n5252 , n295681 );
nor ( n5255 , n295679 , n5254 );
buf ( n295684 , n5255 );
buf ( n295685 , n295684 );
not ( n5258 , n295685 );
buf ( n5259 , n5258 );
not ( n295688 , n5259 );
or ( n5261 , n5097 , n295688 );
not ( n295690 , n5096 );
nand ( n295691 , n295690 , n295684 );
nand ( n5264 , n5261 , n295691 );
nand ( n295693 , n295405 , n5264 );
not ( n5266 , n295693 );
not ( n295695 , n295404 );
nor ( n5268 , n5264 , n295695 );
nor ( n5269 , n5266 , n5268 );
nand ( n295698 , n295208 , n5269 );
not ( n5271 , n295698 );
buf ( n295700 , n294568 );
buf ( n295701 , n294532 );
or ( n295702 , n295700 , n295701 );
buf ( n295703 , n294549 );
nand ( n295704 , n295702 , n295703 );
buf ( n295705 , n295704 );
buf ( n295706 , n295705 );
buf ( n295707 , n294568 );
buf ( n5280 , n294532 );
nand ( n5281 , n295707 , n5280 );
buf ( n295710 , n5281 );
buf ( n295711 , n295710 );
nand ( n5284 , n295706 , n295711 );
buf ( n295713 , n5284 );
buf ( n295714 , n295713 );
not ( n5287 , n295714 );
buf ( n295716 , n5287 );
buf ( n295717 , n295716 );
not ( n5290 , n295717 );
not ( n295719 , n4042 );
not ( n295720 , n294485 );
or ( n5293 , n295719 , n295720 );
or ( n295722 , n4042 , n294485 );
nand ( n295723 , n295722 , n294509 );
nand ( n5296 , n5293 , n295723 );
not ( n5297 , n5296 );
buf ( n295726 , n5297 );
not ( n295727 , n295726 );
or ( n295728 , n5290 , n295727 );
xor ( n5301 , n294420 , n294437 );
and ( n5302 , n5301 , n294455 );
and ( n5303 , n294420 , n294437 );
or ( n295732 , n5302 , n5303 );
buf ( n295733 , n295732 );
buf ( n295734 , n295733 );
nand ( n5307 , n295728 , n295734 );
buf ( n295736 , n5307 );
nand ( n295737 , n295713 , n5296 );
nand ( n5310 , n295736 , n295737 );
not ( n5311 , n5310 );
buf ( n295740 , n294677 );
not ( n295741 , n295740 );
buf ( n295742 , n294663 );
not ( n5315 , n295742 );
or ( n5316 , n295741 , n5315 );
buf ( n295745 , n294677 );
buf ( n295746 , n294663 );
or ( n5319 , n295745 , n295746 );
buf ( n5320 , n4220 );
buf ( n295749 , n5320 );
nand ( n295750 , n5319 , n295749 );
buf ( n295751 , n295750 );
buf ( n295752 , n295751 );
nand ( n5325 , n5316 , n295752 );
buf ( n295754 , n5325 );
not ( n295755 , n295754 );
xor ( n295756 , n295365 , n295377 );
xor ( n5329 , n295756 , n295395 );
not ( n5330 , n5329 );
or ( n5331 , n295755 , n5330 );
buf ( n295760 , n295754 );
buf ( n295761 , n5329 );
or ( n5334 , n295760 , n295761 );
buf ( n295763 , n293454 );
not ( n5336 , n295763 );
buf ( n295765 , n294525 );
not ( n5338 , n295765 );
or ( n5339 , n5336 , n5338 );
buf ( n5340 , n295570 );
buf ( n5341 , n831 );
nand ( n5342 , n5340 , n5341 );
buf ( n5343 , n5342 );
buf ( n295772 , n5343 );
nand ( n5345 , n5339 , n295772 );
buf ( n295774 , n5345 );
buf ( n295775 , n295774 );
not ( n5348 , n4049 );
not ( n295777 , n3539 );
or ( n295778 , n5348 , n295777 );
buf ( n295779 , n2026 );
buf ( n295780 , n295292 );
nand ( n295781 , n295779 , n295780 );
buf ( n295782 , n295781 );
nand ( n295783 , n295778 , n295782 );
buf ( n295784 , n295783 );
xor ( n295785 , n295775 , n295784 );
buf ( n295786 , n4075 );
not ( n5359 , n295786 );
buf ( n295788 , n293058 );
not ( n295789 , n295788 );
or ( n5362 , n5359 , n295789 );
buf ( n295791 , n292841 );
buf ( n295792 , n295253 );
nand ( n5365 , n295791 , n295792 );
buf ( n295794 , n5365 );
buf ( n295795 , n295794 );
nand ( n5368 , n5362 , n295795 );
buf ( n5369 , n5368 );
buf ( n295798 , n5369 );
xor ( n5371 , n295785 , n295798 );
buf ( n295800 , n5371 );
buf ( n295801 , n295800 );
nand ( n5374 , n5334 , n295801 );
buf ( n295803 , n5374 );
nand ( n295804 , n5331 , n295803 );
not ( n295805 , n295804 );
or ( n5378 , n5311 , n295805 );
not ( n295807 , n5310 );
not ( n295808 , n295804 );
nand ( n5381 , n295807 , n295808 );
nand ( n295810 , n5378 , n5381 );
nand ( n5383 , n295516 , n295500 );
not ( n5384 , n5089 );
not ( n295813 , n295503 );
or ( n295814 , n5384 , n295813 );
nand ( n5387 , n295814 , n295485 );
nand ( n295816 , n5383 , n5387 );
xor ( n295817 , n295775 , n295784 );
and ( n5390 , n295817 , n295798 );
and ( n295819 , n295775 , n295784 );
or ( n295820 , n5390 , n295819 );
buf ( n295821 , n295820 );
and ( n295822 , n295816 , n295821 );
not ( n5395 , n295816 );
buf ( n295824 , n295821 );
not ( n5397 , n295824 );
buf ( n295826 , n5397 );
and ( n295827 , n5395 , n295826 );
nor ( n295828 , n295822 , n295827 );
xor ( n5401 , n295422 , n295445 );
and ( n295830 , n5401 , n5034 );
and ( n295831 , n295422 , n295445 );
or ( n5404 , n295830 , n295831 );
buf ( n295833 , n5404 );
not ( n295834 , n295833 );
and ( n5407 , n295828 , n295834 );
not ( n295836 , n295828 );
and ( n295837 , n295836 , n295833 );
nor ( n5410 , n5407 , n295837 );
buf ( n295839 , n5410 );
not ( n295840 , n295839 );
and ( n5413 , n295810 , n295840 );
not ( n295842 , n295810 );
and ( n5415 , n295842 , n295839 );
nor ( n5416 , n5413 , n5415 );
buf ( n5417 , n5416 );
not ( n295846 , n5417 );
buf ( n295847 , n295846 );
not ( n295848 , n295847 );
buf ( n295849 , n295716 );
not ( n5422 , n295849 );
buf ( n295851 , n5296 );
not ( n295852 , n295851 );
and ( n5425 , n5422 , n295852 );
buf ( n295854 , n5296 );
buf ( n295855 , n295716 );
and ( n295856 , n295854 , n295855 );
nor ( n5429 , n5425 , n295856 );
buf ( n295858 , n5429 );
buf ( n295859 , n295733 );
not ( n295860 , n295859 );
buf ( n295861 , n295860 );
and ( n5434 , n295858 , n295861 );
not ( n5435 , n295858 );
and ( n5436 , n5435 , n295733 );
nor ( n5437 , n5434 , n5436 );
buf ( n295866 , n5437 );
not ( n5439 , n295866 );
xor ( n5440 , n295407 , n295463 );
xor ( n5441 , n5440 , n5093 );
buf ( n295870 , n5441 );
not ( n5443 , n295870 );
or ( n5444 , n5439 , n5443 );
buf ( n295873 , n5441 );
buf ( n295874 , n5437 );
or ( n5447 , n295873 , n295874 );
xor ( n5448 , n295754 , n295800 );
xor ( n5449 , n5448 , n5329 );
buf ( n295878 , n5449 );
nand ( n5451 , n5447 , n295878 );
buf ( n295880 , n5451 );
buf ( n295881 , n295880 );
nand ( n5454 , n5444 , n295881 );
buf ( n295883 , n5454 );
xor ( n5456 , n295166 , n295175 );
and ( n5457 , n5456 , n295187 );
and ( n5458 , n295166 , n295175 );
or ( n5459 , n5457 , n5458 );
buf ( n295888 , n5459 );
buf ( n295889 , n295888 );
not ( n5462 , n295889 );
buf ( n295891 , n5462 );
and ( n5464 , n295883 , n295891 );
not ( n295893 , n295883 );
and ( n5466 , n295893 , n295888 );
nor ( n5467 , n5464 , n5466 );
not ( n5468 , n5467 );
or ( n295897 , n295848 , n5468 );
not ( n295898 , n5467 );
not ( n5471 , n295847 );
nand ( n5472 , n295898 , n5471 );
nand ( n5473 , n295897 , n5472 );
not ( n5474 , n5473 );
or ( n5475 , n5271 , n5474 );
or ( n5476 , n5264 , n295695 );
nand ( n5477 , n5476 , n295693 );
nand ( n5478 , n4779 , n5477 );
nand ( n5479 , n5475 , n5478 );
buf ( n295908 , n5479 );
xor ( n5481 , n295153 , n295908 );
buf ( n295910 , n295555 );
not ( n295911 , n295910 );
buf ( n295912 , n291835 );
not ( n5485 , n295912 );
or ( n5486 , n295911 , n5485 );
buf ( n295915 , n777 );
buf ( n5488 , n824 );
xor ( n5489 , n295915 , n5488 );
buf ( n295918 , n5489 );
buf ( n295919 , n295918 );
buf ( n295920 , n1613 );
nand ( n295921 , n295919 , n295920 );
buf ( n295922 , n295921 );
buf ( n295923 , n295922 );
nand ( n5496 , n5486 , n295923 );
buf ( n295925 , n5496 );
not ( n295926 , n295925 );
not ( n5499 , n295926 );
buf ( n295928 , n799 );
xor ( n295929 , n803 , n804 );
buf ( n295930 , n295929 );
nand ( n295931 , n295928 , n295930 );
buf ( n295932 , n295931 );
buf ( n5505 , n295932 );
not ( n295934 , n5505 );
buf ( n295935 , n295934 );
not ( n5508 , n295935 );
buf ( n295937 , n4918 );
not ( n295938 , n295937 );
buf ( n295939 , n294329 );
not ( n5512 , n295939 );
or ( n295941 , n295938 , n5512 );
buf ( n295942 , n1508 );
xor ( n5515 , n828 , n773 );
buf ( n295944 , n5515 );
nand ( n295945 , n295942 , n295944 );
buf ( n295946 , n295945 );
buf ( n295947 , n295946 );
nand ( n295948 , n295941 , n295947 );
buf ( n295949 , n295948 );
not ( n5522 , n295949 );
not ( n295951 , n5522 );
or ( n295952 , n5508 , n295951 );
buf ( n295953 , n295949 );
buf ( n295954 , n295932 );
nand ( n295955 , n295953 , n295954 );
buf ( n295956 , n295955 );
nand ( n5529 , n295952 , n295956 );
not ( n295958 , n5529 );
or ( n295959 , n5499 , n295958 );
nand ( n295960 , n295935 , n5522 );
nand ( n295961 , n295960 , n295956 , n295925 );
nand ( n5534 , n295959 , n295961 );
not ( n295963 , n4890 );
not ( n295964 , n4798 );
or ( n5537 , n295963 , n295964 );
buf ( n295966 , n291988 );
not ( n5539 , n818 );
nand ( n5540 , n783 , n5539 );
not ( n295969 , n783 );
nand ( n295970 , n295969 , n818 );
nand ( n5543 , n5540 , n295970 );
buf ( n295972 , n5543 );
nand ( n295973 , n295966 , n295972 );
buf ( n295974 , n295973 );
nand ( n295975 , n5537 , n295974 );
buf ( n295976 , n5238 );
not ( n295977 , n295976 );
buf ( n295978 , n804 );
buf ( n295979 , n805 );
xnor ( n295980 , n295978 , n295979 );
buf ( n295981 , n295980 );
xor ( n5554 , n805 , n806 );
nor ( n295983 , n295981 , n5554 );
buf ( n295984 , n295983 );
not ( n5557 , n295984 );
or ( n295986 , n295977 , n5557 );
buf ( n295987 , n5554 );
buf ( n295988 , n797 );
buf ( n295989 , n804 );
xor ( n295990 , n295988 , n295989 );
buf ( n295991 , n295990 );
buf ( n295992 , n295991 );
nand ( n295993 , n295987 , n295992 );
buf ( n295994 , n295993 );
buf ( n295995 , n295994 );
nand ( n295996 , n295986 , n295995 );
buf ( n295997 , n295996 );
buf ( n295998 , n295997 );
not ( n5571 , n295998 );
buf ( n296000 , n5571 );
xor ( n296001 , n295975 , n296000 );
buf ( n296002 , n295650 );
not ( n5575 , n296002 );
buf ( n296004 , n291880 );
not ( n5577 , n296004 );
or ( n296006 , n5575 , n5577 );
buf ( n296007 , n293402 );
buf ( n296008 , n775 );
buf ( n296009 , n826 );
xor ( n296010 , n296008 , n296009 );
buf ( n296011 , n296010 );
buf ( n296012 , n296011 );
nand ( n296013 , n296007 , n296012 );
buf ( n296014 , n296013 );
buf ( n296015 , n296014 );
nand ( n296016 , n296006 , n296015 );
buf ( n296017 , n296016 );
xor ( n5590 , n296001 , n296017 );
xor ( n296019 , n5534 , n5590 );
not ( n5592 , n295579 );
not ( n296021 , n1933 );
or ( n296022 , n5592 , n296021 );
not ( n5595 , n771 );
not ( n5596 , n292367 );
or ( n5597 , n5595 , n5596 );
not ( n5598 , n771 );
nand ( n296027 , n5598 , n830 );
nand ( n296028 , n5597 , n296027 );
buf ( n296029 , n296028 );
buf ( n296030 , n831 );
nand ( n5603 , n296029 , n296030 );
buf ( n296032 , n5603 );
nand ( n296033 , n296022 , n296032 );
not ( n5606 , n296033 );
buf ( n296035 , n295264 );
not ( n296036 , n296035 );
buf ( n296037 , n3041 );
not ( n296038 , n296037 );
or ( n296039 , n296036 , n296038 );
buf ( n296040 , n295259 );
buf ( n296041 , n791 );
buf ( n5614 , n810 );
xor ( n5615 , n296041 , n5614 );
buf ( n5616 , n5615 );
buf ( n5617 , n5616 );
nand ( n5618 , n296040 , n5617 );
buf ( n5619 , n5618 );
buf ( n296048 , n5619 );
nand ( n5621 , n296039 , n296048 );
buf ( n296050 , n5621 );
not ( n296051 , n296050 );
not ( n5624 , n296051 );
or ( n296053 , n5606 , n5624 );
not ( n5626 , n296033 );
nand ( n5627 , n5626 , n296050 );
nand ( n5628 , n296053 , n5627 );
not ( n5629 , n295302 );
not ( n296058 , n3539 );
or ( n296059 , n5629 , n296058 );
xor ( n296060 , n789 , n812 );
nand ( n5633 , n294479 , n296060 );
nand ( n296062 , n296059 , n5633 );
xor ( n296063 , n5628 , n296062 );
buf ( n5636 , n296063 );
not ( n296065 , n5636 );
and ( n5638 , n296019 , n296065 );
not ( n5639 , n296019 );
and ( n296068 , n5639 , n5636 );
nor ( n296069 , n5638 , n296068 );
xor ( n5642 , n4821 , n295312 );
and ( n296071 , n5642 , n295402 );
and ( n296072 , n4821 , n295312 );
or ( n5645 , n296071 , n296072 );
xor ( n296074 , n296069 , n5645 );
not ( n296075 , n295804 );
not ( n5648 , n5410 );
not ( n5649 , n5648 );
or ( n296078 , n296075 , n5649 );
not ( n5651 , n295808 );
not ( n296080 , n5410 );
or ( n5653 , n5651 , n296080 );
buf ( n5654 , n5310 );
nand ( n296083 , n5653 , n5654 );
nand ( n296084 , n296078 , n296083 );
xor ( n5657 , n296074 , n296084 );
buf ( n296086 , n5657 );
not ( n296087 , n295847 );
not ( n5660 , n295888 );
or ( n296089 , n296087 , n5660 );
not ( n296090 , n5416 );
not ( n5663 , n295891 );
or ( n5664 , n296090 , n5663 );
nand ( n5665 , n5664 , n295883 );
nand ( n296094 , n296089 , n5665 );
buf ( n5667 , n296094 );
xor ( n5668 , n296086 , n5667 );
buf ( n296097 , n295637 );
not ( n296098 , n296097 );
and ( n5671 , n808 , n807 );
not ( n296100 , n808 );
and ( n296101 , n296100 , n295427 );
nor ( n5674 , n5671 , n296101 );
not ( n296103 , n5003 );
nor ( n5676 , n5674 , n296103 );
buf ( n296105 , n5676 );
not ( n296106 , n296105 );
or ( n296107 , n296098 , n296106 );
not ( n5680 , n5001 );
not ( n296109 , n5680 );
buf ( n296110 , n795 );
buf ( n296111 , n806 );
xor ( n296112 , n296110 , n296111 );
buf ( n296113 , n296112 );
nand ( n296114 , n296109 , n296113 );
buf ( n296115 , n296114 );
nand ( n296116 , n296107 , n296115 );
buf ( n296117 , n296116 );
not ( n5690 , n295615 );
not ( n296119 , n292668 );
or ( n5692 , n5690 , n296119 );
buf ( n296121 , n781 );
buf ( n296122 , n820 );
xor ( n296123 , n296121 , n296122 );
buf ( n296124 , n296123 );
nand ( n5697 , n291969 , n296124 );
nand ( n296126 , n5692 , n5697 );
buf ( n296127 , n296126 );
not ( n5700 , n296127 );
not ( n296129 , n295597 );
not ( n5702 , n4983 );
or ( n5703 , n296129 , n5702 );
xor ( n296132 , n808 , n793 );
buf ( n296133 , n296132 );
buf ( n296134 , n3114 );
nand ( n296135 , n296133 , n296134 );
buf ( n296136 , n296135 );
nand ( n5709 , n5703 , n296136 );
buf ( n296138 , n5709 );
not ( n5711 , n296138 );
buf ( n296140 , n5711 );
buf ( n296141 , n296140 );
not ( n296142 , n296141 );
or ( n5715 , n5700 , n296142 );
buf ( n296144 , n296140 );
buf ( n296145 , n296126 );
or ( n5718 , n296144 , n296145 );
nand ( n296147 , n5715 , n5718 );
buf ( n296148 , n296147 );
xor ( n5721 , n296117 , n296148 );
not ( n296150 , n295322 );
nand ( n296151 , n296150 , n295356 );
and ( n296152 , n295398 , n296151 );
not ( n296153 , n295322 );
nor ( n5726 , n296153 , n295356 );
nor ( n296155 , n296152 , n5726 );
not ( n296156 , n296155 );
xor ( n5729 , n5721 , n296156 );
not ( n296158 , n5404 );
not ( n296159 , n295821 );
or ( n5732 , n296158 , n296159 );
not ( n5733 , n5387 );
not ( n5734 , n5383 );
or ( n296163 , n5733 , n5734 );
or ( n296164 , n295821 , n5404 );
nand ( n5737 , n296163 , n296164 );
nand ( n5738 , n5732 , n5737 );
not ( n5739 , n5738 );
xnor ( n296168 , n5729 , n5739 );
buf ( n296169 , n296168 );
not ( n5742 , n295629 );
buf ( n296171 , n295671 );
not ( n5744 , n296171 );
buf ( n296173 , n5744 );
not ( n296174 , n296173 );
or ( n5747 , n5742 , n296174 );
not ( n5748 , n295671 );
not ( n296177 , n5196 );
or ( n296178 , n5748 , n296177 );
nand ( n5751 , n296178 , n5138 );
nand ( n5752 , n5747 , n5751 );
buf ( n296181 , n5102 );
not ( n296182 , n296181 );
buf ( n296183 , n3977 );
not ( n5756 , n296183 );
or ( n5757 , n296182 , n5756 );
buf ( n296186 , n1712 );
xor ( n5759 , n816 , n785 );
buf ( n296188 , n5759 );
nand ( n296189 , n296186 , n296188 );
buf ( n296190 , n296189 );
buf ( n296191 , n296190 );
nand ( n296192 , n5757 , n296191 );
buf ( n296193 , n296192 );
buf ( n296194 , n296193 );
buf ( n296195 , n295542 );
not ( n5768 , n296195 );
buf ( n296197 , n2078 );
not ( n296198 , n296197 );
or ( n296199 , n5768 , n296198 );
xor ( n5772 , n787 , n814 );
and ( n296201 , n816 , n815 );
not ( n296202 , n816 );
and ( n5775 , n296202 , n2086 );
nor ( n296204 , n296201 , n5775 );
nand ( n296205 , n5772 , n296204 );
buf ( n296206 , n296205 );
nand ( n296207 , n296199 , n296206 );
buf ( n296208 , n296207 );
buf ( n296209 , n296208 );
xor ( n296210 , n296194 , n296209 );
buf ( n296211 , n295284 );
not ( n296212 , n296211 );
buf ( n296213 , n292631 );
not ( n5786 , n296213 );
or ( n296215 , n296212 , n5786 );
buf ( n296216 , n1600 );
buf ( n296217 , n779 );
buf ( n296218 , n822 );
xor ( n5791 , n296217 , n296218 );
buf ( n296220 , n5791 );
buf ( n296221 , n296220 );
nand ( n296222 , n296216 , n296221 );
buf ( n296223 , n296222 );
buf ( n296224 , n296223 );
nand ( n296225 , n296215 , n296224 );
buf ( n296226 , n296225 );
buf ( n296227 , n296226 );
xor ( n296228 , n296210 , n296227 );
buf ( n296229 , n296228 );
buf ( n296230 , n296229 );
not ( n5803 , n296230 );
buf ( n296232 , n5803 );
not ( n5805 , n296232 );
buf ( n296234 , n295586 );
not ( n296235 , n296234 );
buf ( n296236 , n296235 );
buf ( n296237 , n296236 );
not ( n296238 , n296237 );
buf ( n296239 , n4990 );
not ( n5812 , n296239 );
buf ( n296241 , n3408 );
not ( n296242 , n296241 );
or ( n5815 , n5812 , n296242 );
buf ( n296244 , n295600 );
nand ( n296245 , n5815 , n296244 );
buf ( n296246 , n296245 );
buf ( n5819 , n296246 );
not ( n296248 , n5819 );
buf ( n296249 , n296248 );
buf ( n296250 , n296249 );
not ( n296251 , n296250 );
or ( n5824 , n296238 , n296251 );
buf ( n296253 , n295621 );
nand ( n296254 , n5824 , n296253 );
buf ( n296255 , n296254 );
buf ( n296256 , n296236 );
not ( n5829 , n296256 );
buf ( n296258 , n296246 );
nand ( n296259 , n5829 , n296258 );
buf ( n296260 , n296259 );
nand ( n5833 , n296255 , n296260 );
not ( n5834 , n5833 );
buf ( n296263 , n295641 );
not ( n5836 , n296263 );
buf ( n296265 , n295652 );
not ( n5838 , n296265 );
or ( n5839 , n5836 , n5838 );
or ( n5840 , n295652 , n295641 );
nand ( n5841 , n5840 , n5240 );
buf ( n296270 , n5841 );
nand ( n5843 , n5839 , n296270 );
buf ( n296272 , n5843 );
and ( n5845 , n5834 , n296272 );
not ( n296274 , n5834 );
not ( n5847 , n296272 );
and ( n5848 , n296274 , n5847 );
nor ( n5849 , n5845 , n5848 );
not ( n296278 , n5849 );
not ( n296279 , n296278 );
or ( n5852 , n5805 , n296279 );
nand ( n5853 , n5849 , n296229 );
nand ( n5854 , n5852 , n5853 );
and ( n296283 , n5752 , n5854 );
not ( n296284 , n5752 );
not ( n5857 , n5854 );
and ( n5858 , n296284 , n5857 );
nor ( n5859 , n296283 , n5858 );
and ( n296288 , n295338 , n295352 );
not ( n296289 , n5136 );
not ( n5862 , n5104 );
or ( n5863 , n296289 , n5862 );
or ( n5864 , n5136 , n5104 );
nand ( n296293 , n5864 , n295548 );
nand ( n296294 , n5863 , n296293 );
xor ( n5867 , n296288 , n296294 );
buf ( n296296 , n4860 );
not ( n5869 , n296296 );
buf ( n296298 , n295308 );
not ( n5871 , n296298 );
or ( n5872 , n5869 , n5871 );
buf ( n296301 , n295308 );
buf ( n296302 , n4860 );
or ( n296303 , n296301 , n296302 );
buf ( n296304 , n4842 );
nand ( n296305 , n296303 , n296304 );
buf ( n296306 , n296305 );
buf ( n296307 , n296306 );
nand ( n5880 , n5872 , n296307 );
buf ( n5881 , n5880 );
xnor ( n296310 , n5867 , n5881 );
buf ( n296311 , n296310 );
buf ( n296312 , n296311 );
buf ( n296313 , n296312 );
buf ( n296314 , n296313 );
not ( n296315 , n296314 );
buf ( n296316 , n296315 );
and ( n5889 , n5859 , n296316 );
not ( n296318 , n5859 );
and ( n296319 , n296318 , n296313 );
nor ( n5892 , n5889 , n296319 );
buf ( n296321 , n5892 );
xor ( n5894 , n296169 , n296321 );
buf ( n296323 , n4975 );
buf ( n296324 , n5096 );
or ( n5897 , n296323 , n296324 );
buf ( n296326 , n5259 );
nand ( n5899 , n5897 , n296326 );
buf ( n296328 , n5899 );
buf ( n296329 , n296328 );
buf ( n5902 , n5096 );
buf ( n296331 , n4975 );
nand ( n5904 , n5902 , n296331 );
buf ( n296333 , n5904 );
buf ( n296334 , n296333 );
nand ( n5907 , n296329 , n296334 );
buf ( n296336 , n5907 );
buf ( n296337 , n296336 );
xor ( n296338 , n5894 , n296337 );
buf ( n296339 , n296338 );
buf ( n296340 , n296339 );
xor ( n296341 , n5668 , n296340 );
buf ( n296342 , n296341 );
buf ( n296343 , n296342 );
and ( n5916 , n5481 , n296343 );
and ( n296345 , n295153 , n295908 );
or ( n296346 , n5916 , n296345 );
buf ( n296347 , n296346 );
buf ( n296348 , n296347 );
not ( n5921 , n296348 );
or ( n296350 , n295152 , n5921 );
buf ( n296351 , n831 );
not ( n296352 , n296351 );
buf ( n296353 , n867 );
buf ( n296354 , n5479 );
xor ( n296355 , n296353 , n296354 );
buf ( n296356 , n296342 );
and ( n296357 , n296355 , n296356 );
and ( n5930 , n296353 , n296354 );
or ( n296359 , n296357 , n5930 );
buf ( n296360 , n296359 );
buf ( n296361 , n296360 );
nand ( n296362 , n296352 , n296361 );
buf ( n296363 , n296362 );
buf ( n296364 , n296363 );
nand ( n296365 , n296350 , n296364 );
buf ( n296366 , n296365 );
buf ( n5939 , n296366 );
buf ( n296368 , n5939 );
not ( n296369 , n831 );
buf ( n296370 , n840 );
xor ( n296371 , n293298 , n293304 );
and ( n5944 , n296371 , n293573 );
and ( n296373 , n293298 , n293304 );
or ( n5946 , n5944 , n296373 );
buf ( n296375 , n5946 );
buf ( n296376 , n296375 );
xor ( n5949 , n296370 , n296376 );
xor ( n296378 , n293282 , n293288 );
and ( n296379 , n296378 , n293295 );
and ( n5952 , n293282 , n293288 );
or ( n296381 , n296379 , n5952 );
buf ( n296382 , n296381 );
buf ( n296383 , n296382 );
xor ( n296384 , n3019 , n293563 );
and ( n5957 , n296384 , n293570 );
and ( n296386 , n3019 , n293563 );
or ( n5959 , n5957 , n296386 );
buf ( n296388 , n5959 );
buf ( n296389 , n296388 );
xor ( n5962 , n296383 , n296389 );
xor ( n296391 , n294283 , n294301 );
xor ( n296392 , n296391 , n294306 );
buf ( n296393 , n296392 );
buf ( n296394 , n296393 );
xor ( n296395 , n5962 , n296394 );
buf ( n296396 , n296395 );
buf ( n296397 , n296396 );
and ( n5970 , n5949 , n296397 );
and ( n5971 , n296370 , n296376 );
or ( n296400 , n5970 , n5971 );
buf ( n296401 , n296400 );
not ( n296402 , n296401 );
or ( n5975 , n296369 , n296402 );
xor ( n296404 , n872 , n296375 );
and ( n296405 , n296404 , n296396 );
and ( n5978 , n872 , n296375 );
or ( n296407 , n296405 , n5978 );
not ( n5980 , n831 );
nand ( n296409 , n296407 , n5980 );
nand ( n5982 , n5975 , n296409 );
buf ( n296411 , n5982 );
not ( n296412 , n831 );
not ( n5985 , n296412 );
buf ( n296414 , n768 );
buf ( n296415 , n816 );
xor ( n5988 , n296414 , n296415 );
buf ( n5989 , n5988 );
buf ( n296418 , n5989 );
not ( n296419 , n296418 );
buf ( n296420 , n2118 );
not ( n5993 , n296420 );
or ( n296422 , n296419 , n5993 );
buf ( n296423 , n1712 );
buf ( n296424 , n296423 );
buf ( n296425 , n816 );
nand ( n5998 , n296424 , n296425 );
buf ( n296427 , n5998 );
buf ( n296428 , n296427 );
nand ( n6001 , n296422 , n296428 );
buf ( n296430 , n6001 );
buf ( n6003 , n296430 );
buf ( n296432 , n779 );
buf ( n296433 , n804 );
xor ( n296434 , n296432 , n296433 );
buf ( n296435 , n296434 );
buf ( n296436 , n296435 );
not ( n296437 , n296436 );
and ( n6010 , n295658 , n295657 );
buf ( n296439 , n6010 );
buf ( n296440 , n296439 );
buf ( n296441 , n296440 );
buf ( n296442 , n296441 );
not ( n296443 , n296442 );
or ( n296444 , n296437 , n296443 );
buf ( n6017 , n295361 );
buf ( n296446 , n6017 );
buf ( n6019 , n296446 );
buf ( n6020 , n778 );
buf ( n6021 , n804 );
xor ( n6022 , n6020 , n6021 );
buf ( n6023 , n6022 );
buf ( n296452 , n6023 );
nand ( n6025 , n6019 , n296452 );
buf ( n296454 , n6025 );
buf ( n296455 , n296454 );
nand ( n6028 , n296444 , n296455 );
buf ( n296457 , n6028 );
buf ( n6030 , n296457 );
xor ( n6031 , n6003 , n6030 );
buf ( n296460 , n800 );
buf ( n296461 , n784 );
xor ( n6034 , n296460 , n296461 );
buf ( n296463 , n6034 );
buf ( n296464 , n296463 );
not ( n6037 , n296464 );
buf ( n296466 , n801 );
buf ( n296467 , n802 );
xor ( n6040 , n296466 , n296467 );
buf ( n296469 , n6040 );
not ( n296470 , n296469 );
and ( n6043 , n800 , n801 );
not ( n296472 , n800 );
not ( n296473 , n801 );
and ( n6046 , n296472 , n296473 );
nor ( n296475 , n6043 , n6046 );
nand ( n6048 , n296470 , n296475 );
not ( n6049 , n6048 );
buf ( n296478 , n6049 );
buf ( n6051 , n296478 );
buf ( n296480 , n6051 );
buf ( n296481 , n296480 );
not ( n296482 , n296481 );
or ( n6055 , n6037 , n296482 );
xor ( n6056 , n801 , n802 );
buf ( n6057 , n6056 );
buf ( n296486 , n6057 );
xor ( n6059 , n783 , n800 );
buf ( n296488 , n6059 );
nand ( n6061 , n296486 , n296488 );
buf ( n296490 , n6061 );
buf ( n296491 , n296490 );
nand ( n6064 , n6055 , n296491 );
buf ( n296493 , n6064 );
not ( n296494 , n296493 );
buf ( n296495 , n782 );
buf ( n296496 , n802 );
xor ( n6069 , n296495 , n296496 );
buf ( n296498 , n6069 );
buf ( n296499 , n296498 );
not ( n296500 , n296499 );
nor ( n296501 , n803 , n804 );
not ( n296502 , n296501 );
not ( n6075 , n802 );
or ( n6076 , n296502 , n6075 );
not ( n296505 , n802 );
nand ( n6078 , n296505 , n804 , n803 );
nand ( n6079 , n6076 , n6078 );
buf ( n296508 , n6079 );
buf ( n296509 , n296508 );
not ( n6082 , n296509 );
or ( n6083 , n296500 , n6082 );
buf ( n296512 , n295929 );
not ( n6085 , n296512 );
buf ( n296514 , n6085 );
buf ( n296515 , n296514 );
not ( n296516 , n296515 );
buf ( n296517 , n296516 );
buf ( n296518 , n296517 );
buf ( n296519 , n781 );
buf ( n296520 , n802 );
xor ( n296521 , n296519 , n296520 );
buf ( n296522 , n296521 );
buf ( n6095 , n296522 );
nand ( n6096 , n296518 , n6095 );
buf ( n6097 , n6096 );
buf ( n6098 , n6097 );
nand ( n6099 , n6083 , n6098 );
buf ( n6100 , n6099 );
not ( n6101 , n6100 );
or ( n6102 , n296494 , n6101 );
buf ( n296531 , n296493 );
buf ( n296532 , n6100 );
nor ( n296533 , n296531 , n296532 );
buf ( n296534 , n296533 );
buf ( n296535 , n774 );
buf ( n296536 , n810 );
xor ( n296537 , n296535 , n296536 );
buf ( n296538 , n296537 );
buf ( n296539 , n296538 );
not ( n296540 , n296539 );
buf ( n296541 , n293058 );
not ( n296542 , n296541 );
or ( n6115 , n296540 , n296542 );
buf ( n6116 , n295259 );
buf ( n296545 , n773 );
buf ( n296546 , n810 );
xor ( n296547 , n296545 , n296546 );
buf ( n296548 , n296547 );
buf ( n296549 , n296548 );
nand ( n6122 , n6116 , n296549 );
buf ( n296551 , n6122 );
buf ( n296552 , n296551 );
nand ( n6125 , n6115 , n296552 );
buf ( n296554 , n6125 );
buf ( n6127 , n296554 );
not ( n296556 , n6127 );
buf ( n296557 , n296556 );
or ( n296558 , n296534 , n296557 );
nand ( n296559 , n6102 , n296558 );
buf ( n296560 , n296559 );
and ( n296561 , n6031 , n296560 );
and ( n6134 , n6003 , n6030 );
or ( n6135 , n296561 , n6134 );
buf ( n296564 , n6135 );
buf ( n296565 , n296564 );
and ( n6138 , n785 , n800 );
not ( n6139 , n6138 );
buf ( n296568 , n770 );
buf ( n296569 , n814 );
xor ( n6142 , n296568 , n296569 );
buf ( n296571 , n6142 );
not ( n6144 , n296571 );
not ( n6145 , n2893 );
or ( n6146 , n6144 , n6145 );
buf ( n296575 , n2089 );
buf ( n296576 , n814 );
buf ( n296577 , n769 );
xor ( n6150 , n296576 , n296577 );
buf ( n296579 , n6150 );
buf ( n296580 , n296579 );
nand ( n6153 , n296575 , n296580 );
buf ( n296582 , n6153 );
nand ( n6155 , n6146 , n296582 );
not ( n6156 , n6155 );
or ( n6157 , n6139 , n6156 );
nand ( n6158 , n2893 , n296571 );
not ( n296587 , n296582 );
nor ( n6160 , n296587 , n6138 );
nand ( n296589 , n6158 , n6160 );
xor ( n6162 , n808 , n776 );
not ( n6163 , n6162 );
buf ( n296592 , n293655 );
buf ( n6165 , n296592 );
buf ( n296594 , n6165 );
not ( n6167 , n296594 );
or ( n296596 , n6163 , n6167 );
buf ( n296597 , n294557 );
xor ( n6170 , n808 , n775 );
buf ( n296599 , n6170 );
nand ( n6172 , n296597 , n296599 );
buf ( n296601 , n6172 );
nand ( n296602 , n296596 , n296601 );
nand ( n6175 , n296589 , n296602 );
nand ( n6176 , n6157 , n6175 );
buf ( n296605 , n6176 );
and ( n296606 , n296460 , n296461 );
buf ( n296607 , n296606 );
buf ( n296608 , n296607 );
buf ( n296609 , n777 );
buf ( n296610 , n806 );
xor ( n296611 , n296609 , n296610 );
buf ( n296612 , n296611 );
buf ( n296613 , n296612 );
not ( n6186 , n296613 );
buf ( n296615 , n295433 );
buf ( n296616 , n296615 );
buf ( n296617 , n296616 );
buf ( n296618 , n296617 );
not ( n6191 , n296618 );
or ( n6192 , n6186 , n6191 );
buf ( n296621 , n295437 );
buf ( n296622 , n776 );
buf ( n296623 , n806 );
xor ( n296624 , n296622 , n296623 );
buf ( n296625 , n296624 );
buf ( n296626 , n296625 );
nand ( n6199 , n296621 , n296626 );
buf ( n296628 , n6199 );
buf ( n296629 , n296628 );
nand ( n6202 , n6192 , n296629 );
buf ( n296631 , n6202 );
buf ( n296632 , n296631 );
xor ( n6205 , n296608 , n296632 );
xor ( n6206 , n812 , n771 );
buf ( n296635 , n6206 );
not ( n296636 , n296635 );
buf ( n6209 , n2376 );
buf ( n296638 , n6209 );
not ( n296639 , n296638 );
or ( n6212 , n296636 , n296639 );
buf ( n296641 , n2383 );
xor ( n296642 , n812 , n770 );
buf ( n296643 , n296642 );
nand ( n296644 , n296641 , n296643 );
buf ( n296645 , n296644 );
buf ( n296646 , n296645 );
nand ( n296647 , n6212 , n296646 );
buf ( n296648 , n296647 );
buf ( n296649 , n296648 );
xor ( n296650 , n6205 , n296649 );
buf ( n296651 , n296650 );
buf ( n296652 , n296651 );
xor ( n296653 , n296605 , n296652 );
buf ( n6226 , n780 );
buf ( n296655 , n804 );
xor ( n296656 , n6226 , n296655 );
buf ( n296657 , n296656 );
buf ( n296658 , n296657 );
not ( n6231 , n296658 );
buf ( n296660 , n296441 );
not ( n6233 , n296660 );
or ( n6234 , n6231 , n6233 );
buf ( n296663 , n295361 );
buf ( n296664 , n296663 );
buf ( n296665 , n296664 );
buf ( n296666 , n296435 );
nand ( n6239 , n296665 , n296666 );
buf ( n296668 , n6239 );
buf ( n296669 , n296668 );
nand ( n296670 , n6234 , n296669 );
buf ( n296671 , n296670 );
buf ( n296672 , n296671 );
buf ( n296673 , n778 );
buf ( n296674 , n806 );
xor ( n296675 , n296673 , n296674 );
buf ( n296676 , n296675 );
buf ( n296677 , n296676 );
not ( n296678 , n296677 );
buf ( n296679 , n296617 );
not ( n6252 , n296679 );
or ( n296681 , n296678 , n6252 );
buf ( n296682 , n295437 );
buf ( n296683 , n296612 );
nand ( n296684 , n296682 , n296683 );
buf ( n296685 , n296684 );
buf ( n296686 , n296685 );
nand ( n296687 , n296681 , n296686 );
buf ( n296688 , n296687 );
buf ( n296689 , n296688 );
xor ( n296690 , n296672 , n296689 );
buf ( n296691 , n772 );
buf ( n296692 , n812 );
xor ( n296693 , n296691 , n296692 );
buf ( n296694 , n296693 );
buf ( n296695 , n296694 );
not ( n296696 , n296695 );
buf ( n296697 , n6209 );
not ( n6270 , n296697 );
or ( n296699 , n296696 , n6270 );
not ( n296700 , n2383 );
not ( n6273 , n296700 );
nand ( n296702 , n6273 , n6206 );
buf ( n296703 , n296702 );
nand ( n6276 , n296699 , n296703 );
buf ( n296705 , n6276 );
buf ( n296706 , n296705 );
and ( n296707 , n296690 , n296706 );
and ( n296708 , n296672 , n296689 );
or ( n6281 , n296707 , n296708 );
buf ( n296710 , n6281 );
buf ( n296711 , n296710 );
and ( n296712 , n296653 , n296711 );
and ( n296713 , n296605 , n296652 );
or ( n6286 , n296712 , n296713 );
buf ( n296715 , n6286 );
buf ( n296716 , n296715 );
xor ( n296717 , n296565 , n296716 );
xor ( n296718 , n296608 , n296632 );
and ( n6291 , n296718 , n296649 );
and ( n6292 , n296608 , n296632 );
or ( n296721 , n6291 , n6292 );
buf ( n296722 , n296721 );
buf ( n296723 , n296722 );
buf ( n296724 , n6170 );
not ( n6297 , n296724 );
buf ( n296726 , n296594 );
not ( n296727 , n296726 );
or ( n6300 , n6297 , n296727 );
xor ( n6301 , n809 , n810 );
buf ( n296730 , n6301 );
buf ( n296731 , n774 );
buf ( n6304 , n808 );
xor ( n6305 , n296731 , n6304 );
buf ( n296734 , n6305 );
buf ( n296735 , n296734 );
nand ( n296736 , n296730 , n296735 );
buf ( n296737 , n296736 );
buf ( n296738 , n296737 );
nand ( n6311 , n6300 , n296738 );
buf ( n296740 , n6311 );
buf ( n296741 , n296740 );
buf ( n296742 , n296522 );
not ( n6315 , n296742 );
buf ( n296744 , n296508 );
not ( n6317 , n296744 );
or ( n296746 , n6315 , n6317 );
buf ( n296747 , n295929 );
buf ( n6320 , n296747 );
buf ( n296749 , n6320 );
buf ( n296750 , n296749 );
xor ( n296751 , n802 , n780 );
buf ( n6324 , n296751 );
nand ( n6325 , n296750 , n6324 );
buf ( n6326 , n6325 );
buf ( n296755 , n6326 );
nand ( n6328 , n296746 , n296755 );
buf ( n6329 , n6328 );
buf ( n296758 , n6329 );
xor ( n6331 , n296741 , n296758 );
buf ( n296760 , n6059 );
not ( n296761 , n296760 );
buf ( n296762 , n296480 );
not ( n6335 , n296762 );
or ( n6336 , n296761 , n6335 );
buf ( n296765 , n6057 );
buf ( n296766 , n800 );
buf ( n296767 , n782 );
xor ( n6340 , n296766 , n296767 );
buf ( n296769 , n6340 );
buf ( n296770 , n296769 );
nand ( n296771 , n296765 , n296770 );
buf ( n296772 , n296771 );
buf ( n296773 , n296772 );
nand ( n296774 , n6336 , n296773 );
buf ( n296775 , n296774 );
buf ( n296776 , n296775 );
and ( n296777 , n6331 , n296776 );
and ( n296778 , n296741 , n296758 );
or ( n6351 , n296777 , n296778 );
buf ( n296780 , n6351 );
buf ( n296781 , n296780 );
xor ( n6354 , n296723 , n296781 );
buf ( n296783 , n296579 );
not ( n6356 , n296783 );
buf ( n296785 , n2893 );
not ( n296786 , n296785 );
or ( n296787 , n6356 , n296786 );
buf ( n296788 , n292518 );
xor ( n6361 , n814 , n768 );
buf ( n296790 , n6361 );
nand ( n296791 , n296788 , n296790 );
buf ( n296792 , n296791 );
buf ( n296793 , n296792 );
nand ( n296794 , n296787 , n296793 );
buf ( n296795 , n296794 );
buf ( n296796 , n296795 );
buf ( n296797 , n296423 );
not ( n6370 , n296797 );
buf ( n296799 , n6370 );
buf ( n296800 , n296799 );
not ( n6373 , n296800 );
buf ( n296802 , n292543 );
not ( n6375 , n296802 );
or ( n6376 , n6373 , n6375 );
buf ( n296805 , n816 );
nand ( n6378 , n6376 , n296805 );
buf ( n296807 , n6378 );
buf ( n296808 , n296807 );
xor ( n6381 , n296796 , n296808 );
buf ( n296810 , n296548 );
not ( n296811 , n296810 );
buf ( n296812 , n293058 );
not ( n6385 , n296812 );
or ( n296814 , n296811 , n6385 );
buf ( n296815 , n295259 );
buf ( n296816 , n772 );
buf ( n296817 , n810 );
xor ( n296818 , n296816 , n296817 );
buf ( n296819 , n296818 );
buf ( n296820 , n296819 );
nand ( n6393 , n296815 , n296820 );
buf ( n296822 , n6393 );
buf ( n296823 , n296822 );
nand ( n296824 , n296814 , n296823 );
buf ( n296825 , n296824 );
buf ( n296826 , n296825 );
and ( n296827 , n6381 , n296826 );
and ( n6400 , n296796 , n296808 );
or ( n296829 , n296827 , n6400 );
buf ( n296830 , n296829 );
buf ( n296831 , n296830 );
xor ( n296832 , n6354 , n296831 );
buf ( n296833 , n296832 );
buf ( n296834 , n296833 );
xor ( n6407 , n296717 , n296834 );
buf ( n296836 , n6407 );
buf ( n296837 , n296836 );
xor ( n296838 , n296741 , n296758 );
xor ( n296839 , n296838 , n296776 );
buf ( n296840 , n296839 );
buf ( n296841 , n296840 );
xor ( n296842 , n296796 , n296808 );
xor ( n6415 , n296842 , n296826 );
buf ( n296844 , n6415 );
buf ( n296845 , n296844 );
xor ( n296846 , n296841 , n296845 );
xor ( n6419 , n6003 , n6030 );
xor ( n296848 , n6419 , n296560 );
buf ( n296849 , n296848 );
buf ( n296850 , n296849 );
xor ( n296851 , n296846 , n296850 );
buf ( n296852 , n296851 );
buf ( n296853 , n296852 );
buf ( n296854 , n779 );
buf ( n296855 , n806 );
xor ( n6428 , n296854 , n296855 );
buf ( n296857 , n6428 );
buf ( n296858 , n296857 );
not ( n6431 , n296858 );
buf ( n296860 , n295433 );
not ( n296861 , n296860 );
or ( n6434 , n6431 , n296861 );
buf ( n296863 , n295437 );
buf ( n296864 , n296676 );
nand ( n296865 , n296863 , n296864 );
buf ( n296866 , n296865 );
buf ( n296867 , n296866 );
nand ( n296868 , n6434 , n296867 );
buf ( n296869 , n296868 );
buf ( n296870 , n296869 );
buf ( n296871 , n770 );
buf ( n296872 , n816 );
xor ( n6445 , n296871 , n296872 );
buf ( n296874 , n6445 );
buf ( n296875 , n296874 );
not ( n296876 , n296875 );
buf ( n296877 , n2118 );
not ( n296878 , n296877 );
or ( n296879 , n296876 , n296878 );
buf ( n296880 , n296423 );
buf ( n296881 , n769 );
buf ( n6454 , n816 );
xor ( n6455 , n296881 , n6454 );
buf ( n296884 , n6455 );
buf ( n296885 , n296884 );
nand ( n296886 , n296880 , n296885 );
buf ( n296887 , n296886 );
buf ( n296888 , n296887 );
nand ( n296889 , n296879 , n296888 );
buf ( n296890 , n296889 );
buf ( n296891 , n296890 );
xor ( n296892 , n296870 , n296891 );
buf ( n296893 , n777 );
buf ( n296894 , n808 );
xor ( n6467 , n296893 , n296894 );
buf ( n6468 , n6467 );
buf ( n296897 , n6468 );
not ( n6470 , n296897 );
buf ( n296899 , n296594 );
not ( n296900 , n296899 );
or ( n296901 , n6470 , n296900 );
buf ( n296902 , n6301 );
buf ( n296903 , n6162 );
nand ( n6476 , n296902 , n296903 );
buf ( n296905 , n6476 );
buf ( n296906 , n296905 );
nand ( n6479 , n296901 , n296906 );
buf ( n296908 , n6479 );
buf ( n296909 , n296908 );
and ( n296910 , n296892 , n296909 );
and ( n296911 , n296870 , n296891 );
or ( n6484 , n296910 , n296911 );
buf ( n296913 , n6484 );
buf ( n296914 , n296913 );
xor ( n6487 , n296672 , n296689 );
xor ( n6488 , n6487 , n296706 );
buf ( n296917 , n6488 );
buf ( n296918 , n296917 );
xor ( n6491 , n296914 , n296918 );
buf ( n296920 , n786 );
buf ( n296921 , n800 );
xor ( n6494 , n296920 , n296921 );
buf ( n296923 , n6494 );
buf ( n296924 , n296923 );
not ( n6497 , n296924 );
buf ( n296926 , n296480 );
not ( n296927 , n296926 );
or ( n6500 , n6497 , n296927 );
buf ( n296929 , n6057 );
xor ( n6502 , n785 , n800 );
buf ( n296931 , n6502 );
nand ( n296932 , n296929 , n296931 );
buf ( n296933 , n296932 );
buf ( n296934 , n296933 );
nand ( n296935 , n6500 , n296934 );
buf ( n296936 , n296935 );
not ( n6509 , n296936 );
buf ( n296938 , n787 );
buf ( n296939 , n800 );
and ( n296940 , n296938 , n296939 );
buf ( n296941 , n296940 );
not ( n6514 , n296941 );
nand ( n296943 , n6509 , n6514 );
not ( n296944 , n296943 );
buf ( n296945 , n776 );
buf ( n296946 , n810 );
xor ( n6519 , n296945 , n296946 );
buf ( n296948 , n6519 );
buf ( n296949 , n296948 );
not ( n296950 , n296949 );
buf ( n296951 , n293058 );
not ( n296952 , n296951 );
or ( n296953 , n296950 , n296952 );
buf ( n296954 , n295259 );
xor ( n296955 , n810 , n775 );
buf ( n296956 , n296955 );
nand ( n6529 , n296954 , n296956 );
buf ( n296958 , n6529 );
buf ( n296959 , n296958 );
nand ( n296960 , n296953 , n296959 );
buf ( n296961 , n296960 );
not ( n296962 , n296961 );
or ( n6535 , n296944 , n296962 );
buf ( n296964 , n296936 );
nand ( n296965 , n296941 , n296964 );
nand ( n296966 , n6535 , n296965 );
buf ( n296967 , n774 );
buf ( n296968 , n812 );
xor ( n6541 , n296967 , n296968 );
buf ( n296970 , n6541 );
buf ( n296971 , n296970 );
not ( n296972 , n296971 );
buf ( n296973 , n2376 );
not ( n296974 , n296973 );
or ( n6547 , n296972 , n296974 );
buf ( n296976 , n2383 );
buf ( n6549 , n773 );
buf ( n6550 , n812 );
xor ( n6551 , n6549 , n6550 );
buf ( n6552 , n6551 );
buf ( n296981 , n6552 );
nand ( n6554 , n296976 , n296981 );
buf ( n296983 , n6554 );
buf ( n296984 , n296983 );
nand ( n6557 , n6547 , n296984 );
buf ( n296986 , n6557 );
buf ( n296987 , n296986 );
not ( n6560 , n296987 );
buf ( n296989 , n782 );
buf ( n296990 , n804 );
xor ( n296991 , n296989 , n296990 );
buf ( n296992 , n296991 );
buf ( n296993 , n296992 );
not ( n6566 , n296993 );
buf ( n296995 , n6010 );
not ( n6568 , n296995 );
or ( n296997 , n6566 , n6568 );
buf ( n296998 , n296663 );
buf ( n296999 , n781 );
buf ( n297000 , n804 );
xor ( n6573 , n296999 , n297000 );
buf ( n297002 , n6573 );
buf ( n297003 , n297002 );
nand ( n6576 , n296998 , n297003 );
buf ( n6577 , n6576 );
buf ( n297006 , n6577 );
nand ( n6579 , n296997 , n297006 );
buf ( n297008 , n6579 );
buf ( n297009 , n297008 );
not ( n297010 , n297009 );
or ( n6583 , n6560 , n297010 );
or ( n6584 , n296986 , n297008 );
buf ( n297013 , n784 );
buf ( n297014 , n802 );
xor ( n297015 , n297013 , n297014 );
buf ( n297016 , n297015 );
buf ( n297017 , n297016 );
not ( n6590 , n297017 );
buf ( n297019 , n296508 );
not ( n6592 , n297019 );
or ( n6593 , n6590 , n6592 );
buf ( n297022 , n296749 );
buf ( n297023 , n783 );
buf ( n297024 , n802 );
xor ( n6597 , n297023 , n297024 );
buf ( n297026 , n6597 );
buf ( n297027 , n297026 );
nand ( n6600 , n297022 , n297027 );
buf ( n297029 , n6600 );
buf ( n297030 , n297029 );
nand ( n297031 , n6593 , n297030 );
buf ( n297032 , n297031 );
nand ( n6605 , n6584 , n297032 );
buf ( n297034 , n6605 );
nand ( n297035 , n6583 , n297034 );
buf ( n297036 , n297035 );
or ( n297037 , n296966 , n297036 );
buf ( n297038 , n768 );
buf ( n297039 , n818 );
xor ( n297040 , n297038 , n297039 );
buf ( n297041 , n297040 );
buf ( n297042 , n297041 );
not ( n6615 , n297042 );
buf ( n297044 , n292393 );
not ( n297045 , n297044 );
or ( n6618 , n6615 , n297045 );
buf ( n297047 , n291788 );
buf ( n297048 , n818 );
nand ( n6621 , n297047 , n297048 );
buf ( n297050 , n6621 );
buf ( n297051 , n297050 );
nand ( n6624 , n6618 , n297051 );
buf ( n297053 , n6624 );
not ( n6626 , n297053 );
and ( n297055 , n294557 , n6468 );
and ( n297056 , n778 , n294635 );
not ( n6629 , n778 );
and ( n297058 , n6629 , n808 );
nor ( n297059 , n297056 , n297058 );
nor ( n297060 , n297059 , n295410 , n4981 );
nor ( n297061 , n297055 , n297060 );
nand ( n6634 , n6626 , n297061 );
not ( n297063 , n6634 );
buf ( n297064 , n772 );
buf ( n297065 , n814 );
xor ( n297066 , n297064 , n297065 );
buf ( n297067 , n297066 );
buf ( n297068 , n297067 );
not ( n297069 , n297068 );
buf ( n297070 , n2893 );
not ( n6643 , n297070 );
or ( n297072 , n297069 , n6643 );
buf ( n297073 , n2089 );
buf ( n297074 , n771 );
buf ( n297075 , n814 );
xor ( n6648 , n297074 , n297075 );
buf ( n297077 , n6648 );
buf ( n6650 , n297077 );
nand ( n6651 , n297073 , n6650 );
buf ( n6652 , n6651 );
buf ( n297081 , n6652 );
nand ( n6654 , n297072 , n297081 );
buf ( n297083 , n6654 );
not ( n6656 , n297083 );
or ( n6657 , n297063 , n6656 );
not ( n297086 , n297061 );
nand ( n297087 , n297086 , n297053 );
nand ( n6660 , n6657 , n297087 );
nand ( n297089 , n297037 , n6660 );
nand ( n297090 , n297036 , n296966 );
nand ( n6663 , n297089 , n297090 );
buf ( n297092 , n6663 );
and ( n6665 , n6491 , n297092 );
and ( n6666 , n296914 , n296918 );
or ( n297095 , n6665 , n6666 );
buf ( n297096 , n297095 );
buf ( n297097 , n297096 );
xor ( n297098 , n296853 , n297097 );
not ( n297099 , n295230 );
buf ( n297100 , n297099 );
not ( n6673 , n297100 );
buf ( n297102 , n1962 );
not ( n297103 , n297102 );
buf ( n297104 , n297103 );
buf ( n6677 , n297104 );
not ( n6678 , n6677 );
or ( n6679 , n6673 , n6678 );
buf ( n297108 , n818 );
nand ( n297109 , n6679 , n297108 );
buf ( n297110 , n297109 );
not ( n297111 , n2118 );
not ( n297112 , n296884 );
or ( n6685 , n297111 , n297112 );
buf ( n297114 , n296423 );
buf ( n297115 , n5989 );
nand ( n6688 , n297114 , n297115 );
buf ( n6689 , n6688 );
nand ( n6690 , n6685 , n6689 );
xor ( n6691 , n297110 , n6690 );
buf ( n297120 , n6552 );
not ( n6693 , n297120 );
buf ( n297122 , n2376 );
not ( n6695 , n297122 );
or ( n6696 , n6693 , n6695 );
buf ( n297125 , n2383 );
buf ( n297126 , n296694 );
nand ( n297127 , n297125 , n297126 );
buf ( n297128 , n297127 );
buf ( n297129 , n297128 );
nand ( n6702 , n6696 , n297129 );
buf ( n297131 , n6702 );
and ( n6704 , n6691 , n297131 );
and ( n6705 , n297110 , n6690 );
or ( n6706 , n6704 , n6705 );
buf ( n297135 , n6706 );
not ( n297136 , n297135 );
buf ( n297137 , n296430 );
not ( n6710 , n297137 );
and ( n297139 , n297136 , n6710 );
buf ( n297140 , n6706 );
buf ( n297141 , n296430 );
and ( n6714 , n297140 , n297141 );
nor ( n6715 , n297139 , n6714 );
buf ( n297144 , n6715 );
buf ( n297145 , n297144 );
buf ( n297146 , n297026 );
not ( n6719 , n297146 );
buf ( n297148 , n296508 );
not ( n297149 , n297148 );
or ( n6722 , n6719 , n297149 );
buf ( n297151 , n296749 );
buf ( n297152 , n296498 );
nand ( n6725 , n297151 , n297152 );
buf ( n297154 , n6725 );
buf ( n297155 , n297154 );
nand ( n297156 , n6722 , n297155 );
buf ( n297157 , n297156 );
buf ( n297158 , n297157 );
buf ( n297159 , n297002 );
not ( n297160 , n297159 );
buf ( n297161 , n296441 );
not ( n6734 , n297161 );
or ( n6735 , n297160 , n6734 );
buf ( n297164 , n296664 );
buf ( n297165 , n296657 );
nand ( n297166 , n297164 , n297165 );
buf ( n297167 , n297166 );
buf ( n297168 , n297167 );
nand ( n6741 , n6735 , n297168 );
buf ( n297170 , n6741 );
buf ( n297171 , n297170 );
xor ( n6744 , n297158 , n297171 );
buf ( n297173 , n296955 );
not ( n6746 , n297173 );
buf ( n297175 , n293058 );
buf ( n297176 , n297175 );
not ( n6749 , n297176 );
or ( n6750 , n6746 , n6749 );
buf ( n297179 , n295259 );
buf ( n297180 , n296538 );
nand ( n297181 , n297179 , n297180 );
buf ( n297182 , n297181 );
buf ( n297183 , n297182 );
nand ( n6756 , n6750 , n297183 );
buf ( n297185 , n6756 );
buf ( n297186 , n297185 );
and ( n6759 , n6744 , n297186 );
and ( n6760 , n297158 , n297171 );
or ( n6761 , n6759 , n6760 );
buf ( n297190 , n6761 );
buf ( n297191 , n297190 );
xor ( n6764 , n297145 , n297191 );
buf ( n297193 , n6764 );
not ( n6766 , n297193 );
buf ( n297195 , n786 );
buf ( n6768 , n800 );
and ( n6769 , n297195 , n6768 );
buf ( n6770 , n6769 );
buf ( n6771 , n6770 );
buf ( n297200 , n6502 );
not ( n6773 , n297200 );
buf ( n297202 , n296480 );
not ( n297203 , n297202 );
or ( n297204 , n6773 , n297203 );
buf ( n297205 , n6057 );
buf ( n297206 , n296463 );
nand ( n297207 , n297205 , n297206 );
buf ( n297208 , n297207 );
buf ( n297209 , n297208 );
nand ( n6782 , n297204 , n297209 );
buf ( n297211 , n6782 );
buf ( n6784 , n297211 );
xor ( n6785 , n6771 , n6784 );
buf ( n6786 , n297077 );
not ( n6787 , n6786 );
buf ( n297216 , n292509 );
not ( n6789 , n297216 );
or ( n297218 , n6787 , n6789 );
buf ( n297219 , n292518 );
buf ( n297220 , n296571 );
nand ( n297221 , n297219 , n297220 );
buf ( n297222 , n297221 );
buf ( n297223 , n297222 );
nand ( n6796 , n297218 , n297223 );
buf ( n6797 , n6796 );
buf ( n297226 , n6797 );
and ( n6799 , n6785 , n297226 );
and ( n6800 , n6771 , n6784 );
or ( n297229 , n6799 , n6800 );
buf ( n297230 , n297229 );
buf ( n297231 , n297230 );
not ( n6804 , n297231 );
buf ( n6805 , n6804 );
buf ( n297234 , n6805 );
not ( n6807 , n297234 );
not ( n6808 , n296463 );
not ( n297237 , n296480 );
or ( n297238 , n6808 , n297237 );
nand ( n6811 , n297238 , n296490 );
xor ( n6812 , n6811 , n296554 );
xnor ( n6813 , n6812 , n6100 );
buf ( n297242 , n6813 );
not ( n297243 , n297242 );
buf ( n297244 , n297243 );
buf ( n297245 , n297244 );
not ( n6818 , n297245 );
or ( n297247 , n6807 , n6818 );
buf ( n6820 , n6813 );
buf ( n297249 , n297230 );
nand ( n6822 , n6820 , n297249 );
buf ( n297251 , n6822 );
buf ( n297252 , n297251 );
nand ( n6825 , n297247 , n297252 );
buf ( n297254 , n6825 );
buf ( n297255 , n6138 );
buf ( n297256 , n296602 );
xor ( n6829 , n297255 , n297256 );
buf ( n297258 , n6155 );
xnor ( n297259 , n6829 , n297258 );
buf ( n297260 , n297259 );
and ( n6833 , n297254 , n297260 );
not ( n6834 , n297254 );
buf ( n297263 , n297260 );
not ( n297264 , n297263 );
buf ( n297265 , n297264 );
and ( n6838 , n6834 , n297265 );
nor ( n6839 , n6833 , n6838 );
not ( n6840 , n6839 );
or ( n297269 , n6766 , n6840 );
xor ( n297270 , n6771 , n6784 );
xor ( n6843 , n297270 , n297226 );
buf ( n297272 , n6843 );
buf ( n297273 , n297272 );
xor ( n297274 , n297110 , n6690 );
xor ( n297275 , n297274 , n297131 );
buf ( n297276 , n297275 );
xor ( n6849 , n297273 , n297276 );
xor ( n6850 , n297158 , n297171 );
xor ( n297279 , n6850 , n297186 );
buf ( n297280 , n297279 );
buf ( n297281 , n297280 );
and ( n297282 , n6849 , n297281 );
and ( n297283 , n297273 , n297276 );
or ( n6856 , n297282 , n297283 );
buf ( n297285 , n6856 );
nand ( n297286 , n297269 , n297285 );
buf ( n297287 , n297286 );
buf ( n297288 , n297193 );
not ( n297289 , n297288 );
not ( n6862 , n6839 );
buf ( n297291 , n6862 );
nand ( n297292 , n297289 , n297291 );
buf ( n297293 , n297292 );
buf ( n297294 , n297293 );
nand ( n297295 , n297287 , n297294 );
buf ( n297296 , n297295 );
buf ( n297297 , n297296 );
and ( n297298 , n297098 , n297297 );
and ( n6871 , n296853 , n297097 );
or ( n297300 , n297298 , n6871 );
buf ( n297301 , n297300 );
buf ( n297302 , n297301 );
xor ( n6875 , n296837 , n297302 );
xor ( n6876 , n296841 , n296845 );
and ( n297305 , n6876 , n296850 );
and ( n6878 , n296841 , n296845 );
or ( n297307 , n297305 , n6878 );
buf ( n297308 , n297307 );
buf ( n297309 , n297308 );
and ( n6882 , n783 , n800 );
not ( n297311 , n6882 );
not ( n6884 , n297311 );
buf ( n297313 , n296734 );
not ( n6886 , n297313 );
buf ( n297315 , n296594 );
not ( n6888 , n297315 );
or ( n6889 , n6886 , n6888 );
buf ( n297318 , n6301 );
buf ( n6891 , n808 );
buf ( n297320 , n773 );
xor ( n6893 , n6891 , n297320 );
buf ( n297322 , n6893 );
buf ( n297323 , n297322 );
nand ( n297324 , n297318 , n297323 );
buf ( n297325 , n297324 );
buf ( n297326 , n297325 );
nand ( n6899 , n6889 , n297326 );
buf ( n297328 , n6899 );
not ( n6901 , n297328 );
buf ( n297330 , n296769 );
not ( n297331 , n297330 );
buf ( n297332 , n296480 );
not ( n297333 , n297332 );
or ( n6906 , n297331 , n297333 );
buf ( n297335 , n6057 );
buf ( n6908 , n800 );
buf ( n6909 , n781 );
xor ( n6910 , n6908 , n6909 );
buf ( n297339 , n6910 );
buf ( n297340 , n297339 );
nand ( n297341 , n297335 , n297340 );
buf ( n297342 , n297341 );
buf ( n297343 , n297342 );
nand ( n297344 , n6906 , n297343 );
buf ( n297345 , n297344 );
not ( n6918 , n297345 );
nand ( n297347 , n6884 , n6901 , n6918 );
nand ( n6920 , n6918 , n297311 );
not ( n6921 , n6920 );
nand ( n297350 , n6921 , n297328 );
not ( n297351 , n297345 );
nor ( n6924 , n297351 , n6882 );
nand ( n297353 , n6901 , n6924 );
not ( n297354 , n6918 );
nand ( n6927 , n297328 , n297354 , n6882 );
nand ( n297356 , n297347 , n297350 , n297353 , n6927 );
buf ( n297357 , n296751 );
not ( n6930 , n297357 );
buf ( n297359 , n296508 );
not ( n6932 , n297359 );
or ( n6933 , n6930 , n6932 );
buf ( n297362 , n296749 );
buf ( n297363 , n802 );
buf ( n297364 , n779 );
xor ( n6937 , n297363 , n297364 );
buf ( n297366 , n6937 );
buf ( n297367 , n297366 );
nand ( n297368 , n297362 , n297367 );
buf ( n297369 , n297368 );
buf ( n297370 , n297369 );
nand ( n297371 , n6933 , n297370 );
buf ( n297372 , n297371 );
buf ( n297373 , n297372 );
buf ( n297374 , n6023 );
not ( n6947 , n297374 );
buf ( n297376 , n296441 );
not ( n6949 , n297376 );
or ( n297378 , n6947 , n6949 );
buf ( n297379 , n804 );
not ( n297380 , n297379 );
buf ( n297381 , n777 );
nor ( n6954 , n297380 , n297381 );
buf ( n6955 , n6954 );
buf ( n297384 , n6955 );
buf ( n297385 , n777 );
not ( n297386 , n297385 );
buf ( n6959 , n804 );
nor ( n6960 , n297386 , n6959 );
buf ( n6961 , n6960 );
buf ( n297390 , n6961 );
nor ( n6963 , n297384 , n297390 );
buf ( n297392 , n6963 );
buf ( n297393 , n297392 );
not ( n6966 , n297393 );
buf ( n297395 , n6017 );
buf ( n6968 , n297395 );
nand ( n6969 , n6966 , n6968 );
buf ( n6970 , n6969 );
buf ( n6971 , n6970 );
nand ( n6972 , n297378 , n6971 );
buf ( n6973 , n6972 );
buf ( n297402 , n6973 );
xor ( n6975 , n297373 , n297402 );
buf ( n297404 , n6361 );
not ( n297405 , n297404 );
buf ( n297406 , n2893 );
not ( n6979 , n297406 );
or ( n297408 , n297405 , n6979 );
buf ( n297409 , n292518 );
buf ( n297410 , n814 );
nand ( n297411 , n297409 , n297410 );
buf ( n297412 , n297411 );
buf ( n297413 , n297412 );
nand ( n297414 , n297408 , n297413 );
buf ( n297415 , n297414 );
buf ( n297416 , n297415 );
not ( n297417 , n297416 );
buf ( n297418 , n297417 );
buf ( n297419 , n297418 );
xor ( n297420 , n6975 , n297419 );
buf ( n297421 , n297420 );
not ( n6994 , n297421 );
xor ( n297423 , n297356 , n6994 );
buf ( n297424 , n296642 );
not ( n6997 , n297424 );
buf ( n297426 , n2376 );
not ( n297427 , n297426 );
or ( n7000 , n6997 , n297427 );
buf ( n297429 , n2383 );
xor ( n7002 , n812 , n769 );
buf ( n297431 , n7002 );
nand ( n297432 , n297429 , n297431 );
buf ( n297433 , n297432 );
buf ( n297434 , n297433 );
nand ( n297435 , n7000 , n297434 );
buf ( n297436 , n297435 );
buf ( n297437 , n297436 );
buf ( n297438 , n775 );
buf ( n297439 , n806 );
xor ( n7012 , n297438 , n297439 );
buf ( n297441 , n7012 );
buf ( n297442 , n297441 );
not ( n7015 , n297442 );
buf ( n297444 , n295437 );
not ( n297445 , n297444 );
or ( n7018 , n7015 , n297445 );
buf ( n7019 , n296617 );
buf ( n297448 , n296625 );
nand ( n297449 , n7019 , n297448 );
buf ( n297450 , n297449 );
buf ( n297451 , n297450 );
nand ( n7024 , n7018 , n297451 );
buf ( n297453 , n7024 );
buf ( n297454 , n297453 );
xor ( n7027 , n297437 , n297454 );
buf ( n297456 , n296819 );
not ( n297457 , n297456 );
buf ( n297458 , n297175 );
not ( n297459 , n297458 );
or ( n7032 , n297457 , n297459 );
buf ( n297461 , n292841 );
buf ( n7034 , n810 );
buf ( n297463 , n771 );
xor ( n297464 , n7034 , n297463 );
buf ( n297465 , n297464 );
buf ( n297466 , n297465 );
nand ( n7039 , n297461 , n297466 );
buf ( n7040 , n7039 );
buf ( n297469 , n7040 );
nand ( n297470 , n7032 , n297469 );
buf ( n297471 , n297470 );
buf ( n297472 , n297471 );
xor ( n297473 , n7027 , n297472 );
buf ( n297474 , n297473 );
not ( n7047 , n297474 );
xor ( n297476 , n297423 , n7047 );
buf ( n297477 , n297476 );
xor ( n7050 , n297309 , n297477 );
buf ( n297479 , n6706 );
buf ( n297480 , n296430 );
not ( n7053 , n297480 );
buf ( n7054 , n7053 );
buf ( n297483 , n7054 );
or ( n7056 , n297479 , n297483 );
buf ( n297485 , n297190 );
nand ( n297486 , n7056 , n297485 );
buf ( n297487 , n297486 );
buf ( n297488 , n297487 );
buf ( n297489 , n6706 );
buf ( n297490 , n7054 );
nand ( n7063 , n297489 , n297490 );
buf ( n297492 , n7063 );
buf ( n7065 , n297492 );
nand ( n7066 , n297488 , n7065 );
buf ( n297495 , n7066 );
buf ( n297496 , n297495 );
buf ( n297497 , n297265 );
not ( n7070 , n297497 );
buf ( n297499 , n297244 );
not ( n297500 , n297499 );
or ( n297501 , n7070 , n297500 );
buf ( n297502 , n297260 );
not ( n7075 , n297502 );
buf ( n297504 , n6813 );
not ( n297505 , n297504 );
or ( n7078 , n7075 , n297505 );
buf ( n297507 , n297230 );
nand ( n297508 , n7078 , n297507 );
buf ( n297509 , n297508 );
buf ( n297510 , n297509 );
nand ( n297511 , n297501 , n297510 );
buf ( n297512 , n297511 );
buf ( n297513 , n297512 );
xor ( n7086 , n297496 , n297513 );
xor ( n7087 , n296605 , n296652 );
xor ( n297516 , n7087 , n296711 );
buf ( n297517 , n297516 );
buf ( n297518 , n297517 );
and ( n7091 , n7086 , n297518 );
and ( n7092 , n297496 , n297513 );
or ( n297521 , n7091 , n7092 );
buf ( n297522 , n297521 );
buf ( n297523 , n297522 );
xor ( n7096 , n7050 , n297523 );
buf ( n297525 , n7096 );
buf ( n297526 , n297525 );
xor ( n7099 , n6875 , n297526 );
buf ( n297528 , n7099 );
buf ( n7101 , n297528 );
xor ( n7102 , n297496 , n297513 );
xor ( n7103 , n7102 , n297518 );
buf ( n7104 , n7103 );
buf ( n297533 , n7104 );
xor ( n7106 , n296853 , n297097 );
xor ( n7107 , n7106 , n297297 );
buf ( n7108 , n7107 );
buf ( n297537 , n7108 );
xor ( n7110 , n297533 , n297537 );
xor ( n7111 , n296914 , n296918 );
xor ( n7112 , n7111 , n297092 );
buf ( n297541 , n7112 );
buf ( n297542 , n297541 );
xor ( n7115 , n296870 , n296891 );
xor ( n7116 , n7115 , n296909 );
buf ( n297545 , n7116 );
buf ( n297546 , n297545 );
buf ( n297547 , n780 );
buf ( n297548 , n806 );
xor ( n7121 , n297547 , n297548 );
buf ( n297550 , n7121 );
buf ( n297551 , n297550 );
not ( n297552 , n297551 );
buf ( n297553 , n296617 );
not ( n7126 , n297553 );
or ( n7127 , n297552 , n7126 );
buf ( n297556 , n295437 );
buf ( n7129 , n296857 );
nand ( n7130 , n297556 , n7129 );
buf ( n297559 , n7130 );
buf ( n297560 , n297559 );
nand ( n297561 , n7127 , n297560 );
buf ( n297562 , n297561 );
buf ( n297563 , n297562 );
buf ( n297564 , n296890 );
not ( n7137 , n297564 );
buf ( n297566 , n7137 );
buf ( n7139 , n297566 );
xor ( n7140 , n297563 , n7139 );
buf ( n297569 , n787 );
buf ( n297570 , n800 );
xor ( n7143 , n297569 , n297570 );
buf ( n297572 , n7143 );
buf ( n297573 , n297572 );
not ( n297574 , n297573 );
buf ( n297575 , n296480 );
not ( n7148 , n297575 );
or ( n297577 , n297574 , n7148 );
buf ( n297578 , n6057 );
buf ( n297579 , n296923 );
nand ( n297580 , n297578 , n297579 );
buf ( n297581 , n297580 );
buf ( n297582 , n297581 );
nand ( n7155 , n297577 , n297582 );
buf ( n297584 , n7155 );
buf ( n297585 , n297584 );
buf ( n297586 , n785 );
buf ( n297587 , n802 );
xor ( n297588 , n297586 , n297587 );
buf ( n297589 , n297588 );
buf ( n297590 , n297589 );
not ( n297591 , n297590 );
buf ( n297592 , n296508 );
not ( n7165 , n297592 );
or ( n297594 , n297591 , n7165 );
buf ( n297595 , n296517 );
buf ( n297596 , n297016 );
nand ( n297597 , n297595 , n297596 );
buf ( n297598 , n297597 );
buf ( n297599 , n297598 );
nand ( n297600 , n297594 , n297599 );
buf ( n297601 , n297600 );
buf ( n297602 , n297601 );
or ( n297603 , n297585 , n297602 );
not ( n7176 , n296423 );
not ( n297605 , n296874 );
or ( n7178 , n7176 , n297605 );
and ( n7179 , n816 , n771 );
not ( n297608 , n816 );
and ( n297609 , n297608 , n5598 );
nor ( n7182 , n7179 , n297609 );
nand ( n297611 , n2118 , n7182 );
nand ( n297612 , n7178 , n297611 );
buf ( n297613 , n297612 );
nand ( n297614 , n297603 , n297613 );
buf ( n297615 , n297614 );
buf ( n297616 , n297615 );
buf ( n297617 , n297584 );
buf ( n297618 , n297601 );
nand ( n7191 , n297617 , n297618 );
buf ( n7192 , n7191 );
buf ( n297621 , n7192 );
nand ( n297622 , n297616 , n297621 );
buf ( n297623 , n297622 );
buf ( n297624 , n297623 );
and ( n297625 , n7140 , n297624 );
and ( n297626 , n297563 , n7139 );
or ( n297627 , n297625 , n297626 );
buf ( n297628 , n297627 );
buf ( n297629 , n297628 );
xor ( n7202 , n297546 , n297629 );
buf ( n297631 , n788 );
buf ( n297632 , n800 );
and ( n7205 , n297631 , n297632 );
buf ( n297634 , n7205 );
buf ( n297635 , n297634 );
buf ( n7208 , n779 );
buf ( n7209 , n808 );
xor ( n7210 , n7208 , n7209 );
buf ( n7211 , n7210 );
buf ( n297640 , n7211 );
not ( n297641 , n297640 );
buf ( n297642 , n293655 );
not ( n297643 , n297642 );
or ( n7216 , n297641 , n297643 );
not ( n7217 , n297059 );
nand ( n7218 , n7217 , n294557 );
buf ( n297647 , n7218 );
nand ( n297648 , n7216 , n297647 );
buf ( n297649 , n297648 );
buf ( n297650 , n297649 );
xor ( n7223 , n297635 , n297650 );
buf ( n297652 , n777 );
buf ( n297653 , n810 );
xor ( n297654 , n297652 , n297653 );
buf ( n297655 , n297654 );
buf ( n297656 , n297655 );
not ( n297657 , n297656 );
buf ( n297658 , n293058 );
not ( n7231 , n297658 );
or ( n297660 , n297657 , n7231 );
buf ( n297661 , n292841 );
buf ( n297662 , n296948 );
nand ( n297663 , n297661 , n297662 );
buf ( n297664 , n297663 );
buf ( n297665 , n297664 );
nand ( n7238 , n297660 , n297665 );
buf ( n297667 , n7238 );
buf ( n297668 , n297667 );
and ( n7241 , n7223 , n297668 );
and ( n297670 , n297635 , n297650 );
or ( n7243 , n7241 , n297670 );
buf ( n297672 , n7243 );
buf ( n297673 , n297672 );
xor ( n7246 , n812 , n775 );
buf ( n297675 , n7246 );
not ( n7248 , n297675 );
buf ( n297677 , n2376 );
not ( n7250 , n297677 );
or ( n297679 , n7248 , n7250 );
buf ( n297680 , n2383 );
buf ( n297681 , n296970 );
nand ( n297682 , n297680 , n297681 );
buf ( n297683 , n297682 );
buf ( n297684 , n297683 );
nand ( n7257 , n297679 , n297684 );
buf ( n297686 , n7257 );
buf ( n7259 , n297686 );
buf ( n297688 , n7259 );
not ( n297689 , n297688 );
buf ( n297690 , n781 );
buf ( n297691 , n806 );
xor ( n297692 , n297690 , n297691 );
buf ( n297693 , n297692 );
buf ( n297694 , n297693 );
not ( n297695 , n297694 );
buf ( n297696 , n296617 );
not ( n7269 , n297696 );
or ( n297698 , n297695 , n7269 );
buf ( n297699 , n295437 );
buf ( n297700 , n297550 );
nand ( n297701 , n297699 , n297700 );
buf ( n297702 , n297701 );
buf ( n297703 , n297702 );
nand ( n297704 , n297698 , n297703 );
buf ( n297705 , n297704 );
buf ( n297706 , n297705 );
not ( n297707 , n297706 );
or ( n7280 , n297689 , n297707 );
buf ( n297709 , n297705 );
buf ( n297710 , n297686 );
or ( n7283 , n297709 , n297710 );
buf ( n297712 , n783 );
buf ( n297713 , n804 );
xor ( n7286 , n297712 , n297713 );
buf ( n297715 , n7286 );
buf ( n297716 , n297715 );
not ( n7289 , n297716 );
buf ( n297718 , n296441 );
not ( n297719 , n297718 );
or ( n7292 , n7289 , n297719 );
buf ( n297721 , n6017 );
buf ( n297722 , n296992 );
nand ( n297723 , n297721 , n297722 );
buf ( n297724 , n297723 );
buf ( n297725 , n297724 );
nand ( n297726 , n7292 , n297725 );
buf ( n297727 , n297726 );
buf ( n297728 , n297727 );
nand ( n7301 , n7283 , n297728 );
buf ( n297730 , n7301 );
buf ( n297731 , n297730 );
nand ( n7304 , n7280 , n297731 );
buf ( n297733 , n7304 );
buf ( n297734 , n297733 );
xor ( n7307 , n297673 , n297734 );
buf ( n297736 , n769 );
buf ( n297737 , n818 );
xor ( n297738 , n297736 , n297737 );
buf ( n297739 , n297738 );
buf ( n297740 , n297739 );
not ( n297741 , n297740 );
buf ( n297742 , n291984 );
not ( n7315 , n297742 );
or ( n297744 , n297741 , n7315 );
buf ( n297745 , n291989 );
buf ( n297746 , n297041 );
nand ( n297747 , n297745 , n297746 );
buf ( n297748 , n297747 );
buf ( n297749 , n297748 );
nand ( n297750 , n297744 , n297749 );
buf ( n297751 , n297750 );
buf ( n297752 , n297751 );
buf ( n297753 , n291968 );
buf ( n297754 , n291722 );
or ( n7327 , n297753 , n297754 );
buf ( n297756 , n820 );
nand ( n297757 , n7327 , n297756 );
buf ( n297758 , n297757 );
buf ( n297759 , n297758 );
or ( n7332 , n297752 , n297759 );
buf ( n297761 , n773 );
buf ( n297762 , n814 );
xor ( n7335 , n297761 , n297762 );
buf ( n297764 , n7335 );
buf ( n297765 , n297764 );
not ( n7338 , n297765 );
buf ( n297767 , n2893 );
not ( n7340 , n297767 );
or ( n7341 , n7338 , n7340 );
buf ( n297770 , n292518 );
buf ( n297771 , n297067 );
nand ( n297772 , n297770 , n297771 );
buf ( n297773 , n297772 );
buf ( n297774 , n297773 );
nand ( n297775 , n7341 , n297774 );
buf ( n297776 , n297775 );
buf ( n297777 , n297776 );
nand ( n7350 , n7332 , n297777 );
buf ( n7351 , n7350 );
buf ( n297780 , n7351 );
buf ( n7353 , n297758 );
buf ( n297782 , n297751 );
nand ( n297783 , n7353 , n297782 );
buf ( n297784 , n297783 );
buf ( n297785 , n297784 );
nand ( n7358 , n297780 , n297785 );
buf ( n297787 , n7358 );
buf ( n297788 , n297787 );
and ( n7361 , n7307 , n297788 );
and ( n297790 , n297673 , n297734 );
or ( n7363 , n7361 , n297790 );
buf ( n297792 , n7363 );
buf ( n297793 , n297792 );
and ( n7366 , n7202 , n297793 );
and ( n297795 , n297546 , n297629 );
or ( n7368 , n7366 , n297795 );
buf ( n297797 , n7368 );
buf ( n297798 , n297797 );
xor ( n297799 , n297542 , n297798 );
xor ( n7372 , n297273 , n297276 );
xor ( n297801 , n7372 , n297281 );
buf ( n297802 , n297801 );
not ( n7375 , n297802 );
not ( n297804 , n297036 );
not ( n297805 , n297804 );
buf ( n7378 , n296966 );
nand ( n297807 , n297805 , n6660 , n7378 );
not ( n7380 , n7378 );
nand ( n297809 , n297804 , n6660 , n7380 );
not ( n7382 , n6660 );
nand ( n7383 , n297804 , n7378 , n7382 );
nand ( n297812 , n7382 , n297805 , n7380 );
nand ( n297813 , n297807 , n297809 , n7383 , n297812 );
not ( n7386 , n297813 );
or ( n7387 , n7375 , n7386 );
xor ( n297816 , n296966 , n297036 );
xor ( n297817 , n297816 , n7382 );
not ( n7390 , n297817 );
buf ( n297819 , n7390 );
buf ( n297820 , n297802 );
or ( n297821 , n297819 , n297820 );
buf ( n297822 , n296986 );
not ( n297823 , n297822 );
buf ( n297824 , n297823 );
xor ( n7397 , n297008 , n297824 );
xnor ( n297826 , n7397 , n297032 );
not ( n297827 , n297826 );
not ( n7400 , n297827 );
buf ( n297829 , n7400 );
not ( n7402 , n297829 );
xor ( n7403 , n297061 , n297083 );
not ( n297832 , n297053 );
xor ( n297833 , n7403 , n297832 );
buf ( n297834 , n297833 );
not ( n297835 , n297834 );
or ( n297836 , n7402 , n297835 );
not ( n7409 , n297833 );
not ( n297838 , n7409 );
not ( n297839 , n297827 );
or ( n7412 , n297838 , n297839 );
not ( n297841 , n296965 );
buf ( n297842 , n296961 );
nand ( n7415 , n297841 , n297842 );
not ( n297844 , n296943 );
nand ( n7417 , n297844 , n297842 );
not ( n7418 , n297842 );
nand ( n297847 , n7418 , n296964 , n6514 );
nor ( n297848 , n296964 , n6514 );
nand ( n7421 , n7418 , n297848 );
nand ( n297850 , n7415 , n7417 , n297847 , n7421 );
nand ( n7423 , n7412 , n297850 );
buf ( n297852 , n7423 );
nand ( n7425 , n297836 , n297852 );
buf ( n297854 , n7425 );
buf ( n297855 , n297854 );
nand ( n7428 , n297821 , n297855 );
buf ( n297857 , n7428 );
nand ( n7430 , n7387 , n297857 );
buf ( n297859 , n7430 );
and ( n7432 , n297799 , n297859 );
and ( n7433 , n297542 , n297798 );
or ( n7434 , n7432 , n7433 );
buf ( n297863 , n7434 );
buf ( n297864 , n297863 );
and ( n7437 , n7110 , n297864 );
and ( n7438 , n297533 , n297537 );
or ( n7439 , n7437 , n7438 );
buf ( n297868 , n7439 );
buf ( n297869 , n297868 );
and ( n7442 , n7101 , n297869 );
buf ( n297871 , n7442 );
not ( n7444 , n297871 );
or ( n7445 , n5985 , n7444 );
nand ( n7446 , n297528 , n297868 , n831 );
nand ( n297875 , n7445 , n7446 );
buf ( n7448 , n297875 );
not ( n7449 , n831 );
buf ( n297878 , n843 );
buf ( n297879 , n2376 );
buf ( n297880 , n2378 );
and ( n7453 , n297879 , n297880 );
buf ( n297882 , n2383 );
buf ( n297883 , n292813 );
and ( n297884 , n297882 , n297883 );
nor ( n297885 , n7453 , n297884 );
buf ( n297886 , n297885 );
xor ( n297887 , n297886 , n292787 );
xnor ( n7460 , n297887 , n2342 );
buf ( n297889 , n7460 );
xor ( n7462 , n292443 , n2066 );
xnor ( n297891 , n7462 , n2150 );
buf ( n297892 , n297891 );
xor ( n297893 , n297889 , n297892 );
buf ( n297894 , n292649 );
not ( n7467 , n297894 );
buf ( n297896 , n291788 );
not ( n297897 , n297896 );
or ( n297898 , n7467 , n297897 );
buf ( n297899 , n292393 );
xor ( n297900 , n818 , n794 );
buf ( n297901 , n297900 );
nand ( n7474 , n297899 , n297901 );
buf ( n297903 , n7474 );
buf ( n297904 , n297903 );
nand ( n7477 , n297898 , n297904 );
buf ( n297906 , n7477 );
buf ( n297907 , n297906 );
not ( n297908 , n297907 );
not ( n7481 , n292450 );
not ( n297910 , n831 );
or ( n7483 , n7481 , n297910 );
buf ( n297912 , n783 );
buf ( n297913 , n830 );
xor ( n7486 , n297912 , n297913 );
buf ( n297915 , n7486 );
buf ( n297916 , n297915 );
not ( n7489 , n297916 );
buf ( n297918 , n7489 );
or ( n297919 , n297918 , n291653 );
nand ( n297920 , n7483 , n297919 );
buf ( n297921 , n297920 );
buf ( n297922 , n799 );
buf ( n297923 , n815 );
nand ( n7496 , n297922 , n297923 );
buf ( n297925 , n7496 );
or ( n7498 , n799 , n815 );
nand ( n7499 , n7498 , n816 );
and ( n297928 , n297925 , n814 , n7499 );
buf ( n7501 , n297928 );
nand ( n7502 , n297921 , n7501 );
buf ( n7503 , n7502 );
buf ( n297932 , n7503 );
nand ( n7505 , n297908 , n297932 );
buf ( n7506 , n7505 );
buf ( n297935 , n7506 );
not ( n7508 , n297935 );
buf ( n297937 , n292529 );
not ( n297938 , n297937 );
buf ( n297939 , n296423 );
not ( n7512 , n297939 );
or ( n297941 , n297938 , n7512 );
buf ( n297942 , n292892 );
xor ( n297943 , n816 , n797 );
buf ( n7516 , n297943 );
nand ( n7517 , n297942 , n7516 );
buf ( n7518 , n7517 );
buf ( n297947 , n7518 );
nand ( n7520 , n297941 , n297947 );
buf ( n7521 , n7520 );
not ( n297950 , n7521 );
xor ( n7523 , n824 , n789 );
not ( n297952 , n7523 );
nand ( n297953 , n292464 , n292471 , n1402 );
not ( n7526 , n297953 );
not ( n297955 , n7526 );
or ( n297956 , n297952 , n297955 );
nand ( n7529 , n292461 , n1613 );
nand ( n297958 , n297956 , n7529 );
not ( n7531 , n297958 );
or ( n7532 , n297950 , n7531 );
buf ( n297961 , n7521 );
buf ( n297962 , n297958 );
nor ( n7535 , n297961 , n297962 );
buf ( n297964 , n7535 );
buf ( n297965 , n799 );
buf ( n297966 , n814 );
xor ( n297967 , n297965 , n297966 );
buf ( n297968 , n297967 );
buf ( n297969 , n297968 );
not ( n297970 , n297969 );
buf ( n297971 , n292509 );
not ( n7544 , n297971 );
or ( n297973 , n297970 , n7544 );
buf ( n297974 , n2089 );
buf ( n297975 , n292500 );
nand ( n297976 , n297974 , n297975 );
buf ( n297977 , n297976 );
buf ( n297978 , n297977 );
nand ( n7551 , n297973 , n297978 );
buf ( n297980 , n7551 );
buf ( n297981 , n297980 );
not ( n7554 , n297981 );
buf ( n297983 , n7554 );
or ( n297984 , n297964 , n297983 );
nand ( n7557 , n7532 , n297984 );
buf ( n297986 , n7557 );
not ( n297987 , n297986 );
or ( n7560 , n7508 , n297987 );
buf ( n297989 , n7503 );
not ( n7562 , n297989 );
buf ( n297991 , n297906 );
nand ( n297992 , n7562 , n297991 );
buf ( n297993 , n297992 );
buf ( n297994 , n297993 );
nand ( n297995 , n7560 , n297994 );
buf ( n297996 , n297995 );
buf ( n297997 , n297996 );
xor ( n297998 , n297893 , n297997 );
buf ( n297999 , n297998 );
buf ( n298000 , n297999 );
and ( n298001 , n292725 , n799 );
buf ( n298002 , n784 );
buf ( n298003 , n830 );
xor ( n298004 , n298002 , n298003 );
buf ( n298005 , n298004 );
buf ( n298006 , n298005 );
not ( n7579 , n298006 );
buf ( n298008 , n291656 );
not ( n298009 , n298008 );
or ( n298010 , n7579 , n298009 );
buf ( n298011 , n297915 );
buf ( n298012 , n831 );
nand ( n298013 , n298011 , n298012 );
buf ( n298014 , n298013 );
buf ( n298015 , n298014 );
nand ( n7588 , n298010 , n298015 );
buf ( n298017 , n7588 );
or ( n298018 , n298001 , n298017 );
buf ( n298019 , n786 );
buf ( n298020 , n828 );
xor ( n298021 , n298019 , n298020 );
buf ( n298022 , n298021 );
buf ( n298023 , n298022 );
not ( n298024 , n298023 );
buf ( n298025 , n291808 );
not ( n298026 , n298025 );
or ( n7599 , n298024 , n298026 );
buf ( n298028 , n291939 );
buf ( n298029 , n785 );
buf ( n298030 , n828 );
xor ( n298031 , n298029 , n298030 );
buf ( n298032 , n298031 );
buf ( n298033 , n298032 );
nand ( n298034 , n298028 , n298033 );
buf ( n298035 , n298034 );
buf ( n298036 , n298035 );
nand ( n298037 , n7599 , n298036 );
buf ( n298038 , n298037 );
nand ( n7611 , n298018 , n298038 );
buf ( n298040 , n7611 );
buf ( n298041 , n292725 );
buf ( n298042 , n799 );
nand ( n7615 , n298041 , n298042 );
buf ( n7616 , n7615 );
buf ( n298045 , n7616 );
not ( n7618 , n298045 );
buf ( n298047 , n298017 );
nand ( n298048 , n7618 , n298047 );
buf ( n298049 , n298048 );
buf ( n298050 , n298049 );
nand ( n298051 , n298040 , n298050 );
buf ( n298052 , n298051 );
buf ( n298053 , n298052 );
buf ( n7626 , n796 );
buf ( n298055 , n818 );
xor ( n298056 , n7626 , n298055 );
buf ( n298057 , n298056 );
buf ( n298058 , n298057 );
not ( n7631 , n298058 );
buf ( n298060 , n292393 );
not ( n298061 , n298060 );
or ( n7634 , n7631 , n298061 );
buf ( n298063 , n291788 );
xor ( n298064 , n818 , n795 );
buf ( n298065 , n298064 );
nand ( n298066 , n298063 , n298065 );
buf ( n298067 , n298066 );
buf ( n298068 , n298067 );
nand ( n298069 , n7634 , n298068 );
buf ( n298070 , n298069 );
buf ( n298071 , n298070 );
not ( n7644 , n298071 );
buf ( n298073 , n788 );
buf ( n298074 , n826 );
xor ( n298075 , n298073 , n298074 );
buf ( n298076 , n298075 );
not ( n7649 , n298076 );
not ( n298078 , n291880 );
or ( n298079 , n7649 , n298078 );
buf ( n298080 , n291886 );
buf ( n298081 , n787 );
buf ( n298082 , n826 );
xor ( n7655 , n298081 , n298082 );
buf ( n298084 , n7655 );
buf ( n298085 , n298084 );
nand ( n7658 , n298080 , n298085 );
buf ( n298087 , n7658 );
nand ( n7660 , n298079 , n298087 );
buf ( n298089 , n7660 );
not ( n7662 , n298089 );
or ( n7663 , n7644 , n7662 );
or ( n7664 , n298070 , n7660 );
buf ( n7665 , n794 );
buf ( n7666 , n820 );
xor ( n7667 , n7665 , n7666 );
buf ( n7668 , n7667 );
not ( n298097 , n7668 );
not ( n7670 , n291719 );
nor ( n298099 , n7670 , n291714 );
not ( n298100 , n298099 );
or ( n7673 , n298097 , n298100 );
buf ( n298102 , n1995 );
buf ( n7675 , n793 );
buf ( n7676 , n820 );
xor ( n7677 , n7675 , n7676 );
buf ( n7678 , n7677 );
buf ( n298107 , n7678 );
nand ( n298108 , n298102 , n298107 );
buf ( n298109 , n298108 );
nand ( n7682 , n7673 , n298109 );
nand ( n298111 , n7664 , n7682 );
buf ( n298112 , n298111 );
nand ( n298113 , n7663 , n298112 );
buf ( n298114 , n298113 );
buf ( n298115 , n298114 );
xor ( n7688 , n298053 , n298115 );
xor ( n298117 , n824 , n790 );
buf ( n298118 , n298117 );
not ( n298119 , n298118 );
buf ( n298120 , n291835 );
not ( n7693 , n298120 );
or ( n7694 , n298119 , n7693 );
buf ( n7695 , n1613 );
buf ( n298124 , n7523 );
nand ( n7697 , n7695 , n298124 );
buf ( n7698 , n7697 );
buf ( n7699 , n7698 );
nand ( n7700 , n7694 , n7699 );
buf ( n7701 , n7700 );
buf ( n298130 , n7701 );
buf ( n298131 , n792 );
buf ( n298132 , n822 );
xor ( n7705 , n298131 , n298132 );
buf ( n298134 , n7705 );
buf ( n298135 , n298134 );
not ( n7708 , n298135 );
buf ( n298137 , n291761 );
not ( n7710 , n298137 );
or ( n7711 , n7708 , n7710 );
buf ( n298140 , n292105 );
xor ( n298141 , n822 , n791 );
buf ( n298142 , n298141 );
nand ( n7715 , n298140 , n298142 );
buf ( n298144 , n7715 );
buf ( n298145 , n298144 );
nand ( n7718 , n7711 , n298145 );
buf ( n298147 , n7718 );
buf ( n298148 , n298147 );
xor ( n298149 , n298130 , n298148 );
buf ( n298150 , n798 );
buf ( n298151 , n816 );
xor ( n298152 , n298150 , n298151 );
buf ( n298153 , n298152 );
buf ( n298154 , n298153 );
not ( n298155 , n298154 );
buf ( n298156 , n2118 );
not ( n298157 , n298156 );
or ( n7730 , n298155 , n298157 );
buf ( n298159 , n296423 );
buf ( n298160 , n297943 );
nand ( n7733 , n298159 , n298160 );
buf ( n298162 , n7733 );
buf ( n7735 , n298162 );
nand ( n298164 , n7730 , n7735 );
buf ( n298165 , n298164 );
buf ( n298166 , n298165 );
and ( n298167 , n298149 , n298166 );
and ( n7740 , n298130 , n298148 );
or ( n7741 , n298167 , n7740 );
buf ( n298170 , n7741 );
buf ( n298171 , n298170 );
and ( n7744 , n7688 , n298171 );
and ( n298173 , n298053 , n298115 );
or ( n7746 , n7744 , n298173 );
buf ( n298175 , n7746 );
not ( n298176 , n292455 );
not ( n298177 , n292488 );
or ( n298178 , n298176 , n298177 );
not ( n7751 , n292452 );
nand ( n298180 , n7751 , n2026 , n799 );
nand ( n298181 , n298178 , n298180 );
xor ( n298182 , n298181 , n292484 );
buf ( n298183 , n298141 );
not ( n298184 , n298183 );
buf ( n298185 , n291761 );
not ( n298186 , n298185 );
or ( n298187 , n298184 , n298186 );
buf ( n298188 , n1600 );
buf ( n298189 , n292626 );
nand ( n298190 , n298188 , n298189 );
buf ( n298191 , n298190 );
buf ( n298192 , n298191 );
nand ( n7765 , n298187 , n298192 );
buf ( n298194 , n7765 );
not ( n298195 , n298194 );
not ( n298196 , n298084 );
not ( n7769 , n1453 );
or ( n298198 , n298196 , n7769 );
buf ( n298199 , n291886 );
buf ( n298200 , n292603 );
nand ( n298201 , n298199 , n298200 );
buf ( n298202 , n298201 );
nand ( n7775 , n298198 , n298202 );
not ( n298204 , n7775 );
or ( n298205 , n298195 , n298204 );
not ( n298206 , n298194 );
not ( n7779 , n298206 );
not ( n298208 , n7775 );
not ( n298209 , n298208 );
or ( n7782 , n7779 , n298209 );
nand ( n298211 , n298032 , n291808 );
buf ( n298212 , n291939 );
buf ( n298213 , n292561 );
nand ( n298214 , n298212 , n298213 );
buf ( n298215 , n298214 );
nand ( n7788 , n298211 , n298215 );
nand ( n298217 , n7782 , n7788 );
nand ( n298218 , n298205 , n298217 );
xor ( n7791 , n298182 , n298218 );
not ( n298220 , n292599 );
not ( n7793 , n292645 );
not ( n7794 , n7793 );
or ( n7795 , n298220 , n7794 );
not ( n7796 , n292599 );
nand ( n7797 , n292645 , n7796 );
nand ( n298226 , n7795 , n7797 );
and ( n298227 , n298226 , n2187 );
not ( n7800 , n298226 );
not ( n298229 , n2187 );
and ( n7802 , n7800 , n298229 );
nor ( n7803 , n298227 , n7802 );
xor ( n7804 , n7791 , n7803 );
xor ( n7805 , n298175 , n7804 );
not ( n7806 , n297900 );
not ( n7807 , n291989 );
or ( n298236 , n7806 , n7807 );
not ( n298237 , n1355 );
nand ( n7810 , n298237 , n298064 , n2997 );
nand ( n298239 , n298236 , n7810 );
buf ( n298240 , n298239 );
not ( n7813 , n2155 );
not ( n298242 , n291906 );
or ( n7815 , n7813 , n298242 );
nand ( n7816 , n7678 , n291722 );
nand ( n298245 , n7815 , n7816 );
buf ( n7818 , n298245 );
xor ( n7819 , n298240 , n7818 );
xor ( n298248 , n297928 , n297920 );
buf ( n298249 , n298248 );
xor ( n7822 , n7819 , n298249 );
buf ( n298251 , n7822 );
buf ( n298252 , n298251 );
not ( n7825 , n298252 );
not ( n7826 , n291939 );
not ( n298255 , n292561 );
or ( n298256 , n7826 , n298255 );
nand ( n7829 , n298256 , n298211 );
xor ( n298258 , n7829 , n298194 );
and ( n298259 , n298258 , n298208 );
not ( n7832 , n298258 );
and ( n298261 , n7832 , n7775 );
or ( n7834 , n298259 , n298261 );
buf ( n298263 , n7834 );
not ( n298264 , n298263 );
or ( n298265 , n7825 , n298264 );
buf ( n298266 , n7834 );
buf ( n298267 , n298251 );
or ( n298268 , n298266 , n298267 );
not ( n7841 , n7521 );
nand ( n298270 , n7841 , n297958 , n297983 );
not ( n298271 , n297983 );
nand ( n7844 , n298271 , n297958 , n7521 );
nor ( n7845 , n7841 , n297958 );
nand ( n7846 , n297983 , n7845 );
nand ( n7847 , n297980 , n297964 );
nand ( n298276 , n298270 , n7844 , n7846 , n7847 );
buf ( n298277 , n298276 );
nand ( n7850 , n298268 , n298277 );
buf ( n7851 , n7850 );
buf ( n298280 , n7851 );
nand ( n298281 , n298265 , n298280 );
buf ( n298282 , n298281 );
and ( n298283 , n7805 , n298282 );
and ( n298284 , n298175 , n7804 );
or ( n7857 , n298283 , n298284 );
buf ( n298286 , n7857 );
xor ( n298287 , n298000 , n298286 );
xor ( n7860 , n298182 , n298218 );
and ( n298289 , n7860 , n7803 );
and ( n7862 , n298182 , n298218 );
or ( n7863 , n298289 , n7862 );
xor ( n298292 , n298240 , n7818 );
and ( n298293 , n298292 , n298249 );
and ( n7866 , n298240 , n7818 );
or ( n298295 , n298293 , n7866 );
buf ( n298296 , n298295 );
not ( n7869 , n298296 );
not ( n298298 , n292527 );
not ( n298299 , n292557 );
not ( n7872 , n2145 );
or ( n298301 , n298299 , n7872 );
or ( n298302 , n2145 , n292557 );
nand ( n298303 , n298301 , n298302 );
not ( n298304 , n298303 );
or ( n7877 , n298298 , n298304 );
or ( n298306 , n298303 , n292527 );
nand ( n298307 , n7877 , n298306 );
not ( n7880 , n298307 );
nand ( n298309 , n7869 , n7880 );
not ( n7882 , n298309 );
and ( n7883 , n297906 , n7503 );
not ( n7884 , n297906 );
and ( n298313 , n297920 , n297928 );
and ( n7886 , n7884 , n298313 );
or ( n7887 , n7883 , n7886 );
xor ( n7888 , n7887 , n7557 );
not ( n7889 , n7888 );
or ( n7890 , n7882 , n7889 );
nand ( n7891 , n298296 , n298307 );
nand ( n7892 , n7890 , n7891 );
xor ( n7893 , n7863 , n7892 );
buf ( n298322 , n2315 );
nor ( n7895 , n2219 , n2262 );
nand ( n7896 , n298322 , n7895 );
and ( n298325 , n2262 , n2219 );
nand ( n7898 , n298322 , n298325 );
not ( n298327 , n292747 );
buf ( n7900 , n292744 );
nand ( n298329 , n298327 , n7900 );
not ( n298330 , n2263 );
nand ( n7903 , n7900 , n298330 );
nand ( n7904 , n7896 , n7898 , n298329 , n7903 );
xor ( n7905 , n7893 , n7904 );
buf ( n298334 , n7905 );
and ( n7907 , n298287 , n298334 );
and ( n7908 , n298000 , n298286 );
or ( n7909 , n7907 , n7908 );
buf ( n298338 , n7909 );
buf ( n298339 , n298338 );
xor ( n298340 , n297878 , n298339 );
xor ( n7913 , n297889 , n297892 );
and ( n7914 , n7913 , n297997 );
and ( n7915 , n297889 , n297892 );
or ( n7916 , n7914 , n7915 );
buf ( n298345 , n7916 );
buf ( n298346 , n298345 );
xor ( n7919 , n7863 , n7892 );
and ( n7920 , n7919 , n7904 );
and ( n7921 , n7863 , n7892 );
or ( n7922 , n7920 , n7921 );
buf ( n298351 , n7922 );
xor ( n7924 , n298346 , n298351 );
xor ( n7925 , n292837 , n293001 );
xor ( n298354 , n7925 , n293006 );
buf ( n298355 , n298354 );
buf ( n298356 , n298355 );
xor ( n7929 , n7924 , n298356 );
buf ( n298358 , n7929 );
buf ( n298359 , n298358 );
and ( n7932 , n298340 , n298359 );
and ( n7933 , n297878 , n298339 );
or ( n298362 , n7932 , n7933 );
buf ( n298363 , n298362 );
not ( n7936 , n298363 );
or ( n298365 , n7449 , n7936 );
buf ( n298366 , n831 );
not ( n7939 , n298366 );
buf ( n298368 , n875 );
buf ( n298369 , n298338 );
xor ( n7942 , n298368 , n298369 );
buf ( n298371 , n298358 );
and ( n7944 , n7942 , n298371 );
and ( n7945 , n298368 , n298369 );
or ( n7946 , n7944 , n7945 );
buf ( n298375 , n7946 );
buf ( n7948 , n298375 );
nand ( n7949 , n7939 , n7948 );
buf ( n298378 , n7949 );
nand ( n7951 , n298365 , n298378 );
buf ( n298380 , n7951 );
buf ( n298381 , n831 );
not ( n7954 , n298381 );
xor ( n7955 , n802 , n794 );
not ( n298384 , n7955 );
not ( n7957 , n296501 );
not ( n7958 , n802 );
or ( n7959 , n7957 , n7958 );
nand ( n7960 , n7959 , n6078 );
not ( n298389 , n7960 );
or ( n298390 , n298384 , n298389 );
xor ( n7963 , n802 , n793 );
nand ( n298392 , n296749 , n7963 );
nand ( n7965 , n298390 , n298392 );
buf ( n298394 , n7965 );
not ( n298395 , n298394 );
buf ( n298396 , n298395 );
not ( n7969 , n298396 );
xor ( n7970 , n816 , n780 );
buf ( n298399 , n7970 );
not ( n298400 , n298399 );
buf ( n298401 , n292892 );
not ( n298402 , n298401 );
or ( n7975 , n298400 , n298402 );
and ( n7976 , n779 , n292885 );
not ( n298405 , n779 );
and ( n7978 , n298405 , n816 );
or ( n7979 , n7976 , n7978 );
nand ( n298408 , n7979 , n1712 );
buf ( n298409 , n298408 );
nand ( n298410 , n7975 , n298409 );
buf ( n298411 , n298410 );
not ( n7984 , n298411 );
or ( n298413 , n7969 , n7984 );
buf ( n298414 , n298411 );
not ( n7987 , n298414 );
buf ( n298416 , n7965 );
nand ( n7989 , n7987 , n298416 );
buf ( n298418 , n7989 );
nand ( n298419 , n298413 , n298418 );
not ( n298420 , n6049 );
buf ( n298421 , n800 );
not ( n298422 , n298421 );
buf ( n298423 , n298422 );
and ( n7996 , n796 , n298423 );
not ( n298425 , n796 );
and ( n298426 , n298425 , n800 );
or ( n7999 , n7996 , n298426 );
not ( n298428 , n7999 );
or ( n298429 , n298420 , n298428 );
buf ( n298430 , n6057 );
buf ( n8003 , n795 );
buf ( n8004 , n800 );
xor ( n8005 , n8003 , n8004 );
buf ( n8006 , n8005 );
buf ( n298435 , n8006 );
nand ( n298436 , n298430 , n298435 );
buf ( n298437 , n298436 );
nand ( n8010 , n298429 , n298437 );
and ( n298439 , n298419 , n8010 );
not ( n298440 , n298419 );
not ( n8013 , n8010 );
and ( n298442 , n298440 , n8013 );
nor ( n8015 , n298439 , n298442 );
not ( n8016 , n8015 );
not ( n298445 , n8016 );
buf ( n298446 , n784 );
buf ( n298447 , n812 );
xor ( n298448 , n298446 , n298447 );
buf ( n298449 , n298448 );
buf ( n298450 , n298449 );
not ( n298451 , n298450 );
buf ( n298452 , n2373 );
not ( n8025 , n298452 );
or ( n298454 , n298451 , n8025 );
buf ( n298455 , n292810 );
buf ( n298456 , n783 );
buf ( n298457 , n812 );
xor ( n298458 , n298456 , n298457 );
buf ( n298459 , n298458 );
buf ( n298460 , n298459 );
nand ( n8033 , n298455 , n298460 );
buf ( n298462 , n8033 );
buf ( n298463 , n298462 );
nand ( n298464 , n298454 , n298463 );
buf ( n298465 , n298464 );
buf ( n298466 , n298465 );
not ( n298467 , n298466 );
xor ( n8040 , n814 , n782 );
buf ( n298469 , n8040 );
not ( n298470 , n298469 );
buf ( n298471 , n2893 );
not ( n8044 , n298471 );
or ( n8045 , n298470 , n8044 );
buf ( n298474 , n2089 );
buf ( n298475 , n781 );
buf ( n298476 , n814 );
xor ( n8049 , n298475 , n298476 );
buf ( n298478 , n8049 );
buf ( n298479 , n298478 );
nand ( n298480 , n298474 , n298479 );
buf ( n298481 , n298480 );
buf ( n298482 , n298481 );
nand ( n298483 , n8045 , n298482 );
buf ( n298484 , n298483 );
buf ( n8057 , n298484 );
not ( n298486 , n8057 );
buf ( n298487 , n298486 );
buf ( n298488 , n298487 );
not ( n8061 , n298488 );
or ( n8062 , n298467 , n8061 );
buf ( n298491 , n298465 );
buf ( n298492 , n298487 );
or ( n298493 , n298491 , n298492 );
nand ( n8066 , n8062 , n298493 );
buf ( n8067 , n8066 );
buf ( n298496 , n8067 );
xor ( n8069 , n776 , n820 );
buf ( n298498 , n8069 );
not ( n298499 , n298498 );
buf ( n298500 , n291722 );
not ( n298501 , n298500 );
or ( n8074 , n298499 , n298501 );
buf ( n298503 , n291906 );
buf ( n298504 , n775 );
buf ( n298505 , n820 );
xor ( n298506 , n298504 , n298505 );
buf ( n298507 , n298506 );
buf ( n298508 , n298507 );
nand ( n8081 , n298503 , n298508 );
buf ( n298510 , n8081 );
buf ( n298511 , n298510 );
nand ( n8084 , n8074 , n298511 );
buf ( n298513 , n8084 );
buf ( n298514 , n298513 );
xnor ( n8087 , n298496 , n298514 );
buf ( n298516 , n8087 );
not ( n8089 , n298516 );
or ( n298518 , n298445 , n8089 );
xor ( n298519 , n804 , n793 );
buf ( n298520 , n298519 );
not ( n8093 , n298520 );
not ( n298522 , n5231 );
buf ( n298523 , n298522 );
not ( n8096 , n298523 );
or ( n298525 , n8093 , n8096 );
xor ( n298526 , n805 , n806 );
buf ( n298527 , n298526 );
buf ( n298528 , n792 );
buf ( n298529 , n804 );
xor ( n8102 , n298528 , n298529 );
buf ( n298531 , n8102 );
buf ( n298532 , n298531 );
nand ( n8105 , n298527 , n298532 );
buf ( n298534 , n8105 );
buf ( n298535 , n298534 );
nand ( n298536 , n298525 , n298535 );
buf ( n298537 , n298536 );
buf ( n298538 , n298537 );
buf ( n298539 , n779 );
buf ( n298540 , n818 );
xor ( n8113 , n298539 , n298540 );
buf ( n298542 , n8113 );
buf ( n298543 , n298542 );
not ( n298544 , n298543 );
buf ( n298545 , n292393 );
not ( n8118 , n298545 );
or ( n298547 , n298544 , n8118 );
buf ( n298548 , n291989 );
xor ( n8121 , n818 , n778 );
buf ( n298550 , n8121 );
nand ( n8123 , n298548 , n298550 );
buf ( n298552 , n8123 );
buf ( n298553 , n298552 );
nand ( n8126 , n298547 , n298553 );
buf ( n298555 , n8126 );
buf ( n298556 , n298555 );
xor ( n298557 , n298538 , n298556 );
buf ( n298558 , n791 );
buf ( n298559 , n806 );
xor ( n298560 , n298558 , n298559 );
buf ( n298561 , n298560 );
buf ( n298562 , n298561 );
not ( n8135 , n298562 );
buf ( n298564 , n296617 );
not ( n298565 , n298564 );
or ( n298566 , n8135 , n298565 );
buf ( n298567 , n295437 );
xor ( n298568 , n806 , n790 );
buf ( n298569 , n298568 );
nand ( n8142 , n298567 , n298569 );
buf ( n8143 , n8142 );
buf ( n298572 , n8143 );
nand ( n298573 , n298566 , n298572 );
buf ( n298574 , n298573 );
buf ( n298575 , n298574 );
and ( n298576 , n298557 , n298575 );
and ( n8149 , n298538 , n298556 );
or ( n298578 , n298576 , n8149 );
buf ( n298579 , n298578 );
nand ( n8152 , n298518 , n298579 );
or ( n8153 , n298516 , n8016 );
nand ( n298582 , n8152 , n8153 );
not ( n298583 , n298582 );
buf ( n298584 , n772 );
buf ( n298585 , n824 );
xor ( n8158 , n298584 , n298585 );
buf ( n298587 , n8158 );
not ( n298588 , n298587 );
not ( n8161 , n291835 );
or ( n8162 , n298588 , n8161 );
buf ( n298591 , n291842 );
buf ( n298592 , n771 );
buf ( n298593 , n824 );
xor ( n298594 , n298592 , n298593 );
buf ( n298595 , n298594 );
buf ( n298596 , n298595 );
nand ( n8169 , n298591 , n298596 );
buf ( n298598 , n8169 );
nand ( n298599 , n8162 , n298598 );
buf ( n8172 , n298599 );
buf ( n8173 , n786 );
buf ( n8174 , n810 );
xor ( n8175 , n8173 , n8174 );
buf ( n8176 , n8175 );
buf ( n8177 , n8176 );
not ( n8178 , n8177 );
buf ( n8179 , n3041 );
not ( n8180 , n8179 );
or ( n8181 , n8178 , n8180 );
buf ( n8182 , n295259 );
buf ( n298611 , n785 );
buf ( n298612 , n810 );
xor ( n298613 , n298611 , n298612 );
buf ( n298614 , n298613 );
buf ( n298615 , n298614 );
nand ( n298616 , n8182 , n298615 );
buf ( n298617 , n298616 );
buf ( n298618 , n298617 );
nand ( n298619 , n8181 , n298618 );
buf ( n298620 , n298619 );
buf ( n298621 , n298620 );
xor ( n8194 , n8172 , n298621 );
buf ( n298623 , n788 );
buf ( n298624 , n808 );
xor ( n298625 , n298623 , n298624 );
buf ( n298626 , n298625 );
buf ( n298627 , n298626 );
not ( n298628 , n298627 );
buf ( n298629 , n293655 );
not ( n298630 , n298629 );
or ( n8203 , n298628 , n298630 );
buf ( n298632 , n6301 );
buf ( n8205 , n787 );
buf ( n298634 , n808 );
xor ( n298635 , n8205 , n298634 );
buf ( n298636 , n298635 );
buf ( n298637 , n298636 );
nand ( n298638 , n298632 , n298637 );
buf ( n298639 , n298638 );
buf ( n298640 , n298639 );
nand ( n298641 , n8203 , n298640 );
buf ( n298642 , n298641 );
buf ( n298643 , n298642 );
and ( n8216 , n8194 , n298643 );
and ( n8217 , n8172 , n298621 );
or ( n298646 , n8216 , n8217 );
buf ( n298647 , n298646 );
not ( n8220 , n298647 );
buf ( n298649 , n298531 );
not ( n298650 , n298649 );
buf ( n298651 , n295660 );
not ( n298652 , n298651 );
or ( n298653 , n298650 , n298652 );
buf ( n298654 , n295361 );
buf ( n298655 , n791 );
buf ( n298656 , n804 );
xor ( n298657 , n298655 , n298656 );
buf ( n298658 , n298657 );
buf ( n298659 , n298658 );
nand ( n298660 , n298654 , n298659 );
buf ( n298661 , n298660 );
buf ( n298662 , n298661 );
nand ( n298663 , n298653 , n298662 );
buf ( n298664 , n298663 );
buf ( n298665 , n298664 );
buf ( n298666 , n298568 );
not ( n298667 , n298666 );
buf ( n298668 , n5676 );
not ( n298669 , n298668 );
or ( n298670 , n298667 , n298669 );
buf ( n298671 , n295437 );
buf ( n298672 , n789 );
buf ( n298673 , n806 );
xor ( n8246 , n298672 , n298673 );
buf ( n8247 , n8246 );
buf ( n298676 , n8247 );
nand ( n8249 , n298671 , n298676 );
buf ( n298678 , n8249 );
buf ( n298679 , n298678 );
nand ( n8252 , n298670 , n298679 );
buf ( n8253 , n8252 );
buf ( n298682 , n8253 );
xor ( n8255 , n298665 , n298682 );
buf ( n298684 , n8121 );
not ( n298685 , n298684 );
buf ( n298686 , n292393 );
not ( n8259 , n298686 );
or ( n298688 , n298685 , n8259 );
buf ( n298689 , n291788 );
buf ( n298690 , n777 );
buf ( n298691 , n818 );
xor ( n8264 , n298690 , n298691 );
buf ( n298693 , n8264 );
buf ( n298694 , n298693 );
nand ( n298695 , n298689 , n298694 );
buf ( n298696 , n298695 );
buf ( n298697 , n298696 );
nand ( n8270 , n298688 , n298697 );
buf ( n298699 , n8270 );
buf ( n298700 , n298699 );
and ( n298701 , n8255 , n298700 );
and ( n8274 , n298665 , n298682 );
or ( n298703 , n298701 , n8274 );
buf ( n298704 , n298703 );
and ( n8277 , n8220 , n298704 );
not ( n298706 , n8220 );
not ( n298707 , n298704 );
and ( n8280 , n298706 , n298707 );
nor ( n8281 , n8277 , n8280 );
not ( n298710 , n298484 );
or ( n8283 , n298465 , n298513 );
not ( n298712 , n8283 );
or ( n8285 , n298710 , n298712 );
buf ( n298714 , n298513 );
buf ( n298715 , n298465 );
nand ( n298716 , n298714 , n298715 );
buf ( n298717 , n298716 );
nand ( n298718 , n8285 , n298717 );
and ( n298719 , n8281 , n298718 );
not ( n8292 , n8281 );
not ( n298721 , n298718 );
and ( n298722 , n8292 , n298721 );
nor ( n8295 , n298719 , n298722 );
not ( n8296 , n8295 );
not ( n298725 , n8296 );
or ( n298726 , n298583 , n298725 );
xnor ( n8299 , n8281 , n298718 );
or ( n298728 , n8299 , n298582 );
xor ( n298729 , n8172 , n298621 );
xor ( n8302 , n298729 , n298643 );
buf ( n298731 , n8302 );
buf ( n298732 , n797 );
buf ( n298733 , n800 );
and ( n298734 , n298732 , n298733 );
buf ( n298735 , n298734 );
buf ( n298736 , n770 );
buf ( n298737 , n826 );
xor ( n298738 , n298736 , n298737 );
buf ( n298739 , n298738 );
buf ( n298740 , n298739 );
not ( n298741 , n298740 );
buf ( n298742 , n295643 );
not ( n298743 , n298742 );
or ( n298744 , n298741 , n298743 );
not ( n8317 , n291885 );
not ( n298746 , n8317 );
buf ( n298747 , n298746 );
buf ( n298748 , n769 );
buf ( n298749 , n826 );
xor ( n8322 , n298748 , n298749 );
buf ( n298751 , n8322 );
buf ( n298752 , n298751 );
nand ( n8325 , n298747 , n298752 );
buf ( n298754 , n8325 );
buf ( n298755 , n298754 );
nand ( n8328 , n298744 , n298755 );
buf ( n298757 , n8328 );
xor ( n298758 , n298735 , n298757 );
buf ( n298759 , n774 );
buf ( n298760 , n822 );
xor ( n8333 , n298759 , n298760 );
buf ( n298762 , n8333 );
buf ( n298763 , n298762 );
not ( n298764 , n298763 );
not ( n8337 , n291757 );
and ( n298766 , n824 , n823 );
not ( n298767 , n824 );
not ( n8340 , n823 );
and ( n298769 , n298767 , n8340 );
nor ( n8342 , n298766 , n298769 );
nor ( n298771 , n8337 , n8342 );
buf ( n298772 , n298771 );
not ( n8345 , n298772 );
or ( n298774 , n298764 , n8345 );
buf ( n298775 , n292104 );
and ( n8348 , n773 , n822 );
not ( n298777 , n773 );
and ( n8350 , n298777 , n1299 );
nor ( n8351 , n8348 , n8350 );
buf ( n298780 , n8351 );
nand ( n8353 , n298775 , n298780 );
buf ( n8354 , n8353 );
buf ( n298783 , n8354 );
nand ( n298784 , n298774 , n298783 );
buf ( n298785 , n298784 );
xor ( n298786 , n298758 , n298785 );
or ( n298787 , n298731 , n298786 );
xor ( n8360 , n298665 , n298682 );
xor ( n298789 , n8360 , n298700 );
buf ( n298790 , n298789 );
nand ( n8363 , n298787 , n298790 );
nand ( n8364 , n298731 , n298786 );
nand ( n298793 , n8363 , n8364 );
nand ( n298794 , n298728 , n298793 );
nand ( n8367 , n298726 , n298794 );
nand ( n298796 , n795 , n800 );
buf ( n298797 , n794 );
buf ( n298798 , n800 );
xor ( n298799 , n298797 , n298798 );
buf ( n298800 , n298799 );
not ( n8373 , n298800 );
not ( n298802 , n296480 );
or ( n298803 , n8373 , n298802 );
buf ( n298804 , n6057 );
buf ( n298805 , n793 );
buf ( n298806 , n800 );
xor ( n8379 , n298805 , n298806 );
buf ( n8380 , n8379 );
buf ( n298809 , n8380 );
nand ( n8382 , n298804 , n298809 );
buf ( n298811 , n8382 );
nand ( n8384 , n298803 , n298811 );
xor ( n8385 , n298796 , n8384 );
xor ( n8386 , n826 , n768 );
not ( n298815 , n8386 );
not ( n8388 , n1453 );
or ( n8389 , n298815 , n8388 );
buf ( n298818 , n1580 );
buf ( n298819 , n826 );
nand ( n298820 , n298818 , n298819 );
buf ( n298821 , n298820 );
nand ( n8394 , n8389 , n298821 );
xnor ( n8395 , n8385 , n8394 );
xor ( n298824 , n828 , n768 );
buf ( n298825 , n298824 );
not ( n8398 , n298825 );
buf ( n298827 , n292168 );
not ( n8400 , n298827 );
or ( n298829 , n8398 , n8400 );
buf ( n298830 , n291812 );
buf ( n298831 , n828 );
nand ( n8404 , n298830 , n298831 );
buf ( n298833 , n8404 );
buf ( n298834 , n298833 );
nand ( n298835 , n298829 , n298834 );
buf ( n298836 , n298835 );
buf ( n298837 , n298836 );
buf ( n298838 , n8006 );
not ( n298839 , n298838 );
buf ( n298840 , n296480 );
not ( n8413 , n298840 );
or ( n298842 , n298839 , n8413 );
buf ( n298843 , n6057 );
buf ( n298844 , n298800 );
nand ( n8417 , n298843 , n298844 );
buf ( n298846 , n8417 );
buf ( n298847 , n298846 );
nand ( n298848 , n298842 , n298847 );
buf ( n298849 , n298848 );
buf ( n298850 , n298849 );
xor ( n298851 , n298837 , n298850 );
xor ( n298852 , n298735 , n298757 );
and ( n8425 , n298852 , n298785 );
and ( n298854 , n298735 , n298757 );
or ( n8427 , n8425 , n298854 );
buf ( n298856 , n8427 );
and ( n298857 , n298851 , n298856 );
and ( n8430 , n298837 , n298850 );
or ( n8431 , n298857 , n8430 );
buf ( n298860 , n8431 );
buf ( n298861 , n298860 );
not ( n8434 , n298861 );
buf ( n298863 , n8434 );
and ( n8436 , n8395 , n298863 );
not ( n8437 , n8395 );
and ( n8438 , n8437 , n298860 );
or ( n8439 , n8436 , n8438 );
not ( n298868 , n298707 );
not ( n8441 , n8220 );
and ( n8442 , n298868 , n8441 );
nand ( n8443 , n298707 , n8220 );
and ( n8444 , n298718 , n8443 );
nor ( n8445 , n8442 , n8444 );
and ( n8446 , n8439 , n8445 );
not ( n298875 , n8439 );
not ( n298876 , n8445 );
and ( n8449 , n298875 , n298876 );
or ( n298878 , n8446 , n8449 );
and ( n298879 , n8367 , n298878 );
not ( n8452 , n8367 );
not ( n298881 , n298878 );
and ( n8454 , n8452 , n298881 );
nor ( n8455 , n298879 , n8454 );
not ( n298884 , n293525 );
not ( n298885 , n291802 );
or ( n8458 , n298884 , n298885 );
nand ( n298887 , n8458 , n828 );
not ( n298888 , n8351 );
not ( n8461 , n4031 );
or ( n298890 , n298888 , n8461 );
xor ( n298891 , n772 , n822 );
nand ( n298892 , n292104 , n298891 );
nand ( n298893 , n298890 , n298892 );
xor ( n8466 , n298887 , n298893 );
not ( n298895 , n298751 );
not ( n298896 , n291880 );
or ( n8469 , n298895 , n298896 );
buf ( n298898 , n291886 );
buf ( n298899 , n8386 );
nand ( n8472 , n298898 , n298899 );
buf ( n298901 , n8472 );
nand ( n8474 , n8469 , n298901 );
xor ( n298903 , n8466 , n8474 );
buf ( n298904 , n298903 );
or ( n298905 , n8010 , n7965 );
nand ( n298906 , n298905 , n298411 );
nand ( n8479 , n7965 , n8010 );
nand ( n298908 , n298906 , n8479 );
buf ( n298909 , n298908 );
xor ( n8482 , n298904 , n298909 );
buf ( n298911 , n796 );
buf ( n298912 , n800 );
and ( n8485 , n298911 , n298912 );
buf ( n298914 , n8485 );
buf ( n298915 , n298914 );
buf ( n298916 , n298459 );
not ( n298917 , n298916 );
buf ( n298918 , n2373 );
not ( n298919 , n298918 );
or ( n8492 , n298917 , n298919 );
buf ( n298921 , n2026 );
buf ( n298922 , n782 );
buf ( n298923 , n812 );
xor ( n8496 , n298922 , n298923 );
buf ( n8497 , n8496 );
buf ( n8498 , n8497 );
nand ( n8499 , n298921 , n8498 );
buf ( n8500 , n8499 );
buf ( n298929 , n8500 );
nand ( n8502 , n8492 , n298929 );
buf ( n298931 , n8502 );
buf ( n8504 , n298931 );
xor ( n8505 , n298915 , n8504 );
buf ( n298934 , n298478 );
not ( n298935 , n298934 );
buf ( n298936 , n2893 );
not ( n298937 , n298936 );
or ( n8510 , n298935 , n298937 );
buf ( n298939 , n5051 );
buf ( n8512 , n780 );
buf ( n8513 , n814 );
xor ( n8514 , n8512 , n8513 );
buf ( n8515 , n8514 );
buf ( n298944 , n8515 );
nand ( n298945 , n298939 , n298944 );
buf ( n298946 , n298945 );
buf ( n298947 , n298946 );
nand ( n298948 , n8510 , n298947 );
buf ( n298949 , n298948 );
buf ( n298950 , n298949 );
xor ( n298951 , n8505 , n298950 );
buf ( n298952 , n298951 );
buf ( n298953 , n298952 );
and ( n8526 , n8482 , n298953 );
and ( n298955 , n298904 , n298909 );
or ( n298956 , n8526 , n298955 );
buf ( n298957 , n298956 );
buf ( n298958 , n298957 );
xor ( n8531 , n298887 , n298893 );
and ( n8532 , n8531 , n8474 );
and ( n298961 , n298887 , n298893 );
or ( n298962 , n8532 , n298961 );
buf ( n298963 , n298962 );
xor ( n8536 , n298915 , n8504 );
and ( n298965 , n8536 , n298950 );
and ( n298966 , n298915 , n8504 );
or ( n8539 , n298965 , n298966 );
buf ( n298968 , n8539 );
buf ( n298969 , n298968 );
xor ( n8542 , n298963 , n298969 );
buf ( n298971 , n298507 );
not ( n298972 , n298971 );
buf ( n298973 , n298099 );
not ( n298974 , n298973 );
or ( n298975 , n298972 , n298974 );
buf ( n298976 , n291969 );
buf ( n298977 , n774 );
buf ( n298978 , n820 );
xor ( n8551 , n298977 , n298978 );
buf ( n298980 , n8551 );
buf ( n298981 , n298980 );
nand ( n8554 , n298976 , n298981 );
buf ( n298983 , n8554 );
buf ( n298984 , n298983 );
nand ( n298985 , n298975 , n298984 );
buf ( n298986 , n298985 );
not ( n298987 , n298986 );
buf ( n298988 , n298636 );
not ( n8561 , n298988 );
nor ( n298990 , n4981 , n295410 );
buf ( n298991 , n298990 );
not ( n8564 , n298991 );
or ( n298993 , n8561 , n8564 );
buf ( n298994 , n6301 );
buf ( n298995 , n786 );
buf ( n298996 , n808 );
xor ( n8569 , n298995 , n298996 );
buf ( n298998 , n8569 );
buf ( n298999 , n298998 );
nand ( n8572 , n298994 , n298999 );
buf ( n299001 , n8572 );
buf ( n299002 , n299001 );
nand ( n299003 , n298993 , n299002 );
buf ( n299004 , n299003 );
not ( n8577 , n299004 );
or ( n8578 , n298987 , n8577 );
buf ( n299007 , n298986 );
buf ( n299008 , n299004 );
nor ( n8581 , n299007 , n299008 );
buf ( n299010 , n8581 );
buf ( n299011 , n298614 );
not ( n299012 , n299011 );
buf ( n299013 , n293058 );
not ( n299014 , n299013 );
or ( n8587 , n299012 , n299014 );
buf ( n299016 , n292841 );
buf ( n299017 , n784 );
buf ( n8590 , n810 );
xor ( n8591 , n299017 , n8590 );
buf ( n299020 , n8591 );
buf ( n299021 , n299020 );
nand ( n8594 , n299016 , n299021 );
buf ( n299023 , n8594 );
buf ( n299024 , n299023 );
nand ( n299025 , n8587 , n299024 );
buf ( n299026 , n299025 );
buf ( n299027 , n299026 );
not ( n299028 , n299027 );
buf ( n299029 , n299028 );
or ( n8602 , n299010 , n299029 );
nand ( n299031 , n8578 , n8602 );
buf ( n299032 , n299031 );
xor ( n8605 , n8542 , n299032 );
buf ( n299034 , n8605 );
buf ( n299035 , n299034 );
xor ( n299036 , n298958 , n299035 );
nand ( n299037 , n7960 , n7963 );
xor ( n8610 , n802 , n792 );
nand ( n299039 , n296517 , n8610 );
nand ( n299040 , n299037 , n299039 );
not ( n299041 , n299040 );
not ( n8614 , n298658 );
not ( n299043 , n298522 );
or ( n8616 , n8614 , n299043 );
buf ( n299045 , n298526 );
xor ( n299046 , n804 , n790 );
buf ( n8619 , n299046 );
nand ( n8620 , n299045 , n8619 );
buf ( n8621 , n8620 );
nand ( n299050 , n8616 , n8621 );
not ( n8623 , n299050 );
or ( n299052 , n299041 , n8623 );
nand ( n299053 , n299037 , n299039 );
or ( n8626 , n299053 , n299050 );
xor ( n299055 , n816 , n778 );
not ( n8628 , n299055 );
not ( n299057 , n296423 );
or ( n8630 , n8628 , n299057 );
nand ( n8631 , n7979 , n292892 );
nand ( n299060 , n8630 , n8631 );
nand ( n299061 , n8626 , n299060 );
nand ( n8634 , n299052 , n299061 );
buf ( n299063 , n8634 );
buf ( n299064 , n8247 );
not ( n8637 , n299064 );
buf ( n299066 , n295433 );
not ( n299067 , n299066 );
or ( n8640 , n8637 , n299067 );
xor ( n8641 , n806 , n788 );
not ( n8642 , n5680 );
nand ( n299071 , n8641 , n8642 );
buf ( n299072 , n299071 );
nand ( n8645 , n8640 , n299072 );
buf ( n299074 , n8645 );
buf ( n299075 , n299074 );
buf ( n299076 , n298693 );
not ( n8649 , n299076 );
buf ( n299078 , n291984 );
not ( n299079 , n299078 );
or ( n299080 , n8649 , n299079 );
buf ( n299081 , n295230 );
buf ( n299082 , n776 );
buf ( n299083 , n818 );
xor ( n8656 , n299082 , n299083 );
buf ( n8657 , n8656 );
buf ( n299086 , n8657 );
nand ( n299087 , n299081 , n299086 );
buf ( n299088 , n299087 );
buf ( n299089 , n299088 );
nand ( n299090 , n299080 , n299089 );
buf ( n299091 , n299090 );
buf ( n299092 , n299091 );
xor ( n299093 , n299075 , n299092 );
buf ( n299094 , n298595 );
not ( n8667 , n299094 );
buf ( n299096 , n291838 );
not ( n299097 , n299096 );
or ( n8670 , n8667 , n299097 );
buf ( n299099 , n1613 );
and ( n299100 , n770 , n824 );
not ( n8673 , n770 );
and ( n299102 , n8673 , n4959 );
nor ( n299103 , n299100 , n299102 );
buf ( n299104 , n299103 );
nand ( n299105 , n299099 , n299104 );
buf ( n299106 , n299105 );
buf ( n299107 , n299106 );
nand ( n8680 , n8670 , n299107 );
buf ( n299109 , n8680 );
buf ( n299110 , n299109 );
and ( n299111 , n299093 , n299110 );
and ( n8684 , n299075 , n299092 );
or ( n299113 , n299111 , n8684 );
buf ( n299114 , n299113 );
buf ( n299115 , n299114 );
xor ( n299116 , n299063 , n299115 );
not ( n299117 , n291842 );
buf ( n299118 , n769 );
buf ( n299119 , n824 );
xor ( n8692 , n299118 , n299119 );
buf ( n299121 , n8692 );
not ( n299122 , n299121 );
or ( n8695 , n299117 , n299122 );
nand ( n8696 , n299103 , n295562 , n5133 );
nand ( n8697 , n8695 , n8696 );
buf ( n299126 , n8697 );
buf ( n299127 , n8497 );
not ( n8700 , n299127 );
buf ( n299129 , n2373 );
not ( n299130 , n299129 );
or ( n8703 , n8700 , n299130 );
buf ( n299132 , n294479 );
buf ( n299133 , n781 );
buf ( n299134 , n812 );
xor ( n299135 , n299133 , n299134 );
buf ( n299136 , n299135 );
buf ( n299137 , n299136 );
nand ( n8710 , n299132 , n299137 );
buf ( n299139 , n8710 );
buf ( n299140 , n299139 );
nand ( n8713 , n8703 , n299140 );
buf ( n299142 , n8713 );
buf ( n299143 , n299142 );
xor ( n299144 , n299126 , n299143 );
buf ( n299145 , n298980 );
not ( n8718 , n299145 );
buf ( n299147 , n291722 );
not ( n8720 , n299147 );
or ( n8721 , n8718 , n8720 );
buf ( n299150 , n291969 );
buf ( n299151 , n773 );
buf ( n299152 , n820 );
xor ( n299153 , n299151 , n299152 );
buf ( n299154 , n299153 );
buf ( n299155 , n299154 );
nand ( n8728 , n299150 , n299155 );
buf ( n299157 , n8728 );
buf ( n299158 , n299157 );
nand ( n299159 , n8721 , n299158 );
buf ( n299160 , n299159 );
buf ( n299161 , n299160 );
xor ( n8734 , n299144 , n299161 );
buf ( n299163 , n8734 );
buf ( n299164 , n299163 );
xor ( n299165 , n299116 , n299164 );
buf ( n299166 , n299165 );
buf ( n299167 , n299166 );
xor ( n8740 , n299036 , n299167 );
buf ( n299169 , n8740 );
not ( n299170 , n299169 );
and ( n299171 , n8455 , n299170 );
not ( n8744 , n8455 );
and ( n299173 , n8744 , n299169 );
nor ( n299174 , n299171 , n299173 );
buf ( n299175 , n299174 );
xor ( n299176 , n298786 , n298731 );
xor ( n299177 , n299176 , n298790 );
not ( n8750 , n8016 );
not ( n8751 , n298579 );
not ( n8752 , n8751 );
or ( n299181 , n8750 , n8752 );
nand ( n299182 , n8015 , n298579 );
nand ( n8755 , n299181 , n299182 );
and ( n8756 , n8755 , n298516 );
not ( n8757 , n8755 );
not ( n8758 , n298516 );
and ( n299187 , n8757 , n8758 );
nor ( n299188 , n8756 , n299187 );
xor ( n8761 , n299177 , n299188 );
buf ( n299190 , n830 );
buf ( n299191 , n795 );
buf ( n299192 , n802 );
xor ( n8765 , n299191 , n299192 );
buf ( n299194 , n8765 );
buf ( n299195 , n299194 );
not ( n8768 , n299195 );
buf ( n299197 , n296508 );
not ( n299198 , n299197 );
or ( n8771 , n8768 , n299198 );
buf ( n299200 , n296749 );
buf ( n299201 , n7955 );
nand ( n8774 , n299200 , n299201 );
buf ( n299203 , n8774 );
buf ( n299204 , n299203 );
nand ( n299205 , n8771 , n299204 );
buf ( n299206 , n299205 );
buf ( n299207 , n299206 );
xor ( n8780 , n299190 , n299207 );
buf ( n299209 , n799 );
buf ( n299210 , n800 );
and ( n299211 , n299209 , n299210 );
buf ( n299212 , n299211 );
buf ( n299213 , n299212 );
buf ( n299214 , n768 );
buf ( n299215 , n830 );
xor ( n299216 , n299214 , n299215 );
buf ( n299217 , n299216 );
buf ( n299218 , n299217 );
not ( n299219 , n299218 );
buf ( n299220 , n1271 );
not ( n8793 , n299220 );
or ( n299222 , n299219 , n8793 );
buf ( n299223 , n830 );
buf ( n299224 , n831 );
nand ( n299225 , n299223 , n299224 );
buf ( n299226 , n299225 );
buf ( n299227 , n299226 );
nand ( n8800 , n299222 , n299227 );
buf ( n299229 , n8800 );
buf ( n299230 , n299229 );
xor ( n299231 , n299213 , n299230 );
buf ( n299232 , n770 );
buf ( n299233 , n828 );
xor ( n299234 , n299232 , n299233 );
buf ( n299235 , n299234 );
buf ( n8808 , n299235 );
not ( n8809 , n8808 );
buf ( n299238 , n292168 );
not ( n299239 , n299238 );
or ( n8812 , n8809 , n299239 );
buf ( n299241 , n291812 );
buf ( n299242 , n769 );
not ( n8815 , n299242 );
buf ( n299244 , n8815 );
and ( n299245 , n828 , n299244 );
not ( n8818 , n828 );
and ( n299247 , n8818 , n769 );
or ( n8820 , n299245 , n299247 );
buf ( n299249 , n8820 );
nand ( n8822 , n299241 , n299249 );
buf ( n299251 , n8822 );
buf ( n299252 , n299251 );
nand ( n8825 , n8812 , n299252 );
buf ( n299254 , n8825 );
buf ( n299255 , n299254 );
and ( n299256 , n299231 , n299255 );
and ( n299257 , n299213 , n299230 );
or ( n8830 , n299256 , n299257 );
buf ( n299259 , n8830 );
buf ( n299260 , n299259 );
xor ( n8833 , n8780 , n299260 );
buf ( n299262 , n8833 );
buf ( n299263 , n299262 );
buf ( n8836 , n292104 );
xor ( n299265 , n822 , n775 );
buf ( n299266 , n299265 );
nand ( n299267 , n8836 , n299266 );
buf ( n299268 , n299267 );
xor ( n8841 , n822 , n776 );
nand ( n299270 , n8841 , n1338 , n291757 );
and ( n299271 , n299268 , n299270 );
buf ( n299272 , n784 );
buf ( n299273 , n814 );
xor ( n299274 , n299272 , n299273 );
buf ( n299275 , n299274 );
not ( n299276 , n299275 );
buf ( n299277 , n814 );
buf ( n299278 , n815 );
xnor ( n299279 , n299277 , n299278 );
buf ( n299280 , n299279 );
nor ( n8853 , n299280 , n292502 );
not ( n299282 , n8853 );
or ( n8855 , n299276 , n299282 );
buf ( n299284 , n783 );
buf ( n299285 , n814 );
xor ( n299286 , n299284 , n299285 );
buf ( n299287 , n299286 );
nand ( n8860 , n5051 , n299287 );
nand ( n299289 , n8855 , n8860 );
nand ( n8862 , n299271 , n299289 );
not ( n299291 , n8862 );
not ( n8864 , n299271 );
not ( n299293 , n299289 );
nand ( n8866 , n8864 , n299293 );
not ( n8867 , n8866 );
or ( n299296 , n299291 , n8867 );
xor ( n8869 , n812 , n786 );
buf ( n299298 , n8869 );
not ( n299299 , n299298 );
buf ( n299300 , n2373 );
not ( n299301 , n299300 );
or ( n8874 , n299299 , n299301 );
buf ( n299303 , n294479 );
xor ( n299304 , n812 , n785 );
buf ( n299305 , n299304 );
nand ( n8878 , n299303 , n299305 );
buf ( n299307 , n8878 );
buf ( n299308 , n299307 );
nand ( n299309 , n8874 , n299308 );
buf ( n299310 , n299309 );
buf ( n299311 , n299310 );
not ( n8884 , n299311 );
buf ( n299313 , n8884 );
not ( n299314 , n299313 );
nand ( n8887 , n299296 , n299314 );
nand ( n299316 , n8866 , n8862 , n299313 );
nand ( n299317 , n8887 , n299316 );
buf ( n299318 , n299317 );
not ( n299319 , n299318 );
buf ( n299320 , n299319 );
buf ( n299321 , n299320 );
not ( n299322 , n299321 );
buf ( n299323 , n790 );
buf ( n299324 , n808 );
xor ( n299325 , n299323 , n299324 );
buf ( n299326 , n299325 );
buf ( n299327 , n299326 );
not ( n8900 , n299327 );
buf ( n299329 , n3408 );
not ( n299330 , n299329 );
or ( n299331 , n8900 , n299330 );
buf ( n8904 , n3114 );
buf ( n299333 , n789 );
buf ( n299334 , n808 );
xor ( n299335 , n299333 , n299334 );
buf ( n299336 , n299335 );
buf ( n299337 , n299336 );
nand ( n8910 , n8904 , n299337 );
buf ( n299339 , n8910 );
buf ( n299340 , n299339 );
nand ( n8913 , n299331 , n299340 );
buf ( n299342 , n8913 );
buf ( n299343 , n299342 );
buf ( n299344 , n792 );
buf ( n299345 , n806 );
xor ( n299346 , n299344 , n299345 );
buf ( n299347 , n299346 );
buf ( n299348 , n299347 );
not ( n299349 , n299348 );
buf ( n299350 , n294637 );
not ( n8923 , n299350 );
or ( n299352 , n299349 , n8923 );
buf ( n299353 , n293902 );
buf ( n299354 , n298561 );
nand ( n299355 , n299353 , n299354 );
buf ( n299356 , n299355 );
buf ( n299357 , n299356 );
nand ( n299358 , n299352 , n299357 );
buf ( n299359 , n299358 );
buf ( n299360 , n299359 );
xor ( n299361 , n299343 , n299360 );
buf ( n8934 , n780 );
buf ( n299363 , n818 );
xor ( n299364 , n8934 , n299363 );
buf ( n299365 , n299364 );
buf ( n299366 , n299365 );
not ( n8939 , n299366 );
buf ( n299368 , n1962 );
not ( n299369 , n299368 );
or ( n299370 , n8939 , n299369 );
buf ( n299371 , n295230 );
buf ( n299372 , n298542 );
nand ( n299373 , n299371 , n299372 );
buf ( n299374 , n299373 );
buf ( n299375 , n299374 );
nand ( n299376 , n299370 , n299375 );
buf ( n299377 , n299376 );
buf ( n299378 , n299377 );
xor ( n8951 , n299361 , n299378 );
buf ( n299380 , n8951 );
buf ( n299381 , n299380 );
not ( n8954 , n299381 );
or ( n299383 , n299322 , n8954 );
buf ( n299384 , n299320 );
buf ( n299385 , n299380 );
or ( n8958 , n299384 , n299385 );
buf ( n299387 , n778 );
buf ( n299388 , n820 );
xor ( n8961 , n299387 , n299388 );
buf ( n299390 , n8961 );
not ( n8963 , n299390 );
not ( n299392 , n292668 );
or ( n299393 , n8963 , n299392 );
buf ( n299394 , n777 );
buf ( n299395 , n820 );
xor ( n8968 , n299394 , n299395 );
buf ( n299397 , n8968 );
buf ( n299398 , n299397 );
buf ( n299399 , n1995 );
nand ( n8972 , n299398 , n299399 );
buf ( n299401 , n8972 );
nand ( n299402 , n299393 , n299401 );
buf ( n299403 , n772 );
buf ( n299404 , n826 );
xor ( n8977 , n299403 , n299404 );
buf ( n299406 , n8977 );
buf ( n299407 , n299406 );
not ( n8980 , n299407 );
buf ( n299409 , n291880 );
not ( n8982 , n299409 );
or ( n299411 , n8980 , n8982 );
buf ( n299412 , n1579 );
buf ( n299413 , n771 );
buf ( n299414 , n826 );
xor ( n8987 , n299413 , n299414 );
buf ( n299416 , n8987 );
buf ( n8989 , n299416 );
nand ( n8990 , n299412 , n8989 );
buf ( n8991 , n8990 );
buf ( n299420 , n8991 );
nand ( n8993 , n299411 , n299420 );
buf ( n299422 , n8993 );
xor ( n299423 , n299402 , n299422 );
buf ( n8996 , n788 );
buf ( n299425 , n810 );
xor ( n8998 , n8996 , n299425 );
buf ( n299427 , n8998 );
buf ( n299428 , n299427 );
not ( n299429 , n299428 );
buf ( n299430 , n293058 );
not ( n299431 , n299430 );
or ( n9004 , n299429 , n299431 );
buf ( n299433 , n292841 );
buf ( n9006 , n787 );
buf ( n299435 , n810 );
xor ( n299436 , n9006 , n299435 );
buf ( n299437 , n299436 );
buf ( n299438 , n299437 );
nand ( n299439 , n299433 , n299438 );
buf ( n299440 , n299439 );
buf ( n299441 , n299440 );
nand ( n9014 , n9004 , n299441 );
buf ( n299443 , n9014 );
xor ( n299444 , n299423 , n299443 );
buf ( n299445 , n299444 );
nand ( n9018 , n8958 , n299445 );
buf ( n9019 , n9018 );
buf ( n9020 , n9019 );
nand ( n9021 , n299383 , n9020 );
buf ( n9022 , n9021 );
buf ( n9023 , n9022 );
xor ( n9024 , n299263 , n9023 );
or ( n299453 , n8864 , n299310 );
nand ( n299454 , n299453 , n299289 );
buf ( n299455 , n299454 );
nand ( n299456 , n299310 , n8864 );
buf ( n299457 , n299456 );
nand ( n9030 , n299455 , n299457 );
buf ( n299459 , n9030 );
buf ( n299460 , n299459 );
xor ( n9033 , n299343 , n299360 );
and ( n299462 , n9033 , n299378 );
and ( n299463 , n299343 , n299360 );
or ( n9036 , n299462 , n299463 );
buf ( n299465 , n9036 );
buf ( n299466 , n299465 );
xor ( n9039 , n299460 , n299466 );
buf ( n299468 , n798 );
buf ( n299469 , n800 );
xor ( n9042 , n299468 , n299469 );
buf ( n299471 , n9042 );
buf ( n299472 , n299471 );
not ( n299473 , n299472 );
buf ( n299474 , n6049 );
not ( n299475 , n299474 );
or ( n299476 , n299473 , n299475 );
buf ( n299477 , n6057 );
xor ( n299478 , n800 , n797 );
buf ( n299479 , n299478 );
nand ( n9052 , n299477 , n299479 );
buf ( n299481 , n9052 );
buf ( n299482 , n299481 );
nand ( n9055 , n299476 , n299482 );
buf ( n299484 , n9055 );
buf ( n299485 , n299484 );
buf ( n299486 , n774 );
buf ( n299487 , n824 );
xor ( n299488 , n299486 , n299487 );
buf ( n299489 , n299488 );
buf ( n299490 , n299489 );
not ( n299491 , n299490 );
buf ( n299492 , n291838 );
not ( n299493 , n299492 );
or ( n9066 , n299491 , n299493 );
buf ( n299495 , n1613 );
buf ( n299496 , n773 );
buf ( n299497 , n824 );
xor ( n299498 , n299496 , n299497 );
buf ( n299499 , n299498 );
buf ( n299500 , n299499 );
nand ( n299501 , n299495 , n299500 );
buf ( n299502 , n299501 );
buf ( n299503 , n299502 );
nand ( n299504 , n9066 , n299503 );
buf ( n299505 , n299504 );
buf ( n299506 , n299505 );
xor ( n299507 , n299485 , n299506 );
buf ( n299508 , n782 );
buf ( n299509 , n816 );
xor ( n299510 , n299508 , n299509 );
buf ( n299511 , n299510 );
buf ( n299512 , n299511 );
not ( n9085 , n299512 );
buf ( n299514 , n2118 );
not ( n299515 , n299514 );
or ( n299516 , n9085 , n299515 );
buf ( n299517 , n296423 );
xor ( n9090 , n816 , n781 );
buf ( n299519 , n9090 );
nand ( n299520 , n299517 , n299519 );
buf ( n299521 , n299520 );
buf ( n299522 , n299521 );
nand ( n299523 , n299516 , n299522 );
buf ( n299524 , n299523 );
buf ( n299525 , n299524 );
and ( n299526 , n299507 , n299525 );
and ( n299527 , n299485 , n299506 );
or ( n9100 , n299526 , n299527 );
buf ( n299529 , n9100 );
buf ( n299530 , n299529 );
xor ( n299531 , n9039 , n299530 );
buf ( n299532 , n299531 );
buf ( n299533 , n299532 );
and ( n9106 , n9024 , n299533 );
and ( n9107 , n299263 , n9023 );
or ( n299536 , n9106 , n9107 );
buf ( n299537 , n299536 );
and ( n9110 , n8761 , n299537 );
and ( n9111 , n299177 , n299188 );
or ( n9112 , n9110 , n9111 );
xor ( n299541 , n298904 , n298909 );
xor ( n299542 , n299541 , n298953 );
buf ( n299543 , n299542 );
buf ( n299544 , n299543 );
not ( n9117 , n299053 );
and ( n299546 , n299050 , n9117 );
not ( n299547 , n299050 );
and ( n9120 , n299547 , n299040 );
nor ( n9121 , n299546 , n9120 );
not ( n9122 , n299060 );
xor ( n299551 , n9121 , n9122 );
buf ( n299552 , n299551 );
xor ( n9125 , n299075 , n299092 );
xor ( n9126 , n9125 , n299110 );
buf ( n299555 , n9126 );
buf ( n299556 , n299555 );
xor ( n299557 , n299552 , n299556 );
xor ( n9130 , n298986 , n299004 );
buf ( n299559 , n9130 );
buf ( n299560 , n299026 );
and ( n299561 , n299559 , n299560 );
not ( n299562 , n299559 );
buf ( n299563 , n299029 );
and ( n299564 , n299562 , n299563 );
nor ( n299565 , n299561 , n299564 );
buf ( n299566 , n299565 );
buf ( n299567 , n299566 );
xor ( n299568 , n299557 , n299567 );
buf ( n299569 , n299568 );
buf ( n299570 , n299569 );
xor ( n299571 , n299544 , n299570 );
buf ( n299572 , n292367 );
buf ( n9145 , n298836 );
not ( n9146 , n9145 );
buf ( n299575 , n9146 );
buf ( n299576 , n299575 );
xor ( n299577 , n299572 , n299576 );
buf ( n9150 , n798 );
buf ( n9151 , n800 );
and ( n9152 , n9150 , n9151 );
buf ( n9153 , n9152 );
buf ( n299582 , n9153 );
buf ( n299583 , n299478 );
not ( n299584 , n299583 );
buf ( n299585 , n296475 );
not ( n9158 , n299585 );
buf ( n299587 , n296469 );
nor ( n299588 , n9158 , n299587 );
buf ( n299589 , n299588 );
buf ( n299590 , n299589 );
not ( n299591 , n299590 );
or ( n9164 , n299584 , n299591 );
nand ( n299593 , n6056 , n7999 );
buf ( n299594 , n299593 );
nand ( n9167 , n9164 , n299594 );
buf ( n299596 , n9167 );
buf ( n299597 , n299596 );
xor ( n9170 , n299582 , n299597 );
buf ( n299599 , n9090 );
not ( n9172 , n299599 );
buf ( n299601 , n2118 );
not ( n299602 , n299601 );
or ( n299603 , n9172 , n299602 );
buf ( n299604 , n1712 );
buf ( n299605 , n7970 );
nand ( n299606 , n299604 , n299605 );
buf ( n299607 , n299606 );
buf ( n299608 , n299607 );
nand ( n9181 , n299603 , n299608 );
buf ( n9182 , n9181 );
buf ( n299611 , n9182 );
and ( n9184 , n9170 , n299611 );
and ( n299613 , n299582 , n299597 );
or ( n299614 , n9184 , n299613 );
buf ( n299615 , n299614 );
buf ( n299616 , n299615 );
and ( n299617 , n299577 , n299616 );
and ( n299618 , n299572 , n299576 );
or ( n9191 , n299617 , n299618 );
buf ( n299620 , n9191 );
buf ( n299621 , n299620 );
xor ( n9194 , n298837 , n298850 );
xor ( n299623 , n9194 , n298856 );
buf ( n299624 , n299623 );
buf ( n299625 , n299624 );
xor ( n299626 , n299621 , n299625 );
buf ( n299627 , n299499 );
not ( n9200 , n299627 );
buf ( n299629 , n292473 );
not ( n299630 , n299629 );
or ( n9203 , n9200 , n299630 );
buf ( n299632 , n1613 );
buf ( n299633 , n298587 );
nand ( n9206 , n299632 , n299633 );
buf ( n9207 , n9206 );
buf ( n299636 , n9207 );
nand ( n299637 , n9203 , n299636 );
buf ( n299638 , n299637 );
not ( n299639 , n299638 );
buf ( n299640 , n8820 );
not ( n9213 , n299640 );
buf ( n299642 , n294329 );
not ( n299643 , n299642 );
or ( n9216 , n9213 , n299643 );
buf ( n299645 , n1508 );
buf ( n299646 , n298824 );
nand ( n9219 , n299645 , n299646 );
buf ( n9220 , n9219 );
buf ( n299649 , n9220 );
nand ( n9222 , n9216 , n299649 );
buf ( n299651 , n9222 );
not ( n9224 , n299651 );
or ( n9225 , n299639 , n9224 );
buf ( n9226 , n299638 );
buf ( n9227 , n299651 );
nor ( n9228 , n9226 , n9227 );
buf ( n9229 , n9228 );
buf ( n299658 , n299287 );
not ( n9231 , n299658 );
buf ( n299660 , n2078 );
not ( n9233 , n299660 );
or ( n299662 , n9231 , n9233 );
buf ( n299663 , n2089 );
buf ( n299664 , n8040 );
nand ( n9237 , n299663 , n299664 );
buf ( n299666 , n9237 );
buf ( n299667 , n299666 );
nand ( n9240 , n299662 , n299667 );
buf ( n299669 , n9240 );
not ( n9242 , n299669 );
or ( n299671 , n9229 , n9242 );
nand ( n299672 , n9225 , n299671 );
buf ( n299673 , n299397 );
not ( n9246 , n299673 );
buf ( n299675 , n2787 );
not ( n299676 , n299675 );
or ( n299677 , n9246 , n299676 );
nand ( n9250 , n291734 , n8069 );
buf ( n299679 , n9250 );
nand ( n9252 , n299677 , n299679 );
buf ( n299681 , n9252 );
buf ( n299682 , n299681 );
buf ( n299683 , n299416 );
not ( n9256 , n299683 );
buf ( n299685 , n291880 );
not ( n299686 , n299685 );
or ( n9259 , n9256 , n299686 );
buf ( n299688 , n293402 );
buf ( n299689 , n298739 );
nand ( n9262 , n299688 , n299689 );
buf ( n299691 , n9262 );
buf ( n299692 , n299691 );
nand ( n299693 , n9259 , n299692 );
buf ( n299694 , n299693 );
buf ( n299695 , n299694 );
xor ( n299696 , n299682 , n299695 );
not ( n299697 , n299336 );
not ( n299698 , n293655 );
or ( n299699 , n299697 , n299698 );
nand ( n9272 , n294557 , n298626 );
nand ( n299701 , n299699 , n9272 );
buf ( n299702 , n299701 );
and ( n9275 , n299696 , n299702 );
and ( n299704 , n299682 , n299695 );
or ( n9277 , n9275 , n299704 );
buf ( n299706 , n9277 );
xor ( n299707 , n299672 , n299706 );
buf ( n299708 , n299265 );
not ( n9281 , n299708 );
buf ( n299710 , n298771 );
not ( n299711 , n299710 );
or ( n9284 , n9281 , n299711 );
buf ( n299713 , n292104 );
buf ( n299714 , n298762 );
nand ( n299715 , n299713 , n299714 );
buf ( n299716 , n299715 );
buf ( n299717 , n299716 );
nand ( n299718 , n9284 , n299717 );
buf ( n299719 , n299718 );
buf ( n9292 , n299719 );
not ( n299721 , n9292 );
buf ( n299722 , n299721 );
buf ( n299723 , n299722 );
not ( n299724 , n299723 );
buf ( n299725 , n299304 );
not ( n299726 , n299725 );
buf ( n299727 , n2373 );
not ( n9300 , n299727 );
or ( n299729 , n299726 , n9300 );
buf ( n299730 , n294479 );
buf ( n299731 , n298449 );
nand ( n299732 , n299730 , n299731 );
buf ( n299733 , n299732 );
buf ( n299734 , n299733 );
nand ( n299735 , n299729 , n299734 );
buf ( n299736 , n299735 );
buf ( n299737 , n299736 );
not ( n9310 , n299737 );
buf ( n299739 , n9310 );
buf ( n299740 , n299739 );
not ( n299741 , n299740 );
or ( n9314 , n299724 , n299741 );
buf ( n299743 , n299437 );
not ( n299744 , n299743 );
buf ( n299745 , n293058 );
not ( n9318 , n299745 );
or ( n299747 , n299744 , n9318 );
buf ( n299748 , n295259 );
buf ( n299749 , n8176 );
nand ( n299750 , n299748 , n299749 );
buf ( n299751 , n299750 );
buf ( n299752 , n299751 );
nand ( n9325 , n299747 , n299752 );
buf ( n299754 , n9325 );
buf ( n299755 , n299754 );
nand ( n299756 , n9314 , n299755 );
buf ( n299757 , n299756 );
buf ( n299758 , n299736 );
buf ( n299759 , n299719 );
nand ( n299760 , n299758 , n299759 );
buf ( n299761 , n299760 );
nand ( n9334 , n299757 , n299761 );
and ( n299763 , n299707 , n9334 );
and ( n299764 , n299672 , n299706 );
or ( n9337 , n299763 , n299764 );
buf ( n299766 , n9337 );
xor ( n299767 , n299626 , n299766 );
buf ( n299768 , n299767 );
buf ( n299769 , n299768 );
xor ( n9342 , n299571 , n299769 );
buf ( n299771 , n9342 );
xor ( n299772 , n9112 , n299771 );
xor ( n299773 , n299190 , n299207 );
and ( n9346 , n299773 , n299260 );
and ( n9347 , n299190 , n299207 );
or ( n9348 , n9346 , n9347 );
buf ( n299777 , n9348 );
xor ( n299778 , n299460 , n299466 );
and ( n9351 , n299778 , n299530 );
and ( n9352 , n299460 , n299466 );
or ( n9353 , n9351 , n9352 );
buf ( n9354 , n9353 );
xor ( n299783 , n299777 , n9354 );
xor ( n9356 , n299672 , n299706 );
xor ( n9357 , n9356 , n9334 );
xor ( n9358 , n299783 , n9357 );
xor ( n299787 , n299572 , n299576 );
xor ( n299788 , n299787 , n299616 );
buf ( n299789 , n299788 );
buf ( n299790 , n299651 );
not ( n9363 , n299790 );
not ( n299792 , n299669 );
buf ( n299793 , n299792 );
not ( n9366 , n299793 );
or ( n299795 , n9363 , n9366 );
buf ( n299796 , n299651 );
not ( n299797 , n299796 );
buf ( n299798 , n299669 );
nand ( n299799 , n299797 , n299798 );
buf ( n299800 , n299799 );
buf ( n299801 , n299800 );
nand ( n9374 , n299795 , n299801 );
buf ( n299803 , n9374 );
buf ( n299804 , n299638 );
not ( n299805 , n299804 );
buf ( n299806 , n299805 );
and ( n299807 , n299803 , n299806 );
not ( n299808 , n299803 );
buf ( n299809 , n299638 );
and ( n299810 , n299808 , n299809 );
nor ( n9383 , n299807 , n299810 );
not ( n299812 , n9383 );
not ( n299813 , n299812 );
xor ( n9386 , n299722 , n299736 );
xor ( n299815 , n9386 , n299754 );
buf ( n299816 , n299815 );
not ( n9389 , n299816 );
buf ( n299818 , n9389 );
not ( n299819 , n299818 );
or ( n9392 , n299813 , n299819 );
not ( n299821 , n299815 );
not ( n299822 , n9383 );
or ( n9395 , n299821 , n299822 );
xor ( n299824 , n299682 , n299695 );
xor ( n299825 , n299824 , n299702 );
buf ( n299826 , n299825 );
nand ( n299827 , n9395 , n299826 );
nand ( n9400 , n9392 , n299827 );
xor ( n299829 , n299789 , n9400 );
not ( n9402 , n299443 );
buf ( n299831 , n299402 );
not ( n299832 , n299831 );
or ( n299833 , n9402 , n299832 );
or ( n299834 , n299831 , n299443 );
nand ( n9407 , n299834 , n299422 );
nand ( n299836 , n299833 , n9407 );
buf ( n299837 , n299836 );
xor ( n299838 , n299582 , n299597 );
xor ( n9411 , n299838 , n299611 );
buf ( n299840 , n9411 );
buf ( n299841 , n299840 );
xor ( n9414 , n299837 , n299841 );
xor ( n299843 , n298538 , n298556 );
xor ( n299844 , n299843 , n298575 );
buf ( n299845 , n299844 );
buf ( n299846 , n299845 );
and ( n299847 , n9414 , n299846 );
and ( n9420 , n299837 , n299841 );
or ( n299849 , n299847 , n9420 );
buf ( n299850 , n299849 );
xor ( n9423 , n299829 , n299850 );
nand ( n299852 , n9358 , n9423 );
or ( n299853 , n9358 , n9423 );
not ( n9426 , n7960 );
buf ( n299855 , n796 );
buf ( n299856 , n802 );
xor ( n9429 , n299855 , n299856 );
buf ( n299858 , n9429 );
not ( n299859 , n299858 );
or ( n9432 , n9426 , n299859 );
buf ( n299861 , n296517 );
buf ( n299862 , n299194 );
nand ( n9435 , n299861 , n299862 );
buf ( n9436 , n9435 );
nand ( n299865 , n9432 , n9436 );
buf ( n299866 , n299865 );
buf ( n299867 , n794 );
buf ( n299868 , n804 );
xor ( n9441 , n299867 , n299868 );
buf ( n299870 , n9441 );
buf ( n299871 , n299870 );
not ( n299872 , n299871 );
buf ( n299873 , n6010 );
not ( n299874 , n299873 );
or ( n299875 , n299872 , n299874 );
buf ( n299876 , n296663 );
buf ( n299877 , n298519 );
nand ( n9450 , n299876 , n299877 );
buf ( n299879 , n9450 );
buf ( n299880 , n299879 );
nand ( n9453 , n299875 , n299880 );
buf ( n9454 , n9453 );
buf ( n299883 , n9454 );
xor ( n9456 , n299866 , n299883 );
buf ( n299885 , n799 );
buf ( n299886 , n801 );
or ( n299887 , n299885 , n299886 );
buf ( n299888 , n802 );
nand ( n299889 , n299887 , n299888 );
buf ( n299890 , n299889 );
buf ( n299891 , n299890 );
buf ( n299892 , n799 );
buf ( n299893 , n801 );
nand ( n9466 , n299892 , n299893 );
buf ( n9467 , n9466 );
buf ( n299896 , n9467 );
buf ( n299897 , n800 );
and ( n9470 , n299891 , n299896 , n299897 );
buf ( n299899 , n9470 );
buf ( n299900 , n299899 );
buf ( n299901 , n769 );
buf ( n9474 , n830 );
xor ( n9475 , n299901 , n9474 );
buf ( n9476 , n9475 );
buf ( n299905 , n9476 );
not ( n9478 , n299905 );
buf ( n299907 , n1271 );
not ( n299908 , n299907 );
or ( n9481 , n9478 , n299908 );
buf ( n299910 , n299217 );
buf ( n299911 , n831 );
nand ( n299912 , n299910 , n299911 );
buf ( n299913 , n299912 );
buf ( n299914 , n299913 );
nand ( n9487 , n9481 , n299914 );
buf ( n299916 , n9487 );
buf ( n299917 , n299916 );
and ( n299918 , n299900 , n299917 );
buf ( n299919 , n299918 );
buf ( n299920 , n299919 );
and ( n299921 , n9456 , n299920 );
and ( n9494 , n299866 , n299883 );
or ( n9495 , n299921 , n9494 );
buf ( n299924 , n9495 );
buf ( n299925 , n299924 );
buf ( n299926 , n791 );
buf ( n299927 , n808 );
xor ( n9500 , n299926 , n299927 );
buf ( n299929 , n9500 );
not ( n299930 , n299929 );
not ( n299931 , n4983 );
or ( n9504 , n299930 , n299931 );
buf ( n299933 , n3114 );
buf ( n299934 , n299326 );
nand ( n299935 , n299933 , n299934 );
buf ( n299936 , n299935 );
nand ( n9509 , n9504 , n299936 );
not ( n299938 , n9509 );
buf ( n9511 , n793 );
buf ( n299940 , n806 );
xor ( n299941 , n9511 , n299940 );
buf ( n299942 , n299941 );
buf ( n299943 , n299942 );
not ( n299944 , n299943 );
buf ( n299945 , n295433 );
not ( n9518 , n299945 );
or ( n299947 , n299944 , n9518 );
buf ( n299948 , n293902 );
buf ( n299949 , n299347 );
nand ( n9522 , n299948 , n299949 );
buf ( n299951 , n9522 );
buf ( n299952 , n299951 );
nand ( n299953 , n299947 , n299952 );
buf ( n299954 , n299953 );
not ( n9527 , n299954 );
or ( n299956 , n299938 , n9527 );
or ( n9529 , n299954 , n9509 );
xor ( n299958 , n820 , n779 );
not ( n299959 , n299958 );
not ( n9532 , n2787 );
or ( n9533 , n299959 , n9532 );
buf ( n299962 , n291969 );
buf ( n299963 , n299390 );
nand ( n9536 , n299962 , n299963 );
buf ( n9537 , n9536 );
nand ( n299966 , n9533 , n9537 );
nand ( n299967 , n9529 , n299966 );
nand ( n9540 , n299956 , n299967 );
xor ( n9541 , n299213 , n299230 );
xor ( n299970 , n9541 , n299255 );
buf ( n299971 , n299970 );
xor ( n299972 , n9540 , n299971 );
buf ( n299973 , n781 );
buf ( n299974 , n818 );
xor ( n299975 , n299973 , n299974 );
buf ( n299976 , n299975 );
buf ( n299977 , n299976 );
not ( n299978 , n299977 );
buf ( n299979 , n1553 );
not ( n9552 , n299979 );
or ( n299981 , n299978 , n9552 );
buf ( n299982 , n1357 );
buf ( n299983 , n299365 );
nand ( n299984 , n299982 , n299983 );
buf ( n299985 , n299984 );
buf ( n299986 , n299985 );
nand ( n299987 , n299981 , n299986 );
buf ( n299988 , n299987 );
buf ( n299989 , n299988 );
buf ( n299990 , n795 );
buf ( n299991 , n804 );
xor ( n299992 , n299990 , n299991 );
buf ( n299993 , n299992 );
buf ( n299994 , n299993 );
not ( n299995 , n299994 );
buf ( n299996 , n295983 );
not ( n9569 , n299996 );
or ( n299998 , n299995 , n9569 );
buf ( n299999 , n298526 );
buf ( n300000 , n299870 );
nand ( n300001 , n299999 , n300000 );
buf ( n300002 , n300001 );
buf ( n300003 , n300002 );
nand ( n300004 , n299998 , n300003 );
buf ( n300005 , n300004 );
buf ( n300006 , n300005 );
xor ( n300007 , n299989 , n300006 );
buf ( n300008 , n797 );
buf ( n300009 , n802 );
xor ( n300010 , n300008 , n300009 );
buf ( n300011 , n300010 );
buf ( n300012 , n300011 );
not ( n300013 , n300012 );
buf ( n300014 , n7960 );
not ( n9587 , n300014 );
or ( n300016 , n300013 , n9587 );
buf ( n300017 , n296517 );
buf ( n300018 , n299858 );
nand ( n300019 , n300017 , n300018 );
buf ( n300020 , n300019 );
buf ( n300021 , n300020 );
nand ( n300022 , n300016 , n300021 );
buf ( n300023 , n300022 );
buf ( n300024 , n300023 );
and ( n300025 , n300007 , n300024 );
and ( n9598 , n299989 , n300006 );
or ( n300027 , n300025 , n9598 );
buf ( n300028 , n300027 );
and ( n9601 , n299972 , n300028 );
and ( n300030 , n9540 , n299971 );
or ( n300031 , n9601 , n300030 );
buf ( n300032 , n300031 );
xor ( n9605 , n299925 , n300032 );
buf ( n9606 , n773 );
buf ( n9607 , n826 );
xor ( n9608 , n9606 , n9607 );
buf ( n9609 , n9608 );
buf ( n300038 , n9609 );
not ( n9611 , n300038 );
buf ( n300040 , n291880 );
not ( n9613 , n300040 );
or ( n300042 , n9611 , n9613 );
buf ( n300043 , n293402 );
buf ( n300044 , n299406 );
nand ( n9617 , n300043 , n300044 );
buf ( n300046 , n9617 );
buf ( n300047 , n300046 );
nand ( n300048 , n300042 , n300047 );
buf ( n300049 , n300048 );
buf ( n300050 , n787 );
buf ( n300051 , n812 );
xor ( n300052 , n300050 , n300051 );
buf ( n300053 , n300052 );
buf ( n300054 , n300053 );
not ( n300055 , n300054 );
buf ( n300056 , n2373 );
not ( n9629 , n300056 );
or ( n300058 , n300055 , n9629 );
buf ( n9631 , n294479 );
buf ( n300060 , n8869 );
nand ( n300061 , n9631 , n300060 );
buf ( n300062 , n300061 );
buf ( n300063 , n300062 );
nand ( n300064 , n300058 , n300063 );
buf ( n300065 , n300064 );
or ( n9638 , n300049 , n300065 );
buf ( n300067 , n789 );
buf ( n300068 , n810 );
xor ( n9641 , n300067 , n300068 );
buf ( n9642 , n9641 );
buf ( n300071 , n9642 );
not ( n300072 , n300071 );
buf ( n300073 , n293055 );
not ( n300074 , n300073 );
or ( n300075 , n300072 , n300074 );
buf ( n300076 , n295259 );
buf ( n300077 , n299427 );
nand ( n300078 , n300076 , n300077 );
buf ( n300079 , n300078 );
buf ( n300080 , n300079 );
nand ( n300081 , n300075 , n300080 );
buf ( n300082 , n300081 );
nand ( n300083 , n9638 , n300082 );
buf ( n300084 , n300049 );
buf ( n300085 , n300065 );
nand ( n300086 , n300084 , n300085 );
buf ( n300087 , n300086 );
nand ( n9660 , n300083 , n300087 );
buf ( n9661 , n9660 );
buf ( n300090 , n799 );
buf ( n300091 , n800 );
xor ( n300092 , n300090 , n300091 );
buf ( n300093 , n300092 );
buf ( n300094 , n300093 );
not ( n300095 , n300094 );
buf ( n9668 , n299589 );
not ( n9669 , n9668 );
or ( n9670 , n300095 , n9669 );
buf ( n300099 , n299471 );
buf ( n300100 , n6057 );
nand ( n300101 , n300099 , n300100 );
buf ( n300102 , n300101 );
buf ( n300103 , n300102 );
nand ( n300104 , n9670 , n300103 );
buf ( n300105 , n300104 );
buf ( n300106 , n300105 );
buf ( n9679 , n771 );
buf ( n9680 , n828 );
xor ( n9681 , n9679 , n9680 );
buf ( n9682 , n9681 );
buf ( n9683 , n9682 );
not ( n9684 , n9683 );
buf ( n9685 , n291805 );
not ( n9686 , n9685 );
or ( n9687 , n9684 , n9686 );
buf ( n9688 , n291812 );
buf ( n9689 , n299235 );
nand ( n9690 , n9688 , n9689 );
buf ( n9691 , n9690 );
buf ( n9692 , n9691 );
nand ( n9693 , n9687 , n9692 );
buf ( n9694 , n9693 );
buf ( n300123 , n9694 );
xor ( n9696 , n300106 , n300123 );
buf ( n300125 , n775 );
buf ( n300126 , n824 );
xor ( n9699 , n300125 , n300126 );
buf ( n9700 , n9699 );
buf ( n300129 , n9700 );
not ( n9702 , n300129 );
buf ( n300131 , n292473 );
not ( n300132 , n300131 );
or ( n9705 , n9702 , n300132 );
buf ( n300134 , n292870 );
buf ( n300135 , n299489 );
nand ( n300136 , n300134 , n300135 );
buf ( n300137 , n300136 );
buf ( n300138 , n300137 );
nand ( n300139 , n9705 , n300138 );
buf ( n300140 , n300139 );
buf ( n300141 , n300140 );
and ( n300142 , n9696 , n300141 );
and ( n300143 , n300106 , n300123 );
or ( n9716 , n300142 , n300143 );
buf ( n300145 , n9716 );
buf ( n300146 , n300145 );
xor ( n9719 , n9661 , n300146 );
buf ( n300148 , n785 );
buf ( n9721 , n814 );
xor ( n9722 , n300148 , n9721 );
buf ( n300151 , n9722 );
buf ( n300152 , n300151 );
not ( n300153 , n300152 );
buf ( n300154 , n8853 );
not ( n9727 , n300154 );
or ( n9728 , n300153 , n9727 );
xor ( n9729 , n784 , n814 );
nand ( n300158 , n9729 , n295478 );
buf ( n300159 , n300158 );
nand ( n9732 , n9728 , n300159 );
buf ( n300161 , n9732 );
buf ( n300162 , n300161 );
buf ( n300163 , n783 );
buf ( n300164 , n816 );
xor ( n300165 , n300163 , n300164 );
buf ( n300166 , n300165 );
buf ( n300167 , n300166 );
not ( n9740 , n300167 );
buf ( n300169 , n3977 );
not ( n300170 , n300169 );
or ( n300171 , n9740 , n300170 );
buf ( n300172 , n1712 );
buf ( n300173 , n299511 );
nand ( n300174 , n300172 , n300173 );
buf ( n300175 , n300174 );
buf ( n300176 , n300175 );
nand ( n300177 , n300171 , n300176 );
buf ( n300178 , n300177 );
buf ( n9751 , n300178 );
xor ( n9752 , n300162 , n9751 );
buf ( n300181 , n777 );
buf ( n9754 , n822 );
xor ( n300183 , n300181 , n9754 );
buf ( n300184 , n300183 );
buf ( n300185 , n300184 );
not ( n300186 , n300185 );
buf ( n300187 , n298771 );
not ( n300188 , n300187 );
or ( n9761 , n300186 , n300188 );
buf ( n300190 , n1600 );
buf ( n300191 , n8841 );
nand ( n9764 , n300190 , n300191 );
buf ( n300193 , n9764 );
buf ( n300194 , n300193 );
nand ( n9767 , n9761 , n300194 );
buf ( n300196 , n9767 );
buf ( n300197 , n300196 );
and ( n9770 , n9752 , n300197 );
and ( n300199 , n300162 , n9751 );
or ( n300200 , n9770 , n300199 );
buf ( n300201 , n300200 );
buf ( n300202 , n300201 );
and ( n300203 , n9719 , n300202 );
and ( n9776 , n9661 , n300146 );
or ( n300205 , n300203 , n9776 );
buf ( n300206 , n300205 );
buf ( n300207 , n300206 );
and ( n9780 , n9605 , n300207 );
and ( n300209 , n299925 , n300032 );
or ( n300210 , n9780 , n300209 );
buf ( n300211 , n300210 );
nand ( n300212 , n299853 , n300211 );
nand ( n9785 , n299852 , n300212 );
and ( n9786 , n299772 , n9785 );
and ( n300215 , n9112 , n299771 );
or ( n300216 , n9786 , n300215 );
buf ( n300217 , n300216 );
xor ( n300218 , n299175 , n300217 );
xor ( n300219 , n299544 , n299570 );
and ( n9792 , n300219 , n299769 );
and ( n300221 , n299544 , n299570 );
or ( n9794 , n9792 , n300221 );
buf ( n300223 , n9794 );
not ( n9796 , n300223 );
xor ( n9797 , n299552 , n299556 );
and ( n9798 , n9797 , n299567 );
and ( n9799 , n299552 , n299556 );
or ( n300228 , n9798 , n9799 );
buf ( n300229 , n300228 );
buf ( n300230 , n300229 );
buf ( n9803 , n299046 );
not ( n9804 , n9803 );
buf ( n300233 , n295983 );
not ( n9806 , n300233 );
or ( n300235 , n9804 , n9806 );
buf ( n300236 , n295361 );
xor ( n300237 , n804 , n789 );
buf ( n300238 , n300237 );
nand ( n9811 , n300236 , n300238 );
buf ( n300240 , n9811 );
buf ( n300241 , n300240 );
nand ( n9814 , n300235 , n300241 );
buf ( n300243 , n9814 );
buf ( n300244 , n8610 );
not ( n9817 , n300244 );
buf ( n300246 , n7960 );
not ( n300247 , n300246 );
or ( n9820 , n9817 , n300247 );
buf ( n300249 , n295929 );
xor ( n9822 , n802 , n791 );
buf ( n300251 , n9822 );
nand ( n9824 , n300249 , n300251 );
buf ( n9825 , n9824 );
buf ( n300254 , n9825 );
nand ( n9827 , n9820 , n300254 );
buf ( n300256 , n9827 );
xor ( n300257 , n300243 , n300256 );
buf ( n300258 , n8515 );
not ( n9831 , n300258 );
buf ( n300260 , n2078 );
not ( n9833 , n300260 );
or ( n300262 , n9831 , n9833 );
buf ( n300263 , n2089 );
buf ( n300264 , n779 );
buf ( n300265 , n814 );
xor ( n300266 , n300264 , n300265 );
buf ( n300267 , n300266 );
buf ( n300268 , n300267 );
nand ( n300269 , n300263 , n300268 );
buf ( n300270 , n300269 );
buf ( n300271 , n300270 );
nand ( n9844 , n300262 , n300271 );
buf ( n300273 , n9844 );
not ( n9846 , n300273 );
and ( n300275 , n300257 , n9846 );
not ( n9848 , n300257 );
and ( n300277 , n9848 , n300273 );
nor ( n300278 , n300275 , n300277 );
not ( n9851 , n300278 );
buf ( n300280 , n8641 );
not ( n9853 , n300280 );
buf ( n300282 , n294637 );
not ( n300283 , n300282 );
or ( n9856 , n9853 , n300283 );
buf ( n300285 , n293902 );
xor ( n300286 , n806 , n787 );
buf ( n9859 , n300286 );
nand ( n9860 , n300285 , n9859 );
buf ( n300289 , n9860 );
buf ( n300290 , n300289 );
nand ( n9863 , n9856 , n300290 );
buf ( n9864 , n9863 );
buf ( n9865 , n9864 );
not ( n9866 , n9865 );
buf ( n300295 , n9866 );
not ( n300296 , n300295 );
not ( n300297 , n298891 );
not ( n300298 , n298771 );
or ( n300299 , n300297 , n300298 );
buf ( n300300 , n1600 );
xor ( n9873 , n822 , n771 );
buf ( n300302 , n9873 );
nand ( n300303 , n300300 , n300302 );
buf ( n300304 , n300303 );
nand ( n300305 , n300299 , n300304 );
not ( n9878 , n300305 );
or ( n9879 , n300296 , n9878 );
not ( n300308 , n300305 );
buf ( n300309 , n300308 );
buf ( n300310 , n9864 );
nand ( n300311 , n300309 , n300310 );
buf ( n300312 , n300311 );
nand ( n9885 , n9879 , n300312 );
buf ( n300314 , n299055 );
not ( n300315 , n300314 );
buf ( n300316 , n2118 );
not ( n300317 , n300316 );
or ( n300318 , n300315 , n300317 );
buf ( n300319 , n1712 );
buf ( n9892 , n777 );
buf ( n9893 , n816 );
xor ( n9894 , n9892 , n9893 );
buf ( n9895 , n9894 );
buf ( n300324 , n9895 );
nand ( n9897 , n300319 , n300324 );
buf ( n300326 , n9897 );
buf ( n300327 , n300326 );
nand ( n9900 , n300318 , n300327 );
buf ( n300329 , n9900 );
not ( n300330 , n300329 );
and ( n9903 , n9885 , n300330 );
not ( n300332 , n9885 );
and ( n300333 , n300332 , n300329 );
nor ( n9906 , n9903 , n300333 );
not ( n300335 , n9906 );
and ( n300336 , n9851 , n300335 );
not ( n9909 , n9851 );
and ( n9910 , n9909 , n9906 );
nor ( n9911 , n300336 , n9910 );
buf ( n300340 , n8657 );
not ( n300341 , n300340 );
buf ( n300342 , n292393 );
not ( n9915 , n300342 );
or ( n9916 , n300341 , n9915 );
buf ( n300345 , n291788 );
buf ( n300346 , n775 );
buf ( n300347 , n818 );
xor ( n9920 , n300346 , n300347 );
buf ( n300349 , n9920 );
buf ( n9922 , n300349 );
nand ( n9923 , n300345 , n9922 );
buf ( n9924 , n9923 );
buf ( n300353 , n9924 );
nand ( n9926 , n9916 , n300353 );
buf ( n300355 , n9926 );
buf ( n300356 , n298998 );
not ( n300357 , n300356 );
buf ( n300358 , n298990 );
not ( n300359 , n300358 );
or ( n300360 , n300357 , n300359 );
buf ( n300361 , n294557 );
buf ( n300362 , n785 );
buf ( n300363 , n808 );
xor ( n9936 , n300362 , n300363 );
buf ( n300365 , n9936 );
buf ( n300366 , n300365 );
nand ( n9939 , n300361 , n300366 );
buf ( n300368 , n9939 );
buf ( n300369 , n300368 );
nand ( n9942 , n300360 , n300369 );
buf ( n9943 , n9942 );
xor ( n300372 , n300355 , n9943 );
buf ( n300373 , n300372 );
buf ( n300374 , n299020 );
not ( n9947 , n300374 );
buf ( n300376 , n293058 );
not ( n300377 , n300376 );
or ( n9950 , n9947 , n300377 );
buf ( n300379 , n292841 );
buf ( n9952 , n783 );
buf ( n300381 , n810 );
xor ( n300382 , n9952 , n300381 );
buf ( n300383 , n300382 );
buf ( n300384 , n300383 );
nand ( n300385 , n300379 , n300384 );
buf ( n300386 , n300385 );
buf ( n300387 , n300386 );
nand ( n9960 , n9950 , n300387 );
buf ( n9961 , n9960 );
buf ( n300390 , n9961 );
xor ( n9963 , n300373 , n300390 );
buf ( n300392 , n9963 );
and ( n300393 , n9911 , n300392 );
not ( n300394 , n9911 );
buf ( n300395 , n300392 );
not ( n300396 , n300395 );
buf ( n300397 , n300396 );
and ( n9970 , n300394 , n300397 );
nor ( n300399 , n300393 , n9970 );
buf ( n300400 , n300399 );
xor ( n9973 , n300230 , n300400 );
xor ( n300402 , n299621 , n299625 );
and ( n300403 , n300402 , n299766 );
and ( n9976 , n299621 , n299625 );
or ( n300405 , n300403 , n9976 );
buf ( n300406 , n300405 );
buf ( n300407 , n300406 );
xor ( n300408 , n9973 , n300407 );
buf ( n300409 , n300408 );
not ( n9982 , n300409 );
not ( n300411 , n9982 );
or ( n9984 , n9796 , n300411 );
not ( n300413 , n300223 );
nand ( n9986 , n300409 , n300413 );
nand ( n9987 , n9984 , n9986 );
xor ( n9988 , n299777 , n9354 );
and ( n300417 , n9988 , n9357 );
and ( n300418 , n299777 , n9354 );
or ( n9991 , n300417 , n300418 );
not ( n9992 , n9991 );
xor ( n9993 , n299789 , n9400 );
and ( n300422 , n9993 , n299850 );
and ( n300423 , n299789 , n9400 );
or ( n9996 , n300422 , n300423 );
not ( n300425 , n9996 );
nand ( n300426 , n9992 , n300425 );
not ( n9999 , n300426 );
nand ( n300428 , n8152 , n8153 );
xor ( n300429 , n298793 , n300428 );
xnor ( n10002 , n300429 , n8295 );
not ( n300431 , n10002 );
or ( n300432 , n9999 , n300431 );
nand ( n10005 , n9991 , n9996 );
nand ( n300434 , n300432 , n10005 );
and ( n300435 , n9987 , n300434 );
not ( n10008 , n9987 );
not ( n300437 , n300434 );
and ( n300438 , n10008 , n300437 );
nor ( n300439 , n300435 , n300438 );
buf ( n300440 , n300439 );
and ( n300441 , n300218 , n300440 );
and ( n10014 , n299175 , n300217 );
or ( n300443 , n300441 , n10014 );
buf ( n300444 , n300443 );
buf ( n300445 , n298863 );
buf ( n300446 , n8395 );
nand ( n300447 , n300445 , n300446 );
buf ( n300448 , n300447 );
not ( n10021 , n300448 );
not ( n300450 , n298876 );
or ( n300451 , n10021 , n300450 );
buf ( n300452 , n8395 );
not ( n300453 , n300452 );
buf ( n300454 , n298860 );
nand ( n10027 , n300453 , n300454 );
buf ( n10028 , n10027 );
nand ( n300457 , n300451 , n10028 );
xor ( n300458 , n298958 , n299035 );
and ( n300459 , n300458 , n299167 );
and ( n10032 , n298958 , n299035 );
or ( n300461 , n300459 , n10032 );
buf ( n300462 , n300461 );
xor ( n300463 , n300457 , n300462 );
xor ( n300464 , n299063 , n299115 );
and ( n300465 , n300464 , n299164 );
and ( n300466 , n299063 , n299115 );
or ( n10039 , n300465 , n300466 );
buf ( n300468 , n10039 );
buf ( n300469 , n8394 );
xor ( n300470 , n299126 , n299143 );
and ( n10043 , n300470 , n299161 );
and ( n300472 , n299126 , n299143 );
or ( n300473 , n10043 , n300472 );
buf ( n300474 , n300473 );
buf ( n300475 , n300474 );
xor ( n300476 , n300469 , n300475 );
buf ( n300477 , n9943 );
buf ( n300478 , n300355 );
or ( n300479 , n300477 , n300478 );
buf ( n300480 , n9961 );
nand ( n10053 , n300479 , n300480 );
buf ( n300482 , n10053 );
buf ( n300483 , n300482 );
buf ( n300484 , n9943 );
buf ( n300485 , n300355 );
nand ( n10058 , n300484 , n300485 );
buf ( n300487 , n10058 );
buf ( n300488 , n300487 );
nand ( n10061 , n300483 , n300488 );
buf ( n300490 , n10061 );
buf ( n300491 , n300490 );
xor ( n300492 , n300476 , n300491 );
buf ( n300493 , n300492 );
and ( n300494 , n300468 , n300493 );
not ( n300495 , n300468 );
buf ( n300496 , n300493 );
not ( n10069 , n300496 );
buf ( n300498 , n10069 );
and ( n300499 , n300495 , n300498 );
nor ( n300500 , n300494 , n300499 );
buf ( n300501 , n300256 );
not ( n300502 , n300501 );
buf ( n300503 , n300243 );
not ( n300504 , n300503 );
or ( n300505 , n300502 , n300504 );
buf ( n300506 , n300243 );
buf ( n300507 , n300256 );
or ( n10080 , n300506 , n300507 );
buf ( n300509 , n300273 );
nand ( n300510 , n10080 , n300509 );
buf ( n300511 , n300510 );
buf ( n300512 , n300511 );
nand ( n300513 , n300505 , n300512 );
buf ( n300514 , n300513 );
not ( n10087 , n300329 );
nand ( n300516 , n300295 , n300308 );
not ( n300517 , n300516 );
or ( n10090 , n10087 , n300517 );
nand ( n300519 , n300305 , n9864 );
nand ( n10092 , n10090 , n300519 );
xor ( n300521 , n300514 , n10092 );
buf ( n300522 , n299136 );
not ( n10095 , n300522 );
buf ( n300524 , n3539 );
not ( n300525 , n300524 );
or ( n300526 , n10095 , n300525 );
buf ( n300527 , n780 );
buf ( n300528 , n812 );
xor ( n300529 , n300527 , n300528 );
buf ( n300530 , n300529 );
buf ( n300531 , n300530 );
buf ( n300532 , n292810 );
nand ( n300533 , n300531 , n300532 );
buf ( n300534 , n300533 );
buf ( n300535 , n300534 );
nand ( n300536 , n300526 , n300535 );
buf ( n300537 , n300536 );
buf ( n300538 , n300537 );
buf ( n300539 , n300383 );
not ( n300540 , n300539 );
buf ( n300541 , n3041 );
not ( n10114 , n300541 );
or ( n300543 , n300540 , n10114 );
buf ( n300544 , n295259 );
buf ( n300545 , n782 );
buf ( n300546 , n810 );
xor ( n10119 , n300545 , n300546 );
buf ( n300548 , n10119 );
buf ( n10121 , n300548 );
nand ( n10122 , n300544 , n10121 );
buf ( n10123 , n10122 );
buf ( n300552 , n10123 );
nand ( n10125 , n300543 , n300552 );
buf ( n300554 , n10125 );
buf ( n300555 , n300554 );
xor ( n300556 , n300538 , n300555 );
buf ( n300557 , n300349 );
not ( n300558 , n300557 );
buf ( n300559 , n1553 );
not ( n300560 , n300559 );
or ( n300561 , n300558 , n300560 );
buf ( n300562 , n291989 );
buf ( n300563 , n774 );
buf ( n10136 , n818 );
xor ( n300565 , n300563 , n10136 );
buf ( n300566 , n300565 );
buf ( n300567 , n300566 );
nand ( n300568 , n300562 , n300567 );
buf ( n300569 , n300568 );
buf ( n300570 , n300569 );
nand ( n300571 , n300561 , n300570 );
buf ( n300572 , n300571 );
buf ( n300573 , n300572 );
xor ( n300574 , n300556 , n300573 );
buf ( n300575 , n300574 );
xor ( n300576 , n300521 , n300575 );
and ( n300577 , n300500 , n300576 );
not ( n300578 , n300500 );
not ( n10151 , n300576 );
and ( n300580 , n300578 , n10151 );
nor ( n300581 , n300577 , n300580 );
xor ( n300582 , n300463 , n300581 );
buf ( n300583 , n300582 );
not ( n10156 , n300223 );
not ( n300585 , n9982 );
not ( n300586 , n300585 );
or ( n10159 , n10156 , n300586 );
or ( n300588 , n300585 , n300223 );
nand ( n300589 , n300588 , n300434 );
nand ( n300590 , n10159 , n300589 );
buf ( n300591 , n300590 );
xor ( n10164 , n300583 , n300591 );
xor ( n300593 , n300230 , n300400 );
and ( n10166 , n300593 , n300407 );
and ( n10167 , n300230 , n300400 );
or ( n300596 , n10166 , n10167 );
buf ( n300597 , n300596 );
buf ( n300598 , n794 );
buf ( n300599 , n800 );
and ( n300600 , n300598 , n300599 );
buf ( n300601 , n300600 );
buf ( n300602 , n8380 );
not ( n300603 , n300602 );
buf ( n300604 , n299589 );
not ( n300605 , n300604 );
or ( n300606 , n300603 , n300605 );
buf ( n300607 , n6057 );
buf ( n300608 , n792 );
buf ( n300609 , n800 );
xor ( n10182 , n300608 , n300609 );
buf ( n300611 , n10182 );
buf ( n300612 , n300611 );
nand ( n10185 , n300607 , n300612 );
buf ( n300614 , n10185 );
buf ( n300615 , n300614 );
nand ( n10188 , n300606 , n300615 );
buf ( n10189 , n10188 );
xor ( n300618 , n300601 , n10189 );
buf ( n300619 , n778 );
buf ( n300620 , n814 );
xor ( n300621 , n300619 , n300620 );
buf ( n300622 , n300621 );
not ( n300623 , n300622 );
not ( n300624 , n292725 );
or ( n10197 , n300623 , n300624 );
nand ( n300626 , n292509 , n300267 );
nand ( n10199 , n10197 , n300626 );
xor ( n10200 , n300618 , n10199 );
buf ( n300629 , n10200 );
buf ( n300630 , n299121 );
not ( n10203 , n300630 );
buf ( n300632 , n292473 );
not ( n300633 , n300632 );
or ( n10206 , n10203 , n300633 );
buf ( n10207 , n1613 );
buf ( n300636 , n768 );
buf ( n300637 , n824 );
xor ( n300638 , n300636 , n300637 );
buf ( n300639 , n300638 );
buf ( n300640 , n300639 );
nand ( n300641 , n10207 , n300640 );
buf ( n300642 , n300641 );
buf ( n300643 , n300642 );
nand ( n10216 , n10206 , n300643 );
buf ( n300645 , n10216 );
buf ( n10218 , n300645 );
not ( n10219 , n10218 );
buf ( n300648 , n10219 );
buf ( n300649 , n300648 );
not ( n10222 , n300649 );
buf ( n300651 , n299154 );
not ( n300652 , n300651 );
buf ( n300653 , n292668 );
not ( n300654 , n300653 );
or ( n300655 , n300652 , n300654 );
buf ( n300656 , n291969 );
buf ( n300657 , n772 );
buf ( n300658 , n820 );
xor ( n10231 , n300657 , n300658 );
buf ( n300660 , n10231 );
buf ( n300661 , n300660 );
nand ( n300662 , n300656 , n300661 );
buf ( n300663 , n300662 );
buf ( n300664 , n300663 );
nand ( n10237 , n300655 , n300664 );
buf ( n10238 , n10237 );
nand ( n10239 , n8317 , n2965 );
not ( n300668 , n10239 );
not ( n10241 , n291886 );
not ( n300670 , n10241 );
or ( n300671 , n300668 , n300670 );
nand ( n300672 , n300671 , n826 );
xor ( n10245 , n10238 , n300672 );
buf ( n300674 , n10245 );
not ( n300675 , n300674 );
or ( n10248 , n10222 , n300675 );
buf ( n300677 , n10245 );
buf ( n300678 , n300648 );
or ( n10251 , n300677 , n300678 );
nand ( n300680 , n10248 , n10251 );
buf ( n300681 , n300680 );
buf ( n300682 , n300681 );
xor ( n300683 , n300629 , n300682 );
buf ( n300684 , n300237 );
not ( n300685 , n300684 );
buf ( n300686 , n295983 );
not ( n300687 , n300686 );
or ( n10260 , n300685 , n300687 );
buf ( n300689 , n5554 );
buf ( n300690 , n788 );
buf ( n300691 , n804 );
xor ( n300692 , n300690 , n300691 );
buf ( n300693 , n300692 );
buf ( n300694 , n300693 );
nand ( n300695 , n300689 , n300694 );
buf ( n300696 , n300695 );
buf ( n300697 , n300696 );
nand ( n300698 , n10260 , n300697 );
buf ( n300699 , n300698 );
buf ( n300700 , n300699 );
buf ( n300701 , n9895 );
not ( n10274 , n300701 );
buf ( n300703 , n292892 );
not ( n300704 , n300703 );
or ( n300705 , n10274 , n300704 );
buf ( n300706 , n1712 );
buf ( n300707 , n776 );
buf ( n300708 , n816 );
xor ( n300709 , n300707 , n300708 );
buf ( n300710 , n300709 );
buf ( n300711 , n300710 );
nand ( n300712 , n300706 , n300711 );
buf ( n300713 , n300712 );
buf ( n300714 , n300713 );
nand ( n10287 , n300705 , n300714 );
buf ( n10288 , n10287 );
buf ( n300717 , n10288 );
xor ( n10290 , n300700 , n300717 );
buf ( n300719 , n9822 );
not ( n300720 , n300719 );
buf ( n300721 , n6079 );
not ( n300722 , n300721 );
or ( n300723 , n300720 , n300722 );
buf ( n300724 , n296749 );
buf ( n300725 , n790 );
buf ( n300726 , n802 );
xor ( n10299 , n300725 , n300726 );
buf ( n10300 , n10299 );
buf ( n300729 , n10300 );
nand ( n10302 , n300724 , n300729 );
buf ( n10303 , n10302 );
buf ( n300732 , n10303 );
nand ( n10305 , n300723 , n300732 );
buf ( n10306 , n10305 );
buf ( n300735 , n10306 );
xor ( n300736 , n10290 , n300735 );
buf ( n300737 , n300736 );
buf ( n300738 , n300737 );
xor ( n300739 , n300683 , n300738 );
buf ( n300740 , n300739 );
not ( n10313 , n9851 );
not ( n300742 , n300335 );
or ( n300743 , n10313 , n300742 );
not ( n300744 , n9906 );
not ( n300745 , n300278 );
or ( n10318 , n300744 , n300745 );
nand ( n300747 , n10318 , n300392 );
nand ( n300748 , n300743 , n300747 );
not ( n10321 , n300748 );
xor ( n300750 , n300740 , n10321 );
or ( n300751 , n8394 , n298796 );
not ( n10324 , n298796 );
not ( n300753 , n8394 );
or ( n300754 , n10324 , n300753 );
nand ( n10327 , n300754 , n8384 );
nand ( n300756 , n300751 , n10327 );
buf ( n300757 , n300756 );
buf ( n300758 , n300365 );
not ( n10331 , n300758 );
buf ( n300760 , n293655 );
not ( n300761 , n300760 );
or ( n10334 , n10331 , n300761 );
buf ( n300763 , n294557 );
buf ( n300764 , n784 );
buf ( n300765 , n808 );
xor ( n10338 , n300764 , n300765 );
buf ( n300767 , n10338 );
buf ( n300768 , n300767 );
nand ( n300769 , n300763 , n300768 );
buf ( n300770 , n300769 );
buf ( n300771 , n300770 );
nand ( n300772 , n10334 , n300771 );
buf ( n300773 , n300772 );
buf ( n300774 , n300773 );
not ( n300775 , n300774 );
buf ( n300776 , n300775 );
buf ( n300777 , n300286 );
not ( n10350 , n300777 );
buf ( n300779 , n5676 );
not ( n300780 , n300779 );
or ( n10353 , n10350 , n300780 );
buf ( n300782 , n295437 );
and ( n10355 , n786 , n806 );
not ( n10356 , n786 );
not ( n300785 , n806 );
and ( n10358 , n10356 , n300785 );
nor ( n300787 , n10355 , n10358 );
buf ( n300788 , n300787 );
nand ( n10361 , n300782 , n300788 );
buf ( n10362 , n10361 );
buf ( n300791 , n10362 );
nand ( n10364 , n10353 , n300791 );
buf ( n300793 , n10364 );
xor ( n10366 , n300776 , n300793 );
buf ( n300795 , n9873 );
not ( n10368 , n300795 );
buf ( n300797 , n292631 );
not ( n300798 , n300797 );
or ( n10371 , n10368 , n300798 );
buf ( n300800 , n1600 );
buf ( n300801 , n770 );
buf ( n300802 , n822 );
xor ( n300803 , n300801 , n300802 );
buf ( n300804 , n300803 );
buf ( n300805 , n300804 );
nand ( n300806 , n300800 , n300805 );
buf ( n300807 , n300806 );
buf ( n300808 , n300807 );
nand ( n300809 , n10371 , n300808 );
buf ( n300810 , n300809 );
buf ( n300811 , n300810 );
not ( n300812 , n300811 );
buf ( n300813 , n300812 );
xor ( n10386 , n10366 , n300813 );
buf ( n300815 , n10386 );
xor ( n10388 , n300757 , n300815 );
xor ( n10389 , n298963 , n298969 );
and ( n300818 , n10389 , n299032 );
and ( n300819 , n298963 , n298969 );
or ( n10392 , n300818 , n300819 );
buf ( n300821 , n10392 );
buf ( n300822 , n300821 );
xor ( n10395 , n10388 , n300822 );
buf ( n300824 , n10395 );
xnor ( n10397 , n300750 , n300824 );
xor ( n300826 , n300597 , n10397 );
buf ( n300827 , n298881 );
not ( n10400 , n300827 );
buf ( n300829 , n299169 );
not ( n300830 , n300829 );
or ( n10403 , n10400 , n300830 );
or ( n300832 , n299169 , n298881 );
nand ( n10405 , n300832 , n8367 );
buf ( n10406 , n10405 );
nand ( n10407 , n10403 , n10406 );
buf ( n10408 , n10407 );
xor ( n300837 , n300826 , n10408 );
buf ( n300838 , n300837 );
xor ( n300839 , n10164 , n300838 );
buf ( n300840 , n300839 );
and ( n10413 , n300444 , n300840 );
buf ( n300842 , n10413 );
not ( n300843 , n300842 );
or ( n10416 , n7954 , n300843 );
buf ( n300845 , n831 );
not ( n300846 , n300845 );
buf ( n300847 , n300840 );
buf ( n300848 , n300444 );
and ( n300849 , n300847 , n300848 );
buf ( n300850 , n300849 );
buf ( n300851 , n300850 );
nand ( n300852 , n300846 , n300851 );
buf ( n300853 , n300852 );
buf ( n300854 , n300853 );
nand ( n300855 , n10416 , n300854 );
buf ( n300856 , n300855 );
buf ( n10429 , n300856 );
buf ( n300858 , n831 );
not ( n300859 , n300858 );
buf ( n300860 , n847 );
not ( n10433 , n292288 );
not ( n10434 , n292277 );
not ( n300863 , n10434 );
or ( n10436 , n10433 , n300863 );
nand ( n300865 , n10436 , n1877 );
not ( n300866 , n292288 );
nand ( n10439 , n300866 , n292277 );
nand ( n300868 , n300865 , n10439 );
buf ( n10441 , n300868 );
buf ( n300870 , n292176 );
not ( n300871 , n300870 );
buf ( n300872 , n292168 );
not ( n300873 , n300872 );
or ( n300874 , n300871 , n300873 );
buf ( n300875 , n291812 );
buf ( n300876 , n298022 );
nand ( n10449 , n300875 , n300876 );
buf ( n300878 , n10449 );
buf ( n300879 , n300878 );
nand ( n10452 , n300874 , n300879 );
buf ( n300881 , n10452 );
not ( n10454 , n292283 );
not ( n300883 , n7526 );
or ( n300884 , n10454 , n300883 );
buf ( n300885 , n1613 );
buf ( n300886 , n298117 );
nand ( n300887 , n300885 , n300886 );
buf ( n300888 , n300887 );
nand ( n300889 , n300884 , n300888 );
xor ( n300890 , n300881 , n300889 );
buf ( n300891 , n799 );
buf ( n300892 , n816 );
xor ( n300893 , n300891 , n300892 );
buf ( n300894 , n300893 );
buf ( n300895 , n300894 );
not ( n10468 , n300895 );
buf ( n300897 , n2118 );
not ( n300898 , n300897 );
or ( n300899 , n10468 , n300898 );
buf ( n300900 , n1712 );
buf ( n300901 , n298153 );
nand ( n300902 , n300900 , n300901 );
buf ( n300903 , n300902 );
buf ( n300904 , n300903 );
nand ( n300905 , n300899 , n300904 );
buf ( n300906 , n300905 );
xor ( n300907 , n300890 , n300906 );
buf ( n300908 , n300907 );
xor ( n10481 , n10441 , n300908 );
buf ( n300910 , n292255 );
not ( n300911 , n300910 );
buf ( n300912 , n291722 );
not ( n300913 , n300912 );
or ( n10486 , n300911 , n300913 );
buf ( n300915 , n291969 );
buf ( n300916 , n7668 );
nand ( n10489 , n300915 , n300916 );
buf ( n300918 , n10489 );
buf ( n300919 , n300918 );
nand ( n10492 , n10486 , n300919 );
buf ( n300921 , n10492 );
buf ( n300922 , n292273 );
not ( n10495 , n300922 );
buf ( n300924 , n1453 );
not ( n300925 , n300924 );
or ( n10498 , n10495 , n300925 );
buf ( n300927 , n291886 );
buf ( n300928 , n298076 );
nand ( n300929 , n300927 , n300928 );
buf ( n300930 , n300929 );
buf ( n300931 , n300930 );
nand ( n300932 , n10498 , n300931 );
buf ( n300933 , n300932 );
buf ( n300934 , n300933 );
not ( n300935 , n300934 );
buf ( n300936 , n300935 );
xor ( n300937 , n300921 , n300936 );
buf ( n300938 , n292301 );
not ( n10511 , n300938 );
buf ( n300940 , n291761 );
not ( n300941 , n300940 );
or ( n300942 , n10511 , n300941 );
buf ( n300943 , n292104 );
buf ( n300944 , n298134 );
nand ( n300945 , n300943 , n300944 );
buf ( n300946 , n300945 );
buf ( n300947 , n300946 );
nand ( n300948 , n300942 , n300947 );
buf ( n300949 , n300948 );
xnor ( n300950 , n300937 , n300949 );
buf ( n300951 , n300950 );
xor ( n10524 , n10481 , n300951 );
buf ( n300953 , n10524 );
buf ( n10526 , n300953 );
xor ( n300955 , n1799 , n292244 );
and ( n300956 , n300955 , n292262 );
and ( n10529 , n1799 , n292244 );
or ( n300958 , n300956 , n10529 );
buf ( n300959 , n300958 );
buf ( n300960 , n300959 );
buf ( n300961 , n292237 );
not ( n10534 , n300961 );
buf ( n300963 , n291984 );
not ( n300964 , n300963 );
or ( n300965 , n10534 , n300964 );
buf ( n300966 , n291989 );
buf ( n300967 , n298057 );
nand ( n300968 , n300966 , n300967 );
buf ( n300969 , n300968 );
buf ( n300970 , n300969 );
nand ( n300971 , n300965 , n300970 );
buf ( n300972 , n300971 );
buf ( n300973 , n300972 );
buf ( n300974 , n799 );
buf ( n300975 , n817 );
or ( n10548 , n300974 , n300975 );
buf ( n300977 , n818 );
nand ( n300978 , n10548 , n300977 );
buf ( n300979 , n300978 );
buf ( n300980 , n300979 );
buf ( n300981 , n799 );
buf ( n300982 , n817 );
nand ( n300983 , n300981 , n300982 );
buf ( n300984 , n300983 );
buf ( n300985 , n300984 );
buf ( n300986 , n816 );
and ( n300987 , n300980 , n300985 , n300986 );
buf ( n300988 , n300987 );
buf ( n300989 , n300988 );
buf ( n300990 , n292154 );
not ( n300991 , n300990 );
buf ( n300992 , n291656 );
not ( n300993 , n300992 );
or ( n300994 , n300991 , n300993 );
buf ( n300995 , n298005 );
buf ( n300996 , n831 );
nand ( n300997 , n300995 , n300996 );
buf ( n300998 , n300997 );
buf ( n300999 , n300998 );
nand ( n10572 , n300994 , n300999 );
buf ( n301001 , n10572 );
buf ( n301002 , n301001 );
xor ( n10575 , n300989 , n301002 );
buf ( n301004 , n10575 );
buf ( n301005 , n301004 );
xor ( n301006 , n300973 , n301005 );
xor ( n301007 , n292145 , n292162 );
and ( n10580 , n301007 , n292183 );
and ( n301009 , n292145 , n292162 );
or ( n301010 , n10580 , n301009 );
buf ( n301011 , n301010 );
buf ( n301012 , n301011 );
xor ( n301013 , n301006 , n301012 );
buf ( n301014 , n301013 );
buf ( n301015 , n301014 );
xor ( n10588 , n300960 , n301015 );
xor ( n10589 , n1758 , n292205 );
and ( n301018 , n10589 , n292212 );
and ( n301019 , n1758 , n292205 );
or ( n301020 , n301018 , n301019 );
buf ( n301021 , n301020 );
buf ( n301022 , n301021 );
xor ( n301023 , n10588 , n301022 );
buf ( n301024 , n301023 );
buf ( n301025 , n301024 );
xor ( n301026 , n10526 , n301025 );
xor ( n10599 , n292265 , n292310 );
and ( n301028 , n10599 , n292317 );
and ( n301029 , n292265 , n292310 );
or ( n10602 , n301028 , n301029 );
buf ( n301031 , n10602 );
buf ( n301032 , n301031 );
and ( n10605 , n301026 , n301032 );
and ( n10606 , n10526 , n301025 );
or ( n301035 , n10605 , n10606 );
buf ( n301036 , n301035 );
buf ( n301037 , n301036 );
xor ( n301038 , n300860 , n301037 );
xor ( n10611 , n298017 , n7616 );
xor ( n10612 , n10611 , n298038 );
not ( n301041 , n7682 );
not ( n10614 , n7660 );
or ( n10615 , n301041 , n10614 );
or ( n301044 , n7682 , n7660 );
nand ( n301045 , n10615 , n301044 );
buf ( n301046 , n301045 );
buf ( n301047 , n298070 );
buf ( n10620 , n301047 );
and ( n10621 , n301046 , n10620 );
not ( n301050 , n301046 );
not ( n301051 , n301047 );
buf ( n301052 , n301051 );
and ( n301053 , n301050 , n301052 );
nor ( n10626 , n10621 , n301053 );
buf ( n301055 , n10626 );
buf ( n10628 , n301055 );
not ( n301057 , n10628 );
buf ( n301058 , n301057 );
xor ( n10631 , n10612 , n301058 );
xor ( n301060 , n298130 , n298148 );
xor ( n301061 , n301060 , n298166 );
buf ( n301062 , n301061 );
xnor ( n301063 , n10631 , n301062 );
buf ( n301064 , n301063 );
xor ( n10637 , n300960 , n301015 );
and ( n301066 , n10637 , n301022 );
and ( n301067 , n300960 , n301015 );
or ( n10640 , n301066 , n301067 );
buf ( n301069 , n10640 );
buf ( n301070 , n301069 );
xor ( n10643 , n301064 , n301070 );
xor ( n301072 , n300973 , n301005 );
and ( n301073 , n301072 , n301012 );
and ( n301074 , n300973 , n301005 );
or ( n301075 , n301073 , n301074 );
buf ( n301076 , n301075 );
buf ( n301077 , n301076 );
and ( n301078 , n300989 , n301002 );
buf ( n301079 , n301078 );
buf ( n301080 , n301079 );
buf ( n301081 , n300881 );
not ( n10654 , n301081 );
buf ( n301083 , n300889 );
not ( n301084 , n301083 );
or ( n301085 , n10654 , n301084 );
buf ( n301086 , n300889 );
buf ( n301087 , n300881 );
or ( n301088 , n301086 , n301087 );
buf ( n301089 , n300906 );
nand ( n301090 , n301088 , n301089 );
buf ( n301091 , n301090 );
buf ( n301092 , n301091 );
nand ( n301093 , n301085 , n301092 );
buf ( n301094 , n301093 );
buf ( n10667 , n301094 );
xor ( n10668 , n301080 , n10667 );
not ( n301097 , n300933 );
not ( n301098 , n300921 );
or ( n10671 , n301097 , n301098 );
buf ( n10672 , n300933 );
buf ( n301101 , n300921 );
nor ( n301102 , n10672 , n301101 );
buf ( n301103 , n301102 );
buf ( n301104 , n300949 );
not ( n10677 , n301104 );
buf ( n301106 , n10677 );
or ( n301107 , n301103 , n301106 );
nand ( n301108 , n10671 , n301107 );
buf ( n301109 , n301108 );
xor ( n301110 , n10668 , n301109 );
buf ( n301111 , n301110 );
buf ( n301112 , n301111 );
xor ( n301113 , n301077 , n301112 );
xor ( n301114 , n10441 , n300908 );
and ( n10687 , n301114 , n300951 );
and ( n301116 , n10441 , n300908 );
or ( n10689 , n10687 , n301116 );
buf ( n301118 , n10689 );
buf ( n301119 , n301118 );
xor ( n10692 , n301113 , n301119 );
buf ( n301121 , n10692 );
buf ( n301122 , n301121 );
xor ( n10695 , n10643 , n301122 );
buf ( n301124 , n10695 );
buf ( n301125 , n301124 );
and ( n10698 , n301038 , n301125 );
and ( n301127 , n300860 , n301037 );
or ( n301128 , n10698 , n301127 );
buf ( n301129 , n301128 );
buf ( n301130 , n301129 );
not ( n301131 , n301130 );
or ( n301132 , n300859 , n301131 );
buf ( n301133 , n879 );
buf ( n301134 , n301036 );
xor ( n301135 , n301133 , n301134 );
buf ( n301136 , n301124 );
and ( n301137 , n301135 , n301136 );
and ( n10710 , n301133 , n301134 );
or ( n301139 , n301137 , n10710 );
buf ( n301140 , n301139 );
buf ( n301141 , n301140 );
buf ( n301142 , n5980 );
nand ( n10715 , n301141 , n301142 );
buf ( n301144 , n10715 );
buf ( n301145 , n301144 );
nand ( n301146 , n301132 , n301145 );
buf ( n301147 , n301146 );
buf ( n10720 , n301147 );
not ( n301149 , n831 );
xor ( n301150 , n297635 , n297650 );
xor ( n10723 , n301150 , n297668 );
buf ( n301152 , n10723 );
buf ( n301153 , n301152 );
buf ( n301154 , n788 );
buf ( n301155 , n800 );
xor ( n301156 , n301154 , n301155 );
buf ( n301157 , n301156 );
buf ( n301158 , n301157 );
not ( n301159 , n301158 );
buf ( n301160 , n296480 );
not ( n10733 , n301160 );
or ( n301162 , n301159 , n10733 );
buf ( n301163 , n6057 );
buf ( n301164 , n297572 );
nand ( n301165 , n301163 , n301164 );
buf ( n301166 , n301165 );
buf ( n301167 , n301166 );
nand ( n301168 , n301162 , n301167 );
buf ( n301169 , n301168 );
buf ( n301170 , n301169 );
buf ( n301171 , n786 );
buf ( n301172 , n802 );
xor ( n301173 , n301171 , n301172 );
buf ( n301174 , n301173 );
buf ( n301175 , n301174 );
not ( n301176 , n301175 );
buf ( n301177 , n296508 );
not ( n301178 , n301177 );
or ( n10751 , n301176 , n301178 );
buf ( n301180 , n296749 );
buf ( n10753 , n297589 );
nand ( n10754 , n301180 , n10753 );
buf ( n10755 , n10754 );
buf ( n10756 , n10755 );
nand ( n10757 , n10751 , n10756 );
buf ( n10758 , n10757 );
buf ( n10759 , n10758 );
xor ( n10760 , n301170 , n10759 );
xor ( n301189 , n812 , n776 );
buf ( n301190 , n301189 );
not ( n10763 , n301190 );
buf ( n301192 , n2376 );
not ( n301193 , n301192 );
or ( n10766 , n10763 , n301193 );
buf ( n301195 , n2383 );
buf ( n301196 , n7246 );
nand ( n10769 , n301195 , n301196 );
buf ( n301198 , n10769 );
buf ( n301199 , n301198 );
nand ( n301200 , n10766 , n301199 );
buf ( n301201 , n301200 );
buf ( n301202 , n301201 );
and ( n301203 , n10760 , n301202 );
and ( n10776 , n301170 , n10759 );
or ( n301205 , n301203 , n10776 );
buf ( n301206 , n301205 );
buf ( n301207 , n301206 );
xor ( n10780 , n301153 , n301207 );
xor ( n10781 , n297601 , n297612 );
xor ( n301210 , n10781 , n297584 );
buf ( n301211 , n301210 );
and ( n10784 , n10780 , n301211 );
and ( n301213 , n301153 , n301207 );
or ( n301214 , n10784 , n301213 );
buf ( n301215 , n301214 );
buf ( n301216 , n301215 );
buf ( n301217 , n780 );
buf ( n301218 , n808 );
xor ( n301219 , n301217 , n301218 );
buf ( n301220 , n301219 );
not ( n301221 , n301220 );
not ( n301222 , n293655 );
or ( n10795 , n301221 , n301222 );
buf ( n301224 , n294557 );
buf ( n301225 , n7211 );
nand ( n301226 , n301224 , n301225 );
buf ( n301227 , n301226 );
nand ( n301228 , n10795 , n301227 );
not ( n301229 , n291788 );
not ( n10802 , n297739 );
or ( n301231 , n301229 , n10802 );
buf ( n10804 , n770 );
buf ( n301233 , n818 );
xor ( n10806 , n10804 , n301233 );
buf ( n301235 , n10806 );
nand ( n10808 , n291984 , n301235 );
nand ( n10809 , n301231 , n10808 );
not ( n301238 , n10809 );
or ( n301239 , n301228 , n301238 );
not ( n301240 , n293058 );
buf ( n301241 , n778 );
buf ( n301242 , n810 );
xor ( n301243 , n301241 , n301242 );
buf ( n301244 , n301243 );
not ( n301245 , n301244 );
or ( n301246 , n301240 , n301245 );
buf ( n301247 , n295259 );
buf ( n301248 , n297655 );
nand ( n301249 , n301247 , n301248 );
buf ( n301250 , n301249 );
nand ( n301251 , n301246 , n301250 );
nand ( n10824 , n301239 , n301251 );
nand ( n301253 , n301228 , n301238 );
nand ( n10826 , n10824 , n301253 );
buf ( n301255 , n10826 );
buf ( n10828 , n297705 );
not ( n301257 , n10828 );
buf ( n301258 , n301257 );
xor ( n10831 , n297727 , n301258 );
xnor ( n301260 , n10831 , n7259 );
buf ( n10833 , n301260 );
xor ( n10834 , n301255 , n10833 );
xor ( n301263 , n297751 , n297758 );
xor ( n301264 , n301263 , n297776 );
buf ( n301265 , n301264 );
and ( n301266 , n10834 , n301265 );
and ( n301267 , n301255 , n10833 );
or ( n10840 , n301266 , n301267 );
buf ( n301269 , n10840 );
buf ( n301270 , n301269 );
xor ( n10843 , n301216 , n301270 );
not ( n301272 , n297850 );
buf ( n301273 , n297833 );
not ( n10846 , n301273 );
and ( n301275 , n301272 , n10846 );
not ( n301276 , n301272 );
and ( n301277 , n301276 , n301273 );
nor ( n10850 , n301275 , n301277 );
buf ( n301279 , n7400 );
and ( n301280 , n10850 , n301279 );
not ( n10853 , n10850 );
not ( n301282 , n301279 );
and ( n10855 , n10853 , n301282 );
nor ( n10856 , n301280 , n10855 );
buf ( n301285 , n10856 );
xor ( n10858 , n10843 , n301285 );
buf ( n301287 , n10858 );
buf ( n10860 , n301287 );
buf ( n301289 , n790 );
buf ( n301290 , n800 );
and ( n301291 , n301289 , n301290 );
buf ( n301292 , n301291 );
buf ( n301293 , n301292 );
buf ( n301294 , n789 );
buf ( n301295 , n800 );
xor ( n301296 , n301294 , n301295 );
buf ( n301297 , n301296 );
buf ( n301298 , n301297 );
not ( n301299 , n301298 );
buf ( n301300 , n299589 );
not ( n10873 , n301300 );
or ( n301302 , n301299 , n10873 );
buf ( n301303 , n6057 );
buf ( n301304 , n301157 );
nand ( n10877 , n301303 , n301304 );
buf ( n301306 , n10877 );
buf ( n301307 , n301306 );
nand ( n10880 , n301302 , n301307 );
buf ( n301309 , n10880 );
buf ( n301310 , n301309 );
xor ( n301311 , n301293 , n301310 );
buf ( n301312 , n777 );
buf ( n301313 , n812 );
xor ( n301314 , n301312 , n301313 );
buf ( n301315 , n301314 );
buf ( n301316 , n301315 );
not ( n301317 , n301316 );
buf ( n301318 , n2373 );
not ( n301319 , n301318 );
or ( n10892 , n301317 , n301319 );
buf ( n301321 , n2383 );
buf ( n301322 , n301189 );
nand ( n10895 , n301321 , n301322 );
buf ( n10896 , n10895 );
buf ( n301325 , n10896 );
nand ( n10898 , n10892 , n301325 );
buf ( n301327 , n10898 );
buf ( n301328 , n301327 );
and ( n10901 , n301311 , n301328 );
and ( n301330 , n301293 , n301310 );
or ( n301331 , n10901 , n301330 );
buf ( n301332 , n301331 );
buf ( n301333 , n301332 );
xor ( n301334 , n802 , n787 );
buf ( n301335 , n301334 );
not ( n301336 , n301335 );
buf ( n301337 , n7960 );
not ( n301338 , n301337 );
or ( n10911 , n301336 , n301338 );
buf ( n301340 , n295929 );
buf ( n301341 , n301174 );
nand ( n301342 , n301340 , n301341 );
buf ( n301343 , n301342 );
buf ( n301344 , n301343 );
nand ( n301345 , n10911 , n301344 );
buf ( n301346 , n301345 );
buf ( n301347 , n301346 );
xor ( n301348 , n804 , n785 );
buf ( n301349 , n301348 );
not ( n301350 , n301349 );
buf ( n10923 , n6010 );
not ( n10924 , n10923 );
or ( n10925 , n301350 , n10924 );
buf ( n10926 , n298526 );
xor ( n301355 , n804 , n784 );
buf ( n10928 , n301355 );
nand ( n10929 , n10926 , n10928 );
buf ( n10930 , n10929 );
buf ( n301359 , n10930 );
nand ( n10932 , n10925 , n301359 );
buf ( n10933 , n10932 );
buf ( n301362 , n10933 );
xor ( n10935 , n301347 , n301362 );
buf ( n301364 , n771 );
buf ( n301365 , n818 );
xor ( n301366 , n301364 , n301365 );
buf ( n301367 , n301366 );
buf ( n301368 , n301367 );
not ( n301369 , n301368 );
buf ( n301370 , n292393 );
not ( n10943 , n301370 );
or ( n301372 , n301369 , n10943 );
buf ( n301373 , n291788 );
buf ( n301374 , n301235 );
nand ( n301375 , n301373 , n301374 );
buf ( n301376 , n301375 );
buf ( n301377 , n301376 );
nand ( n301378 , n301372 , n301377 );
buf ( n301379 , n301378 );
buf ( n301380 , n301379 );
and ( n301381 , n10935 , n301380 );
and ( n301382 , n301347 , n301362 );
or ( n10955 , n301381 , n301382 );
buf ( n301384 , n10955 );
buf ( n10957 , n301384 );
xor ( n10958 , n301333 , n10957 );
buf ( n301387 , n1597 );
not ( n301388 , n301387 );
buf ( n301389 , n1330 );
not ( n301390 , n301389 );
or ( n10963 , n301388 , n301390 );
buf ( n301392 , n822 );
nand ( n301393 , n10963 , n301392 );
buf ( n301394 , n301393 );
buf ( n301395 , n301394 );
not ( n301396 , n301395 );
buf ( n301397 , n301396 );
buf ( n301398 , n301397 );
not ( n10971 , n301398 );
buf ( n301400 , n769 );
buf ( n301401 , n820 );
xor ( n10974 , n301400 , n301401 );
buf ( n10975 , n10974 );
buf ( n301404 , n10975 );
not ( n10977 , n301404 );
buf ( n301406 , n298099 );
not ( n10979 , n301406 );
or ( n301408 , n10977 , n10979 );
buf ( n301409 , n291906 );
buf ( n301410 , n768 );
buf ( n301411 , n820 );
xor ( n301412 , n301410 , n301411 );
buf ( n301413 , n301412 );
buf ( n10986 , n301413 );
nand ( n10987 , n301409 , n10986 );
buf ( n301416 , n10987 );
buf ( n301417 , n301416 );
nand ( n301418 , n301408 , n301417 );
buf ( n301419 , n301418 );
buf ( n301420 , n301419 );
not ( n301421 , n301420 );
buf ( n301422 , n301421 );
buf ( n301423 , n301422 );
not ( n301424 , n301423 );
or ( n10997 , n10971 , n301424 );
buf ( n301426 , n773 );
buf ( n10999 , n816 );
xor ( n11000 , n301426 , n10999 );
buf ( n11001 , n11000 );
buf ( n301430 , n11001 );
not ( n11003 , n301430 );
buf ( n301432 , n2118 );
not ( n11005 , n301432 );
or ( n301434 , n11003 , n11005 );
buf ( n301435 , n1712 );
xor ( n11008 , n816 , n772 );
buf ( n301437 , n11008 );
nand ( n301438 , n301435 , n301437 );
buf ( n301439 , n301438 );
buf ( n301440 , n301439 );
nand ( n11013 , n301434 , n301440 );
buf ( n301442 , n11013 );
buf ( n301443 , n301442 );
nand ( n301444 , n10997 , n301443 );
buf ( n301445 , n301444 );
buf ( n301446 , n301445 );
buf ( n301447 , n301419 );
buf ( n301448 , n301394 );
nand ( n301449 , n301447 , n301448 );
buf ( n301450 , n301449 );
buf ( n301451 , n301450 );
nand ( n301452 , n301446 , n301451 );
buf ( n301453 , n301452 );
buf ( n301454 , n301453 );
and ( n301455 , n10958 , n301454 );
and ( n11028 , n301333 , n10957 );
or ( n301457 , n301455 , n11028 );
buf ( n301458 , n301457 );
buf ( n301459 , n301458 );
not ( n301460 , n301238 );
buf ( n301461 , n789 );
buf ( n301462 , n800 );
and ( n11035 , n301461 , n301462 );
buf ( n301464 , n11035 );
buf ( n11037 , n301464 );
not ( n11038 , n11008 );
not ( n301467 , n2118 );
or ( n11040 , n11038 , n301467 );
nand ( n301469 , n7182 , n1712 );
nand ( n301470 , n11040 , n301469 );
buf ( n301471 , n301470 );
xor ( n301472 , n11037 , n301471 );
buf ( n301473 , n301413 );
not ( n301474 , n301473 );
buf ( n301475 , n298099 );
not ( n301476 , n301475 );
or ( n11049 , n301474 , n301476 );
buf ( n301478 , n291969 );
buf ( n301479 , n820 );
nand ( n11052 , n301478 , n301479 );
buf ( n301481 , n11052 );
buf ( n301482 , n301481 );
nand ( n11055 , n11049 , n301482 );
buf ( n301484 , n11055 );
buf ( n301485 , n301484 );
and ( n301486 , n301472 , n301485 );
and ( n301487 , n11037 , n301471 );
or ( n11060 , n301486 , n301487 );
buf ( n301489 , n11060 );
xor ( n301490 , n301460 , n301489 );
buf ( n301491 , n782 );
buf ( n301492 , n806 );
xor ( n11065 , n301491 , n301492 );
buf ( n301494 , n11065 );
buf ( n301495 , n301494 );
not ( n301496 , n301495 );
buf ( n301497 , n5676 );
not ( n301498 , n301497 );
or ( n11071 , n301496 , n301498 );
buf ( n301500 , n295437 );
buf ( n301501 , n297693 );
nand ( n11074 , n301500 , n301501 );
buf ( n301503 , n11074 );
buf ( n301504 , n301503 );
nand ( n301505 , n11071 , n301504 );
buf ( n301506 , n301505 );
buf ( n301507 , n301506 );
buf ( n301508 , n774 );
buf ( n11081 , n814 );
xor ( n11082 , n301508 , n11081 );
buf ( n301511 , n11082 );
buf ( n301512 , n301511 );
not ( n301513 , n301512 );
buf ( n301514 , n292719 );
not ( n11087 , n301514 );
or ( n301516 , n301513 , n11087 );
buf ( n11089 , n292725 );
buf ( n11090 , n297764 );
nand ( n11091 , n11089 , n11090 );
buf ( n11092 , n11091 );
buf ( n301521 , n11092 );
nand ( n11094 , n301516 , n301521 );
buf ( n11095 , n11094 );
buf ( n301524 , n11095 );
xor ( n11097 , n301507 , n301524 );
buf ( n301526 , n301355 );
not ( n301527 , n301526 );
buf ( n301528 , n296441 );
not ( n11101 , n301528 );
or ( n11102 , n301527 , n11101 );
buf ( n301531 , n296664 );
buf ( n301532 , n297715 );
nand ( n11105 , n301531 , n301532 );
buf ( n301534 , n11105 );
buf ( n301535 , n301534 );
nand ( n301536 , n11102 , n301535 );
buf ( n301537 , n301536 );
buf ( n301538 , n301537 );
and ( n11111 , n11097 , n301538 );
and ( n301540 , n301507 , n301524 );
or ( n11113 , n11111 , n301540 );
buf ( n301542 , n11113 );
xor ( n301543 , n301490 , n301542 );
buf ( n301544 , n301543 );
xor ( n301545 , n301459 , n301544 );
not ( n11118 , n301494 );
not ( n301547 , n295437 );
or ( n301548 , n11118 , n301547 );
xor ( n11121 , n806 , n783 );
not ( n301550 , n5674 );
nand ( n301551 , n11121 , n301550 , n5003 );
nand ( n11124 , n301548 , n301551 );
buf ( n301553 , n11124 );
buf ( n301554 , n775 );
buf ( n301555 , n814 );
xor ( n11128 , n301554 , n301555 );
buf ( n301557 , n11128 );
not ( n301558 , n301557 );
not ( n301559 , n292719 );
or ( n11132 , n301558 , n301559 );
buf ( n301561 , n292725 );
buf ( n301562 , n301511 );
nand ( n301563 , n301561 , n301562 );
buf ( n301564 , n301563 );
nand ( n301565 , n11132 , n301564 );
buf ( n301566 , n301565 );
xor ( n11139 , n301553 , n301566 );
buf ( n301568 , n781 );
buf ( n301569 , n808 );
xor ( n301570 , n301568 , n301569 );
buf ( n301571 , n301570 );
buf ( n11144 , n301571 );
not ( n11145 , n11144 );
buf ( n11146 , n298990 );
not ( n11147 , n11146 );
or ( n11148 , n11145 , n11147 );
buf ( n11149 , n294557 );
buf ( n301578 , n301220 );
nand ( n301579 , n11149 , n301578 );
buf ( n301580 , n301579 );
buf ( n301581 , n301580 );
nand ( n301582 , n11148 , n301581 );
buf ( n301583 , n301582 );
buf ( n301584 , n301583 );
and ( n301585 , n11139 , n301584 );
and ( n11158 , n301553 , n301566 );
or ( n301587 , n301585 , n11158 );
buf ( n301588 , n301587 );
buf ( n301589 , n301588 );
xor ( n11162 , n11037 , n301471 );
xor ( n11163 , n11162 , n301485 );
buf ( n301592 , n11163 );
buf ( n301593 , n301592 );
xor ( n301594 , n301589 , n301593 );
xor ( n11167 , n301507 , n301524 );
xor ( n301596 , n11167 , n301538 );
buf ( n301597 , n301596 );
buf ( n301598 , n301597 );
and ( n301599 , n301594 , n301598 );
and ( n11172 , n301589 , n301593 );
or ( n11173 , n301599 , n11172 );
buf ( n301602 , n11173 );
buf ( n301603 , n301602 );
and ( n301604 , n301545 , n301603 );
and ( n11177 , n301459 , n301544 );
or ( n301606 , n301604 , n11177 );
buf ( n301607 , n301606 );
buf ( n301608 , n301607 );
xor ( n301609 , n297563 , n7139 );
xor ( n301610 , n301609 , n297624 );
buf ( n301611 , n301610 );
buf ( n301612 , n301611 );
not ( n11185 , n301542 );
buf ( n301614 , n301489 );
not ( n11187 , n301614 );
or ( n11188 , n11185 , n11187 );
nor ( n301617 , n301614 , n301542 );
or ( n301618 , n301617 , n301238 );
nand ( n11191 , n11188 , n301618 );
buf ( n301620 , n11191 );
xor ( n11193 , n301612 , n301620 );
xor ( n11194 , n297673 , n297734 );
xor ( n11195 , n11194 , n297788 );
buf ( n301624 , n11195 );
buf ( n301625 , n301624 );
xor ( n11198 , n11193 , n301625 );
buf ( n301627 , n11198 );
buf ( n301628 , n301627 );
xor ( n11201 , n301608 , n301628 );
xor ( n301630 , n301153 , n301207 );
xor ( n301631 , n301630 , n301211 );
buf ( n301632 , n301631 );
buf ( n301633 , n301632 );
not ( n301634 , n301633 );
not ( n11207 , n301251 );
not ( n11208 , n301238 );
or ( n301637 , n11207 , n11208 );
or ( n11210 , n301238 , n301251 );
nand ( n301639 , n301637 , n11210 );
not ( n11212 , n301228 );
and ( n301641 , n301639 , n11212 );
not ( n301642 , n301639 );
and ( n11215 , n301642 , n301228 );
nor ( n301644 , n301641 , n11215 );
xor ( n301645 , n301170 , n10759 );
xor ( n11218 , n301645 , n301202 );
buf ( n301647 , n11218 );
xor ( n11220 , n301644 , n301647 );
buf ( n301649 , n768 );
buf ( n301650 , n822 );
xor ( n11223 , n301649 , n301650 );
buf ( n301652 , n11223 );
buf ( n301653 , n301652 );
not ( n301654 , n301653 );
buf ( n301655 , n292631 );
not ( n301656 , n301655 );
or ( n301657 , n301654 , n301656 );
buf ( n301658 , n292105 );
buf ( n301659 , n822 );
nand ( n301660 , n301658 , n301659 );
buf ( n301661 , n301660 );
buf ( n301662 , n301661 );
nand ( n301663 , n301657 , n301662 );
buf ( n301664 , n301663 );
buf ( n301665 , n301664 );
not ( n301666 , n301665 );
buf ( n301667 , n778 );
buf ( n301668 , n812 );
xor ( n301669 , n301667 , n301668 );
buf ( n301670 , n301669 );
buf ( n301671 , n301670 );
not ( n11244 , n301671 );
buf ( n301673 , n2373 );
not ( n301674 , n301673 );
or ( n11247 , n11244 , n301674 );
buf ( n11248 , n2026 );
buf ( n301677 , n301315 );
nand ( n11250 , n11248 , n301677 );
buf ( n301679 , n11250 );
buf ( n301680 , n301679 );
nand ( n11253 , n11247 , n301680 );
buf ( n301682 , n11253 );
buf ( n301683 , n301682 );
not ( n301684 , n301683 );
or ( n11257 , n301666 , n301684 );
buf ( n301686 , n301682 );
buf ( n301687 , n301664 );
or ( n11260 , n301686 , n301687 );
buf ( n301689 , n790 );
buf ( n301690 , n800 );
xor ( n11263 , n301689 , n301690 );
buf ( n11264 , n11263 );
buf ( n301693 , n11264 );
not ( n11266 , n301693 );
buf ( n301695 , n296480 );
not ( n11268 , n301695 );
or ( n301697 , n11266 , n11268 );
buf ( n301698 , n6057 );
buf ( n301699 , n301297 );
nand ( n11272 , n301698 , n301699 );
buf ( n301701 , n11272 );
buf ( n301702 , n301701 );
nand ( n301703 , n301697 , n301702 );
buf ( n301704 , n301703 );
buf ( n301705 , n301704 );
nand ( n11278 , n11260 , n301705 );
buf ( n301707 , n11278 );
buf ( n301708 , n301707 );
nand ( n11281 , n11257 , n301708 );
buf ( n301710 , n11281 );
buf ( n301711 , n791 );
buf ( n11284 , n800 );
and ( n11285 , n301711 , n11284 );
buf ( n11286 , n11285 );
buf ( n301715 , n11286 );
xor ( n11288 , n810 , n779 );
not ( n301717 , n11288 );
buf ( n301718 , n2410 );
not ( n11291 , n301718 );
or ( n11292 , n301717 , n11291 );
not ( n11293 , n293468 );
not ( n301722 , n2410 );
xor ( n301723 , n810 , n780 );
nand ( n11296 , n11293 , n301722 , n301723 );
nand ( n11297 , n11292 , n11296 );
buf ( n301726 , n11297 );
xor ( n11299 , n301715 , n301726 );
buf ( n301728 , n772 );
buf ( n301729 , n818 );
xor ( n301730 , n301728 , n301729 );
buf ( n301731 , n301730 );
buf ( n301732 , n301731 );
not ( n11305 , n301732 );
buf ( n301734 , n1962 );
not ( n11307 , n301734 );
or ( n11308 , n11305 , n11307 );
buf ( n301737 , n291989 );
buf ( n301738 , n301367 );
nand ( n301739 , n301737 , n301738 );
buf ( n301740 , n301739 );
buf ( n301741 , n301740 );
nand ( n11314 , n11308 , n301741 );
buf ( n301743 , n11314 );
buf ( n301744 , n301743 );
and ( n301745 , n11299 , n301744 );
and ( n301746 , n301715 , n301726 );
or ( n11319 , n301745 , n301746 );
buf ( n301748 , n11319 );
or ( n301749 , n301710 , n301748 );
not ( n11322 , n301749 );
buf ( n301751 , n784 );
buf ( n301752 , n806 );
xor ( n11325 , n301751 , n301752 );
buf ( n11326 , n11325 );
buf ( n301755 , n11326 );
not ( n301756 , n301755 );
buf ( n301757 , n5676 );
not ( n301758 , n301757 );
or ( n11331 , n301756 , n301758 );
buf ( n301760 , n295437 );
buf ( n301761 , n11121 );
nand ( n301762 , n301760 , n301761 );
buf ( n301763 , n301762 );
buf ( n301764 , n301763 );
nand ( n301765 , n11331 , n301764 );
buf ( n301766 , n301765 );
buf ( n301767 , n301766 );
buf ( n301768 , n782 );
buf ( n301769 , n808 );
xor ( n11342 , n301768 , n301769 );
buf ( n11343 , n11342 );
buf ( n301772 , n11343 );
not ( n11345 , n301772 );
buf ( n301774 , n298990 );
not ( n11347 , n301774 );
or ( n11348 , n11345 , n11347 );
buf ( n301777 , n294557 );
buf ( n301778 , n301571 );
nand ( n301779 , n301777 , n301778 );
buf ( n301780 , n301779 );
buf ( n301781 , n301780 );
nand ( n301782 , n11348 , n301781 );
buf ( n301783 , n301782 );
buf ( n301784 , n301783 );
xor ( n301785 , n301767 , n301784 );
xor ( n11358 , n816 , n774 );
buf ( n301787 , n11358 );
not ( n11360 , n301787 );
buf ( n301789 , n2118 );
not ( n301790 , n301789 );
or ( n11363 , n11360 , n301790 );
buf ( n301792 , n296423 );
buf ( n301793 , n11001 );
nand ( n11366 , n301792 , n301793 );
buf ( n301795 , n11366 );
buf ( n301796 , n301795 );
nand ( n301797 , n11363 , n301796 );
buf ( n301798 , n301797 );
buf ( n301799 , n301798 );
and ( n301800 , n301785 , n301799 );
and ( n11373 , n301767 , n301784 );
or ( n301802 , n301800 , n11373 );
buf ( n301803 , n301802 );
not ( n11376 , n301803 );
or ( n301805 , n11322 , n11376 );
buf ( n301806 , n301748 );
buf ( n301807 , n301710 );
nand ( n301808 , n301806 , n301807 );
buf ( n301809 , n301808 );
nand ( n301810 , n301805 , n301809 );
and ( n11383 , n11220 , n301810 );
and ( n11384 , n301644 , n301647 );
or ( n301813 , n11383 , n11384 );
buf ( n301814 , n301813 );
not ( n301815 , n301814 );
or ( n11388 , n301634 , n301815 );
buf ( n301817 , n301632 );
buf ( n301818 , n301813 );
or ( n11391 , n301817 , n301818 );
xor ( n301820 , n301255 , n10833 );
xor ( n301821 , n301820 , n301265 );
buf ( n301822 , n301821 );
buf ( n301823 , n301822 );
nand ( n301824 , n11391 , n301823 );
buf ( n301825 , n301824 );
buf ( n301826 , n301825 );
nand ( n301827 , n11388 , n301826 );
buf ( n301828 , n301827 );
buf ( n301829 , n301828 );
xor ( n11402 , n11201 , n301829 );
buf ( n301831 , n11402 );
buf ( n301832 , n301831 );
xor ( n301833 , n10860 , n301832 );
buf ( n301834 , n770 );
buf ( n301835 , n820 );
xor ( n301836 , n301834 , n301835 );
buf ( n301837 , n301836 );
buf ( n301838 , n301837 );
not ( n301839 , n301838 );
buf ( n301840 , n291722 );
not ( n11413 , n301840 );
or ( n301842 , n301839 , n11413 );
buf ( n301843 , n291906 );
buf ( n301844 , n10975 );
nand ( n301845 , n301843 , n301844 );
buf ( n301846 , n301845 );
buf ( n301847 , n301846 );
nand ( n301848 , n301842 , n301847 );
buf ( n301849 , n301848 );
buf ( n301850 , n301849 );
buf ( n11423 , n11288 );
not ( n11424 , n11423 );
buf ( n11425 , n293058 );
not ( n11426 , n11425 );
or ( n11427 , n11424 , n11426 );
buf ( n11428 , n295259 );
buf ( n301857 , n301244 );
nand ( n301858 , n11428 , n301857 );
buf ( n301859 , n301858 );
buf ( n301860 , n301859 );
nand ( n301861 , n11427 , n301860 );
buf ( n301862 , n301861 );
buf ( n301863 , n301862 );
xor ( n301864 , n301850 , n301863 );
buf ( n301865 , n786 );
buf ( n301866 , n804 );
xor ( n301867 , n301865 , n301866 );
buf ( n301868 , n301867 );
not ( n11441 , n301868 );
not ( n301870 , n298522 );
or ( n11443 , n11441 , n301870 );
buf ( n301872 , n298526 );
buf ( n301873 , n301348 );
nand ( n301874 , n301872 , n301873 );
buf ( n301875 , n301874 );
nand ( n11448 , n11443 , n301875 );
not ( n301877 , n11448 );
buf ( n301878 , n788 );
buf ( n301879 , n802 );
xor ( n301880 , n301878 , n301879 );
buf ( n301881 , n301880 );
not ( n11454 , n301881 );
not ( n301883 , n296508 );
or ( n301884 , n11454 , n301883 );
buf ( n301885 , n296749 );
buf ( n301886 , n301334 );
nand ( n11459 , n301885 , n301886 );
buf ( n301888 , n11459 );
nand ( n11461 , n301884 , n301888 );
not ( n11462 , n11461 );
or ( n301891 , n301877 , n11462 );
buf ( n11464 , n776 );
buf ( n11465 , n814 );
xor ( n11466 , n11464 , n11465 );
buf ( n11467 , n11466 );
buf ( n301896 , n11467 );
not ( n11469 , n301896 );
buf ( n301898 , n292509 );
not ( n301899 , n301898 );
or ( n11472 , n11469 , n301899 );
buf ( n301901 , n5051 );
buf ( n301902 , n301557 );
nand ( n11475 , n301901 , n301902 );
buf ( n301904 , n11475 );
buf ( n301905 , n301904 );
nand ( n11478 , n11472 , n301905 );
buf ( n301907 , n11478 );
buf ( n301908 , n301907 );
not ( n301909 , n301908 );
buf ( n301910 , n301909 );
nor ( n301911 , n11461 , n11448 );
or ( n301912 , n301910 , n301911 );
nand ( n11485 , n301891 , n301912 );
buf ( n301914 , n11485 );
and ( n301915 , n301864 , n301914 );
and ( n301916 , n301850 , n301863 );
or ( n11489 , n301915 , n301916 );
buf ( n301918 , n11489 );
buf ( n301919 , n301918 );
xor ( n301920 , n301333 , n10957 );
xor ( n11493 , n301920 , n301454 );
buf ( n301922 , n11493 );
buf ( n301923 , n301922 );
xor ( n11496 , n301919 , n301923 );
xor ( n11497 , n301347 , n301362 );
xor ( n11498 , n11497 , n301380 );
buf ( n301927 , n11498 );
buf ( n301928 , n301927 );
xor ( n11501 , n301553 , n301566 );
xor ( n11502 , n11501 , n301584 );
buf ( n301931 , n11502 );
buf ( n301932 , n301931 );
xor ( n11505 , n301928 , n301932 );
xor ( n11506 , n301442 , n301397 );
xnor ( n11507 , n11506 , n301419 );
buf ( n301936 , n11507 );
and ( n301937 , n11505 , n301936 );
and ( n11510 , n301928 , n301932 );
or ( n301939 , n301937 , n11510 );
buf ( n301940 , n301939 );
buf ( n301941 , n301940 );
and ( n301942 , n11496 , n301941 );
and ( n301943 , n301919 , n301923 );
or ( n11516 , n301942 , n301943 );
buf ( n301945 , n11516 );
buf ( n301946 , n301945 );
xor ( n11519 , n301459 , n301544 );
xor ( n11520 , n11519 , n301603 );
buf ( n11521 , n11520 );
buf ( n301950 , n11521 );
xor ( n11523 , n301946 , n301950 );
xor ( n11524 , n301589 , n301593 );
xor ( n11525 , n11524 , n301598 );
buf ( n301954 , n11525 );
buf ( n301955 , n301954 );
xor ( n301956 , n301644 , n301647 );
xor ( n11529 , n301956 , n301810 );
buf ( n301958 , n11529 );
xor ( n301959 , n301955 , n301958 );
xor ( n11532 , n301293 , n301310 );
xor ( n301961 , n11532 , n301328 );
buf ( n301962 , n301961 );
buf ( n301963 , n301962 );
xor ( n11536 , n301850 , n301863 );
xor ( n301965 , n11536 , n301914 );
buf ( n301966 , n301965 );
buf ( n301967 , n301966 );
xor ( n301968 , n301963 , n301967 );
buf ( n301969 , n301849 );
not ( n301970 , n301969 );
buf ( n301971 , n301970 );
buf ( n301972 , n301971 );
not ( n301973 , n293902 );
not ( n11546 , n11326 );
or ( n301975 , n301973 , n11546 );
and ( n301976 , n785 , n806 );
not ( n11549 , n785 );
and ( n301978 , n11549 , n300785 );
nor ( n301979 , n301976 , n301978 );
nand ( n11552 , n5680 , n301979 , n294634 );
nand ( n301981 , n301975 , n11552 );
not ( n301982 , n301981 );
buf ( n301983 , n771 );
buf ( n301984 , n820 );
xor ( n301985 , n301983 , n301984 );
buf ( n301986 , n301985 );
buf ( n301987 , n301986 );
not ( n301988 , n301987 );
buf ( n301989 , n291722 );
not ( n11562 , n301989 );
or ( n301991 , n301988 , n11562 );
buf ( n301992 , n291969 );
buf ( n301993 , n301837 );
nand ( n301994 , n301992 , n301993 );
buf ( n301995 , n301994 );
buf ( n301996 , n301995 );
nand ( n301997 , n301991 , n301996 );
buf ( n301998 , n301997 );
not ( n11571 , n301998 );
or ( n302000 , n301982 , n11571 );
not ( n302001 , n301981 );
not ( n11574 , n302001 );
buf ( n302003 , n301998 );
not ( n11576 , n302003 );
buf ( n302005 , n11576 );
not ( n11578 , n302005 );
or ( n11579 , n11574 , n11578 );
buf ( n11580 , n787 );
buf ( n11581 , n804 );
xor ( n11582 , n11580 , n11581 );
buf ( n11583 , n11582 );
buf ( n302012 , n11583 );
not ( n11585 , n302012 );
buf ( n302014 , n295660 );
not ( n302015 , n302014 );
or ( n11588 , n11585 , n302015 );
buf ( n302017 , n295361 );
buf ( n302018 , n301868 );
nand ( n302019 , n302017 , n302018 );
buf ( n302020 , n302019 );
buf ( n302021 , n302020 );
nand ( n11594 , n11588 , n302021 );
buf ( n302023 , n11594 );
nand ( n11596 , n11579 , n302023 );
nand ( n302025 , n302000 , n11596 );
buf ( n302026 , n302025 );
xor ( n302027 , n301972 , n302026 );
buf ( n302028 , n781 );
buf ( n302029 , n810 );
xor ( n302030 , n302028 , n302029 );
buf ( n302031 , n302030 );
buf ( n302032 , n302031 );
not ( n302033 , n302032 );
buf ( n302034 , n293058 );
not ( n11607 , n302034 );
or ( n11608 , n302033 , n11607 );
buf ( n302037 , n292841 );
buf ( n11610 , n301723 );
nand ( n11611 , n302037 , n11610 );
buf ( n302040 , n11611 );
buf ( n302041 , n302040 );
nand ( n302042 , n11608 , n302041 );
buf ( n302043 , n302042 );
buf ( n302044 , n302043 );
buf ( n11617 , n775 );
buf ( n11618 , n816 );
xor ( n11619 , n11617 , n11618 );
buf ( n11620 , n11619 );
buf ( n302049 , n11620 );
not ( n11622 , n302049 );
buf ( n302051 , n292892 );
not ( n302052 , n302051 );
or ( n302053 , n11622 , n302052 );
buf ( n302054 , n296423 );
buf ( n302055 , n11358 );
nand ( n11628 , n302054 , n302055 );
buf ( n302057 , n11628 );
buf ( n302058 , n302057 );
nand ( n302059 , n302053 , n302058 );
buf ( n302060 , n302059 );
buf ( n302061 , n302060 );
xor ( n302062 , n302044 , n302061 );
buf ( n302063 , n298990 );
not ( n302064 , n302063 );
buf ( n302065 , n302064 );
buf ( n302066 , n302065 );
and ( n302067 , n783 , n808 );
not ( n11640 , n783 );
and ( n302069 , n11640 , n294635 );
nor ( n11642 , n302067 , n302069 );
buf ( n302071 , n11642 );
not ( n302072 , n302071 );
buf ( n302073 , n302072 );
buf ( n302074 , n302073 );
or ( n302075 , n302066 , n302074 );
buf ( n302076 , n6301 );
not ( n11649 , n302076 );
buf ( n11650 , n11649 );
buf ( n11651 , n11650 );
buf ( n302080 , n11343 );
not ( n302081 , n302080 );
buf ( n302082 , n302081 );
buf ( n302083 , n302082 );
or ( n11656 , n11651 , n302083 );
nand ( n302085 , n302075 , n11656 );
buf ( n302086 , n302085 );
buf ( n302087 , n302086 );
and ( n302088 , n302062 , n302087 );
and ( n11661 , n302044 , n302061 );
or ( n302090 , n302088 , n11661 );
buf ( n302091 , n302090 );
buf ( n302092 , n302091 );
and ( n302093 , n302027 , n302092 );
and ( n302094 , n301972 , n302026 );
or ( n11667 , n302093 , n302094 );
buf ( n302096 , n11667 );
buf ( n302097 , n302096 );
and ( n11670 , n301968 , n302097 );
and ( n302099 , n301963 , n301967 );
or ( n11672 , n11670 , n302099 );
buf ( n302101 , n11672 );
buf ( n302102 , n302101 );
and ( n302103 , n301959 , n302102 );
and ( n11676 , n301955 , n301958 );
or ( n11677 , n302103 , n11676 );
buf ( n302106 , n11677 );
buf ( n302107 , n302106 );
and ( n11680 , n11523 , n302107 );
and ( n302109 , n301946 , n301950 );
or ( n302110 , n11680 , n302109 );
buf ( n302111 , n302110 );
buf ( n302112 , n302111 );
and ( n11685 , n301833 , n302112 );
and ( n11686 , n10860 , n301832 );
or ( n11687 , n11685 , n11686 );
buf ( n302116 , n11687 );
buf ( n302117 , n302116 );
xor ( n302118 , n301216 , n301270 );
and ( n11691 , n302118 , n301285 );
and ( n11692 , n301216 , n301270 );
or ( n302121 , n11691 , n11692 );
buf ( n302122 , n302121 );
buf ( n302123 , n302122 );
xor ( n302124 , n301608 , n301628 );
and ( n302125 , n302124 , n301829 );
and ( n11698 , n301608 , n301628 );
or ( n302127 , n302125 , n11698 );
buf ( n302128 , n302127 );
buf ( n302129 , n302128 );
xor ( n302130 , n302123 , n302129 );
xor ( n11703 , n297546 , n297629 );
xor ( n302132 , n11703 , n297793 );
buf ( n302133 , n302132 );
buf ( n302134 , n302133 );
xor ( n11707 , n301612 , n301620 );
and ( n11708 , n11707 , n301625 );
and ( n302137 , n301612 , n301620 );
or ( n11710 , n11708 , n302137 );
buf ( n302139 , n11710 );
buf ( n302140 , n302139 );
xor ( n302141 , n302134 , n302140 );
buf ( n302142 , n297802 );
not ( n11715 , n302142 );
and ( n302144 , n297817 , n297854 );
not ( n302145 , n297817 );
not ( n302146 , n297854 );
and ( n11719 , n302145 , n302146 );
nor ( n302148 , n302144 , n11719 );
buf ( n302149 , n302148 );
not ( n11722 , n302149 );
or ( n302151 , n11715 , n11722 );
buf ( n302152 , n302148 );
buf ( n302153 , n297802 );
or ( n302154 , n302152 , n302153 );
nand ( n302155 , n302151 , n302154 );
buf ( n302156 , n302155 );
buf ( n302157 , n302156 );
xor ( n302158 , n302141 , n302157 );
buf ( n302159 , n302158 );
buf ( n302160 , n302159 );
xor ( n11733 , n302130 , n302160 );
buf ( n302162 , n11733 );
buf ( n302163 , n302162 );
and ( n11736 , n302117 , n302163 );
buf ( n302165 , n11736 );
not ( n302166 , n302165 );
or ( n11739 , n301149 , n302166 );
buf ( n302168 , n831 );
not ( n302169 , n302168 );
buf ( n302170 , n302116 );
buf ( n302171 , n302162 );
and ( n302172 , n302170 , n302171 );
buf ( n302173 , n302172 );
buf ( n302174 , n302173 );
nand ( n11747 , n302169 , n302174 );
buf ( n302176 , n11747 );
nand ( n302177 , n11739 , n302176 );
buf ( n11750 , n302177 );
xor ( n302179 , n297373 , n297402 );
and ( n302180 , n302179 , n297419 );
and ( n302181 , n297373 , n297402 );
or ( n302182 , n302180 , n302181 );
buf ( n302183 , n302182 );
buf ( n302184 , n302183 );
buf ( n302185 , n297415 );
not ( n11758 , n297328 );
not ( n302187 , n6920 );
or ( n302188 , n11758 , n302187 );
nand ( n11761 , n297354 , n6882 );
nand ( n11762 , n302188 , n11761 );
buf ( n302191 , n11762 );
xor ( n302192 , n302185 , n302191 );
xor ( n302193 , n297437 , n297454 );
and ( n11766 , n302193 , n297472 );
and ( n302195 , n297437 , n297454 );
or ( n302196 , n11766 , n302195 );
buf ( n302197 , n302196 );
buf ( n302198 , n302197 );
xor ( n11771 , n302192 , n302198 );
buf ( n302200 , n11771 );
buf ( n11773 , n302200 );
xor ( n11774 , n302184 , n11773 );
xor ( n302203 , n296723 , n296781 );
and ( n302204 , n302203 , n296831 );
and ( n11777 , n296723 , n296781 );
or ( n11778 , n302204 , n11777 );
buf ( n302207 , n11778 );
buf ( n302208 , n302207 );
xor ( n11781 , n11774 , n302208 );
buf ( n302210 , n11781 );
xor ( n11783 , n297309 , n297477 );
and ( n302212 , n11783 , n297523 );
and ( n11785 , n297309 , n297477 );
or ( n302214 , n302212 , n11785 );
buf ( n302215 , n302214 );
xor ( n302216 , n302210 , n302215 );
not ( n11789 , n6994 );
not ( n11790 , n7047 );
or ( n11791 , n11789 , n11790 );
nand ( n302220 , n11791 , n297356 );
not ( n302221 , n6994 );
nand ( n302222 , n302221 , n297474 );
nand ( n11795 , n302220 , n302222 );
buf ( n302224 , n11795 );
and ( n302225 , n296766 , n296767 );
buf ( n302226 , n302225 );
buf ( n302227 , n302226 );
buf ( n302228 , n297339 );
not ( n302229 , n302228 );
buf ( n302230 , n296480 );
not ( n302231 , n302230 );
or ( n302232 , n302229 , n302231 );
buf ( n302233 , n6057 );
buf ( n11806 , n800 );
buf ( n302235 , n780 );
xor ( n302236 , n11806 , n302235 );
buf ( n302237 , n302236 );
buf ( n302238 , n302237 );
nand ( n11811 , n302233 , n302238 );
buf ( n302240 , n11811 );
buf ( n302241 , n302240 );
nand ( n302242 , n302232 , n302241 );
buf ( n302243 , n302242 );
buf ( n302244 , n302243 );
xor ( n302245 , n302227 , n302244 );
buf ( n302246 , n297441 );
not ( n302247 , n302246 );
buf ( n302248 , n296617 );
not ( n11821 , n302248 );
or ( n302250 , n302247 , n11821 );
buf ( n302251 , n295437 );
xor ( n302252 , n806 , n774 );
buf ( n302253 , n302252 );
nand ( n11826 , n302251 , n302253 );
buf ( n302255 , n11826 );
buf ( n302256 , n302255 );
nand ( n302257 , n302250 , n302256 );
buf ( n302258 , n302257 );
buf ( n302259 , n302258 );
xor ( n302260 , n302245 , n302259 );
buf ( n302261 , n302260 );
buf ( n302262 , n302261 );
buf ( n302263 , n297322 );
not ( n11836 , n302263 );
buf ( n302265 , n296594 );
not ( n11838 , n302265 );
or ( n11839 , n11836 , n11838 );
buf ( n302268 , n294557 );
xor ( n11841 , n808 , n772 );
buf ( n302270 , n11841 );
nand ( n11843 , n302268 , n302270 );
buf ( n302272 , n11843 );
buf ( n302273 , n302272 );
nand ( n302274 , n11839 , n302273 );
buf ( n302275 , n302274 );
buf ( n11848 , n2089 );
not ( n302277 , n11848 );
buf ( n302278 , n302277 );
buf ( n302279 , n302278 );
not ( n11852 , n302279 );
buf ( n302281 , n2892 );
not ( n302282 , n302281 );
or ( n11855 , n11852 , n302282 );
buf ( n302284 , n814 );
nand ( n11857 , n11855 , n302284 );
buf ( n302286 , n11857 );
xor ( n11859 , n302275 , n302286 );
buf ( n302288 , n7002 );
not ( n11861 , n302288 );
buf ( n302290 , n2376 );
not ( n302291 , n302290 );
or ( n302292 , n11861 , n302291 );
buf ( n302293 , n2383 );
xor ( n11866 , n812 , n768 );
buf ( n302295 , n11866 );
nand ( n302296 , n302293 , n302295 );
buf ( n302297 , n302296 );
buf ( n302298 , n302297 );
nand ( n302299 , n302292 , n302298 );
buf ( n302300 , n302299 );
xor ( n302301 , n11859 , n302300 );
buf ( n302302 , n302301 );
xor ( n11875 , n302262 , n302302 );
buf ( n11876 , n297366 );
not ( n11877 , n11876 );
buf ( n11878 , n296508 );
not ( n11879 , n11878 );
or ( n11880 , n11877 , n11879 );
buf ( n302309 , n296749 );
buf ( n302310 , n802 );
buf ( n302311 , n778 );
xor ( n302312 , n302310 , n302311 );
buf ( n302313 , n302312 );
buf ( n302314 , n302313 );
nand ( n11887 , n302309 , n302314 );
buf ( n302316 , n11887 );
buf ( n302317 , n302316 );
nand ( n302318 , n11880 , n302317 );
buf ( n302319 , n302318 );
buf ( n302320 , n302319 );
buf ( n302321 , n297465 );
not ( n302322 , n302321 );
buf ( n302323 , n293058 );
not ( n302324 , n302323 );
or ( n302325 , n302322 , n302324 );
buf ( n302326 , n295259 );
buf ( n302327 , n770 );
buf ( n302328 , n810 );
xor ( n302329 , n302327 , n302328 );
buf ( n302330 , n302329 );
buf ( n302331 , n302330 );
nand ( n302332 , n302326 , n302331 );
buf ( n302333 , n302332 );
buf ( n302334 , n302333 );
nand ( n302335 , n302325 , n302334 );
buf ( n302336 , n302335 );
buf ( n11909 , n302336 );
xor ( n11910 , n302320 , n11909 );
buf ( n302339 , n296441 );
not ( n302340 , n302339 );
buf ( n302341 , n302340 );
buf ( n302342 , n302341 );
buf ( n302343 , n297392 );
or ( n11916 , n302342 , n302343 );
not ( n302345 , n296446 );
buf ( n302346 , n302345 );
buf ( n302347 , n804 );
buf ( n302348 , n776 );
xnor ( n302349 , n302347 , n302348 );
buf ( n302350 , n302349 );
buf ( n302351 , n302350 );
or ( n302352 , n302346 , n302351 );
nand ( n11925 , n11916 , n302352 );
buf ( n302354 , n11925 );
buf ( n302355 , n302354 );
xor ( n11928 , n11910 , n302355 );
buf ( n302357 , n11928 );
buf ( n302358 , n302357 );
xor ( n11931 , n11875 , n302358 );
buf ( n302360 , n11931 );
buf ( n302361 , n302360 );
xor ( n11934 , n302224 , n302361 );
xor ( n302363 , n296565 , n296716 );
and ( n302364 , n302363 , n296834 );
and ( n302365 , n296565 , n296716 );
or ( n11938 , n302364 , n302365 );
buf ( n302367 , n11938 );
buf ( n302368 , n302367 );
xor ( n11941 , n11934 , n302368 );
buf ( n302370 , n11941 );
xor ( n302371 , n302216 , n302370 );
not ( n302372 , n302371 );
xor ( n11945 , n296837 , n297302 );
and ( n302374 , n11945 , n297526 );
and ( n302375 , n296837 , n297302 );
or ( n11948 , n302374 , n302375 );
buf ( n302377 , n11948 );
not ( n302378 , n302377 );
nor ( n11951 , n302372 , n302378 );
and ( n302380 , n831 , n11951 );
not ( n302381 , n831 );
buf ( n302382 , n302377 );
buf ( n302383 , n302371 );
and ( n11956 , n302382 , n302383 );
buf ( n302385 , n11956 );
and ( n302386 , n302381 , n302385 );
or ( n11959 , n302380 , n302386 );
buf ( n302388 , n11959 );
xor ( n11961 , n301813 , n301822 );
xor ( n302390 , n11961 , n301632 );
buf ( n302391 , n302390 );
xor ( n11964 , n301919 , n301923 );
xor ( n302393 , n11964 , n301941 );
buf ( n302394 , n302393 );
buf ( n302395 , n302394 );
xor ( n11968 , n301715 , n301726 );
xor ( n302397 , n11968 , n301744 );
buf ( n302398 , n302397 );
buf ( n302399 , n302398 );
buf ( n11972 , n789 );
buf ( n302401 , n802 );
xor ( n302402 , n11972 , n302401 );
buf ( n302403 , n302402 );
buf ( n302404 , n302403 );
not ( n302405 , n302404 );
buf ( n302406 , n7960 );
not ( n302407 , n302406 );
or ( n11980 , n302405 , n302407 );
buf ( n302409 , n296517 );
buf ( n302410 , n301881 );
nand ( n11983 , n302409 , n302410 );
buf ( n302412 , n11983 );
buf ( n302413 , n302412 );
nand ( n11986 , n11980 , n302413 );
buf ( n302415 , n11986 );
buf ( n302416 , n302415 );
buf ( n302417 , n791 );
buf ( n302418 , n800 );
xor ( n302419 , n302417 , n302418 );
buf ( n302420 , n302419 );
buf ( n302421 , n302420 );
not ( n302422 , n302421 );
buf ( n302423 , n6049 );
not ( n11996 , n302423 );
or ( n11997 , n302422 , n11996 );
buf ( n302426 , n6057 );
buf ( n302427 , n11264 );
nand ( n12000 , n302426 , n302427 );
buf ( n302429 , n12000 );
buf ( n302430 , n302429 );
nand ( n302431 , n11997 , n302430 );
buf ( n302432 , n302431 );
buf ( n302433 , n302432 );
xor ( n12006 , n302416 , n302433 );
buf ( n302435 , n777 );
buf ( n302436 , n814 );
xor ( n12009 , n302435 , n302436 );
buf ( n302438 , n12009 );
buf ( n302439 , n302438 );
not ( n12012 , n302439 );
buf ( n302441 , n292509 );
not ( n302442 , n302441 );
or ( n12015 , n12012 , n302442 );
buf ( n302444 , n5051 );
buf ( n302445 , n11467 );
nand ( n302446 , n302444 , n302445 );
buf ( n302447 , n302446 );
buf ( n302448 , n302447 );
nand ( n12021 , n12015 , n302448 );
buf ( n302450 , n12021 );
buf ( n302451 , n302450 );
and ( n302452 , n12006 , n302451 );
and ( n12025 , n302416 , n302433 );
or ( n302454 , n302452 , n12025 );
buf ( n302455 , n302454 );
buf ( n302456 , n302455 );
xor ( n302457 , n302399 , n302456 );
buf ( n302458 , n769 );
buf ( n302459 , n822 );
xor ( n302460 , n302458 , n302459 );
buf ( n302461 , n302460 );
buf ( n302462 , n302461 );
not ( n12035 , n302462 );
buf ( n302464 , n291761 );
not ( n302465 , n302464 );
or ( n302466 , n12035 , n302465 );
buf ( n302467 , n1600 );
buf ( n302468 , n301652 );
nand ( n302469 , n302467 , n302468 );
buf ( n302470 , n302469 );
buf ( n302471 , n302470 );
nand ( n302472 , n302466 , n302471 );
buf ( n302473 , n302472 );
buf ( n302474 , n302473 );
or ( n12047 , n292870 , n7526 );
nand ( n302476 , n12047 , n824 );
buf ( n302477 , n302476 );
xor ( n12050 , n302474 , n302477 );
buf ( n302479 , n773 );
buf ( n302480 , n818 );
xor ( n302481 , n302479 , n302480 );
buf ( n302482 , n302481 );
buf ( n302483 , n302482 );
not ( n12056 , n302483 );
buf ( n302485 , n297104 );
not ( n12058 , n302485 );
buf ( n302487 , n12058 );
buf ( n302488 , n302487 );
not ( n302489 , n302488 );
or ( n12062 , n12056 , n302489 );
not ( n302491 , n297099 );
buf ( n302492 , n302491 );
buf ( n302493 , n301731 );
nand ( n302494 , n302492 , n302493 );
buf ( n302495 , n302494 );
buf ( n302496 , n302495 );
nand ( n302497 , n12062 , n302496 );
buf ( n302498 , n302497 );
buf ( n302499 , n302498 );
and ( n302500 , n12050 , n302499 );
and ( n12073 , n302474 , n302477 );
or ( n12074 , n302500 , n12073 );
buf ( n302503 , n12074 );
buf ( n302504 , n302503 );
and ( n302505 , n302457 , n302504 );
and ( n12078 , n302399 , n302456 );
or ( n302507 , n302505 , n12078 );
buf ( n302508 , n302507 );
buf ( n302509 , n302508 );
not ( n12082 , n301710 );
xor ( n302511 , n301748 , n12082 );
xnor ( n12084 , n302511 , n301803 );
buf ( n302513 , n12084 );
xor ( n302514 , n302509 , n302513 );
xor ( n302515 , n301767 , n301784 );
xor ( n12088 , n302515 , n301799 );
buf ( n302517 , n12088 );
buf ( n302518 , n302517 );
and ( n12091 , n11448 , n301910 );
not ( n302520 , n11448 );
and ( n302521 , n302520 , n301907 );
or ( n12094 , n12091 , n302521 );
and ( n12095 , n12094 , n11461 );
not ( n302524 , n12094 );
not ( n302525 , n11461 );
and ( n12098 , n302524 , n302525 );
nor ( n302527 , n12095 , n12098 );
buf ( n302528 , n302527 );
xor ( n302529 , n302518 , n302528 );
xor ( n12102 , n301664 , n301682 );
xor ( n12103 , n12102 , n301704 );
buf ( n12104 , n12103 );
and ( n12105 , n302529 , n12104 );
and ( n12106 , n302518 , n302528 );
or ( n12107 , n12105 , n12106 );
buf ( n12108 , n12107 );
buf ( n302537 , n12108 );
and ( n12110 , n302514 , n302537 );
and ( n302539 , n302509 , n302513 );
or ( n302540 , n12110 , n302539 );
buf ( n302541 , n302540 );
buf ( n302542 , n302541 );
xor ( n302543 , n302395 , n302542 );
xor ( n12116 , n301928 , n301932 );
xor ( n302545 , n12116 , n301936 );
buf ( n302546 , n302545 );
buf ( n302547 , n302546 );
xor ( n302548 , n301963 , n301967 );
xor ( n302549 , n302548 , n302097 );
buf ( n302550 , n302549 );
buf ( n302551 , n302550 );
xor ( n302552 , n302547 , n302551 );
buf ( n12125 , n792 );
buf ( n12126 , n800 );
nand ( n12127 , n12125 , n12126 );
buf ( n12128 , n12127 );
buf ( n302557 , n12128 );
not ( n12130 , n302557 );
buf ( n302559 , n779 );
buf ( n302560 , n812 );
xor ( n12133 , n302559 , n302560 );
buf ( n302562 , n12133 );
buf ( n302563 , n302562 );
not ( n12136 , n302563 );
buf ( n302565 , n2373 );
not ( n12138 , n302565 );
or ( n302567 , n12136 , n12138 );
buf ( n302568 , n2026 );
buf ( n302569 , n301670 );
nand ( n302570 , n302568 , n302569 );
buf ( n302571 , n302570 );
buf ( n302572 , n302571 );
nand ( n12145 , n302567 , n302572 );
buf ( n12146 , n12145 );
buf ( n12147 , n12146 );
not ( n302576 , n12147 );
buf ( n302577 , n302576 );
buf ( n302578 , n302577 );
not ( n302579 , n302578 );
or ( n12152 , n12130 , n302579 );
buf ( n302581 , n300804 );
not ( n302582 , n302581 );
buf ( n302583 , n291761 );
not ( n12156 , n302583 );
or ( n302585 , n302582 , n12156 );
buf ( n302586 , n1600 );
buf ( n302587 , n302461 );
nand ( n12160 , n302586 , n302587 );
buf ( n302589 , n12160 );
buf ( n302590 , n302589 );
nand ( n302591 , n302585 , n302590 );
buf ( n302592 , n302591 );
buf ( n302593 , n302592 );
nand ( n12166 , n12152 , n302593 );
buf ( n302595 , n12166 );
buf ( n12168 , n302595 );
buf ( n302597 , n12128 );
not ( n12170 , n302597 );
buf ( n12171 , n12146 );
nand ( n12172 , n12170 , n12171 );
buf ( n302601 , n12172 );
buf ( n302602 , n302601 );
nand ( n302603 , n12168 , n302602 );
buf ( n302604 , n302603 );
buf ( n302605 , n302604 );
not ( n12178 , n301979 );
not ( n12179 , n8642 );
or ( n302608 , n12178 , n12179 );
not ( n302609 , n296103 );
nand ( n12182 , n302609 , n300787 , n301550 );
nand ( n12183 , n302608 , n12182 );
not ( n302612 , n12183 );
not ( n302613 , n300693 );
not ( n12186 , n298522 );
or ( n12187 , n302613 , n12186 );
buf ( n302616 , n298526 );
buf ( n302617 , n11583 );
nand ( n12190 , n302616 , n302617 );
buf ( n302619 , n12190 );
nand ( n302620 , n12187 , n302619 );
not ( n302621 , n302620 );
or ( n12194 , n302612 , n302621 );
buf ( n302623 , n12183 );
buf ( n302624 , n302620 );
nor ( n12197 , n302623 , n302624 );
buf ( n302626 , n12197 );
and ( n12199 , n300710 , n292892 );
and ( n302628 , n296423 , n11620 );
nor ( n12201 , n12199 , n302628 );
or ( n302630 , n302626 , n12201 );
nand ( n302631 , n12194 , n302630 );
buf ( n302632 , n302631 );
not ( n302633 , n10300 );
not ( n12206 , n7960 );
or ( n302635 , n302633 , n12206 );
buf ( n302636 , n296517 );
buf ( n302637 , n302403 );
nand ( n12210 , n302636 , n302637 );
buf ( n302639 , n12210 );
nand ( n302640 , n302635 , n302639 );
buf ( n302641 , n302640 );
not ( n12214 , n302641 );
buf ( n302643 , n300639 );
not ( n12216 , n302643 );
buf ( n302645 , n291838 );
not ( n12218 , n302645 );
or ( n12219 , n12216 , n12218 );
buf ( n302648 , n1613 );
buf ( n302649 , n824 );
nand ( n12222 , n302648 , n302649 );
buf ( n302651 , n12222 );
buf ( n302652 , n302651 );
nand ( n302653 , n12219 , n302652 );
buf ( n302654 , n302653 );
buf ( n302655 , n302654 );
not ( n302656 , n302655 );
or ( n302657 , n12214 , n302656 );
or ( n302658 , n302654 , n302640 );
buf ( n302659 , n300622 );
not ( n302660 , n302659 );
buf ( n302661 , n292509 );
not ( n12234 , n302661 );
or ( n302663 , n302660 , n12234 );
buf ( n302664 , n292725 );
buf ( n302665 , n302438 );
nand ( n12238 , n302664 , n302665 );
buf ( n302667 , n12238 );
buf ( n302668 , n302667 );
nand ( n302669 , n302663 , n302668 );
buf ( n302670 , n302669 );
nand ( n302671 , n302658 , n302670 );
buf ( n302672 , n302671 );
nand ( n12245 , n302657 , n302672 );
buf ( n302674 , n12245 );
buf ( n302675 , n302674 );
xor ( n12248 , n302632 , n302675 );
buf ( n302677 , n300767 );
not ( n12250 , n302677 );
buf ( n302679 , n293655 );
not ( n12252 , n302679 );
or ( n302681 , n12250 , n12252 );
not ( n12254 , n809 );
not ( n12255 , n293537 );
or ( n12256 , n12254 , n12255 );
nand ( n302685 , n12256 , n293541 );
nand ( n302686 , n11642 , n302685 );
buf ( n302687 , n302686 );
nand ( n12260 , n302681 , n302687 );
buf ( n302689 , n12260 );
buf ( n302690 , n302689 );
buf ( n302691 , n300548 );
not ( n12264 , n302691 );
buf ( n302693 , n293058 );
not ( n302694 , n302693 );
or ( n302695 , n12264 , n302694 );
buf ( n302696 , n292841 );
buf ( n302697 , n302031 );
nand ( n302698 , n302696 , n302697 );
buf ( n302699 , n302698 );
buf ( n302700 , n302699 );
nand ( n302701 , n302695 , n302700 );
buf ( n302702 , n302701 );
buf ( n302703 , n302702 );
xor ( n302704 , n302690 , n302703 );
buf ( n302705 , n300566 );
not ( n302706 , n302705 );
buf ( n302707 , n302487 );
not ( n302708 , n302707 );
or ( n12281 , n302706 , n302708 );
buf ( n302710 , n302491 );
buf ( n302711 , n302482 );
nand ( n302712 , n302710 , n302711 );
buf ( n302713 , n302712 );
buf ( n302714 , n302713 );
nand ( n302715 , n12281 , n302714 );
buf ( n302716 , n302715 );
buf ( n302717 , n302716 );
and ( n302718 , n302704 , n302717 );
and ( n302719 , n302690 , n302703 );
or ( n12292 , n302718 , n302719 );
buf ( n302721 , n12292 );
buf ( n302722 , n302721 );
and ( n12295 , n12248 , n302722 );
and ( n302724 , n302632 , n302675 );
or ( n302725 , n12295 , n302724 );
buf ( n302726 , n302725 );
buf ( n302727 , n302726 );
xor ( n12300 , n302605 , n302727 );
xor ( n12301 , n301972 , n302026 );
xor ( n12302 , n12301 , n302092 );
buf ( n302731 , n12302 );
buf ( n302732 , n302731 );
and ( n302733 , n12300 , n302732 );
and ( n12306 , n302605 , n302727 );
or ( n302735 , n302733 , n12306 );
buf ( n302736 , n302735 );
buf ( n302737 , n302736 );
and ( n302738 , n302552 , n302737 );
and ( n12311 , n302547 , n302551 );
or ( n302740 , n302738 , n12311 );
buf ( n302741 , n302740 );
buf ( n302742 , n302741 );
and ( n302743 , n302543 , n302742 );
and ( n302744 , n302395 , n302542 );
or ( n12317 , n302743 , n302744 );
buf ( n302746 , n12317 );
buf ( n302747 , n302746 );
xor ( n12320 , n302391 , n302747 );
xor ( n302749 , n301946 , n301950 );
xor ( n302750 , n302749 , n302107 );
buf ( n302751 , n302750 );
buf ( n302752 , n302751 );
xor ( n12325 , n12320 , n302752 );
buf ( n302754 , n12325 );
buf ( n302755 , n302754 );
xor ( n302756 , n301955 , n301958 );
xor ( n12329 , n302756 , n302102 );
buf ( n302758 , n12329 );
buf ( n302759 , n302758 );
buf ( n12332 , n12128 );
buf ( n302761 , n12146 );
xor ( n302762 , n12332 , n302761 );
buf ( n302763 , n302592 );
not ( n12336 , n302763 );
buf ( n302765 , n12336 );
buf ( n302766 , n302765 );
xnor ( n12339 , n302762 , n302766 );
buf ( n12340 , n12339 );
buf ( n302769 , n12340 );
not ( n302770 , n302769 );
xor ( n302771 , n302416 , n302433 );
xor ( n12344 , n302771 , n302451 );
buf ( n302773 , n12344 );
not ( n302774 , n302773 );
buf ( n302775 , n302774 );
not ( n302776 , n302775 );
or ( n302777 , n302770 , n302776 );
and ( n12350 , n302023 , n302001 );
not ( n12351 , n302023 );
and ( n12352 , n12351 , n301981 );
or ( n302781 , n12350 , n12352 );
and ( n302782 , n302781 , n302005 );
not ( n12355 , n302781 );
and ( n12356 , n12355 , n301998 );
nor ( n12357 , n302782 , n12356 );
buf ( n302786 , n12357 );
not ( n12359 , n302786 );
buf ( n302788 , n12359 );
buf ( n302789 , n302788 );
nand ( n302790 , n302777 , n302789 );
buf ( n302791 , n302790 );
buf ( n302792 , n302791 );
buf ( n302793 , n302774 );
not ( n12366 , n302793 );
buf ( n302795 , n12340 );
not ( n12368 , n302795 );
buf ( n302797 , n12368 );
buf ( n302798 , n302797 );
nand ( n302799 , n12366 , n302798 );
buf ( n302800 , n302799 );
buf ( n302801 , n302800 );
nand ( n302802 , n302792 , n302801 );
buf ( n302803 , n302802 );
buf ( n302804 , n302803 );
xor ( n302805 , n302399 , n302456 );
xor ( n12378 , n302805 , n302504 );
buf ( n302807 , n12378 );
buf ( n302808 , n302807 );
xor ( n302809 , n302804 , n302808 );
buf ( n302810 , n793 );
buf ( n302811 , n800 );
and ( n302812 , n302810 , n302811 );
buf ( n302813 , n302812 );
buf ( n302814 , n302813 );
buf ( n302815 , n300611 );
not ( n12388 , n302815 );
buf ( n302817 , n6049 );
not ( n12390 , n302817 );
or ( n12391 , n12388 , n12390 );
buf ( n302820 , n6057 );
buf ( n302821 , n302420 );
nand ( n302822 , n302820 , n302821 );
buf ( n302823 , n302822 );
buf ( n302824 , n302823 );
nand ( n302825 , n12391 , n302824 );
buf ( n302826 , n302825 );
buf ( n302827 , n302826 );
xor ( n302828 , n302814 , n302827 );
buf ( n302829 , n300660 );
not ( n302830 , n302829 );
buf ( n302831 , n298099 );
not ( n12404 , n302831 );
or ( n302833 , n302830 , n12404 );
buf ( n302834 , n291906 );
buf ( n302835 , n301986 );
nand ( n12408 , n302834 , n302835 );
buf ( n12409 , n12408 );
buf ( n302838 , n12409 );
nand ( n12411 , n302833 , n302838 );
buf ( n302840 , n12411 );
buf ( n302841 , n302840 );
and ( n12414 , n302828 , n302841 );
and ( n302843 , n302814 , n302827 );
or ( n12416 , n12414 , n302843 );
buf ( n302845 , n12416 );
buf ( n302846 , n302845 );
xor ( n12419 , n302474 , n302477 );
xor ( n302848 , n12419 , n302499 );
buf ( n302849 , n302848 );
buf ( n302850 , n302849 );
xor ( n12423 , n302846 , n302850 );
xor ( n12424 , n302044 , n302061 );
xor ( n302853 , n12424 , n302087 );
buf ( n302854 , n302853 );
buf ( n302855 , n302854 );
and ( n302856 , n12423 , n302855 );
and ( n302857 , n302846 , n302850 );
or ( n12430 , n302856 , n302857 );
buf ( n302859 , n12430 );
buf ( n302860 , n302859 );
and ( n302861 , n302809 , n302860 );
and ( n302862 , n302804 , n302808 );
or ( n12435 , n302861 , n302862 );
buf ( n302864 , n12435 );
buf ( n302865 , n302864 );
xor ( n302866 , n302509 , n302513 );
xor ( n12439 , n302866 , n302537 );
buf ( n302868 , n12439 );
buf ( n302869 , n302868 );
xor ( n12442 , n302865 , n302869 );
xor ( n302871 , n302518 , n302528 );
xor ( n302872 , n302871 , n12104 );
buf ( n302873 , n302872 );
buf ( n302874 , n302873 );
buf ( n302875 , n300530 );
not ( n12448 , n302875 );
buf ( n302877 , n2376 );
not ( n12450 , n302877 );
or ( n12451 , n12448 , n12450 );
buf ( n302880 , n2383 );
buf ( n302881 , n302562 );
nand ( n302882 , n302880 , n302881 );
buf ( n302883 , n302882 );
buf ( n302884 , n302883 );
nand ( n302885 , n12451 , n302884 );
buf ( n302886 , n302885 );
buf ( n302887 , n302886 );
buf ( n302888 , n302765 );
xor ( n302889 , n302887 , n302888 );
xor ( n302890 , n300700 , n300717 );
and ( n12463 , n302890 , n300735 );
and ( n302892 , n300700 , n300717 );
or ( n12465 , n12463 , n302892 );
buf ( n302894 , n12465 );
buf ( n302895 , n302894 );
and ( n12468 , n302889 , n302895 );
and ( n12469 , n302887 , n302888 );
or ( n302898 , n12468 , n12469 );
buf ( n302899 , n302898 );
buf ( n302900 , n302899 );
not ( n12473 , n300672 );
not ( n302902 , n10238 );
or ( n12475 , n12473 , n302902 );
buf ( n12476 , n10238 );
buf ( n302905 , n300672 );
nor ( n302906 , n12476 , n302905 );
buf ( n302907 , n302906 );
or ( n12480 , n300648 , n302907 );
nand ( n302909 , n12475 , n12480 );
buf ( n302910 , n302909 );
xor ( n12483 , n300538 , n300555 );
and ( n302912 , n12483 , n300573 );
and ( n12485 , n300538 , n300555 );
or ( n302914 , n302912 , n12485 );
buf ( n302915 , n302914 );
buf ( n302916 , n302915 );
xor ( n302917 , n302910 , n302916 );
not ( n12490 , n300773 );
not ( n302919 , n300810 );
or ( n302920 , n12490 , n302919 );
not ( n12493 , n300813 );
not ( n302922 , n300776 );
or ( n12495 , n12493 , n302922 );
nand ( n302924 , n12495 , n300793 );
nand ( n12497 , n302920 , n302924 );
buf ( n302926 , n12497 );
and ( n12499 , n302917 , n302926 );
and ( n12500 , n302910 , n302916 );
or ( n302929 , n12499 , n12500 );
buf ( n302930 , n302929 );
buf ( n302931 , n302930 );
xor ( n302932 , n302900 , n302931 );
xor ( n302933 , n302632 , n302675 );
xor ( n302934 , n302933 , n302722 );
buf ( n302935 , n302934 );
buf ( n302936 , n302935 );
and ( n302937 , n302932 , n302936 );
and ( n12510 , n302900 , n302931 );
or ( n302939 , n302937 , n12510 );
buf ( n302940 , n302939 );
buf ( n302941 , n302940 );
xor ( n12514 , n302874 , n302941 );
xor ( n12515 , n302605 , n302727 );
xor ( n12516 , n12515 , n302732 );
buf ( n302945 , n12516 );
buf ( n302946 , n302945 );
and ( n302947 , n12514 , n302946 );
and ( n12520 , n302874 , n302941 );
or ( n302949 , n302947 , n12520 );
buf ( n302950 , n302949 );
buf ( n302951 , n302950 );
and ( n302952 , n12442 , n302951 );
and ( n12525 , n302865 , n302869 );
or ( n12526 , n302952 , n12525 );
buf ( n302955 , n12526 );
buf ( n302956 , n302955 );
xor ( n302957 , n302759 , n302956 );
xor ( n302958 , n302395 , n302542 );
xor ( n302959 , n302958 , n302742 );
buf ( n302960 , n302959 );
buf ( n302961 , n302960 );
and ( n302962 , n302957 , n302961 );
and ( n302963 , n302759 , n302956 );
or ( n12536 , n302962 , n302963 );
buf ( n302965 , n12536 );
buf ( n302966 , n302965 );
and ( n12539 , n302755 , n302966 );
buf ( n302968 , n12539 );
nand ( n12541 , n302968 , n831 );
buf ( n302970 , n831 );
not ( n302971 , n302970 );
buf ( n302972 , n302965 );
buf ( n302973 , n302754 );
and ( n12546 , n302972 , n302973 );
buf ( n302975 , n12546 );
buf ( n302976 , n302975 );
nand ( n302977 , n302971 , n302976 );
buf ( n302978 , n302977 );
nand ( n12551 , n12541 , n302978 );
buf ( n302980 , n12551 );
xor ( n302981 , n302547 , n302551 );
xor ( n302982 , n302981 , n302737 );
buf ( n302983 , n302982 );
buf ( n302984 , n302983 );
xor ( n302985 , n302865 , n302869 );
xor ( n12558 , n302985 , n302951 );
buf ( n302987 , n12558 );
buf ( n302988 , n302987 );
xor ( n12561 , n302984 , n302988 );
xor ( n12562 , n300601 , n10189 );
and ( n12563 , n12562 , n10199 );
and ( n12564 , n300601 , n10189 );
or ( n302993 , n12563 , n12564 );
buf ( n302994 , n302993 );
xor ( n12567 , n302814 , n302827 );
xor ( n12568 , n12567 , n302841 );
buf ( n12569 , n12568 );
buf ( n302998 , n12569 );
xor ( n12571 , n302994 , n302998 );
xor ( n12572 , n302690 , n302703 );
xor ( n12573 , n12572 , n302717 );
buf ( n303002 , n12573 );
buf ( n303003 , n303002 );
and ( n12576 , n12571 , n303003 );
and ( n12577 , n302994 , n302998 );
or ( n12578 , n12576 , n12577 );
buf ( n303007 , n12578 );
buf ( n303008 , n302774 );
not ( n303009 , n303008 );
buf ( n303010 , n302788 );
not ( n303011 , n303010 );
or ( n12584 , n303009 , n303011 );
buf ( n303013 , n302773 );
buf ( n303014 , n12357 );
nand ( n12587 , n303013 , n303014 );
buf ( n12588 , n12587 );
buf ( n303017 , n12588 );
nand ( n303018 , n12584 , n303017 );
buf ( n303019 , n303018 );
and ( n303020 , n303019 , n302797 );
not ( n12593 , n303019 );
and ( n12594 , n12593 , n12340 );
nor ( n12595 , n303020 , n12594 );
xor ( n12596 , n303007 , n12595 );
xor ( n12597 , n302846 , n302850 );
xor ( n12598 , n12597 , n302855 );
buf ( n303027 , n12598 );
and ( n303028 , n12596 , n303027 );
and ( n12601 , n303007 , n12595 );
or ( n12602 , n303028 , n12601 );
buf ( n303031 , n12602 );
xor ( n12604 , n302804 , n302808 );
xor ( n303033 , n12604 , n302860 );
buf ( n303034 , n303033 );
buf ( n303035 , n303034 );
xor ( n12608 , n303031 , n303035 );
not ( n12609 , n12201 );
not ( n12610 , n302620 );
not ( n303039 , n12183 );
and ( n12612 , n12610 , n303039 );
and ( n303041 , n12183 , n302620 );
nor ( n303042 , n12612 , n303041 );
not ( n12615 , n303042 );
or ( n12616 , n12609 , n12615 );
or ( n12617 , n303042 , n12201 );
nand ( n12618 , n12616 , n12617 );
buf ( n303047 , n12618 );
buf ( n303048 , n302670 );
not ( n12621 , n303048 );
buf ( n303050 , n302640 );
not ( n12623 , n303050 );
buf ( n303052 , n12623 );
buf ( n303053 , n303052 );
not ( n303054 , n303053 );
and ( n303055 , n12621 , n303054 );
buf ( n303056 , n302670 );
buf ( n303057 , n303052 );
and ( n303058 , n303056 , n303057 );
nor ( n12631 , n303055 , n303058 );
buf ( n303060 , n12631 );
buf ( n12633 , n303060 );
buf ( n303062 , n302654 );
xnor ( n12635 , n12633 , n303062 );
buf ( n12636 , n12635 );
buf ( n303065 , n12636 );
xor ( n12638 , n303047 , n303065 );
xor ( n303067 , n302887 , n302888 );
xor ( n12640 , n303067 , n302895 );
buf ( n303069 , n12640 );
buf ( n303070 , n303069 );
and ( n303071 , n12638 , n303070 );
and ( n12644 , n303047 , n303065 );
or ( n303073 , n303071 , n12644 );
buf ( n303074 , n303073 );
buf ( n303075 , n303074 );
xor ( n12648 , n300514 , n10092 );
and ( n12649 , n12648 , n300575 );
and ( n12650 , n300514 , n10092 );
or ( n303079 , n12649 , n12650 );
xor ( n12652 , n300469 , n300475 );
and ( n303081 , n12652 , n300491 );
and ( n12654 , n300469 , n300475 );
or ( n303083 , n303081 , n12654 );
buf ( n303084 , n303083 );
xor ( n303085 , n303079 , n303084 );
xor ( n303086 , n302910 , n302916 );
xor ( n12659 , n303086 , n302926 );
buf ( n303088 , n12659 );
and ( n303089 , n303085 , n303088 );
and ( n12662 , n303079 , n303084 );
or ( n303091 , n303089 , n12662 );
buf ( n303092 , n303091 );
xor ( n303093 , n303075 , n303092 );
xor ( n303094 , n302900 , n302931 );
xor ( n12667 , n303094 , n302936 );
buf ( n303096 , n12667 );
buf ( n303097 , n303096 );
and ( n12670 , n303093 , n303097 );
and ( n303099 , n303075 , n303092 );
or ( n12672 , n12670 , n303099 );
buf ( n303101 , n12672 );
buf ( n303102 , n303101 );
and ( n12675 , n12608 , n303102 );
and ( n303104 , n303031 , n303035 );
or ( n303105 , n12675 , n303104 );
buf ( n303106 , n303105 );
buf ( n303107 , n303106 );
and ( n303108 , n12561 , n303107 );
and ( n303109 , n302984 , n302988 );
or ( n12682 , n303108 , n303109 );
buf ( n303111 , n12682 );
buf ( n303112 , n303111 );
xor ( n12685 , n302759 , n302956 );
xor ( n303114 , n12685 , n302961 );
buf ( n303115 , n303114 );
buf ( n303116 , n303115 );
and ( n12689 , n303112 , n303116 );
buf ( n303118 , n12689 );
and ( n12691 , n831 , n303118 );
not ( n12692 , n831 );
buf ( n303121 , n303115 );
buf ( n303122 , n303111 );
and ( n12695 , n303121 , n303122 );
buf ( n303124 , n12695 );
and ( n12697 , n12692 , n303124 );
or ( n12698 , n12691 , n12697 );
buf ( n12699 , n12698 );
buf ( n303128 , n831 );
not ( n303129 , n303128 );
not ( n12702 , n5437 );
not ( n12703 , n12702 );
not ( n303132 , n5441 );
or ( n303133 , n12703 , n303132 );
or ( n12706 , n12702 , n5441 );
nand ( n303135 , n303133 , n12706 );
buf ( n303136 , n303135 );
buf ( n12709 , n5449 );
buf ( n303138 , n12709 );
and ( n12711 , n303136 , n303138 );
not ( n12712 , n303136 );
buf ( n303141 , n5449 );
not ( n12714 , n303141 );
buf ( n303143 , n12714 );
buf ( n12716 , n303143 );
and ( n12717 , n12712 , n12716 );
nor ( n303146 , n12711 , n12717 );
buf ( n303147 , n303146 );
buf ( n303148 , n303147 );
xor ( n303149 , n294587 , n4266 );
and ( n303150 , n303149 , n294709 );
and ( n12723 , n294587 , n4266 );
or ( n12724 , n303150 , n12723 );
buf ( n303153 , n12724 );
xor ( n12726 , n303148 , n303153 );
buf ( n303155 , n295205 );
not ( n303156 , n303155 );
buf ( n303157 , n303156 );
and ( n12730 , n4766 , n303157 );
not ( n12731 , n4766 );
and ( n12732 , n12731 , n295205 );
nor ( n12733 , n12730 , n12732 );
buf ( n303162 , n295189 );
not ( n303163 , n303162 );
buf ( n303164 , n303163 );
and ( n303165 , n12733 , n303164 );
not ( n12738 , n12733 );
and ( n303167 , n12738 , n295189 );
nor ( n303168 , n303165 , n303167 );
buf ( n303169 , n303168 );
and ( n12742 , n12726 , n303169 );
and ( n303171 , n303148 , n303153 );
or ( n12744 , n12742 , n303171 );
buf ( n303173 , n12744 );
xor ( n303174 , n836 , n303173 );
and ( n303175 , n4779 , n5269 );
not ( n12748 , n4779 );
and ( n12749 , n12748 , n5477 );
nor ( n303178 , n303175 , n12749 );
not ( n303179 , n5473 );
and ( n12752 , n303178 , n303179 );
not ( n303181 , n303178 );
and ( n303182 , n303181 , n5473 );
nor ( n12755 , n12752 , n303182 );
and ( n12756 , n303174 , n12755 );
and ( n12757 , n836 , n303173 );
or ( n12758 , n12756 , n12757 );
buf ( n303187 , n12758 );
not ( n303188 , n303187 );
or ( n303189 , n303129 , n303188 );
buf ( n303190 , n831 );
not ( n12763 , n303190 );
buf ( n303192 , n868 );
buf ( n303193 , n303173 );
xor ( n303194 , n303192 , n303193 );
buf ( n303195 , n12755 );
and ( n12768 , n303194 , n303195 );
and ( n303197 , n303192 , n303193 );
or ( n12770 , n12768 , n303197 );
buf ( n303199 , n12770 );
buf ( n303200 , n303199 );
nand ( n12773 , n12763 , n303200 );
buf ( n303202 , n12773 );
buf ( n303203 , n303202 );
nand ( n303204 , n303189 , n303203 );
buf ( n303205 , n303204 );
buf ( n12778 , n303205 );
buf ( n12779 , n295136 );
buf ( n303208 , n855 );
xor ( n12781 , n295082 , n295095 );
xor ( n12782 , n12781 , n295112 );
not ( n12783 , n12782 );
xor ( n12784 , n294810 , n294825 );
not ( n12785 , n12784 );
buf ( n12786 , n1613 );
buf ( n303215 , n799 );
and ( n303216 , n12786 , n303215 );
buf ( n303217 , n303216 );
buf ( n303218 , n303217 );
buf ( n303219 , n794 );
buf ( n303220 , n830 );
xor ( n303221 , n303219 , n303220 );
buf ( n303222 , n303221 );
buf ( n303223 , n303222 );
not ( n303224 , n303223 );
buf ( n303225 , n291656 );
not ( n12798 , n303225 );
or ( n303227 , n303224 , n12798 );
buf ( n303228 , n294797 );
buf ( n303229 , n831 );
nand ( n303230 , n303228 , n303229 );
buf ( n303231 , n303230 );
buf ( n303232 , n303231 );
nand ( n303233 , n303227 , n303232 );
buf ( n303234 , n303233 );
buf ( n303235 , n303234 );
xor ( n12808 , n303218 , n303235 );
buf ( n303237 , n796 );
buf ( n303238 , n828 );
xor ( n12811 , n303237 , n303238 );
buf ( n303240 , n12811 );
buf ( n303241 , n303240 );
not ( n12814 , n303241 );
buf ( n303243 , n291808 );
not ( n303244 , n303243 );
or ( n12817 , n12814 , n303244 );
buf ( n303246 , n291939 );
buf ( n303247 , n295100 );
nand ( n303248 , n303246 , n303247 );
buf ( n303249 , n303248 );
buf ( n303250 , n303249 );
nand ( n303251 , n12817 , n303250 );
buf ( n303252 , n303251 );
buf ( n303253 , n303252 );
and ( n303254 , n12808 , n303253 );
and ( n303255 , n303218 , n303235 );
or ( n12828 , n303254 , n303255 );
buf ( n303257 , n12828 );
not ( n303258 , n303257 );
nand ( n12831 , n12785 , n303258 );
not ( n303260 , n12831 );
or ( n303261 , n12783 , n303260 );
nand ( n12834 , n303257 , n12784 );
nand ( n303263 , n303261 , n12834 );
buf ( n303264 , n303263 );
xor ( n12837 , n303208 , n303264 );
nand ( n12838 , n295118 , n4687 , n4693 );
not ( n12839 , n295118 );
not ( n303268 , n4687 );
nand ( n303269 , n12839 , n4693 , n303268 );
not ( n12842 , n295118 );
not ( n303271 , n4693 );
nand ( n303272 , n12842 , n303271 , n4687 );
nand ( n12845 , n303271 , n295118 , n303268 );
nand ( n303274 , n12838 , n303269 , n303272 , n12845 );
buf ( n303275 , n303274 );
and ( n12848 , n12837 , n303275 );
and ( n303277 , n303208 , n303264 );
or ( n303278 , n12848 , n303277 );
buf ( n303279 , n303278 );
buf ( n303280 , n303279 );
buf ( n303281 , n858 );
buf ( n303282 , n1580 );
buf ( n303283 , n799 );
and ( n303284 , n303282 , n303283 );
buf ( n303285 , n303284 );
buf ( n303286 , n303285 );
xor ( n303287 , n830 , n796 );
buf ( n303288 , n303287 );
not ( n12861 , n303288 );
buf ( n303290 , n291656 );
not ( n303291 , n303290 );
or ( n12864 , n12861 , n303291 );
buf ( n303293 , n795 );
buf ( n303294 , n830 );
xor ( n303295 , n303293 , n303294 );
buf ( n303296 , n303295 );
buf ( n303297 , n303296 );
buf ( n303298 , n831 );
nand ( n12871 , n303297 , n303298 );
buf ( n303300 , n12871 );
buf ( n303301 , n303300 );
nand ( n303302 , n12864 , n303301 );
buf ( n303303 , n303302 );
buf ( n303304 , n303303 );
xor ( n303305 , n303286 , n303304 );
buf ( n303306 , n828 );
buf ( n303307 , n798 );
xor ( n303308 , n303306 , n303307 );
buf ( n303309 , n303308 );
buf ( n303310 , n303309 );
not ( n303311 , n303310 );
buf ( n303312 , n291808 );
not ( n303313 , n303312 );
or ( n12886 , n303311 , n303313 );
buf ( n12887 , n291939 );
buf ( n303316 , n828 );
buf ( n303317 , n797 );
xor ( n303318 , n303316 , n303317 );
buf ( n303319 , n303318 );
buf ( n303320 , n303319 );
nand ( n303321 , n12887 , n303320 );
buf ( n303322 , n303321 );
buf ( n303323 , n303322 );
nand ( n12896 , n12886 , n303323 );
buf ( n12897 , n12896 );
buf ( n303326 , n12897 );
and ( n12899 , n303305 , n303326 );
and ( n303328 , n303286 , n303304 );
or ( n303329 , n12899 , n303328 );
buf ( n303330 , n303329 );
buf ( n303331 , n303330 );
xor ( n303332 , n303281 , n303331 );
buf ( n303333 , n799 );
buf ( n303334 , n827 );
or ( n303335 , n303333 , n303334 );
buf ( n303336 , n828 );
nand ( n303337 , n303335 , n303336 );
buf ( n303338 , n303337 );
buf ( n303339 , n303338 );
buf ( n303340 , n799 );
buf ( n303341 , n827 );
nand ( n303342 , n303340 , n303341 );
buf ( n303343 , n303342 );
buf ( n303344 , n303343 );
buf ( n303345 , n826 );
and ( n12918 , n303339 , n303344 , n303345 );
buf ( n303347 , n12918 );
buf ( n12920 , n303347 );
buf ( n303349 , n303296 );
not ( n12922 , n303349 );
buf ( n303351 , n291656 );
not ( n303352 , n303351 );
or ( n12925 , n12922 , n303352 );
buf ( n303354 , n303222 );
buf ( n303355 , n831 );
nand ( n12928 , n303354 , n303355 );
buf ( n12929 , n12928 );
buf ( n303358 , n12929 );
nand ( n12931 , n12925 , n303358 );
buf ( n303360 , n12931 );
buf ( n303361 , n303360 );
xor ( n303362 , n12920 , n303361 );
buf ( n303363 , n303362 );
buf ( n303364 , n303363 );
buf ( n12937 , n799 );
buf ( n12938 , n826 );
xor ( n12939 , n12937 , n12938 );
buf ( n12940 , n12939 );
buf ( n303369 , n12940 );
not ( n12942 , n303369 );
buf ( n303371 , n1453 );
not ( n12944 , n303371 );
or ( n303373 , n12942 , n12944 );
buf ( n303374 , n1580 );
buf ( n303375 , n826 );
buf ( n303376 , n798 );
xor ( n303377 , n303375 , n303376 );
buf ( n303378 , n303377 );
buf ( n303379 , n303378 );
nand ( n303380 , n303374 , n303379 );
buf ( n303381 , n303380 );
buf ( n303382 , n303381 );
nand ( n303383 , n303373 , n303382 );
buf ( n303384 , n303383 );
buf ( n303385 , n303384 );
xor ( n12958 , n303364 , n303385 );
buf ( n303387 , n303319 );
not ( n12960 , n303387 );
buf ( n303389 , n291808 );
not ( n303390 , n303389 );
or ( n12963 , n12960 , n303390 );
buf ( n303392 , n291939 );
buf ( n303393 , n303240 );
nand ( n12966 , n303392 , n303393 );
buf ( n303395 , n12966 );
buf ( n303396 , n303395 );
nand ( n12969 , n12963 , n303396 );
buf ( n303398 , n12969 );
buf ( n303399 , n303398 );
xor ( n12972 , n12958 , n303399 );
buf ( n303401 , n12972 );
buf ( n303402 , n303401 );
and ( n12975 , n303332 , n303402 );
and ( n303404 , n303281 , n303331 );
or ( n303405 , n12975 , n303404 );
buf ( n303406 , n303405 );
buf ( n303407 , n303406 );
buf ( n12980 , n301129 );
buf ( n303409 , n839 );
xor ( n12982 , n296383 , n296389 );
and ( n12983 , n12982 , n296394 );
and ( n303412 , n296383 , n296389 );
or ( n303413 , n12983 , n303412 );
buf ( n303414 , n303413 );
buf ( n303415 , n303414 );
xor ( n12988 , n303409 , n303415 );
xor ( n12989 , n294080 , n294277 );
xor ( n12990 , n12989 , n294310 );
buf ( n303419 , n12990 );
xor ( n12992 , n12988 , n303419 );
buf ( n303421 , n12992 );
buf ( n12994 , n303421 );
buf ( n303423 , n844 );
xor ( n303424 , n298296 , n7880 );
xnor ( n303425 , n303424 , n7888 );
buf ( n303426 , n303425 );
xor ( n12999 , n301080 , n10667 );
and ( n303428 , n12999 , n301109 );
and ( n303429 , n301080 , n10667 );
or ( n13002 , n303428 , n303429 );
buf ( n303431 , n13002 );
buf ( n303432 , n303431 );
buf ( n303433 , n10612 );
not ( n303434 , n303433 );
buf ( n303435 , n301055 );
not ( n303436 , n303435 );
or ( n303437 , n303434 , n303436 );
buf ( n303438 , n301062 );
nand ( n303439 , n303437 , n303438 );
buf ( n303440 , n303439 );
buf ( n303441 , n303440 );
buf ( n303442 , n10612 );
not ( n303443 , n303442 );
buf ( n13016 , n301058 );
nand ( n13017 , n303443 , n13016 );
buf ( n13018 , n13017 );
buf ( n13019 , n13018 );
nand ( n13020 , n303441 , n13019 );
buf ( n13021 , n13020 );
buf ( n303450 , n13021 );
xor ( n13023 , n303432 , n303450 );
xor ( n303452 , n298053 , n298115 );
xor ( n13025 , n303452 , n298171 );
buf ( n303454 , n13025 );
buf ( n303455 , n303454 );
and ( n303456 , n13023 , n303455 );
and ( n303457 , n303432 , n303450 );
or ( n13030 , n303456 , n303457 );
buf ( n303459 , n13030 );
buf ( n303460 , n303459 );
xor ( n13033 , n303426 , n303460 );
xor ( n13034 , n298175 , n7804 );
xor ( n303463 , n13034 , n298282 );
buf ( n303464 , n303463 );
and ( n303465 , n13033 , n303464 );
and ( n13038 , n303426 , n303460 );
or ( n13039 , n303465 , n13038 );
buf ( n303468 , n13039 );
buf ( n303469 , n303468 );
xor ( n303470 , n303423 , n303469 );
xor ( n13043 , n298000 , n298286 );
xor ( n303472 , n13043 , n298334 );
buf ( n303473 , n303472 );
buf ( n303474 , n303473 );
xor ( n303475 , n303470 , n303474 );
buf ( n303476 , n303475 );
buf ( n303477 , n303476 );
xor ( n13050 , n7834 , n298251 );
buf ( n303479 , n13050 );
buf ( n303480 , n298276 );
and ( n303481 , n303479 , n303480 );
not ( n13054 , n303479 );
buf ( n303483 , n298276 );
not ( n303484 , n303483 );
buf ( n303485 , n303484 );
buf ( n303486 , n303485 );
and ( n13059 , n13054 , n303486 );
nor ( n303488 , n303481 , n13059 );
buf ( n303489 , n303488 );
buf ( n303490 , n303489 );
xor ( n303491 , n303432 , n303450 );
xor ( n303492 , n303491 , n303455 );
buf ( n303493 , n303492 );
buf ( n303494 , n303493 );
xor ( n303495 , n303490 , n303494 );
xor ( n303496 , n301077 , n301112 );
and ( n13069 , n303496 , n301119 );
and ( n303498 , n301077 , n301112 );
or ( n13071 , n13069 , n303498 );
buf ( n303500 , n13071 );
buf ( n303501 , n303500 );
and ( n303502 , n303495 , n303501 );
and ( n303503 , n303490 , n303494 );
or ( n13076 , n303502 , n303503 );
buf ( n303505 , n13076 );
xor ( n303506 , n845 , n303505 );
xor ( n13079 , n303426 , n303460 );
xor ( n303508 , n13079 , n303464 );
buf ( n303509 , n303508 );
xor ( n13082 , n303506 , n303509 );
buf ( n303511 , n13082 );
xor ( n303512 , n300860 , n301037 );
xor ( n13085 , n303512 , n301125 );
buf ( n303514 , n13085 );
buf ( n303515 , n303514 );
buf ( n303516 , n850 );
xor ( n303517 , n292083 , n292089 );
xor ( n13090 , n303517 , n292124 );
buf ( n303519 , n13090 );
buf ( n303520 , n303519 );
xor ( n13093 , n294968 , n294981 );
and ( n303522 , n13093 , n294995 );
and ( n13095 , n294968 , n294981 );
or ( n13096 , n303522 , n13095 );
buf ( n303525 , n13096 );
buf ( n303526 , n303525 );
xor ( n303527 , n295020 , n295033 );
and ( n303528 , n303527 , n295047 );
and ( n13101 , n295020 , n295033 );
or ( n303530 , n303528 , n13101 );
buf ( n303531 , n303530 );
buf ( n303532 , n303531 );
xor ( n303533 , n303526 , n303532 );
xor ( n13106 , n292102 , n292110 );
xor ( n303535 , n13106 , n1692 );
buf ( n13108 , n303535 );
and ( n13109 , n303533 , n13108 );
and ( n303538 , n303526 , n303532 );
or ( n303539 , n13109 , n303538 );
buf ( n303540 , n303539 );
buf ( n303541 , n303540 );
xor ( n303542 , n303520 , n303541 );
xor ( n13115 , n291864 , n291868 );
xor ( n13116 , n13115 , n291958 );
buf ( n303545 , n13116 );
buf ( n303546 , n303545 );
and ( n13119 , n303542 , n303546 );
and ( n303548 , n303520 , n303541 );
or ( n13121 , n13119 , n303548 );
buf ( n303550 , n13121 );
buf ( n303551 , n303550 );
xor ( n13124 , n303516 , n303551 );
xor ( n303553 , n291860 , n291963 );
xor ( n303554 , n303553 , n292132 );
buf ( n303555 , n303554 );
buf ( n303556 , n303555 );
xor ( n13129 , n13124 , n303556 );
buf ( n303558 , n13129 );
buf ( n13131 , n303558 );
xor ( n303560 , n294738 , n294954 );
xor ( n303561 , n303560 , n295052 );
buf ( n303562 , n303561 );
buf ( n13135 , n303562 );
xor ( n13136 , n295070 , n295125 );
xor ( n13137 , n13136 , n295132 );
buf ( n303566 , n13137 );
buf ( n303567 , n303566 );
xor ( n13140 , n303208 , n303264 );
xor ( n303569 , n13140 , n303275 );
buf ( n303570 , n303569 );
buf ( n13143 , n303570 );
buf ( n303572 , n10413 );
not ( n303573 , n9991 );
not ( n303574 , n303573 );
not ( n303575 , n300425 );
or ( n13148 , n303574 , n303575 );
nand ( n303577 , n13148 , n10005 );
not ( n13150 , n10002 );
and ( n303579 , n303577 , n13150 );
not ( n303580 , n303577 );
and ( n13153 , n303580 , n10002 );
nor ( n303582 , n303579 , n13153 );
buf ( n13155 , n303582 );
xor ( n303584 , n299837 , n299841 );
xor ( n13157 , n303584 , n299846 );
buf ( n303586 , n13157 );
buf ( n303587 , n303586 );
and ( n13160 , n299826 , n299812 );
not ( n303589 , n299826 );
and ( n13162 , n299803 , n299806 );
not ( n303591 , n299803 );
and ( n13164 , n303591 , n299809 );
nor ( n303593 , n13162 , n13164 );
and ( n303594 , n303589 , n303593 );
nor ( n13167 , n13160 , n303594 );
buf ( n13168 , n299815 );
not ( n303597 , n13168 );
and ( n13170 , n13167 , n303597 );
not ( n303599 , n13167 );
and ( n303600 , n303599 , n13168 );
nor ( n13173 , n13170 , n303600 );
buf ( n303602 , n13173 );
xor ( n303603 , n303587 , n303602 );
xor ( n13176 , n299866 , n299883 );
xor ( n13177 , n13176 , n299920 );
buf ( n303606 , n13177 );
buf ( n303607 , n303606 );
xor ( n13180 , n299485 , n299506 );
xor ( n303609 , n13180 , n299525 );
buf ( n303610 , n303609 );
buf ( n303611 , n303610 );
xor ( n303612 , n303607 , n303611 );
buf ( n303613 , n778 );
buf ( n303614 , n822 );
xor ( n303615 , n303613 , n303614 );
buf ( n303616 , n303615 );
not ( n13189 , n303616 );
not ( n303618 , n4031 );
or ( n303619 , n13189 , n303618 );
buf ( n303620 , n1600 );
buf ( n303621 , n300184 );
nand ( n303622 , n303620 , n303621 );
buf ( n303623 , n303622 );
nand ( n13196 , n303619 , n303623 );
not ( n13197 , n13196 );
buf ( n303626 , n788 );
buf ( n303627 , n812 );
xor ( n303628 , n303626 , n303627 );
buf ( n303629 , n303628 );
buf ( n303630 , n303629 );
not ( n303631 , n303630 );
buf ( n303632 , n3539 );
not ( n13205 , n303632 );
or ( n303634 , n303631 , n13205 );
buf ( n303635 , n292810 );
buf ( n303636 , n300053 );
nand ( n303637 , n303635 , n303636 );
buf ( n303638 , n303637 );
buf ( n303639 , n303638 );
nand ( n13212 , n303634 , n303639 );
buf ( n303641 , n13212 );
not ( n13214 , n303641 );
or ( n303643 , n13197 , n13214 );
not ( n303644 , n13196 );
not ( n13217 , n303644 );
not ( n303646 , n303641 );
not ( n303647 , n303646 );
or ( n13220 , n13217 , n303647 );
buf ( n303649 , n790 );
buf ( n303650 , n810 );
xor ( n13223 , n303649 , n303650 );
buf ( n13224 , n13223 );
buf ( n303653 , n13224 );
not ( n13226 , n303653 );
buf ( n303655 , n293058 );
not ( n303656 , n303655 );
or ( n13229 , n13226 , n303656 );
buf ( n303658 , n292841 );
buf ( n303659 , n9642 );
nand ( n13232 , n303658 , n303659 );
buf ( n303661 , n13232 );
buf ( n303662 , n303661 );
nand ( n13235 , n13229 , n303662 );
buf ( n13236 , n13235 );
nand ( n303665 , n13220 , n13236 );
nand ( n303666 , n303643 , n303665 );
not ( n13239 , n303666 );
buf ( n303668 , n782 );
buf ( n303669 , n818 );
xor ( n13242 , n303668 , n303669 );
buf ( n13243 , n13242 );
buf ( n303672 , n13243 );
not ( n303673 , n303672 );
nor ( n303674 , n2996 , n1961 );
buf ( n303675 , n303674 );
not ( n303676 , n303675 );
or ( n303677 , n303673 , n303676 );
buf ( n303678 , n1357 );
buf ( n303679 , n299976 );
nand ( n303680 , n303678 , n303679 );
buf ( n303681 , n303680 );
buf ( n303682 , n303681 );
nand ( n303683 , n303677 , n303682 );
buf ( n303684 , n303683 );
buf ( n303685 , n303684 );
xor ( n13258 , n796 , n804 );
buf ( n303687 , n13258 );
not ( n303688 , n303687 );
buf ( n303689 , n295983 );
not ( n303690 , n303689 );
or ( n13263 , n303688 , n303690 );
buf ( n303692 , n5554 );
buf ( n303693 , n299993 );
nand ( n13266 , n303692 , n303693 );
buf ( n303695 , n13266 );
buf ( n303696 , n303695 );
nand ( n13269 , n13263 , n303696 );
buf ( n13270 , n13269 );
buf ( n303699 , n13270 );
xor ( n13272 , n303685 , n303699 );
buf ( n303701 , n794 );
buf ( n303702 , n806 );
xor ( n13275 , n303701 , n303702 );
buf ( n13276 , n13275 );
buf ( n303705 , n13276 );
not ( n13278 , n303705 );
buf ( n303707 , n294637 );
not ( n13280 , n303707 );
or ( n13281 , n13278 , n13280 );
buf ( n303710 , n295437 );
buf ( n303711 , n299942 );
nand ( n13284 , n303710 , n303711 );
buf ( n303713 , n13284 );
buf ( n303714 , n303713 );
nand ( n13287 , n13281 , n303714 );
buf ( n303716 , n13287 );
buf ( n303717 , n303716 );
and ( n13290 , n13272 , n303717 );
and ( n303719 , n303685 , n303699 );
or ( n303720 , n13290 , n303719 );
buf ( n303721 , n303720 );
buf ( n303722 , n303721 );
not ( n13295 , n303722 );
buf ( n303724 , n13295 );
nand ( n13297 , n13239 , n303724 );
not ( n303726 , n13297 );
xor ( n13299 , n808 , n792 );
not ( n13300 , n13299 );
not ( n13301 , n4983 );
or ( n13302 , n13300 , n13301 );
buf ( n303731 , n3114 );
buf ( n303732 , n299929 );
nand ( n13305 , n303731 , n303732 );
buf ( n303734 , n13305 );
nand ( n13307 , n13302 , n303734 );
buf ( n303736 , n13307 );
buf ( n13309 , n780 );
buf ( n303738 , n820 );
xor ( n13311 , n13309 , n303738 );
buf ( n303740 , n13311 );
buf ( n303741 , n303740 );
not ( n13314 , n303741 );
buf ( n303743 , n298099 );
not ( n303744 , n303743 );
or ( n303745 , n13314 , n303744 );
buf ( n303746 , n1995 );
buf ( n303747 , n299958 );
nand ( n303748 , n303746 , n303747 );
buf ( n303749 , n303748 );
buf ( n303750 , n303749 );
nand ( n303751 , n303745 , n303750 );
buf ( n303752 , n303751 );
buf ( n303753 , n303752 );
xor ( n303754 , n303736 , n303753 );
buf ( n303755 , n774 );
buf ( n303756 , n826 );
xor ( n303757 , n303755 , n303756 );
buf ( n303758 , n303757 );
buf ( n303759 , n303758 );
not ( n303760 , n303759 );
buf ( n303761 , n291880 );
not ( n303762 , n303761 );
or ( n13335 , n303760 , n303762 );
buf ( n303764 , n291886 );
buf ( n13337 , n9609 );
nand ( n13338 , n303764 , n13337 );
buf ( n13339 , n13338 );
buf ( n13340 , n13339 );
nand ( n13341 , n13335 , n13340 );
buf ( n13342 , n13341 );
buf ( n303771 , n13342 );
and ( n13344 , n303754 , n303771 );
and ( n303773 , n303736 , n303753 );
or ( n303774 , n13344 , n303773 );
buf ( n303775 , n303774 );
not ( n303776 , n303775 );
or ( n303777 , n303726 , n303776 );
nand ( n13350 , n303721 , n303666 );
nand ( n303779 , n303777 , n13350 );
buf ( n303780 , n303779 );
and ( n303781 , n303612 , n303780 );
and ( n303782 , n303607 , n303611 );
or ( n303783 , n303781 , n303782 );
buf ( n303784 , n303783 );
buf ( n303785 , n303784 );
and ( n303786 , n303603 , n303785 );
and ( n303787 , n303587 , n303602 );
or ( n13360 , n303786 , n303787 );
buf ( n303789 , n13360 );
xor ( n303790 , n299177 , n299188 );
xor ( n13363 , n303790 , n299537 );
xor ( n13364 , n303789 , n13363 );
xor ( n303793 , n9540 , n299971 );
xor ( n303794 , n303793 , n300028 );
xor ( n13367 , n299900 , n299917 );
buf ( n13368 , n13367 );
buf ( n303797 , n13368 );
buf ( n303798 , n772 );
buf ( n303799 , n828 );
xor ( n13372 , n303798 , n303799 );
buf ( n303801 , n13372 );
not ( n13374 , n303801 );
not ( n13375 , n294329 );
or ( n303804 , n13374 , n13375 );
buf ( n13377 , n1508 );
buf ( n13378 , n9682 );
nand ( n13379 , n13377 , n13378 );
buf ( n13380 , n13379 );
nand ( n303809 , n303804 , n13380 );
not ( n13382 , n303809 );
buf ( n303811 , n770 );
buf ( n303812 , n830 );
xor ( n13385 , n303811 , n303812 );
buf ( n13386 , n13385 );
buf ( n303815 , n13386 );
not ( n303816 , n303815 );
buf ( n303817 , n293454 );
not ( n303818 , n303817 );
or ( n13391 , n303816 , n303818 );
buf ( n303820 , n9476 );
buf ( n303821 , n831 );
nand ( n303822 , n303820 , n303821 );
buf ( n303823 , n303822 );
buf ( n303824 , n303823 );
nand ( n303825 , n13391 , n303824 );
buf ( n303826 , n303825 );
buf ( n303827 , n303826 );
not ( n303828 , n303827 );
buf ( n303829 , n799 );
buf ( n303830 , n296469 );
nand ( n303831 , n303829 , n303830 );
buf ( n303832 , n303831 );
buf ( n303833 , n303832 );
nand ( n13406 , n303828 , n303833 );
buf ( n303835 , n13406 );
not ( n13408 , n303835 );
or ( n13409 , n13382 , n13408 );
buf ( n303838 , n303832 );
not ( n13411 , n303838 );
buf ( n303840 , n303826 );
nand ( n13413 , n13411 , n303840 );
buf ( n303842 , n13413 );
nand ( n13415 , n13409 , n303842 );
buf ( n303844 , n13415 );
xor ( n13417 , n303797 , n303844 );
buf ( n303846 , n776 );
buf ( n303847 , n824 );
xor ( n13420 , n303846 , n303847 );
buf ( n303849 , n13420 );
buf ( n303850 , n303849 );
not ( n303851 , n303850 );
buf ( n303852 , n292473 );
not ( n303853 , n303852 );
or ( n13426 , n303851 , n303853 );
buf ( n303855 , n1613 );
buf ( n303856 , n9700 );
nand ( n303857 , n303855 , n303856 );
buf ( n303858 , n303857 );
buf ( n303859 , n303858 );
nand ( n303860 , n13426 , n303859 );
buf ( n303861 , n303860 );
buf ( n303862 , n784 );
buf ( n303863 , n816 );
xor ( n303864 , n303862 , n303863 );
buf ( n303865 , n303864 );
buf ( n303866 , n303865 );
not ( n303867 , n303866 );
buf ( n303868 , n292892 );
not ( n13441 , n303868 );
or ( n303870 , n303867 , n13441 );
buf ( n13443 , n1712 );
buf ( n303872 , n300166 );
nand ( n303873 , n13443 , n303872 );
buf ( n303874 , n303873 );
buf ( n303875 , n303874 );
nand ( n303876 , n303870 , n303875 );
buf ( n303877 , n303876 );
or ( n13450 , n303861 , n303877 );
buf ( n303879 , n786 );
buf ( n303880 , n814 );
xor ( n13453 , n303879 , n303880 );
buf ( n303882 , n13453 );
not ( n303883 , n303882 );
not ( n303884 , n2893 );
or ( n13457 , n303883 , n303884 );
buf ( n303886 , n292725 );
buf ( n13459 , n300151 );
nand ( n13460 , n303886 , n13459 );
buf ( n13461 , n13460 );
nand ( n303890 , n13457 , n13461 );
nand ( n13463 , n13450 , n303890 );
buf ( n303892 , n13463 );
buf ( n303893 , n303877 );
buf ( n303894 , n303861 );
nand ( n13467 , n303893 , n303894 );
buf ( n303896 , n13467 );
buf ( n303897 , n303896 );
nand ( n13470 , n303892 , n303897 );
buf ( n303899 , n13470 );
buf ( n303900 , n303899 );
and ( n303901 , n13417 , n303900 );
and ( n13474 , n303797 , n303844 );
or ( n303903 , n303901 , n13474 );
buf ( n303904 , n303903 );
or ( n13477 , n303794 , n303904 );
xor ( n303906 , n300162 , n9751 );
xor ( n303907 , n303906 , n300197 );
buf ( n303908 , n303907 );
buf ( n303909 , n303908 );
xor ( n303910 , n299989 , n300006 );
xor ( n303911 , n303910 , n300024 );
buf ( n303912 , n303911 );
buf ( n303913 , n303912 );
xor ( n303914 , n303909 , n303913 );
xor ( n13487 , n300106 , n300123 );
xor ( n303916 , n13487 , n300141 );
buf ( n303917 , n303916 );
buf ( n303918 , n303917 );
and ( n303919 , n303914 , n303918 );
and ( n13492 , n303909 , n303913 );
or ( n303921 , n303919 , n13492 );
buf ( n303922 , n303921 );
nand ( n13495 , n13477 , n303922 );
nand ( n303924 , n303794 , n303904 );
nand ( n13497 , n13495 , n303924 );
buf ( n303926 , n13497 );
xor ( n13499 , n299925 , n300032 );
xor ( n13500 , n13499 , n300207 );
buf ( n303929 , n13500 );
buf ( n303930 , n303929 );
xor ( n303931 , n303926 , n303930 );
xor ( n13504 , n299263 , n9023 );
xor ( n303933 , n13504 , n299533 );
buf ( n303934 , n303933 );
buf ( n303935 , n303934 );
and ( n303936 , n303931 , n303935 );
and ( n303937 , n303926 , n303930 );
or ( n13510 , n303936 , n303937 );
buf ( n303939 , n13510 );
and ( n303940 , n13364 , n303939 );
and ( n13513 , n303789 , n13363 );
or ( n13514 , n303940 , n13513 );
buf ( n303943 , n13514 );
xor ( n13516 , n13155 , n303943 );
xor ( n303945 , n9112 , n299771 );
xor ( n13518 , n303945 , n9785 );
buf ( n303947 , n13518 );
and ( n13520 , n13516 , n303947 );
and ( n303949 , n13155 , n303943 );
or ( n13522 , n13520 , n303949 );
buf ( n303951 , n13522 );
buf ( n303952 , n303951 );
xor ( n303953 , n299175 , n300217 );
xor ( n13526 , n303953 , n300440 );
buf ( n303955 , n13526 );
buf ( n303956 , n303955 );
and ( n13529 , n303952 , n303956 );
buf ( n303958 , n13529 );
buf ( n303959 , n303958 );
buf ( n303960 , n4288 );
xor ( n13533 , n303409 , n303415 );
and ( n303962 , n13533 , n303419 );
and ( n303963 , n303409 , n303415 );
or ( n13536 , n303962 , n303963 );
buf ( n303965 , n13536 );
buf ( n303966 , n303965 );
buf ( n13539 , n296401 );
xor ( n303968 , n845 , n303505 );
and ( n303969 , n303968 , n303509 );
and ( n13542 , n845 , n303505 );
or ( n303971 , n303969 , n13542 );
buf ( n13544 , n303971 );
buf ( n303973 , n297285 );
not ( n13546 , n303973 );
buf ( n303975 , n297193 );
not ( n13548 , n303975 );
and ( n303977 , n13546 , n13548 );
buf ( n303978 , n297285 );
buf ( n303979 , n297193 );
and ( n13552 , n303978 , n303979 );
nor ( n303981 , n303977 , n13552 );
buf ( n303982 , n303981 );
buf ( n303983 , n6862 );
not ( n13556 , n303983 );
and ( n303985 , n303982 , n13556 );
not ( n13558 , n303982 );
and ( n303987 , n13558 , n303983 );
nor ( n13560 , n303985 , n303987 );
buf ( n303989 , n13560 );
xor ( n303990 , n297542 , n297798 );
xor ( n303991 , n303990 , n297859 );
buf ( n303992 , n303991 );
buf ( n303993 , n303992 );
xor ( n303994 , n303989 , n303993 );
xor ( n303995 , n302134 , n302140 );
and ( n13568 , n303995 , n302157 );
and ( n303997 , n302134 , n302140 );
or ( n303998 , n13568 , n303997 );
buf ( n303999 , n303998 );
buf ( n304000 , n303999 );
and ( n304001 , n303994 , n304000 );
and ( n13574 , n303989 , n303993 );
or ( n304003 , n304001 , n13574 );
buf ( n304004 , n304003 );
buf ( n304005 , n304004 );
xor ( n13578 , n297533 , n297537 );
xor ( n304007 , n13578 , n297864 );
buf ( n304008 , n304007 );
buf ( n304009 , n304008 );
and ( n304010 , n304005 , n304009 );
buf ( n304011 , n304010 );
buf ( n13584 , n304011 );
not ( n304013 , n303809 );
and ( n13586 , n303826 , n303832 );
not ( n13587 , n303826 );
and ( n13588 , n799 , n6056 );
and ( n13589 , n13587 , n13588 );
nor ( n13590 , n13586 , n13589 );
and ( n13591 , n304013 , n13590 );
not ( n304020 , n304013 );
not ( n304021 , n13590 );
and ( n13594 , n304020 , n304021 );
nor ( n13595 , n13591 , n13594 );
buf ( n304024 , n13595 );
xor ( n13597 , n303685 , n303699 );
xor ( n304026 , n13597 , n303717 );
buf ( n304027 , n304026 );
buf ( n304028 , n304027 );
xor ( n13601 , n304024 , n304028 );
xor ( n304030 , n303736 , n303753 );
xor ( n13603 , n304030 , n303771 );
buf ( n304032 , n13603 );
buf ( n304033 , n304032 );
xor ( n13606 , n13601 , n304033 );
buf ( n304035 , n13606 );
buf ( n304036 , n304035 );
buf ( n304037 , n295991 );
not ( n304038 , n304037 );
buf ( n304039 , n295660 );
not ( n13612 , n304039 );
or ( n304041 , n304038 , n13612 );
nand ( n13614 , n298526 , n13258 );
buf ( n304043 , n13614 );
nand ( n304044 , n304041 , n304043 );
buf ( n304045 , n304044 );
not ( n13618 , n304045 );
buf ( n304047 , n799 );
buf ( n304048 , n802 );
xor ( n304049 , n304047 , n304048 );
buf ( n304050 , n304049 );
buf ( n304051 , n304050 );
not ( n304052 , n304051 );
buf ( n304053 , n296508 );
not ( n13626 , n304053 );
or ( n13627 , n304052 , n13626 );
buf ( n304056 , n296749 );
buf ( n304057 , n798 );
buf ( n304058 , n802 );
xor ( n304059 , n304057 , n304058 );
buf ( n304060 , n304059 );
buf ( n304061 , n304060 );
nand ( n304062 , n304056 , n304061 );
buf ( n304063 , n304062 );
buf ( n304064 , n304063 );
nand ( n13637 , n13627 , n304064 );
buf ( n304066 , n13637 );
buf ( n304067 , n304066 );
not ( n13640 , n304067 );
buf ( n304069 , n13640 );
not ( n304070 , n304069 );
or ( n13643 , n13618 , n304070 );
not ( n304072 , n304045 );
nand ( n304073 , n304072 , n304066 );
nand ( n13646 , n13643 , n304073 );
buf ( n304075 , n799 );
buf ( n304076 , n803 );
or ( n13649 , n304075 , n304076 );
buf ( n304078 , n804 );
nand ( n304079 , n13649 , n304078 );
buf ( n304080 , n304079 );
buf ( n304081 , n304080 );
buf ( n304082 , n799 );
buf ( n304083 , n803 );
nand ( n304084 , n304082 , n304083 );
buf ( n304085 , n304084 );
buf ( n304086 , n304085 );
buf ( n304087 , n802 );
and ( n13660 , n304081 , n304086 , n304087 );
buf ( n13661 , n13660 );
buf ( n304090 , n13661 );
buf ( n304091 , n296028 );
not ( n13664 , n304091 );
buf ( n304093 , n291656 );
not ( n304094 , n304093 );
or ( n13667 , n13664 , n304094 );
buf ( n304096 , n13386 );
buf ( n304097 , n831 );
nand ( n13670 , n304096 , n304097 );
buf ( n13671 , n13670 );
buf ( n304100 , n13671 );
nand ( n13673 , n13667 , n304100 );
buf ( n13674 , n13673 );
buf ( n13675 , n13674 );
xor ( n13676 , n304090 , n13675 );
buf ( n304105 , n13676 );
and ( n304106 , n13646 , n304105 );
not ( n13679 , n13646 );
not ( n304108 , n304105 );
and ( n304109 , n13679 , n304108 );
nor ( n13682 , n304106 , n304109 );
not ( n13683 , n296063 );
not ( n13684 , n5534 );
or ( n13685 , n13683 , n13684 );
nor ( n13686 , n5534 , n296063 );
or ( n13687 , n13686 , n5590 );
nand ( n13688 , n13685 , n13687 );
xor ( n13689 , n13682 , n13688 );
not ( n13690 , n296288 );
buf ( n304119 , n4860 );
not ( n13692 , n304119 );
buf ( n304121 , n295308 );
not ( n13694 , n304121 );
or ( n13695 , n13692 , n13694 );
buf ( n304124 , n296306 );
nand ( n13697 , n13695 , n304124 );
buf ( n304126 , n13697 );
not ( n304127 , n304126 );
or ( n13700 , n13690 , n304127 );
buf ( n304129 , n304126 );
buf ( n304130 , n296288 );
nor ( n304131 , n304129 , n304130 );
buf ( n304132 , n304131 );
not ( n13705 , n296294 );
or ( n13706 , n304132 , n13705 );
nand ( n13707 , n13700 , n13706 );
and ( n13708 , n13689 , n13707 );
and ( n13709 , n13682 , n13688 );
or ( n13710 , n13708 , n13709 );
buf ( n304139 , n13710 );
xor ( n13712 , n304036 , n304139 );
nand ( n13713 , n296062 , n296033 );
buf ( n13714 , n13713 );
or ( n13715 , n296062 , n296033 );
nand ( n13716 , n13715 , n296050 );
buf ( n304145 , n13716 );
nand ( n13718 , n13714 , n304145 );
buf ( n304147 , n13718 );
not ( n304148 , n295935 );
not ( n13721 , n295949 );
or ( n304150 , n304148 , n13721 );
or ( n13723 , n295935 , n295949 );
nand ( n304152 , n13723 , n295925 );
nand ( n304153 , n304150 , n304152 );
xor ( n13726 , n304147 , n304153 );
xor ( n304155 , n296194 , n296209 );
and ( n304156 , n304155 , n296227 );
and ( n13729 , n296194 , n296209 );
or ( n304158 , n304156 , n13729 );
buf ( n304159 , n304158 );
xor ( n304160 , n13726 , n304159 );
buf ( n304161 , n304160 );
not ( n304162 , n295975 );
nand ( n13735 , n304162 , n296000 );
not ( n304164 , n13735 );
not ( n304165 , n296017 );
or ( n13738 , n304164 , n304165 );
buf ( n304167 , n296000 );
not ( n304168 , n304167 );
buf ( n13741 , n295975 );
buf ( n304170 , n13741 );
nand ( n304171 , n304168 , n304170 );
buf ( n304172 , n304171 );
nand ( n13745 , n13738 , n304172 );
buf ( n304174 , n13745 );
buf ( n304175 , n5709 );
buf ( n304176 , n296126 );
or ( n304177 , n304175 , n304176 );
buf ( n13750 , n296117 );
nand ( n13751 , n304177 , n13750 );
buf ( n13752 , n13751 );
buf ( n304181 , n13752 );
buf ( n304182 , n5709 );
buf ( n304183 , n296126 );
nand ( n13756 , n304182 , n304183 );
buf ( n304185 , n13756 );
buf ( n304186 , n304185 );
nand ( n304187 , n304181 , n304186 );
buf ( n304188 , n304187 );
buf ( n304189 , n304188 );
xor ( n304190 , n304174 , n304189 );
buf ( n304191 , n5515 );
not ( n13764 , n304191 );
buf ( n304193 , n294329 );
not ( n304194 , n304193 );
or ( n13767 , n13764 , n304194 );
buf ( n304196 , n1508 );
buf ( n304197 , n303801 );
nand ( n13770 , n304196 , n304197 );
buf ( n13771 , n13770 );
buf ( n304200 , n13771 );
nand ( n13773 , n13767 , n304200 );
buf ( n304202 , n13773 );
buf ( n304203 , n304202 );
buf ( n304204 , n5759 );
not ( n304205 , n304204 );
buf ( n304206 , n292892 );
not ( n13779 , n304206 );
or ( n13780 , n304205 , n13779 );
buf ( n304209 , n1712 );
buf ( n304210 , n303865 );
nand ( n304211 , n304209 , n304210 );
buf ( n304212 , n304211 );
buf ( n304213 , n304212 );
nand ( n13786 , n13780 , n304213 );
buf ( n304215 , n13786 );
buf ( n304216 , n304215 );
xor ( n304217 , n304203 , n304216 );
buf ( n304218 , n295918 );
not ( n304219 , n304218 );
buf ( n304220 , n291835 );
not ( n13793 , n304220 );
or ( n304222 , n304219 , n13793 );
buf ( n304223 , n291843 );
buf ( n304224 , n303849 );
nand ( n304225 , n304223 , n304224 );
buf ( n304226 , n304225 );
buf ( n304227 , n304226 );
nand ( n13800 , n304222 , n304227 );
buf ( n304229 , n13800 );
buf ( n304230 , n304229 );
xor ( n304231 , n304217 , n304230 );
buf ( n304232 , n304231 );
buf ( n304233 , n304232 );
xor ( n304234 , n304190 , n304233 );
buf ( n304235 , n304234 );
buf ( n304236 , n304235 );
xor ( n304237 , n304161 , n304236 );
buf ( n304238 , n5833 );
not ( n13811 , n304238 );
not ( n304240 , n13811 );
not ( n304241 , n296232 );
or ( n13814 , n304240 , n304241 );
nand ( n304243 , n13814 , n296272 );
buf ( n13816 , n304243 );
nand ( n304245 , n296229 , n304238 );
buf ( n304246 , n304245 );
nand ( n304247 , n13816 , n304246 );
buf ( n304248 , n304247 );
buf ( n304249 , n304248 );
and ( n304250 , n304237 , n304249 );
and ( n304251 , n304161 , n304236 );
or ( n304252 , n304250 , n304251 );
buf ( n304253 , n304252 );
buf ( n304254 , n304253 );
xor ( n304255 , n13712 , n304254 );
buf ( n304256 , n304255 );
buf ( n304257 , n304256 );
xor ( n304258 , n304161 , n304236 );
xor ( n13831 , n304258 , n304249 );
buf ( n304260 , n13831 );
buf ( n13833 , n304260 );
not ( n13834 , n13833 );
buf ( n13835 , n13834 );
buf ( n304264 , n13835 );
xor ( n13837 , n13682 , n13688 );
xor ( n304266 , n13837 , n13707 );
buf ( n304267 , n304266 );
not ( n304268 , n304267 );
buf ( n304269 , n304268 );
buf ( n304270 , n304269 );
nand ( n304271 , n304264 , n304270 );
buf ( n304272 , n304271 );
buf ( n304273 , n304272 );
not ( n13846 , n304273 );
not ( n304275 , n5616 );
not ( n304276 , n293058 );
or ( n13849 , n304275 , n304276 );
buf ( n304278 , n292841 );
buf ( n304279 , n13224 );
nand ( n13852 , n304278 , n304279 );
buf ( n13853 , n13852 );
nand ( n304282 , n13849 , n13853 );
not ( n13855 , n304282 );
not ( n304284 , n13855 );
buf ( n304285 , n296124 );
not ( n13858 , n304285 );
buf ( n304287 , n292668 );
not ( n304288 , n304287 );
or ( n304289 , n13858 , n304288 );
buf ( n304290 , n303740 );
buf ( n304291 , n291734 );
nand ( n304292 , n304290 , n304291 );
buf ( n304293 , n304292 );
buf ( n304294 , n304293 );
nand ( n304295 , n304289 , n304294 );
buf ( n304296 , n304295 );
buf ( n304297 , n304296 );
buf ( n304298 , n296011 );
not ( n304299 , n304298 );
buf ( n304300 , n293394 );
not ( n13873 , n304300 );
or ( n304302 , n304299 , n13873 );
buf ( n304303 , n298746 );
buf ( n304304 , n303758 );
nand ( n13877 , n304303 , n304304 );
buf ( n13878 , n13877 );
buf ( n304307 , n13878 );
nand ( n13880 , n304302 , n304307 );
buf ( n304309 , n13880 );
buf ( n304310 , n304309 );
xor ( n304311 , n304297 , n304310 );
buf ( n304312 , n304311 );
not ( n13885 , n304312 );
or ( n304314 , n304284 , n13885 );
not ( n304315 , n304282 );
or ( n304316 , n304312 , n304315 );
nand ( n13889 , n304314 , n304316 );
buf ( n304318 , n13889 );
not ( n304319 , n296132 );
not ( n13892 , n293655 );
or ( n304321 , n304319 , n13892 );
buf ( n304322 , n6301 );
buf ( n304323 , n13299 );
nand ( n304324 , n304322 , n304323 );
buf ( n304325 , n304324 );
nand ( n13898 , n304321 , n304325 );
not ( n304327 , n296113 );
not ( n13900 , n295433 );
or ( n13901 , n304327 , n13900 );
buf ( n13902 , n295437 );
buf ( n304331 , n13276 );
nand ( n304332 , n13902 , n304331 );
buf ( n304333 , n304332 );
nand ( n304334 , n13901 , n304333 );
not ( n304335 , n304334 );
and ( n13908 , n13898 , n304335 );
not ( n304337 , n13898 );
and ( n304338 , n304337 , n304334 );
nor ( n13911 , n13908 , n304338 );
not ( n304340 , n5543 );
not ( n13913 , n4798 );
or ( n304342 , n304340 , n13913 );
buf ( n304343 , n295230 );
buf ( n304344 , n13243 );
nand ( n13917 , n304343 , n304344 );
buf ( n304346 , n13917 );
nand ( n304347 , n304342 , n304346 );
not ( n13920 , n304347 );
and ( n304349 , n13911 , n13920 );
not ( n13922 , n13911 );
and ( n304351 , n13922 , n304347 );
nor ( n304352 , n304349 , n304351 );
buf ( n304353 , n304352 );
xor ( n304354 , n304318 , n304353 );
buf ( n304355 , n2026 );
buf ( n304356 , n303629 );
nand ( n13929 , n304355 , n304356 );
buf ( n304358 , n13929 );
not ( n304359 , n2366 );
not ( n13932 , n292799 );
nand ( n13933 , n304359 , n13932 , n296060 );
nand ( n13934 , n304358 , n13933 );
not ( n13935 , n296220 );
not ( n304364 , n291761 );
or ( n304365 , n13935 , n304364 );
buf ( n304366 , n292105 );
buf ( n304367 , n303616 );
nand ( n13940 , n304366 , n304367 );
buf ( n304369 , n13940 );
nand ( n13942 , n304365 , n304369 );
xor ( n304371 , n13934 , n13942 );
buf ( n304372 , n5772 );
not ( n13945 , n304372 );
buf ( n304374 , n292719 );
not ( n13947 , n304374 );
or ( n13948 , n13945 , n13947 );
buf ( n304377 , n292518 );
buf ( n13950 , n303882 );
nand ( n13951 , n304377 , n13950 );
buf ( n304380 , n13951 );
buf ( n304381 , n304380 );
nand ( n304382 , n13948 , n304381 );
buf ( n304383 , n304382 );
xor ( n13956 , n304371 , n304383 );
buf ( n304385 , n13956 );
xor ( n304386 , n304354 , n304385 );
buf ( n304387 , n304386 );
not ( n13960 , n5721 );
not ( n304389 , n296156 );
or ( n304390 , n13960 , n304389 );
not ( n13963 , n5721 );
not ( n304392 , n13963 );
not ( n304393 , n296155 );
or ( n13966 , n304392 , n304393 );
nand ( n304395 , n13966 , n5738 );
nand ( n304396 , n304390 , n304395 );
and ( n13969 , n304387 , n304396 );
not ( n304398 , n304387 );
not ( n304399 , n304396 );
and ( n13972 , n304398 , n304399 );
nor ( n13973 , n13969 , n13972 );
not ( n13974 , n296310 );
not ( n13975 , n296232 );
not ( n304404 , n296278 );
or ( n304405 , n13975 , n304404 );
nand ( n13978 , n304405 , n5853 );
nand ( n13979 , n13974 , n13978 );
not ( n13980 , n296310 );
not ( n13981 , n5857 );
or ( n13982 , n13980 , n13981 );
nand ( n304411 , n13982 , n5752 );
nand ( n304412 , n13979 , n304411 );
and ( n13985 , n13973 , n304412 );
not ( n304414 , n13973 );
not ( n304415 , n304412 );
and ( n13988 , n304414 , n304415 );
nor ( n304417 , n13985 , n13988 );
buf ( n304418 , n304417 );
not ( n13991 , n304418 );
or ( n304420 , n13846 , n13991 );
buf ( n13993 , n13835 );
buf ( n304422 , n304269 );
or ( n13995 , n13993 , n304422 );
buf ( n304424 , n13995 );
buf ( n304425 , n304424 );
nand ( n13998 , n304420 , n304425 );
buf ( n304427 , n13998 );
buf ( n304428 , n304427 );
xor ( n14001 , n304257 , n304428 );
and ( n304430 , n304090 , n13675 );
buf ( n304431 , n304430 );
buf ( n304432 , n304431 );
not ( n304433 , n304060 );
not ( n14006 , n296508 );
or ( n304435 , n304433 , n14006 );
buf ( n304436 , n296517 );
buf ( n304437 , n300011 );
nand ( n14010 , n304436 , n304437 );
buf ( n304439 , n14010 );
nand ( n14012 , n304435 , n304439 );
buf ( n304441 , n14012 );
xor ( n14014 , n304432 , n304441 );
xor ( n14015 , n304203 , n304216 );
and ( n14016 , n14015 , n304230 );
and ( n14017 , n304203 , n304216 );
or ( n14018 , n14016 , n14017 );
buf ( n304447 , n14018 );
buf ( n304448 , n304447 );
xor ( n304449 , n14014 , n304448 );
buf ( n304450 , n304449 );
buf ( n304451 , n304450 );
xor ( n304452 , n304147 , n304153 );
and ( n304453 , n304452 , n304159 );
and ( n14026 , n304147 , n304153 );
or ( n304455 , n304453 , n14026 );
buf ( n304456 , n304455 );
xor ( n304457 , n304451 , n304456 );
xor ( n14030 , n304318 , n304353 );
and ( n304459 , n14030 , n304385 );
and ( n14032 , n304318 , n304353 );
or ( n14033 , n304459 , n14032 );
buf ( n304462 , n14033 );
buf ( n304463 , n304462 );
xor ( n304464 , n304457 , n304463 );
buf ( n304465 , n304464 );
buf ( n304466 , n304465 );
xor ( n304467 , n304174 , n304189 );
and ( n14040 , n304467 , n304233 );
and ( n304469 , n304174 , n304189 );
or ( n304470 , n14040 , n304469 );
buf ( n304471 , n304470 );
buf ( n304472 , n304471 );
buf ( n304473 , n296124 );
not ( n14046 , n304473 );
buf ( n304475 , n292668 );
not ( n14048 , n304475 );
or ( n304477 , n14046 , n14048 );
buf ( n304478 , n304293 );
nand ( n14051 , n304477 , n304478 );
buf ( n304480 , n14051 );
nor ( n304481 , n304480 , n304309 );
or ( n304482 , n304315 , n304481 );
nand ( n14055 , n304480 , n304309 );
nand ( n304484 , n304482 , n14055 );
buf ( n304485 , n304484 );
buf ( n304486 , n13920 );
not ( n304487 , n304486 );
not ( n304488 , n13898 );
buf ( n304489 , n304488 );
not ( n304490 , n304489 );
or ( n304491 , n304487 , n304490 );
not ( n14064 , n304335 );
buf ( n304493 , n14064 );
nand ( n304494 , n304491 , n304493 );
buf ( n304495 , n304494 );
buf ( n304496 , n304495 );
buf ( n304497 , n13898 );
buf ( n304498 , n304347 );
nand ( n14071 , n304497 , n304498 );
buf ( n304500 , n14071 );
buf ( n304501 , n304500 );
nand ( n14074 , n304496 , n304501 );
buf ( n14075 , n14074 );
buf ( n304504 , n14075 );
xor ( n304505 , n304485 , n304504 );
xor ( n304506 , n13934 , n13942 );
and ( n14079 , n304506 , n304383 );
and ( n14080 , n13934 , n13942 );
or ( n304509 , n14079 , n14080 );
buf ( n304510 , n304509 );
xor ( n304511 , n304505 , n304510 );
buf ( n304512 , n304511 );
buf ( n304513 , n304512 );
xor ( n304514 , n304472 , n304513 );
not ( n14087 , n304105 );
not ( n304516 , n304045 );
or ( n304517 , n14087 , n304516 );
buf ( n304518 , n304105 );
buf ( n304519 , n304045 );
nor ( n304520 , n304518 , n304519 );
buf ( n304521 , n304520 );
or ( n14094 , n304521 , n304069 );
nand ( n14095 , n304517 , n14094 );
buf ( n304524 , n14095 );
xor ( n14097 , n13196 , n303641 );
xor ( n304526 , n14097 , n13236 );
buf ( n304527 , n304526 );
xor ( n14100 , n304524 , n304527 );
xor ( n304529 , n303877 , n303890 );
xor ( n14102 , n304529 , n303861 );
buf ( n304531 , n14102 );
xor ( n14104 , n14100 , n304531 );
buf ( n304533 , n14104 );
buf ( n304534 , n304533 );
xor ( n14107 , n304514 , n304534 );
buf ( n304536 , n14107 );
buf ( n304537 , n304536 );
xor ( n14110 , n304466 , n304537 );
not ( n304539 , n304412 );
not ( n14112 , n304387 );
nand ( n304541 , n14112 , n304399 );
not ( n14114 , n304541 );
or ( n14115 , n304539 , n14114 );
nand ( n14116 , n304387 , n304396 );
nand ( n14117 , n14115 , n14116 );
buf ( n304546 , n14117 );
xor ( n304547 , n14110 , n304546 );
buf ( n304548 , n304547 );
buf ( n304549 , n304548 );
and ( n14122 , n14001 , n304549 );
and ( n14123 , n304257 , n304428 );
or ( n14124 , n14122 , n14123 );
buf ( n304553 , n14124 );
buf ( n304554 , n304553 );
xor ( n14127 , n292754 , n2583 );
xor ( n14128 , n14127 , n293262 );
buf ( n304557 , n14128 );
buf ( n14130 , n304557 );
buf ( n304559 , n882 );
buf ( n304560 , n850 );
and ( n304561 , n304559 , n304560 );
not ( n304562 , n304559 );
buf ( n304563 , n850 );
not ( n304564 , n304563 );
buf ( n304565 , n304564 );
buf ( n304566 , n304565 );
and ( n14139 , n304562 , n304566 );
nor ( n14140 , n304561 , n14139 );
buf ( n304569 , n14140 );
buf ( n304570 , n304569 );
not ( n304571 , n304570 );
buf ( n304572 , n883 );
buf ( n304573 , n884 );
xor ( n304574 , n304572 , n304573 );
buf ( n304575 , n304574 );
buf ( n304576 , n304575 );
not ( n304577 , n304576 );
xor ( n14150 , n882 , n883 );
buf ( n304579 , n14150 );
nand ( n14152 , n304577 , n304579 );
buf ( n304581 , n14152 );
buf ( n14154 , n304581 );
not ( n14155 , n14154 );
buf ( n304584 , n14155 );
buf ( n304585 , n304584 );
not ( n304586 , n304585 );
or ( n304587 , n304571 , n304586 );
buf ( n304588 , n882 );
buf ( n304589 , n849 );
xnor ( n14162 , n304588 , n304589 );
buf ( n304591 , n14162 );
buf ( n304592 , n304591 );
not ( n304593 , n304592 );
buf ( n304594 , n304575 );
buf ( n14167 , n304594 );
buf ( n304596 , n14167 );
buf ( n304597 , n304596 );
nand ( n304598 , n304593 , n304597 );
buf ( n304599 , n304598 );
buf ( n304600 , n304599 );
nand ( n304601 , n304587 , n304600 );
buf ( n304602 , n304601 );
buf ( n304603 , n304602 );
buf ( n304604 , n890 );
buf ( n304605 , n842 );
and ( n304606 , n304604 , n304605 );
not ( n14179 , n304604 );
buf ( n304608 , n842 );
not ( n304609 , n304608 );
buf ( n304610 , n304609 );
buf ( n304611 , n304610 );
and ( n14184 , n14179 , n304611 );
nor ( n14185 , n304606 , n14184 );
buf ( n304614 , n14185 );
buf ( n304615 , n304614 );
not ( n14188 , n304615 );
not ( n304617 , n890 );
nand ( n304618 , n304617 , n891 );
not ( n304619 , n304618 );
not ( n14192 , n891 );
nand ( n304621 , n14192 , n890 );
not ( n304622 , n304621 );
or ( n14195 , n304619 , n304622 );
and ( n304624 , n891 , n892 );
not ( n304625 , n891 );
not ( n14198 , n892 );
and ( n304627 , n304625 , n14198 );
nor ( n14200 , n304624 , n304627 );
not ( n304629 , n14200 );
nand ( n304630 , n14195 , n304629 );
buf ( n304631 , n304630 );
not ( n14204 , n304631 );
buf ( n304633 , n14204 );
buf ( n304634 , n304633 );
not ( n304635 , n304634 );
or ( n14208 , n14188 , n304635 );
buf ( n304637 , n890 );
not ( n14210 , n304637 );
buf ( n304639 , n841 );
nor ( n14212 , n14210 , n304639 );
buf ( n304641 , n14212 );
buf ( n14214 , n304641 );
buf ( n304643 , n841 );
not ( n304644 , n304643 );
buf ( n304645 , n890 );
nor ( n304646 , n304644 , n304645 );
buf ( n304647 , n304646 );
buf ( n304648 , n304647 );
nor ( n304649 , n14214 , n304648 );
buf ( n304650 , n304649 );
buf ( n304651 , n304650 );
not ( n304652 , n304651 );
buf ( n304653 , n14200 );
not ( n14226 , n304653 );
buf ( n304655 , n14226 );
buf ( n304656 , n304655 );
not ( n304657 , n304656 );
buf ( n304658 , n304657 );
buf ( n304659 , n304658 );
nand ( n304660 , n304652 , n304659 );
buf ( n304661 , n304660 );
buf ( n304662 , n304661 );
nand ( n14235 , n14208 , n304662 );
buf ( n14236 , n14235 );
buf ( n14237 , n14236 );
xor ( n14238 , n304603 , n14237 );
buf ( n304667 , n863 );
buf ( n304668 , n871 );
or ( n14241 , n304667 , n304668 );
buf ( n304670 , n872 );
nand ( n304671 , n14241 , n304670 );
buf ( n304672 , n304671 );
buf ( n304673 , n304672 );
buf ( n304674 , n863 );
buf ( n304675 , n871 );
nand ( n14248 , n304674 , n304675 );
buf ( n304677 , n14248 );
buf ( n304678 , n304677 );
buf ( n304679 , n870 );
and ( n304680 , n304673 , n304678 , n304679 );
buf ( n304681 , n304680 );
buf ( n304682 , n304681 );
buf ( n304683 , n841 );
buf ( n304684 , n892 );
xor ( n304685 , n304683 , n304684 );
buf ( n304686 , n304685 );
buf ( n304687 , n304686 );
not ( n304688 , n304687 );
buf ( n304689 , n892 );
buf ( n304690 , n893 );
xnor ( n304691 , n304689 , n304690 );
buf ( n304692 , n304691 );
buf ( n304693 , n304692 );
xor ( n304694 , n893 , n894 );
buf ( n304695 , n304694 );
nor ( n304696 , n304693 , n304695 );
buf ( n304697 , n304696 );
buf ( n304698 , n304697 );
buf ( n14271 , n304698 );
buf ( n14272 , n14271 );
buf ( n304701 , n14272 );
not ( n304702 , n304701 );
or ( n14275 , n304688 , n304702 );
buf ( n304704 , n892 );
not ( n14277 , n304704 );
buf ( n304706 , n840 );
nor ( n304707 , n14277 , n304706 );
buf ( n304708 , n304707 );
buf ( n304709 , n304708 );
buf ( n304710 , n840 );
not ( n14283 , n304710 );
buf ( n304712 , n892 );
nor ( n304713 , n14283 , n304712 );
buf ( n304714 , n304713 );
buf ( n14287 , n304714 );
nor ( n14288 , n304709 , n14287 );
buf ( n14289 , n14288 );
buf ( n304718 , n14289 );
not ( n14291 , n304718 );
buf ( n304720 , n304694 );
nand ( n304721 , n14291 , n304720 );
buf ( n304722 , n304721 );
buf ( n304723 , n304722 );
nand ( n304724 , n14275 , n304723 );
buf ( n304725 , n304724 );
buf ( n304726 , n304725 );
and ( n14299 , n304682 , n304726 );
buf ( n304728 , n14299 );
buf ( n304729 , n304728 );
xor ( n14302 , n14238 , n304729 );
buf ( n304731 , n14302 );
buf ( n304732 , n304731 );
buf ( n304733 , n870 );
buf ( n304734 , n862 );
and ( n304735 , n304733 , n304734 );
not ( n304736 , n304733 );
buf ( n14309 , n862 );
not ( n304738 , n14309 );
buf ( n304739 , n304738 );
buf ( n304740 , n304739 );
and ( n304741 , n304736 , n304740 );
nor ( n304742 , n304735 , n304741 );
buf ( n304743 , n304742 );
buf ( n304744 , n304743 );
not ( n14317 , n304744 );
xnor ( n14318 , n871 , n872 );
buf ( n304747 , n14318 );
xor ( n14320 , n870 , n871 );
buf ( n304749 , n14320 );
and ( n14322 , n304747 , n304749 );
buf ( n14323 , n14322 );
buf ( n304752 , n14323 );
buf ( n14325 , n304752 );
buf ( n304754 , n14325 );
buf ( n304755 , n304754 );
not ( n304756 , n304755 );
or ( n14329 , n14317 , n304756 );
buf ( n304758 , n14318 );
buf ( n14331 , n304758 );
buf ( n304760 , n14331 );
buf ( n14333 , n304760 );
not ( n304762 , n14333 );
buf ( n304763 , n304762 );
buf ( n304764 , n304763 );
buf ( n304765 , n870 );
buf ( n304766 , n861 );
and ( n304767 , n304765 , n304766 );
not ( n304768 , n304765 );
buf ( n304769 , n861 );
not ( n304770 , n304769 );
buf ( n304771 , n304770 );
buf ( n304772 , n304771 );
and ( n304773 , n304768 , n304772 );
nor ( n304774 , n304767 , n304773 );
buf ( n304775 , n304774 );
buf ( n304776 , n304775 );
nand ( n14349 , n304764 , n304776 );
buf ( n304778 , n14349 );
buf ( n304779 , n304778 );
nand ( n14352 , n14329 , n304779 );
buf ( n304781 , n14352 );
buf ( n304782 , n304781 );
buf ( n304783 , n884 );
buf ( n304784 , n848 );
not ( n14357 , n304784 );
buf ( n304786 , n14357 );
buf ( n304787 , n304786 );
and ( n14360 , n304783 , n304787 );
not ( n304789 , n304783 );
buf ( n304790 , n848 );
and ( n14363 , n304789 , n304790 );
nor ( n304792 , n14360 , n14363 );
buf ( n304793 , n304792 );
buf ( n304794 , n304793 );
not ( n304795 , n304794 );
buf ( n304796 , n304795 );
buf ( n14369 , n304796 );
not ( n14370 , n14369 );
buf ( n304799 , n884 );
buf ( n304800 , n885 );
xnor ( n14373 , n304799 , n304800 );
buf ( n304802 , n14373 );
buf ( n14375 , n304802 );
buf ( n304804 , n885 );
buf ( n304805 , n886 );
xor ( n304806 , n304804 , n304805 );
buf ( n304807 , n304806 );
buf ( n304808 , n304807 );
nor ( n304809 , n14375 , n304808 );
buf ( n304810 , n304809 );
buf ( n304811 , n304810 );
buf ( n304812 , n304811 );
buf ( n304813 , n304812 );
buf ( n304814 , n304813 );
not ( n304815 , n304814 );
or ( n304816 , n14370 , n304815 );
buf ( n304817 , n304807 );
buf ( n14390 , n304817 );
buf ( n304819 , n14390 );
buf ( n304820 , n304819 );
buf ( n304821 , n847 );
buf ( n304822 , n884 );
and ( n304823 , n304821 , n304822 );
not ( n304824 , n304821 );
buf ( n304825 , n884 );
not ( n14398 , n304825 );
buf ( n304827 , n14398 );
buf ( n304828 , n304827 );
and ( n14401 , n304824 , n304828 );
nor ( n14402 , n304823 , n14401 );
buf ( n14403 , n14402 );
buf ( n304832 , n14403 );
nand ( n14405 , n304820 , n304832 );
buf ( n304834 , n14405 );
buf ( n304835 , n304834 );
nand ( n14408 , n304816 , n304835 );
buf ( n304837 , n14408 );
buf ( n304838 , n304837 );
xor ( n14411 , n304782 , n304838 );
buf ( n304840 , n872 );
buf ( n304841 , n873 );
xnor ( n304842 , n304840 , n304841 );
buf ( n304843 , n304842 );
buf ( n304844 , n304843 );
xor ( n304845 , n873 , n874 );
buf ( n304846 , n304845 );
nor ( n14419 , n304844 , n304846 );
buf ( n14420 , n14419 );
buf ( n14421 , n14420 );
buf ( n14422 , n14421 );
buf ( n304851 , n14422 );
buf ( n304852 , n304851 );
not ( n14425 , n304852 );
buf ( n304854 , n14425 );
buf ( n304855 , n304854 );
buf ( n304856 , n860 );
buf ( n304857 , n872 );
xnor ( n304858 , n304856 , n304857 );
buf ( n304859 , n304858 );
buf ( n304860 , n304859 );
or ( n14433 , n304855 , n304860 );
buf ( n304862 , n304845 );
buf ( n14435 , n304862 );
buf ( n304864 , n14435 );
buf ( n304865 , n304864 );
not ( n14438 , n304865 );
buf ( n14439 , n14438 );
buf ( n304868 , n14439 );
buf ( n304869 , n872 );
buf ( n304870 , n859 );
and ( n304871 , n304869 , n304870 );
not ( n14444 , n304869 );
buf ( n304873 , n859 );
not ( n14446 , n304873 );
buf ( n14447 , n14446 );
buf ( n14448 , n14447 );
and ( n304877 , n14444 , n14448 );
nor ( n304878 , n304871 , n304877 );
buf ( n304879 , n304878 );
buf ( n304880 , n304879 );
not ( n304881 , n304880 );
buf ( n304882 , n304881 );
buf ( n304883 , n304882 );
or ( n304884 , n304868 , n304883 );
nand ( n14457 , n14433 , n304884 );
buf ( n304886 , n14457 );
buf ( n304887 , n304886 );
xor ( n14460 , n14411 , n304887 );
buf ( n304889 , n14460 );
buf ( n304890 , n304889 );
xor ( n304891 , n304732 , n304890 );
buf ( n304892 , n846 );
buf ( n304893 , n886 );
xor ( n304894 , n304892 , n304893 );
buf ( n304895 , n304894 );
buf ( n304896 , n304895 );
not ( n14469 , n304896 );
buf ( n304898 , n887 );
buf ( n304899 , n888 );
xor ( n304900 , n304898 , n304899 );
buf ( n304901 , n304900 );
buf ( n304902 , n304901 );
buf ( n304903 , n886 );
buf ( n304904 , n887 );
xnor ( n14477 , n304903 , n304904 );
buf ( n304906 , n14477 );
buf ( n304907 , n304906 );
nor ( n14480 , n304902 , n304907 );
buf ( n304909 , n14480 );
buf ( n304910 , n304909 );
buf ( n14483 , n304910 );
buf ( n304912 , n14483 );
buf ( n304913 , n304912 );
not ( n14486 , n304913 );
or ( n14487 , n14469 , n14486 );
buf ( n304916 , n886 );
buf ( n304917 , n845 );
xnor ( n14490 , n304916 , n304917 );
buf ( n304919 , n14490 );
buf ( n304920 , n304919 );
not ( n14493 , n304920 );
buf ( n304922 , n304901 );
nand ( n14495 , n14493 , n304922 );
buf ( n304924 , n14495 );
buf ( n304925 , n304924 );
nand ( n304926 , n14487 , n304925 );
buf ( n304927 , n304926 );
buf ( n304928 , n304927 );
buf ( n14501 , n879 );
buf ( n304930 , n880 );
xor ( n304931 , n14501 , n304930 );
buf ( n304932 , n304931 );
buf ( n304933 , n304932 );
not ( n14506 , n304933 );
xor ( n14507 , n879 , n878 );
buf ( n304936 , n14507 );
nand ( n14509 , n14506 , n304936 );
buf ( n304938 , n14509 );
buf ( n304939 , n304938 );
buf ( n14512 , n304939 );
buf ( n304941 , n14512 );
buf ( n304942 , n304941 );
buf ( n304943 , n878 );
buf ( n304944 , n854 );
xnor ( n304945 , n304943 , n304944 );
buf ( n304946 , n304945 );
buf ( n304947 , n304946 );
or ( n304948 , n304942 , n304947 );
buf ( n304949 , n304932 );
not ( n14522 , n304949 );
buf ( n14523 , n14522 );
buf ( n304952 , n14523 );
buf ( n304953 , n878 );
buf ( n304954 , n853 );
not ( n14527 , n304954 );
buf ( n304956 , n14527 );
buf ( n304957 , n304956 );
and ( n14530 , n304953 , n304957 );
not ( n14531 , n304953 );
buf ( n14532 , n853 );
and ( n14533 , n14531 , n14532 );
nor ( n304962 , n14530 , n14533 );
buf ( n304963 , n304962 );
buf ( n304964 , n304963 );
or ( n14537 , n304952 , n304964 );
nand ( n304966 , n304948 , n14537 );
buf ( n304967 , n304966 );
buf ( n304968 , n304967 );
xor ( n304969 , n304928 , n304968 );
buf ( n14542 , n881 );
buf ( n304971 , n882 );
xor ( n304972 , n14542 , n304971 );
buf ( n304973 , n304972 );
buf ( n304974 , n304973 );
not ( n304975 , n304974 );
buf ( n304976 , n304975 );
buf ( n304977 , n304976 );
xor ( n14550 , n881 , n880 );
buf ( n304979 , n14550 );
nand ( n304980 , n304977 , n304979 );
buf ( n304981 , n304980 );
buf ( n304982 , n304981 );
not ( n14555 , n304982 );
buf ( n304984 , n14555 );
buf ( n14557 , n304984 );
not ( n304986 , n14557 );
buf ( n304987 , n304986 );
buf ( n304988 , n304987 );
buf ( n304989 , n852 );
buf ( n14562 , n880 );
xnor ( n14563 , n304989 , n14562 );
buf ( n14564 , n14563 );
buf ( n304993 , n14564 );
or ( n14566 , n304988 , n304993 );
buf ( n304995 , n304973 );
buf ( n304996 , n304995 );
buf ( n304997 , n304996 );
buf ( n304998 , n304997 );
not ( n14571 , n304998 );
buf ( n305000 , n14571 );
buf ( n305001 , n305000 );
buf ( n305002 , n880 );
buf ( n305003 , n851 );
xor ( n305004 , n305002 , n305003 );
buf ( n305005 , n305004 );
buf ( n305006 , n305005 );
not ( n305007 , n305006 );
buf ( n305008 , n305007 );
buf ( n305009 , n305008 );
or ( n14582 , n305001 , n305009 );
nand ( n305011 , n14566 , n14582 );
buf ( n305012 , n305011 );
buf ( n305013 , n305012 );
xor ( n14586 , n304969 , n305013 );
buf ( n305015 , n14586 );
buf ( n305016 , n305015 );
and ( n14589 , n304891 , n305016 );
and ( n305018 , n304732 , n304890 );
or ( n305019 , n14589 , n305018 );
buf ( n305020 , n305019 );
buf ( n305021 , n305020 );
xor ( n305022 , n894 , n837 );
buf ( n305023 , n305022 );
not ( n14596 , n305023 );
buf ( n305025 , n895 );
not ( n305026 , n305025 );
buf ( n305027 , n894 );
nand ( n305028 , n305026 , n305027 );
buf ( n305029 , n305028 );
buf ( n305030 , n305029 );
not ( n305031 , n305030 );
buf ( n305032 , n305031 );
buf ( n305033 , n305032 );
not ( n14606 , n305033 );
or ( n305035 , n14596 , n14606 );
buf ( n305036 , n836 );
buf ( n305037 , n894 );
xor ( n305038 , n305036 , n305037 );
buf ( n305039 , n305038 );
buf ( n305040 , n305039 );
buf ( n305041 , n895 );
nand ( n305042 , n305040 , n305041 );
buf ( n305043 , n305042 );
buf ( n305044 , n305043 );
nand ( n305045 , n305035 , n305044 );
buf ( n305046 , n305045 );
buf ( n305047 , n305046 );
buf ( n305048 , n304879 );
not ( n305049 , n305048 );
buf ( n305050 , n304851 );
not ( n14623 , n305050 );
or ( n305052 , n305049 , n14623 );
buf ( n305053 , n304845 );
buf ( n305054 , n872 );
buf ( n305055 , n858 );
and ( n305056 , n305054 , n305055 );
not ( n305057 , n305054 );
buf ( n305058 , n858 );
not ( n305059 , n305058 );
buf ( n305060 , n305059 );
buf ( n305061 , n305060 );
and ( n305062 , n305057 , n305061 );
nor ( n305063 , n305056 , n305062 );
buf ( n305064 , n305063 );
buf ( n305065 , n305064 );
nand ( n305066 , n305053 , n305065 );
buf ( n305067 , n305066 );
buf ( n305068 , n305067 );
nand ( n14641 , n305052 , n305068 );
buf ( n305070 , n14641 );
buf ( n305071 , n305070 );
xor ( n14644 , n305047 , n305071 );
buf ( n305073 , n14403 );
not ( n305074 , n305073 );
buf ( n305075 , n304813 );
not ( n14648 , n305075 );
or ( n305077 , n305074 , n14648 );
buf ( n305078 , n304819 );
buf ( n305079 , n846 );
buf ( n305080 , n884 );
xor ( n305081 , n305079 , n305080 );
buf ( n305082 , n305081 );
buf ( n305083 , n305082 );
nand ( n305084 , n305078 , n305083 );
buf ( n305085 , n305084 );
buf ( n305086 , n305085 );
nand ( n305087 , n305077 , n305086 );
buf ( n305088 , n305087 );
buf ( n305089 , n305088 );
xor ( n305090 , n14644 , n305089 );
buf ( n305091 , n305090 );
buf ( n305092 , n305091 );
buf ( n305093 , n305005 );
not ( n14666 , n305093 );
buf ( n305095 , n304976 );
buf ( n305096 , n14550 );
and ( n305097 , n305095 , n305096 );
buf ( n305098 , n305097 );
buf ( n305099 , n305098 );
not ( n305100 , n305099 );
or ( n14673 , n14666 , n305100 );
buf ( n305102 , n304997 );
xor ( n305103 , n880 , n850 );
buf ( n305104 , n305103 );
nand ( n305105 , n305102 , n305104 );
buf ( n305106 , n305105 );
buf ( n305107 , n305106 );
nand ( n14680 , n14673 , n305107 );
buf ( n14681 , n14680 );
buf ( n305110 , n14681 );
buf ( n305111 , n888 );
buf ( n305112 , n843 );
and ( n305113 , n305111 , n305112 );
not ( n14686 , n305111 );
buf ( n305115 , n843 );
not ( n305116 , n305115 );
buf ( n305117 , n305116 );
buf ( n305118 , n305117 );
and ( n14691 , n14686 , n305118 );
nor ( n14692 , n305113 , n14691 );
buf ( n305121 , n14692 );
buf ( n305122 , n305121 );
not ( n305123 , n305122 );
buf ( n305124 , n889 );
buf ( n305125 , n890 );
xor ( n305126 , n305124 , n305125 );
buf ( n305127 , n305126 );
buf ( n305128 , n305127 );
not ( n14701 , n305128 );
buf ( n305130 , n14701 );
buf ( n305131 , n305130 );
xor ( n305132 , n889 , n888 );
buf ( n305133 , n305132 );
nand ( n305134 , n305131 , n305133 );
buf ( n305135 , n305134 );
buf ( n305136 , n305135 );
not ( n305137 , n305136 );
buf ( n305138 , n305137 );
buf ( n305139 , n305138 );
not ( n14712 , n305139 );
or ( n14713 , n305123 , n14712 );
buf ( n14714 , n305127 );
buf ( n305143 , n14714 );
buf ( n305144 , n305143 );
buf ( n305145 , n305144 );
buf ( n14718 , n888 );
buf ( n305147 , n842 );
xor ( n14720 , n14718 , n305147 );
buf ( n305149 , n14720 );
buf ( n305150 , n305149 );
nand ( n14723 , n305145 , n305150 );
buf ( n305152 , n14723 );
buf ( n305153 , n305152 );
nand ( n305154 , n14713 , n305153 );
buf ( n305155 , n305154 );
buf ( n305156 , n305155 );
xor ( n305157 , n305110 , n305156 );
buf ( n305158 , n304941 );
buf ( n305159 , n304963 );
or ( n305160 , n305158 , n305159 );
buf ( n305161 , n14523 );
buf ( n305162 , n878 );
buf ( n14735 , n852 );
and ( n14736 , n305162 , n14735 );
not ( n305165 , n305162 );
buf ( n305166 , n852 );
not ( n305167 , n305166 );
buf ( n305168 , n305167 );
buf ( n305169 , n305168 );
and ( n305170 , n305165 , n305169 );
nor ( n305171 , n14736 , n305170 );
buf ( n305172 , n305171 );
buf ( n305173 , n305172 );
not ( n305174 , n305173 );
buf ( n305175 , n305174 );
buf ( n305176 , n305175 );
or ( n305177 , n305161 , n305176 );
nand ( n14750 , n305160 , n305177 );
buf ( n305179 , n14750 );
buf ( n305180 , n305179 );
xor ( n14753 , n305157 , n305180 );
buf ( n305182 , n14753 );
buf ( n305183 , n305182 );
xor ( n14756 , n305092 , n305183 );
buf ( n305185 , n868 );
buf ( n305186 , n863 );
and ( n14759 , n305185 , n305186 );
not ( n14760 , n305185 );
buf ( n305189 , n863 );
not ( n14762 , n305189 );
buf ( n305191 , n14762 );
buf ( n305192 , n305191 );
buf ( n305193 , n305192 );
and ( n14766 , n14760 , n305193 );
nor ( n305195 , n14759 , n14766 );
buf ( n305196 , n305195 );
buf ( n305197 , n305196 );
not ( n305198 , n305197 );
buf ( n305199 , n869 );
buf ( n305200 , n870 );
xor ( n14773 , n305199 , n305200 );
buf ( n305202 , n14773 );
buf ( n305203 , n305202 );
not ( n14776 , n305203 );
buf ( n305205 , n14776 );
buf ( n14778 , n305205 );
xor ( n305207 , n868 , n869 );
buf ( n305208 , n305207 );
nand ( n305209 , n14778 , n305208 );
buf ( n305210 , n305209 );
buf ( n305211 , n305210 );
not ( n305212 , n305211 );
buf ( n305213 , n305212 );
buf ( n305214 , n305213 );
not ( n305215 , n305214 );
or ( n14788 , n305198 , n305215 );
buf ( n305217 , n305202 );
buf ( n14790 , n305217 );
buf ( n305219 , n14790 );
buf ( n305220 , n305219 );
xor ( n14793 , n868 , n862 );
buf ( n305222 , n14793 );
nand ( n305223 , n305220 , n305222 );
buf ( n305224 , n305223 );
buf ( n305225 , n305224 );
nand ( n305226 , n14788 , n305225 );
buf ( n305227 , n305226 );
buf ( n305228 , n305227 );
buf ( n305229 , n304775 );
not ( n305230 , n305229 );
buf ( n305231 , n304754 );
not ( n305232 , n305231 );
or ( n14805 , n305230 , n305232 );
buf ( n305234 , n304763 );
buf ( n305235 , n870 );
buf ( n305236 , n860 );
and ( n14809 , n305235 , n305236 );
not ( n14810 , n305235 );
buf ( n305239 , n860 );
not ( n305240 , n305239 );
buf ( n305241 , n305240 );
buf ( n305242 , n305241 );
and ( n305243 , n14810 , n305242 );
nor ( n305244 , n14809 , n305243 );
buf ( n305245 , n305244 );
buf ( n305246 , n305245 );
nand ( n305247 , n305234 , n305246 );
buf ( n305248 , n305247 );
buf ( n305249 , n305248 );
nand ( n14822 , n14805 , n305249 );
buf ( n305251 , n14822 );
buf ( n305252 , n305251 );
xor ( n14825 , n305228 , n305252 );
buf ( n305254 , n304630 );
buf ( n305255 , n304650 );
or ( n305256 , n305254 , n305255 );
buf ( n305257 , n304655 );
buf ( n305258 , n890 );
buf ( n305259 , n840 );
not ( n14832 , n305259 );
buf ( n305261 , n14832 );
buf ( n14834 , n305261 );
and ( n14835 , n305258 , n14834 );
not ( n14836 , n305258 );
buf ( n305265 , n840 );
and ( n14838 , n14836 , n305265 );
nor ( n14839 , n14835 , n14838 );
buf ( n305268 , n14839 );
buf ( n305269 , n305268 );
or ( n305270 , n305257 , n305269 );
nand ( n305271 , n305256 , n305270 );
buf ( n305272 , n305271 );
buf ( n305273 , n305272 );
xor ( n305274 , n14825 , n305273 );
buf ( n305275 , n305274 );
buf ( n305276 , n305275 );
xor ( n14849 , n14756 , n305276 );
buf ( n305278 , n14849 );
buf ( n305279 , n305278 );
xor ( n305280 , n305021 , n305279 );
xor ( n14853 , n874 , n857 );
buf ( n305282 , n14853 );
not ( n305283 , n305282 );
buf ( n305284 , n874 );
buf ( n305285 , n875 );
xnor ( n305286 , n305284 , n305285 );
buf ( n305287 , n305286 );
buf ( n14860 , n305287 );
xor ( n305289 , n875 , n876 );
buf ( n305290 , n305289 );
nor ( n305291 , n14860 , n305290 );
buf ( n305292 , n305291 );
buf ( n305293 , n305292 );
not ( n305294 , n305293 );
or ( n305295 , n305283 , n305294 );
buf ( n305296 , n305289 );
not ( n305297 , n305296 );
buf ( n305298 , n305297 );
buf ( n14871 , n305298 );
not ( n305300 , n14871 );
buf ( n305301 , n305300 );
buf ( n305302 , n305301 );
buf ( n305303 , n874 );
buf ( n305304 , n856 );
xor ( n305305 , n305303 , n305304 );
buf ( n305306 , n305305 );
buf ( n305307 , n305306 );
nand ( n305308 , n305302 , n305307 );
buf ( n305309 , n305308 );
buf ( n305310 , n305309 );
nand ( n305311 , n305295 , n305310 );
buf ( n305312 , n305311 );
buf ( n305313 , n876 );
buf ( n14886 , n855 );
and ( n14887 , n305313 , n14886 );
not ( n14888 , n305313 );
buf ( n305317 , n855 );
not ( n14890 , n305317 );
buf ( n305319 , n14890 );
buf ( n305320 , n305319 );
and ( n305321 , n14888 , n305320 );
nor ( n14894 , n14887 , n305321 );
buf ( n305323 , n14894 );
buf ( n305324 , n305323 );
not ( n14897 , n305324 );
buf ( n305326 , n876 );
buf ( n305327 , n877 );
xnor ( n14900 , n305326 , n305327 );
buf ( n14901 , n14900 );
buf ( n305330 , n14901 );
buf ( n305331 , n877 );
buf ( n305332 , n878 );
xor ( n305333 , n305331 , n305332 );
buf ( n305334 , n305333 );
buf ( n305335 , n305334 );
nor ( n14908 , n305330 , n305335 );
buf ( n305337 , n14908 );
buf ( n305338 , n305337 );
buf ( n305339 , n305338 );
not ( n305340 , n305339 );
or ( n305341 , n14897 , n305340 );
buf ( n305342 , n305334 );
buf ( n305343 , n305342 );
buf ( n305344 , n305343 );
buf ( n305345 , n305344 );
xor ( n14918 , n876 , n854 );
buf ( n305347 , n14918 );
nand ( n305348 , n305345 , n305347 );
buf ( n305349 , n305348 );
buf ( n305350 , n305349 );
nand ( n305351 , n305341 , n305350 );
buf ( n305352 , n305351 );
xor ( n305353 , n305312 , n305352 );
buf ( n305354 , n304912 );
not ( n305355 , n305354 );
buf ( n305356 , n305355 );
buf ( n305357 , n305356 );
buf ( n305358 , n304919 );
or ( n305359 , n305357 , n305358 );
buf ( n305360 , n887 );
buf ( n305361 , n888 );
xnor ( n305362 , n305360 , n305361 );
buf ( n305363 , n305362 );
buf ( n305364 , n305363 );
buf ( n305365 , n844 );
buf ( n305366 , n886 );
xnor ( n14939 , n305365 , n305366 );
buf ( n305368 , n14939 );
buf ( n305369 , n305368 );
or ( n305370 , n305364 , n305369 );
nand ( n14943 , n305359 , n305370 );
buf ( n14944 , n14943 );
xor ( n305373 , n305353 , n14944 );
xor ( n14946 , n304603 , n14237 );
and ( n305375 , n14946 , n304729 );
and ( n14948 , n304603 , n14237 );
or ( n305377 , n305375 , n14948 );
buf ( n305378 , n305377 );
buf ( n305379 , n304584 );
not ( n305380 , n305379 );
buf ( n305381 , n305380 );
buf ( n305382 , n305381 );
buf ( n305383 , n304591 );
or ( n305384 , n305382 , n305383 );
buf ( n305385 , n304596 );
not ( n14958 , n305385 );
buf ( n14959 , n14958 );
buf ( n14960 , n14959 );
xor ( n14961 , n882 , n848 );
buf ( n305390 , n14961 );
not ( n305391 , n305390 );
buf ( n305392 , n305391 );
buf ( n305393 , n305392 );
or ( n305394 , n14960 , n305393 );
nand ( n14967 , n305384 , n305394 );
buf ( n305396 , n14967 );
buf ( n14969 , n305396 );
buf ( n305398 , n863 );
buf ( n305399 , n869 );
or ( n14972 , n305398 , n305399 );
buf ( n305401 , n870 );
nand ( n305402 , n14972 , n305401 );
buf ( n305403 , n305402 );
buf ( n305404 , n305403 );
buf ( n305405 , n863 );
buf ( n305406 , n869 );
nand ( n305407 , n305405 , n305406 );
buf ( n305408 , n305407 );
buf ( n305409 , n305408 );
buf ( n305410 , n868 );
and ( n14983 , n305404 , n305409 , n305410 );
buf ( n305412 , n14983 );
buf ( n305413 , n305412 );
buf ( n305414 , n892 );
buf ( n305415 , n839 );
and ( n14988 , n305414 , n305415 );
not ( n14989 , n305414 );
buf ( n305418 , n839 );
not ( n14991 , n305418 );
buf ( n14992 , n14991 );
buf ( n305421 , n14992 );
and ( n14994 , n14989 , n305421 );
nor ( n305423 , n14988 , n14994 );
buf ( n305424 , n305423 );
buf ( n305425 , n305424 );
not ( n14998 , n305425 );
buf ( n305427 , n14272 );
not ( n15000 , n305427 );
or ( n305429 , n14998 , n15000 );
xor ( n305430 , n893 , n894 );
buf ( n305431 , n305430 );
buf ( n305432 , n838 );
buf ( n305433 , n892 );
xor ( n15006 , n305432 , n305433 );
buf ( n305435 , n15006 );
buf ( n305436 , n305435 );
nand ( n305437 , n305431 , n305436 );
buf ( n305438 , n305437 );
buf ( n305439 , n305438 );
nand ( n305440 , n305429 , n305439 );
buf ( n305441 , n305440 );
buf ( n305442 , n305441 );
xor ( n15015 , n305413 , n305442 );
buf ( n305444 , n15015 );
buf ( n305445 , n305444 );
xor ( n15018 , n14969 , n305445 );
buf ( n15019 , n305219 );
not ( n305448 , n15019 );
buf ( n305449 , n305448 );
buf ( n305450 , n305449 );
buf ( n305451 , n305192 );
nor ( n305452 , n305450 , n305451 );
buf ( n305453 , n305452 );
buf ( n305454 , n305453 );
buf ( n305455 , n888 );
buf ( n305456 , n844 );
not ( n15029 , n305456 );
buf ( n305458 , n15029 );
buf ( n305459 , n305458 );
and ( n305460 , n305455 , n305459 );
not ( n305461 , n305455 );
buf ( n305462 , n844 );
and ( n15035 , n305461 , n305462 );
nor ( n305464 , n305460 , n15035 );
buf ( n305465 , n305464 );
buf ( n305466 , n305465 );
not ( n305467 , n305466 );
buf ( n305468 , n305467 );
buf ( n305469 , n305468 );
not ( n305470 , n305469 );
buf ( n305471 , n305138 );
not ( n305472 , n305471 );
or ( n305473 , n305470 , n305472 );
buf ( n305474 , n305144 );
buf ( n305475 , n305121 );
nand ( n15048 , n305474 , n305475 );
buf ( n305477 , n15048 );
buf ( n305478 , n305477 );
nand ( n305479 , n305473 , n305478 );
buf ( n305480 , n305479 );
buf ( n305481 , n305480 );
xor ( n305482 , n305454 , n305481 );
buf ( n305483 , n14272 );
not ( n15056 , n305483 );
buf ( n15057 , n15056 );
buf ( n305486 , n15057 );
buf ( n305487 , n14289 );
or ( n305488 , n305486 , n305487 );
not ( n305489 , n305430 );
buf ( n305490 , n305489 );
buf ( n305491 , n305424 );
not ( n15064 , n305491 );
buf ( n15065 , n15064 );
buf ( n305494 , n15065 );
or ( n15067 , n305490 , n305494 );
nand ( n15068 , n305488 , n15067 );
buf ( n305497 , n15068 );
buf ( n305498 , n305497 );
and ( n15071 , n305482 , n305498 );
and ( n305500 , n305454 , n305481 );
or ( n305501 , n15071 , n305500 );
buf ( n305502 , n305501 );
buf ( n305503 , n305502 );
xor ( n305504 , n15018 , n305503 );
buf ( n305505 , n305504 );
xor ( n305506 , n305378 , n305505 );
xor ( n15079 , n305373 , n305506 );
buf ( n305508 , n15079 );
xor ( n15081 , n305280 , n305508 );
buf ( n305510 , n15081 );
buf ( n15083 , n305510 );
buf ( n305512 , n304581 );
buf ( n305513 , n882 );
buf ( n305514 , n305168 );
and ( n305515 , n305513 , n305514 );
not ( n305516 , n305513 );
buf ( n305517 , n852 );
and ( n305518 , n305516 , n305517 );
nor ( n305519 , n305515 , n305518 );
buf ( n305520 , n305519 );
buf ( n305521 , n305520 );
or ( n305522 , n305512 , n305521 );
buf ( n305523 , n14959 );
buf ( n305524 , n882 );
not ( n305525 , n305524 );
buf ( n305526 , n305525 );
buf ( n305527 , n305526 );
buf ( n305528 , n851 );
and ( n15101 , n305527 , n305528 );
buf ( n305530 , n851 );
not ( n305531 , n305530 );
buf ( n305532 , n305531 );
buf ( n305533 , n305532 );
buf ( n305534 , n882 );
and ( n15107 , n305533 , n305534 );
nor ( n15108 , n15101 , n15107 );
buf ( n305537 , n15108 );
buf ( n305538 , n305537 );
or ( n305539 , n305523 , n305538 );
nand ( n15112 , n305522 , n305539 );
buf ( n305541 , n15112 );
buf ( n305542 , n305541 );
buf ( n305543 , n863 );
buf ( n305544 , n873 );
or ( n15117 , n305543 , n305544 );
buf ( n305546 , n874 );
nand ( n305547 , n15117 , n305546 );
buf ( n305548 , n305547 );
buf ( n305549 , n305548 );
buf ( n305550 , n863 );
buf ( n305551 , n873 );
nand ( n15124 , n305550 , n305551 );
buf ( n305553 , n15124 );
buf ( n305554 , n305553 );
buf ( n305555 , n872 );
and ( n15128 , n305549 , n305554 , n305555 );
buf ( n15129 , n15128 );
buf ( n305558 , n15129 );
buf ( n305559 , n14272 );
not ( n305560 , n305559 );
buf ( n305561 , n305560 );
buf ( n305562 , n305561 );
buf ( n305563 , n843 );
buf ( n305564 , n892 );
not ( n15137 , n305564 );
buf ( n305566 , n15137 );
buf ( n305567 , n305566 );
and ( n305568 , n305563 , n305567 );
not ( n15141 , n305563 );
buf ( n305570 , n892 );
and ( n305571 , n15141 , n305570 );
nor ( n15144 , n305568 , n305571 );
buf ( n15145 , n15144 );
buf ( n305574 , n15145 );
or ( n15147 , n305562 , n305574 );
buf ( n305576 , n305489 );
buf ( n305577 , n892 );
buf ( n305578 , n842 );
xnor ( n15151 , n305577 , n305578 );
buf ( n305580 , n15151 );
buf ( n305581 , n305580 );
or ( n15154 , n305576 , n305581 );
nand ( n305583 , n15147 , n15154 );
buf ( n305584 , n305583 );
buf ( n15157 , n305584 );
and ( n15158 , n305558 , n15157 );
buf ( n305587 , n15158 );
buf ( n15160 , n305587 );
xor ( n15161 , n305542 , n15160 );
buf ( n305590 , n886 );
buf ( n305591 , n849 );
and ( n15164 , n305590 , n305591 );
not ( n305593 , n305590 );
buf ( n305594 , n849 );
not ( n305595 , n305594 );
buf ( n305596 , n305595 );
buf ( n305597 , n305596 );
and ( n305598 , n305593 , n305597 );
nor ( n15171 , n15164 , n305598 );
buf ( n305600 , n15171 );
buf ( n305601 , n305600 );
not ( n15174 , n305601 );
buf ( n305603 , n304912 );
not ( n305604 , n305603 );
or ( n15177 , n15174 , n305604 );
buf ( n305606 , n304901 );
buf ( n305607 , n848 );
buf ( n305608 , n886 );
xor ( n15181 , n305607 , n305608 );
buf ( n305610 , n15181 );
buf ( n305611 , n305610 );
nand ( n15184 , n305606 , n305611 );
buf ( n15185 , n15184 );
buf ( n305614 , n15185 );
nand ( n15187 , n15177 , n305614 );
buf ( n305616 , n15187 );
buf ( n305617 , n305616 );
xor ( n305618 , n874 , n861 );
buf ( n305619 , n305618 );
not ( n15192 , n305619 );
buf ( n305621 , n305287 );
buf ( n305622 , n305289 );
nor ( n305623 , n305621 , n305622 );
buf ( n305624 , n305623 );
buf ( n305625 , n305624 );
buf ( n15198 , n305625 );
buf ( n305627 , n15198 );
buf ( n305628 , n305627 );
not ( n15201 , n305628 );
or ( n305630 , n15192 , n15201 );
buf ( n15203 , n305301 );
buf ( n305632 , n874 );
buf ( n305633 , n860 );
and ( n15206 , n305632 , n305633 );
not ( n15207 , n305632 );
buf ( n305636 , n305241 );
and ( n305637 , n15207 , n305636 );
nor ( n305638 , n15206 , n305637 );
buf ( n305639 , n305638 );
buf ( n305640 , n305639 );
nand ( n15213 , n15203 , n305640 );
buf ( n305642 , n15213 );
buf ( n305643 , n305642 );
nand ( n305644 , n305630 , n305643 );
buf ( n305645 , n305644 );
buf ( n305646 , n305645 );
xor ( n15219 , n305617 , n305646 );
buf ( n15220 , n305338 );
not ( n305649 , n15220 );
buf ( n305650 , n305649 );
buf ( n305651 , n305650 );
buf ( n305652 , n876 );
buf ( n15225 , n14447 );
and ( n15226 , n305652 , n15225 );
not ( n305655 , n305652 );
buf ( n305656 , n859 );
and ( n15229 , n305655 , n305656 );
nor ( n305658 , n15226 , n15229 );
buf ( n305659 , n305658 );
buf ( n305660 , n305659 );
or ( n15233 , n305651 , n305660 );
buf ( n305662 , n305334 );
not ( n15235 , n305662 );
buf ( n305664 , n15235 );
buf ( n305665 , n305664 );
buf ( n305666 , n876 );
buf ( n305667 , n305060 );
and ( n305668 , n305666 , n305667 );
not ( n15241 , n305666 );
buf ( n305670 , n858 );
and ( n305671 , n15241 , n305670 );
nor ( n15244 , n305668 , n305671 );
buf ( n15245 , n15244 );
buf ( n305674 , n15245 );
or ( n15247 , n305665 , n305674 );
nand ( n305676 , n15233 , n15247 );
buf ( n305677 , n305676 );
buf ( n305678 , n305677 );
and ( n15251 , n15219 , n305678 );
and ( n15252 , n305617 , n305646 );
or ( n305681 , n15251 , n15252 );
buf ( n305682 , n305681 );
buf ( n305683 , n305682 );
and ( n305684 , n15161 , n305683 );
and ( n305685 , n305542 , n15160 );
or ( n15258 , n305684 , n305685 );
buf ( n305687 , n15258 );
buf ( n305688 , n305687 );
buf ( n305689 , n304763 );
buf ( n305690 , n863 );
and ( n305691 , n305689 , n305690 );
buf ( n305692 , n305691 );
buf ( n305693 , n305692 );
buf ( n305694 , n888 );
buf ( n305695 , n846 );
xor ( n305696 , n305694 , n305695 );
buf ( n305697 , n305696 );
not ( n15270 , n305697 );
not ( n305699 , n305138 );
or ( n305700 , n15270 , n305699 );
buf ( n305701 , n888 );
buf ( n305702 , n845 );
xnor ( n305703 , n305701 , n305702 );
buf ( n305704 , n305703 );
or ( n15277 , n305704 , n305130 );
nand ( n15278 , n305700 , n15277 );
buf ( n305707 , n15278 );
xor ( n305708 , n305693 , n305707 );
buf ( n305709 , n305580 );
not ( n15282 , n305709 );
buf ( n305711 , n15282 );
buf ( n305712 , n305711 );
not ( n305713 , n305712 );
buf ( n305714 , n14272 );
not ( n15287 , n305714 );
or ( n15288 , n305713 , n15287 );
buf ( n305717 , n304686 );
buf ( n305718 , n304694 );
nand ( n305719 , n305717 , n305718 );
buf ( n305720 , n305719 );
buf ( n305721 , n305720 );
nand ( n305722 , n15288 , n305721 );
buf ( n305723 , n305722 );
buf ( n305724 , n305723 );
and ( n305725 , n305708 , n305724 );
and ( n15298 , n305693 , n305707 );
or ( n305727 , n305725 , n15298 );
buf ( n305728 , n305727 );
buf ( n15301 , n305728 );
buf ( n305730 , n304845 );
buf ( n305731 , n872 );
buf ( n305732 , n861 );
and ( n305733 , n305731 , n305732 );
not ( n305734 , n305731 );
buf ( n305735 , n304771 );
and ( n15308 , n305734 , n305735 );
nor ( n15309 , n305733 , n15308 );
buf ( n305738 , n15309 );
buf ( n305739 , n305738 );
nand ( n305740 , n305730 , n305739 );
buf ( n305741 , n305740 );
buf ( n305742 , n872 );
buf ( n305743 , n862 );
and ( n305744 , n305742 , n305743 );
not ( n305745 , n305742 );
buf ( n305746 , n304739 );
and ( n305747 , n305745 , n305746 );
nor ( n305748 , n305744 , n305747 );
buf ( n305749 , n305748 );
nand ( n305750 , n305749 , n304851 );
nand ( n305751 , n305741 , n305750 );
buf ( n305752 , n305751 );
buf ( n305753 , n884 );
buf ( n305754 , n850 );
and ( n15327 , n305753 , n305754 );
not ( n15328 , n305753 );
buf ( n305757 , n304565 );
and ( n15330 , n15328 , n305757 );
nor ( n15331 , n15327 , n15330 );
buf ( n305760 , n15331 );
buf ( n305761 , n305760 );
not ( n305762 , n305761 );
buf ( n305763 , n304813 );
not ( n305764 , n305763 );
or ( n305765 , n305762 , n305764 );
buf ( n305766 , n884 );
buf ( n305767 , n849 );
xnor ( n15340 , n305766 , n305767 );
buf ( n15341 , n15340 );
buf ( n305770 , n15341 );
not ( n305771 , n305770 );
buf ( n15344 , n304807 );
nand ( n15345 , n305771 , n15344 );
buf ( n15346 , n15345 );
buf ( n305775 , n15346 );
nand ( n15348 , n305765 , n305775 );
buf ( n15349 , n15348 );
buf ( n305778 , n15349 );
xor ( n15351 , n305752 , n305778 );
buf ( n305780 , n890 );
buf ( n305781 , n843 );
and ( n15354 , n305780 , n305781 );
not ( n305783 , n305780 );
buf ( n305784 , n305117 );
and ( n15357 , n305783 , n305784 );
nor ( n305786 , n15354 , n15357 );
buf ( n305787 , n305786 );
buf ( n305788 , n305787 );
not ( n305789 , n305788 );
buf ( n305790 , n304658 );
not ( n305791 , n305790 );
or ( n15364 , n305789 , n305791 );
buf ( n305793 , n890 );
not ( n15366 , n305793 );
buf ( n305795 , n844 );
nor ( n305796 , n15366 , n305795 );
buf ( n305797 , n305796 );
buf ( n305798 , n305797 );
buf ( n305799 , n844 );
not ( n305800 , n305799 );
buf ( n15373 , n890 );
nor ( n15374 , n305800 , n15373 );
buf ( n15375 , n15374 );
buf ( n305804 , n15375 );
nor ( n15377 , n305798 , n305804 );
buf ( n15378 , n15377 );
buf ( n305807 , n15378 );
not ( n15380 , n305807 );
buf ( n305809 , n304633 );
nand ( n15382 , n15380 , n305809 );
buf ( n305811 , n15382 );
buf ( n305812 , n305811 );
nand ( n15385 , n15364 , n305812 );
buf ( n305814 , n15385 );
buf ( n305815 , n305814 );
and ( n305816 , n15351 , n305815 );
and ( n15389 , n305752 , n305778 );
or ( n305818 , n305816 , n15389 );
buf ( n305819 , n305818 );
buf ( n305820 , n305819 );
xor ( n305821 , n15301 , n305820 );
buf ( n305822 , n870 );
buf ( n305823 , n863 );
and ( n305824 , n305822 , n305823 );
not ( n305825 , n305822 );
buf ( n305826 , n305192 );
and ( n305827 , n305825 , n305826 );
nor ( n305828 , n305824 , n305827 );
buf ( n305829 , n305828 );
buf ( n305830 , n305829 );
not ( n15403 , n305830 );
buf ( n305832 , n14323 );
not ( n305833 , n305832 );
or ( n305834 , n15403 , n305833 );
buf ( n305835 , n304763 );
buf ( n305836 , n304743 );
nand ( n305837 , n305835 , n305836 );
buf ( n305838 , n305837 );
buf ( n305839 , n305838 );
nand ( n305840 , n305834 , n305839 );
buf ( n305841 , n305840 );
buf ( n305842 , n305841 );
buf ( n305843 , n305787 );
not ( n305844 , n305843 );
buf ( n305845 , n304633 );
not ( n15418 , n305845 );
or ( n305847 , n305844 , n15418 );
buf ( n305848 , n304658 );
buf ( n305849 , n304614 );
nand ( n305850 , n305848 , n305849 );
buf ( n305851 , n305850 );
buf ( n305852 , n305851 );
nand ( n15425 , n305847 , n305852 );
buf ( n15426 , n15425 );
buf ( n15427 , n15426 );
xor ( n15428 , n305842 , n15427 );
buf ( n305857 , n304581 );
buf ( n305858 , n305537 );
or ( n15431 , n305857 , n305858 );
buf ( n305860 , n14959 );
buf ( n305861 , n304569 );
not ( n15434 , n305861 );
buf ( n305863 , n15434 );
buf ( n305864 , n305863 );
or ( n305865 , n305860 , n305864 );
nand ( n15438 , n15431 , n305865 );
buf ( n305867 , n15438 );
buf ( n305868 , n305867 );
xor ( n305869 , n15428 , n305868 );
buf ( n305870 , n305869 );
buf ( n305871 , n305870 );
xor ( n305872 , n305821 , n305871 );
buf ( n305873 , n305872 );
buf ( n305874 , n305873 );
xor ( n305875 , n305688 , n305874 );
xor ( n305876 , n305693 , n305707 );
xor ( n15449 , n305876 , n305724 );
buf ( n305878 , n15449 );
buf ( n305879 , n305878 );
not ( n15452 , n895 );
nand ( n305881 , n15452 , n894 );
buf ( n305882 , n305881 );
buf ( n305883 , n840 );
buf ( n305884 , n894 );
xor ( n305885 , n305883 , n305884 );
buf ( n305886 , n305885 );
buf ( n305887 , n305886 );
not ( n305888 , n305887 );
buf ( n305889 , n305888 );
buf ( n305890 , n305889 );
or ( n15463 , n305882 , n305890 );
xor ( n305892 , n894 , n839 );
buf ( n305893 , n305892 );
not ( n15466 , n305893 );
buf ( n15467 , n15466 );
buf ( n15468 , n15467 );
not ( n15469 , n895 );
buf ( n305898 , n15469 );
or ( n305899 , n15468 , n305898 );
nand ( n305900 , n15463 , n305899 );
buf ( n305901 , n305900 );
buf ( n305902 , n305901 );
buf ( n305903 , n305639 );
not ( n15476 , n305903 );
buf ( n305905 , n305627 );
not ( n305906 , n305905 );
or ( n305907 , n15476 , n305906 );
buf ( n305908 , n874 );
not ( n305909 , n305908 );
buf ( n15482 , n859 );
nor ( n15483 , n305909 , n15482 );
buf ( n15484 , n15483 );
buf ( n305913 , n15484 );
buf ( n305914 , n859 );
not ( n305915 , n305914 );
buf ( n15488 , n874 );
nor ( n15489 , n305915 , n15488 );
buf ( n305918 , n15489 );
buf ( n305919 , n305918 );
nor ( n305920 , n305913 , n305919 );
buf ( n305921 , n305920 );
buf ( n305922 , n305921 );
not ( n305923 , n305922 );
buf ( n15496 , n305301 );
nand ( n15497 , n305923 , n15496 );
buf ( n15498 , n15497 );
buf ( n15499 , n15498 );
nand ( n15500 , n305907 , n15499 );
buf ( n15501 , n15500 );
buf ( n305930 , n15501 );
xor ( n15503 , n305902 , n305930 );
buf ( n305932 , n305650 );
buf ( n305933 , n15245 );
or ( n305934 , n305932 , n305933 );
buf ( n305935 , n305664 );
buf ( n305936 , n876 );
buf ( n15509 , n857 );
not ( n15510 , n15509 );
buf ( n305939 , n15510 );
buf ( n305940 , n305939 );
and ( n15513 , n305936 , n305940 );
not ( n305942 , n305936 );
buf ( n305943 , n857 );
and ( n15516 , n305942 , n305943 );
nor ( n305945 , n15513 , n15516 );
buf ( n305946 , n305945 );
buf ( n305947 , n305946 );
or ( n15520 , n305935 , n305947 );
nand ( n15521 , n305934 , n15520 );
buf ( n305950 , n15521 );
buf ( n305951 , n305950 );
xor ( n305952 , n15503 , n305951 );
buf ( n305953 , n305952 );
buf ( n305954 , n305953 );
xor ( n305955 , n305879 , n305954 );
buf ( n305956 , n880 );
buf ( n305957 , n854 );
xor ( n15530 , n305956 , n305957 );
buf ( n305959 , n15530 );
buf ( n305960 , n305959 );
not ( n305961 , n305960 );
buf ( n305962 , n304984 );
not ( n305963 , n305962 );
or ( n15536 , n305961 , n305963 );
buf ( n305965 , n304997 );
buf ( n305966 , n880 );
buf ( n305967 , n853 );
and ( n305968 , n305966 , n305967 );
not ( n15541 , n305966 );
buf ( n305970 , n304956 );
and ( n305971 , n15541 , n305970 );
nor ( n15544 , n305968 , n305971 );
buf ( n305973 , n15544 );
buf ( n305974 , n305973 );
nand ( n15547 , n305965 , n305974 );
buf ( n305976 , n15547 );
buf ( n305977 , n305976 );
nand ( n15550 , n15536 , n305977 );
buf ( n305979 , n15550 );
buf ( n305980 , n305979 );
buf ( n305981 , n305610 );
not ( n305982 , n305981 );
buf ( n305983 , n304912 );
not ( n305984 , n305983 );
or ( n15557 , n305982 , n305984 );
buf ( n15558 , n304901 );
buf ( n305987 , n847 );
buf ( n305988 , n886 );
and ( n15561 , n305987 , n305988 );
not ( n15562 , n305987 );
buf ( n305991 , n886 );
not ( n305992 , n305991 );
buf ( n305993 , n305992 );
buf ( n305994 , n305993 );
and ( n15567 , n15562 , n305994 );
nor ( n305996 , n15561 , n15567 );
buf ( n305997 , n305996 );
buf ( n15570 , n305997 );
nand ( n15571 , n15558 , n15570 );
buf ( n15572 , n15571 );
buf ( n306001 , n15572 );
nand ( n15574 , n15557 , n306001 );
buf ( n15575 , n15574 );
buf ( n306004 , n15575 );
xor ( n306005 , n305980 , n306004 );
buf ( n306006 , n304941 );
buf ( n306007 , n878 );
buf ( n306008 , n856 );
not ( n15581 , n306008 );
buf ( n15582 , n15581 );
buf ( n306011 , n15582 );
and ( n306012 , n306007 , n306011 );
not ( n306013 , n306007 );
buf ( n306014 , n856 );
and ( n306015 , n306013 , n306014 );
nor ( n306016 , n306012 , n306015 );
buf ( n306017 , n306016 );
buf ( n306018 , n306017 );
or ( n306019 , n306006 , n306018 );
buf ( n306020 , n878 );
buf ( n306021 , n855 );
and ( n15594 , n306020 , n306021 );
not ( n15595 , n306020 );
buf ( n306024 , n305319 );
and ( n306025 , n15595 , n306024 );
nor ( n306026 , n15594 , n306025 );
buf ( n306027 , n306026 );
buf ( n306028 , n306027 );
not ( n306029 , n306028 );
buf ( n306030 , n306029 );
buf ( n306031 , n306030 );
buf ( n306032 , n14523 );
or ( n15605 , n306031 , n306032 );
nand ( n15606 , n306019 , n15605 );
buf ( n306035 , n15606 );
buf ( n306036 , n306035 );
xor ( n306037 , n306005 , n306036 );
buf ( n306038 , n306037 );
buf ( n306039 , n306038 );
and ( n306040 , n305955 , n306039 );
and ( n15613 , n305879 , n305954 );
or ( n306042 , n306040 , n15613 );
buf ( n306043 , n306042 );
buf ( n306044 , n306043 );
and ( n306045 , n305875 , n306044 );
and ( n306046 , n305688 , n305874 );
or ( n15619 , n306045 , n306046 );
buf ( n306048 , n15619 );
buf ( n306049 , n306048 );
buf ( n306050 , n880 );
buf ( n306051 , n855 );
xor ( n15624 , n306050 , n306051 );
buf ( n15625 , n15624 );
buf ( n306054 , n15625 );
not ( n15627 , n306054 );
buf ( n306056 , n305098 );
not ( n306057 , n306056 );
or ( n15630 , n15627 , n306057 );
buf ( n306059 , n304997 );
buf ( n306060 , n305959 );
nand ( n15633 , n306059 , n306060 );
buf ( n306062 , n15633 );
buf ( n306063 , n306062 );
nand ( n306064 , n15630 , n306063 );
buf ( n306065 , n306064 );
buf ( n306066 , n306065 );
buf ( n306067 , n847 );
buf ( n306068 , n888 );
xor ( n306069 , n306067 , n306068 );
buf ( n306070 , n306069 );
buf ( n306071 , n306070 );
not ( n15644 , n306071 );
buf ( n306073 , n305138 );
not ( n15646 , n306073 );
or ( n15647 , n15644 , n15646 );
buf ( n306076 , n305144 );
buf ( n306077 , n305697 );
nand ( n306078 , n306076 , n306077 );
buf ( n306079 , n306078 );
buf ( n306080 , n306079 );
nand ( n15653 , n15647 , n306080 );
buf ( n306082 , n15653 );
buf ( n306083 , n306082 );
xor ( n15656 , n306066 , n306083 );
buf ( n306085 , n304938 );
buf ( n15658 , n878 );
buf ( n306087 , n857 );
xnor ( n15660 , n15658 , n306087 );
buf ( n306089 , n15660 );
buf ( n306090 , n306089 );
or ( n306091 , n306085 , n306090 );
buf ( n306092 , n14523 );
buf ( n306093 , n306017 );
or ( n15666 , n306092 , n306093 );
nand ( n15667 , n306091 , n15666 );
buf ( n306096 , n15667 );
buf ( n306097 , n306096 );
and ( n306098 , n15656 , n306097 );
and ( n306099 , n306066 , n306083 );
or ( n15672 , n306098 , n306099 );
buf ( n306101 , n15672 );
buf ( n306102 , n306101 );
buf ( n15675 , n841 );
buf ( n306104 , n894 );
xor ( n306105 , n15675 , n306104 );
buf ( n306106 , n306105 );
buf ( n306107 , n306106 );
not ( n306108 , n306107 );
buf ( n306109 , n305032 );
not ( n306110 , n306109 );
or ( n15683 , n306108 , n306110 );
buf ( n306112 , n305886 );
buf ( n306113 , n895 );
nand ( n15686 , n306112 , n306113 );
buf ( n306115 , n15686 );
buf ( n306116 , n306115 );
nand ( n306117 , n15683 , n306116 );
buf ( n306118 , n306117 );
buf ( n306119 , n872 );
buf ( n306120 , n863 );
and ( n306121 , n306119 , n306120 );
not ( n15694 , n306119 );
buf ( n306123 , n305192 );
and ( n15696 , n15694 , n306123 );
nor ( n15697 , n306121 , n15696 );
buf ( n306126 , n15697 );
buf ( n306127 , n306126 );
not ( n15700 , n306127 );
buf ( n306129 , n304843 );
buf ( n306130 , n304845 );
nor ( n306131 , n306129 , n306130 );
buf ( n306132 , n306131 );
buf ( n306133 , n306132 );
not ( n306134 , n306133 );
or ( n15707 , n15700 , n306134 );
buf ( n306136 , n304864 );
buf ( n306137 , n305749 );
nand ( n15710 , n306136 , n306137 );
buf ( n306139 , n15710 );
buf ( n306140 , n306139 );
nand ( n306141 , n15707 , n306140 );
buf ( n306142 , n306141 );
xor ( n15715 , n306118 , n306142 );
buf ( n306144 , n845 );
buf ( n15717 , n890 );
xor ( n15718 , n306144 , n15717 );
buf ( n306147 , n15718 );
buf ( n306148 , n306147 );
not ( n15721 , n306148 );
buf ( n306150 , n304630 );
not ( n306151 , n306150 );
buf ( n306152 , n306151 );
buf ( n306153 , n306152 );
not ( n306154 , n306153 );
or ( n306155 , n15721 , n306154 );
buf ( n306156 , n15378 );
not ( n15729 , n306156 );
buf ( n306158 , n304658 );
nand ( n15731 , n15729 , n306158 );
buf ( n306160 , n15731 );
buf ( n306161 , n306160 );
nand ( n15734 , n306155 , n306161 );
buf ( n306163 , n15734 );
and ( n15736 , n15715 , n306163 );
and ( n306165 , n306118 , n306142 );
or ( n15738 , n15736 , n306165 );
buf ( n306167 , n15738 );
xor ( n15740 , n306102 , n306167 );
xor ( n15741 , n305752 , n305778 );
xor ( n15742 , n15741 , n305815 );
buf ( n306171 , n15742 );
buf ( n306172 , n306171 );
and ( n306173 , n15740 , n306172 );
and ( n15746 , n306102 , n306167 );
or ( n15747 , n306173 , n15746 );
buf ( n306176 , n15747 );
buf ( n306177 , n306176 );
xor ( n306178 , n304682 , n304726 );
buf ( n306179 , n306178 );
buf ( n306180 , n306179 );
xor ( n15753 , n305980 , n306004 );
and ( n15754 , n15753 , n306036 );
and ( n15755 , n305980 , n306004 );
or ( n15756 , n15754 , n15755 );
buf ( n15757 , n15756 );
buf ( n306186 , n15757 );
xor ( n15759 , n306180 , n306186 );
xor ( n306188 , n305902 , n305930 );
and ( n306189 , n306188 , n305951 );
and ( n15762 , n305902 , n305930 );
or ( n306191 , n306189 , n15762 );
buf ( n306192 , n306191 );
buf ( n306193 , n306192 );
xor ( n306194 , n15759 , n306193 );
buf ( n306195 , n306194 );
buf ( n306196 , n306195 );
xor ( n15769 , n306177 , n306196 );
buf ( n306198 , n305892 );
not ( n15771 , n306198 );
buf ( n306200 , n305032 );
not ( n306201 , n306200 );
or ( n306202 , n15771 , n306201 );
buf ( n306203 , n838 );
buf ( n306204 , n894 );
xor ( n306205 , n306203 , n306204 );
buf ( n306206 , n306205 );
buf ( n306207 , n306206 );
buf ( n306208 , n895 );
nand ( n306209 , n306207 , n306208 );
buf ( n306210 , n306209 );
buf ( n306211 , n306210 );
nand ( n306212 , n306202 , n306211 );
buf ( n306213 , n306212 );
buf ( n306214 , n306213 );
buf ( n306215 , n305738 );
not ( n306216 , n306215 );
buf ( n306217 , n304851 );
not ( n306218 , n306217 );
or ( n306219 , n306216 , n306218 );
buf ( n306220 , n304859 );
not ( n15793 , n306220 );
buf ( n306222 , n304864 );
nand ( n306223 , n15793 , n306222 );
buf ( n306224 , n306223 );
buf ( n306225 , n306224 );
nand ( n306226 , n306219 , n306225 );
buf ( n306227 , n306226 );
buf ( n306228 , n306227 );
xor ( n306229 , n306214 , n306228 );
buf ( n306230 , n304813 );
not ( n15803 , n306230 );
buf ( n15804 , n15803 );
buf ( n306233 , n15804 );
buf ( n306234 , n15341 );
or ( n306235 , n306233 , n306234 );
buf ( n15808 , n304819 );
not ( n15809 , n15808 );
buf ( n306238 , n15809 );
buf ( n306239 , n306238 );
buf ( n306240 , n304793 );
or ( n306241 , n306239 , n306240 );
nand ( n306242 , n306235 , n306241 );
buf ( n306243 , n306242 );
buf ( n306244 , n306243 );
xor ( n306245 , n306229 , n306244 );
buf ( n306246 , n306245 );
buf ( n306247 , n306246 );
buf ( n306248 , n305973 );
not ( n306249 , n306248 );
buf ( n306250 , n304984 );
not ( n306251 , n306250 );
or ( n306252 , n306249 , n306251 );
buf ( n306253 , n14564 );
not ( n306254 , n306253 );
buf ( n306255 , n304973 );
nand ( n15828 , n306254 , n306255 );
buf ( n306257 , n15828 );
buf ( n306258 , n306257 );
nand ( n306259 , n306252 , n306258 );
buf ( n306260 , n306259 );
buf ( n306261 , n306260 );
buf ( n306262 , n306027 );
not ( n306263 , n306262 );
not ( n15836 , n304941 );
buf ( n306265 , n15836 );
not ( n306266 , n306265 );
or ( n306267 , n306263 , n306266 );
buf ( n306268 , n304946 );
not ( n15841 , n306268 );
buf ( n306270 , n14523 );
not ( n306271 , n306270 );
buf ( n306272 , n306271 );
buf ( n306273 , n306272 );
nand ( n306274 , n15841 , n306273 );
buf ( n306275 , n306274 );
buf ( n306276 , n306275 );
nand ( n15849 , n306267 , n306276 );
buf ( n306278 , n15849 );
buf ( n306279 , n306278 );
xor ( n306280 , n306261 , n306279 );
buf ( n306281 , n305138 );
not ( n306282 , n306281 );
buf ( n306283 , n306282 );
buf ( n306284 , n306283 );
buf ( n306285 , n305704 );
or ( n306286 , n306284 , n306285 );
buf ( n306287 , n305144 );
not ( n15860 , n306287 );
buf ( n15861 , n15860 );
buf ( n306290 , n15861 );
buf ( n306291 , n305465 );
or ( n306292 , n306290 , n306291 );
nand ( n306293 , n306286 , n306292 );
buf ( n306294 , n306293 );
buf ( n306295 , n306294 );
xor ( n306296 , n306280 , n306295 );
buf ( n306297 , n306296 );
buf ( n306298 , n306297 );
xor ( n306299 , n306247 , n306298 );
buf ( n306300 , n305997 );
not ( n306301 , n306300 );
buf ( n15874 , n304912 );
not ( n15875 , n15874 );
or ( n15876 , n306301 , n15875 );
buf ( n15877 , n304901 );
buf ( n306306 , n304895 );
nand ( n306307 , n15877 , n306306 );
buf ( n306308 , n306307 );
buf ( n306309 , n306308 );
nand ( n306310 , n15876 , n306309 );
buf ( n306311 , n306310 );
buf ( n306312 , n306311 );
buf ( n306313 , n305946 );
not ( n15886 , n306313 );
buf ( n15887 , n15886 );
buf ( n306316 , n15887 );
not ( n15889 , n306316 );
buf ( n306318 , n305338 );
not ( n15891 , n306318 );
or ( n306320 , n15889 , n15891 );
buf ( n306321 , n876 );
buf ( n306322 , n856 );
and ( n306323 , n306321 , n306322 );
not ( n306324 , n306321 );
buf ( n306325 , n15582 );
and ( n15898 , n306324 , n306325 );
nor ( n306327 , n306323 , n15898 );
buf ( n306328 , n306327 );
buf ( n306329 , n306328 );
buf ( n306330 , n305344 );
nand ( n306331 , n306329 , n306330 );
buf ( n306332 , n306331 );
buf ( n306333 , n306332 );
nand ( n306334 , n306320 , n306333 );
buf ( n306335 , n306334 );
buf ( n306336 , n306335 );
xor ( n306337 , n306312 , n306336 );
buf ( n306338 , n305627 );
not ( n306339 , n306338 );
buf ( n306340 , n306339 );
buf ( n306341 , n306340 );
buf ( n306342 , n305921 );
or ( n306343 , n306341 , n306342 );
buf ( n306344 , n305289 );
not ( n306345 , n306344 );
buf ( n306346 , n306345 );
buf ( n306347 , n306346 );
buf ( n306348 , n874 );
buf ( n306349 , n858 );
and ( n15922 , n306348 , n306349 );
not ( n306351 , n306348 );
buf ( n306352 , n305060 );
and ( n15925 , n306351 , n306352 );
nor ( n15926 , n15922 , n15925 );
buf ( n306355 , n15926 );
buf ( n15928 , n306355 );
not ( n15929 , n15928 );
buf ( n15930 , n15929 );
buf ( n306359 , n15930 );
or ( n15932 , n306347 , n306359 );
nand ( n306361 , n306343 , n15932 );
buf ( n306362 , n306361 );
buf ( n306363 , n306362 );
xor ( n306364 , n306337 , n306363 );
buf ( n306365 , n306364 );
buf ( n306366 , n306365 );
xor ( n306367 , n306299 , n306366 );
buf ( n306368 , n306367 );
buf ( n306369 , n306368 );
and ( n15942 , n15769 , n306369 );
and ( n15943 , n306177 , n306196 );
or ( n15944 , n15942 , n15943 );
buf ( n306373 , n15944 );
buf ( n306374 , n306373 );
xor ( n306375 , n306049 , n306374 );
xor ( n15948 , n306180 , n306186 );
and ( n306377 , n15948 , n306193 );
and ( n15950 , n306180 , n306186 );
or ( n306379 , n306377 , n15950 );
buf ( n306380 , n306379 );
buf ( n306381 , n306380 );
xor ( n15954 , n15301 , n305820 );
and ( n15955 , n15954 , n305871 );
and ( n306384 , n15301 , n305820 );
or ( n15957 , n15955 , n306384 );
buf ( n306386 , n15957 );
buf ( n306387 , n306386 );
xor ( n15960 , n306381 , n306387 );
xor ( n306389 , n306247 , n306298 );
and ( n306390 , n306389 , n306366 );
and ( n306391 , n306247 , n306298 );
or ( n15964 , n306390 , n306391 );
buf ( n306393 , n15964 );
buf ( n306394 , n306393 );
xor ( n15967 , n15960 , n306394 );
buf ( n306396 , n15967 );
buf ( n306397 , n306396 );
and ( n306398 , n306375 , n306397 );
and ( n15971 , n306049 , n306374 );
or ( n306400 , n306398 , n15971 );
buf ( n306401 , n306400 );
buf ( n306402 , n306401 );
xor ( n306403 , n15083 , n306402 );
xor ( n306404 , n306214 , n306228 );
and ( n15977 , n306404 , n306244 );
and ( n306406 , n306214 , n306228 );
or ( n306407 , n15977 , n306406 );
buf ( n306408 , n306407 );
buf ( n306409 , n306408 );
xor ( n306410 , n306261 , n306279 );
and ( n15983 , n306410 , n306295 );
and ( n15984 , n306261 , n306279 );
or ( n306413 , n15983 , n15984 );
buf ( n306414 , n306413 );
buf ( n15987 , n306414 );
xor ( n15988 , n306409 , n15987 );
xor ( n306417 , n306312 , n306336 );
and ( n306418 , n306417 , n306363 );
and ( n15991 , n306312 , n306336 );
or ( n306420 , n306418 , n15991 );
buf ( n306421 , n306420 );
buf ( n306422 , n306421 );
and ( n306423 , n15988 , n306422 );
and ( n306424 , n306409 , n15987 );
or ( n15997 , n306423 , n306424 );
buf ( n306426 , n15997 );
buf ( n306427 , n306426 );
buf ( n306428 , n306206 );
not ( n306429 , n306428 );
buf ( n306430 , n305032 );
not ( n16003 , n306430 );
or ( n306432 , n306429 , n16003 );
buf ( n306433 , n305022 );
buf ( n306434 , n895 );
nand ( n306435 , n306433 , n306434 );
buf ( n306436 , n306435 );
buf ( n306437 , n306436 );
nand ( n306438 , n306432 , n306437 );
buf ( n306439 , n306438 );
buf ( n306440 , n306439 );
buf ( n306441 , n306355 );
not ( n306442 , n306441 );
buf ( n306443 , n305627 );
not ( n16016 , n306443 );
or ( n306445 , n306442 , n16016 );
buf ( n306446 , n305301 );
buf ( n306447 , n14853 );
nand ( n16020 , n306446 , n306447 );
buf ( n16021 , n16020 );
buf ( n306450 , n16021 );
nand ( n16023 , n306445 , n306450 );
buf ( n306452 , n16023 );
buf ( n16025 , n306452 );
xor ( n16026 , n306440 , n16025 );
buf ( n306455 , n306328 );
not ( n306456 , n306455 );
buf ( n306457 , n305338 );
not ( n306458 , n306457 );
or ( n306459 , n306456 , n306458 );
buf ( n306460 , n305344 );
buf ( n306461 , n305323 );
nand ( n306462 , n306460 , n306461 );
buf ( n306463 , n306462 );
buf ( n306464 , n306463 );
nand ( n306465 , n306459 , n306464 );
buf ( n306466 , n306465 );
buf ( n306467 , n306466 );
xor ( n16040 , n16026 , n306467 );
buf ( n306469 , n16040 );
buf ( n306470 , n306469 );
xor ( n16043 , n305842 , n15427 );
and ( n306472 , n16043 , n305868 );
and ( n306473 , n305842 , n15427 );
or ( n16046 , n306472 , n306473 );
buf ( n306475 , n16046 );
buf ( n16048 , n306475 );
xor ( n16049 , n306470 , n16048 );
xor ( n306478 , n305454 , n305481 );
xor ( n16051 , n306478 , n305498 );
buf ( n306480 , n16051 );
buf ( n306481 , n306480 );
and ( n16054 , n16049 , n306481 );
and ( n306483 , n306470 , n16048 );
or ( n306484 , n16054 , n306483 );
buf ( n306485 , n306484 );
buf ( n306486 , n306485 );
xor ( n306487 , n306427 , n306486 );
xor ( n306488 , n306440 , n16025 );
and ( n16061 , n306488 , n306467 );
and ( n306490 , n306440 , n16025 );
or ( n306491 , n16061 , n306490 );
buf ( n306492 , n306491 );
buf ( n306493 , n306492 );
xor ( n306494 , n304928 , n304968 );
and ( n16067 , n306494 , n305013 );
and ( n306496 , n304928 , n304968 );
or ( n306497 , n16067 , n306496 );
buf ( n306498 , n306497 );
buf ( n306499 , n306498 );
xor ( n306500 , n306493 , n306499 );
xor ( n16073 , n304782 , n304838 );
and ( n306502 , n16073 , n304887 );
and ( n16075 , n304782 , n304838 );
or ( n16076 , n306502 , n16075 );
buf ( n306505 , n16076 );
buf ( n306506 , n306505 );
xor ( n16079 , n306500 , n306506 );
buf ( n306508 , n16079 );
buf ( n306509 , n306508 );
xor ( n16082 , n306487 , n306509 );
buf ( n306511 , n16082 );
buf ( n306512 , n306511 );
xor ( n16085 , n306381 , n306387 );
and ( n306514 , n16085 , n306394 );
and ( n16087 , n306381 , n306387 );
or ( n16088 , n306514 , n16087 );
buf ( n306517 , n16088 );
buf ( n306518 , n306517 );
xor ( n16091 , n306512 , n306518 );
xor ( n306520 , n306409 , n15987 );
xor ( n16093 , n306520 , n306422 );
buf ( n306522 , n16093 );
buf ( n306523 , n306522 );
xor ( n16096 , n306470 , n16048 );
xor ( n306525 , n16096 , n306481 );
buf ( n306526 , n306525 );
buf ( n306527 , n306526 );
xor ( n16100 , n306523 , n306527 );
xor ( n16101 , n304732 , n304890 );
xor ( n16102 , n16101 , n305016 );
buf ( n306531 , n16102 );
buf ( n306532 , n306531 );
and ( n306533 , n16100 , n306532 );
and ( n16106 , n306523 , n306527 );
or ( n16107 , n306533 , n16106 );
buf ( n306536 , n16107 );
buf ( n306537 , n306536 );
xor ( n16110 , n16091 , n306537 );
buf ( n306539 , n16110 );
buf ( n306540 , n306539 );
xor ( n16113 , n306403 , n306540 );
buf ( n306542 , n16113 );
buf ( n306543 , n306542 );
xor ( n306544 , n13155 , n303943 );
xor ( n16117 , n306544 , n303947 );
buf ( n306546 , n16117 );
xor ( n306547 , n300211 , n9358 );
xor ( n16120 , n306547 , n9423 );
buf ( n306549 , n299317 );
not ( n16122 , n306549 );
buf ( n306551 , n299380 );
not ( n16124 , n306551 );
or ( n16125 , n16122 , n16124 );
buf ( n306554 , n299317 );
buf ( n306555 , n299380 );
or ( n16128 , n306554 , n306555 );
nand ( n306557 , n16125 , n16128 );
buf ( n306558 , n306557 );
buf ( n306559 , n306558 );
buf ( n306560 , n299444 );
and ( n306561 , n306559 , n306560 );
not ( n306562 , n306559 );
buf ( n306563 , n299444 );
not ( n306564 , n306563 );
buf ( n306565 , n306564 );
buf ( n306566 , n306565 );
and ( n306567 , n306562 , n306566 );
nor ( n306568 , n306561 , n306567 );
buf ( n306569 , n306568 );
buf ( n306570 , n306569 );
xor ( n306571 , n9661 , n300146 );
xor ( n306572 , n306571 , n300202 );
buf ( n306573 , n306572 );
buf ( n306574 , n306573 );
xor ( n16147 , n306570 , n306574 );
not ( n16148 , n9509 );
and ( n306577 , n16148 , n299954 );
not ( n306578 , n16148 );
not ( n306579 , n299954 );
and ( n16152 , n306578 , n306579 );
nor ( n306581 , n306577 , n16152 );
buf ( n306582 , n299966 );
not ( n16155 , n306582 );
and ( n306584 , n306581 , n16155 );
not ( n306585 , n306581 );
and ( n16158 , n306585 , n306582 );
nor ( n306587 , n306584 , n16158 );
buf ( n306588 , n306587 );
xor ( n16161 , n300082 , n300065 );
xor ( n306590 , n16161 , n300049 );
buf ( n306591 , n306590 );
xor ( n306592 , n306588 , n306591 );
xor ( n16165 , n304485 , n304504 );
and ( n16166 , n16165 , n304510 );
and ( n306595 , n304485 , n304504 );
or ( n306596 , n16166 , n306595 );
buf ( n306597 , n306596 );
buf ( n306598 , n306597 );
and ( n306599 , n306592 , n306598 );
and ( n306600 , n306588 , n306591 );
or ( n16173 , n306599 , n306600 );
buf ( n306602 , n16173 );
buf ( n306603 , n306602 );
and ( n16176 , n16147 , n306603 );
and ( n306605 , n306570 , n306574 );
or ( n306606 , n16176 , n306605 );
buf ( n306607 , n306606 );
buf ( n306608 , n306607 );
xor ( n306609 , n303587 , n303602 );
xor ( n16182 , n306609 , n303785 );
buf ( n306611 , n16182 );
buf ( n306612 , n306611 );
xor ( n16185 , n306608 , n306612 );
xor ( n16186 , n303607 , n303611 );
xor ( n306615 , n16186 , n303780 );
buf ( n306616 , n306615 );
buf ( n306617 , n306616 );
xor ( n306618 , n304432 , n304441 );
and ( n306619 , n306618 , n304448 );
and ( n16192 , n304432 , n304441 );
or ( n16193 , n306619 , n16192 );
buf ( n306622 , n16193 );
buf ( n306623 , n306622 );
xor ( n306624 , n303797 , n303844 );
xor ( n306625 , n306624 , n303900 );
buf ( n306626 , n306625 );
buf ( n306627 , n306626 );
xor ( n16200 , n306623 , n306627 );
and ( n16201 , n13239 , n303775 );
not ( n16202 , n13239 );
not ( n306631 , n303775 );
and ( n306632 , n16202 , n306631 );
nor ( n16205 , n16201 , n306632 );
buf ( n306634 , n16205 );
buf ( n16207 , n303724 );
xor ( n16208 , n306634 , n16207 );
buf ( n306637 , n16208 );
buf ( n306638 , n306637 );
and ( n16211 , n16200 , n306638 );
and ( n16212 , n306623 , n306627 );
or ( n306641 , n16211 , n16212 );
buf ( n306642 , n306641 );
buf ( n306643 , n306642 );
xor ( n306644 , n306617 , n306643 );
xor ( n16217 , n304024 , n304028 );
and ( n306646 , n16217 , n304033 );
and ( n16219 , n304024 , n304028 );
or ( n306648 , n306646 , n16219 );
buf ( n306649 , n306648 );
buf ( n306650 , n306649 );
xor ( n306651 , n303909 , n303913 );
xor ( n306652 , n306651 , n303918 );
buf ( n306653 , n306652 );
buf ( n306654 , n306653 );
xor ( n306655 , n306650 , n306654 );
xor ( n16228 , n304524 , n304527 );
and ( n306657 , n16228 , n304531 );
and ( n306658 , n304524 , n304527 );
or ( n16231 , n306657 , n306658 );
buf ( n306660 , n16231 );
buf ( n306661 , n306660 );
and ( n16234 , n306655 , n306661 );
and ( n306663 , n306650 , n306654 );
or ( n16236 , n16234 , n306663 );
buf ( n306665 , n16236 );
buf ( n306666 , n306665 );
and ( n16239 , n306644 , n306666 );
and ( n306668 , n306617 , n306643 );
or ( n306669 , n16239 , n306668 );
buf ( n306670 , n306669 );
buf ( n306671 , n306670 );
and ( n306672 , n16185 , n306671 );
and ( n16245 , n306608 , n306612 );
or ( n306674 , n306672 , n16245 );
buf ( n306675 , n306674 );
xor ( n16248 , n16120 , n306675 );
xor ( n16249 , n303789 , n13363 );
xor ( n306678 , n16249 , n303939 );
and ( n16251 , n16248 , n306678 );
and ( n306680 , n16120 , n306675 );
or ( n16253 , n16251 , n306680 );
and ( n16254 , n306546 , n16253 );
xor ( n306683 , n303952 , n303956 );
buf ( n306684 , n306683 );
nor ( n306685 , n16254 , n306684 );
not ( n16258 , n306685 );
nand ( n16259 , n16254 , n306684 );
nand ( n306688 , n16258 , n16259 );
not ( n16261 , n306688 );
xor ( n306690 , n306588 , n306591 );
xor ( n16263 , n306690 , n306598 );
buf ( n306692 , n16263 );
buf ( n16265 , n306692 );
xor ( n306694 , n304451 , n304456 );
and ( n16267 , n306694 , n304463 );
and ( n306696 , n304451 , n304456 );
or ( n306697 , n16267 , n306696 );
buf ( n306698 , n306697 );
buf ( n306699 , n306698 );
xor ( n306700 , n16265 , n306699 );
xor ( n16273 , n304472 , n304513 );
and ( n16274 , n16273 , n304534 );
and ( n306703 , n304472 , n304513 );
or ( n306704 , n16274 , n306703 );
buf ( n306705 , n306704 );
buf ( n306706 , n306705 );
xor ( n306707 , n306700 , n306706 );
buf ( n306708 , n306707 );
buf ( n306709 , n306708 );
xor ( n306710 , n304466 , n304537 );
and ( n306711 , n306710 , n304546 );
and ( n16284 , n304466 , n304537 );
or ( n306713 , n306711 , n16284 );
buf ( n306714 , n306713 );
buf ( n306715 , n306714 );
xor ( n306716 , n306709 , n306715 );
xor ( n16289 , n306623 , n306627 );
xor ( n306718 , n16289 , n306638 );
buf ( n306719 , n306718 );
buf ( n306720 , n306719 );
xor ( n16293 , n306650 , n306654 );
xor ( n16294 , n16293 , n306661 );
buf ( n306723 , n16294 );
buf ( n306724 , n306723 );
xor ( n16297 , n306720 , n306724 );
xor ( n16298 , n304036 , n304139 );
and ( n16299 , n16298 , n304254 );
and ( n16300 , n304036 , n304139 );
or ( n16301 , n16299 , n16300 );
buf ( n306730 , n16301 );
buf ( n306731 , n306730 );
xor ( n306732 , n16297 , n306731 );
buf ( n306733 , n306732 );
buf ( n306734 , n306733 );
and ( n306735 , n306716 , n306734 );
and ( n16308 , n306709 , n306715 );
or ( n306737 , n306735 , n16308 );
buf ( n306738 , n306737 );
not ( n16311 , n306738 );
xor ( n16312 , n16265 , n306699 );
and ( n16313 , n16312 , n306706 );
and ( n306742 , n16265 , n306699 );
or ( n16315 , n16313 , n306742 );
buf ( n306744 , n16315 );
buf ( n16317 , n306744 );
xor ( n16318 , n306720 , n306724 );
and ( n306747 , n16318 , n306731 );
and ( n306748 , n306720 , n306724 );
or ( n306749 , n306747 , n306748 );
buf ( n306750 , n306749 );
buf ( n306751 , n306750 );
xor ( n306752 , n16317 , n306751 );
buf ( n16325 , n303794 );
not ( n306754 , n16325 );
buf ( n306755 , n303904 );
not ( n16328 , n306755 );
buf ( n306757 , n16328 );
and ( n16330 , n306757 , n303922 );
not ( n16331 , n306757 );
not ( n16332 , n303922 );
and ( n16333 , n16331 , n16332 );
nor ( n306762 , n16330 , n16333 );
not ( n306763 , n306762 );
or ( n306764 , n306754 , n306763 );
or ( n16337 , n306762 , n16325 );
nand ( n306766 , n306764 , n16337 );
buf ( n306767 , n306766 );
xor ( n16340 , n306570 , n306574 );
xor ( n306769 , n16340 , n306603 );
buf ( n306770 , n306769 );
buf ( n306771 , n306770 );
xor ( n16344 , n306767 , n306771 );
xor ( n306773 , n306617 , n306643 );
xor ( n306774 , n306773 , n306666 );
buf ( n306775 , n306774 );
buf ( n306776 , n306775 );
xor ( n306777 , n16344 , n306776 );
buf ( n306778 , n306777 );
buf ( n306779 , n306778 );
xor ( n306780 , n306752 , n306779 );
buf ( n306781 , n306780 );
not ( n16354 , n306781 );
not ( n306783 , n16354 );
or ( n16356 , n16311 , n306783 );
not ( n16357 , n306738 );
nand ( n16358 , n16357 , n306781 );
nand ( n16359 , n16356 , n16358 );
not ( n306788 , n16359 );
buf ( n306789 , n832 );
buf ( n306790 , n304553 );
xor ( n306791 , n306789 , n306790 );
xor ( n16364 , n306709 , n306715 );
xor ( n306793 , n16364 , n306734 );
buf ( n306794 , n306793 );
buf ( n306795 , n306794 );
and ( n306796 , n306791 , n306795 );
and ( n16369 , n306789 , n306790 );
or ( n306798 , n306796 , n16369 );
buf ( n306799 , n306798 );
not ( n306800 , n306799 );
nand ( n306801 , n306788 , n306800 );
not ( n16374 , n306801 );
xor ( n306803 , n16317 , n306751 );
and ( n306804 , n306803 , n306779 );
and ( n16377 , n16317 , n306751 );
or ( n306806 , n306804 , n16377 );
buf ( n306807 , n306806 );
not ( n16380 , n306807 );
xor ( n306809 , n303926 , n303930 );
xor ( n306810 , n306809 , n303935 );
buf ( n306811 , n306810 );
xor ( n16384 , n306767 , n306771 );
and ( n306813 , n16384 , n306776 );
and ( n306814 , n306767 , n306771 );
or ( n16387 , n306813 , n306814 );
buf ( n306816 , n16387 );
xor ( n306817 , n306811 , n306816 );
xor ( n16390 , n306608 , n306612 );
xor ( n306819 , n16390 , n306671 );
buf ( n306820 , n306819 );
xor ( n16393 , n306817 , n306820 );
not ( n306822 , n16393 );
not ( n306823 , n306822 );
or ( n16396 , n16380 , n306823 );
not ( n16397 , n306807 );
nand ( n306826 , n16397 , n16393 );
nand ( n306827 , n16396 , n306826 );
buf ( n306828 , n306781 );
buf ( n306829 , n306738 );
nand ( n306830 , n306828 , n306829 );
buf ( n306831 , n306830 );
not ( n306832 , n306831 );
nor ( n16405 , n306827 , n306832 );
nor ( n306834 , n16374 , n16405 );
xor ( n16407 , n306811 , n306816 );
and ( n306836 , n16407 , n306820 );
and ( n306837 , n306811 , n306816 );
or ( n16410 , n306836 , n306837 );
not ( n306839 , n16410 );
not ( n306840 , n306839 );
xor ( n16413 , n16120 , n306675 );
xor ( n306842 , n16413 , n306678 );
not ( n306843 , n306842 );
or ( n306844 , n306840 , n306843 );
not ( n306845 , n16410 );
or ( n16418 , n306842 , n306845 );
nand ( n306847 , n306844 , n16418 );
nand ( n306848 , n306807 , n16393 );
not ( n16421 , n306848 );
nor ( n306850 , n306847 , n16421 );
nand ( n16423 , n306842 , n16410 );
not ( n306852 , n16423 );
xor ( n16425 , n306546 , n16253 );
nor ( n16426 , n306852 , n16425 );
nor ( n306855 , n306850 , n16426 );
nand ( n306856 , n306834 , n306855 );
buf ( n16429 , n306856 );
not ( n306858 , n16429 );
not ( n306859 , n306858 );
xor ( n16432 , n838 , n294313 );
xor ( n306861 , n16432 , n294713 );
nor ( n16434 , n303966 , n306861 );
nand ( n16435 , n12994 , n13539 );
or ( n306864 , n16434 , n16435 );
nand ( n16437 , n306861 , n303966 );
nand ( n16438 , n306864 , n16437 );
not ( n16439 , n16438 );
xor ( n16440 , n836 , n303173 );
xor ( n306869 , n16440 , n12755 );
buf ( n306870 , n837 );
xor ( n16443 , n4147 , n294581 );
and ( n16444 , n16443 , n294711 );
and ( n16445 , n4147 , n294581 );
or ( n16446 , n16444 , n16445 );
buf ( n306875 , n16446 );
buf ( n306876 , n306875 );
xor ( n306877 , n306870 , n306876 );
xor ( n16450 , n303148 , n303153 );
xor ( n16451 , n16450 , n303169 );
buf ( n306880 , n16451 );
buf ( n306881 , n306880 );
and ( n306882 , n306877 , n306881 );
and ( n306883 , n306870 , n306876 );
or ( n16456 , n306882 , n306883 );
buf ( n306885 , n16456 );
nor ( n306886 , n306869 , n306885 );
xor ( n16459 , n306870 , n306876 );
xor ( n306888 , n16459 , n306881 );
buf ( n306889 , n306888 );
nor ( n306890 , n306889 , n303960 );
nor ( n16463 , n306886 , n306890 );
not ( n306892 , n16463 );
or ( n16465 , n16439 , n306892 );
not ( n16466 , n306886 );
nand ( n306895 , n306889 , n303960 );
not ( n306896 , n306895 );
and ( n306897 , n16466 , n306896 );
nand ( n16470 , n306885 , n306869 );
not ( n306899 , n16470 );
nor ( n306900 , n306897 , n306899 );
nand ( n16473 , n16465 , n306900 );
not ( n306902 , n16473 );
xor ( n306903 , n296086 , n5667 );
and ( n16476 , n306903 , n296340 );
and ( n306905 , n296086 , n5667 );
or ( n306906 , n16476 , n306905 );
buf ( n306907 , n306906 );
xor ( n306908 , n834 , n306907 );
xor ( n16481 , n296069 , n5645 );
and ( n306910 , n16481 , n296084 );
and ( n16483 , n296069 , n5645 );
or ( n16484 , n306910 , n16483 );
buf ( n306913 , n16484 );
xor ( n306914 , n296169 , n296321 );
and ( n306915 , n306914 , n296337 );
and ( n306916 , n296169 , n296321 );
or ( n16489 , n306915 , n306916 );
buf ( n306918 , n16489 );
buf ( n16491 , n306918 );
xor ( n16492 , n306913 , n16491 );
buf ( n306921 , n304266 );
buf ( n306922 , n13835 );
and ( n16495 , n306921 , n306922 );
not ( n306924 , n306921 );
buf ( n306925 , n304260 );
and ( n16498 , n306924 , n306925 );
nor ( n306927 , n16495 , n16498 );
buf ( n306928 , n306927 );
not ( n16501 , n304417 );
and ( n306930 , n306928 , n16501 );
not ( n306931 , n306928 );
and ( n16504 , n306931 , n304417 );
nor ( n306933 , n306930 , n16504 );
buf ( n306934 , n306933 );
xor ( n306935 , n16492 , n306934 );
buf ( n306936 , n306935 );
xor ( n306937 , n306908 , n306936 );
not ( n16510 , n306937 );
not ( n16511 , n296347 );
nand ( n306940 , n16510 , n16511 );
xor ( n306941 , n295153 , n295908 );
xor ( n306942 , n306941 , n296343 );
buf ( n306943 , n306942 );
not ( n306944 , n306943 );
not ( n306945 , n12758 );
nand ( n16518 , n306944 , n306945 );
and ( n306947 , n306940 , n16518 );
not ( n306948 , n306947 );
xor ( n16521 , n306789 , n306790 );
xor ( n306950 , n16521 , n306795 );
buf ( n306951 , n306950 );
not ( n306952 , n306951 );
xor ( n16525 , n306913 , n16491 );
and ( n306954 , n16525 , n306934 );
and ( n16527 , n306913 , n16491 );
or ( n16528 , n306954 , n16527 );
buf ( n306957 , n16528 );
xor ( n306958 , n833 , n306957 );
xor ( n306959 , n304257 , n304428 );
xor ( n16532 , n306959 , n304549 );
buf ( n306961 , n16532 );
and ( n306962 , n306958 , n306961 );
and ( n16535 , n833 , n306957 );
or ( n306964 , n306962 , n16535 );
not ( n306965 , n306964 );
nand ( n16538 , n306952 , n306965 );
xor ( n306967 , n833 , n306957 );
xor ( n306968 , n306967 , n306961 );
not ( n16541 , n306968 );
xor ( n306970 , n834 , n306907 );
and ( n16543 , n306970 , n306936 );
and ( n306972 , n834 , n306907 );
or ( n16545 , n16543 , n306972 );
not ( n16546 , n16545 );
nand ( n306975 , n16541 , n16546 );
nand ( n306976 , n16538 , n306975 );
nor ( n306977 , n306948 , n306976 );
not ( n16550 , n306977 );
or ( n306979 , n306902 , n16550 );
not ( n306980 , n306976 );
not ( n16553 , n306943 );
nor ( n306982 , n16553 , n306945 );
not ( n306983 , n306982 );
not ( n16556 , n306940 );
or ( n306985 , n306983 , n16556 );
not ( n306986 , n16511 );
buf ( n16559 , n306937 );
nand ( n306988 , n306986 , n16559 );
nand ( n306989 , n306985 , n306988 );
and ( n306990 , n306980 , n306989 );
not ( n16563 , n16538 );
not ( n306992 , n16546 );
nand ( n16565 , n306992 , n306968 );
or ( n16566 , n16563 , n16565 );
nand ( n306995 , n306951 , n306964 );
nand ( n306996 , n16566 , n306995 );
nor ( n306997 , n306990 , n306996 );
nand ( n16570 , n306979 , n306997 );
not ( n306999 , n16570 );
buf ( n307000 , n846 );
xor ( n16573 , n301064 , n301070 );
and ( n307002 , n16573 , n301122 );
and ( n307003 , n301064 , n301070 );
or ( n16576 , n307002 , n307003 );
buf ( n307005 , n16576 );
buf ( n307006 , n307005 );
xor ( n307007 , n307000 , n307006 );
xor ( n307008 , n303490 , n303494 );
xor ( n16581 , n307008 , n303501 );
buf ( n307010 , n16581 );
buf ( n307011 , n307010 );
xor ( n307012 , n307007 , n307011 );
buf ( n307013 , n307012 );
buf ( n16586 , n307013 );
nor ( n307015 , n16586 , n12980 );
buf ( n307016 , n848 );
xor ( n307017 , n292215 , n292221 );
and ( n16590 , n307017 , n292320 );
and ( n16591 , n292215 , n292221 );
or ( n307020 , n16590 , n16591 );
buf ( n307021 , n307020 );
buf ( n307022 , n307021 );
xor ( n307023 , n307016 , n307022 );
xor ( n307024 , n10526 , n301025 );
xor ( n307025 , n307024 , n301032 );
buf ( n307026 , n307025 );
buf ( n307027 , n307026 );
and ( n307028 , n307023 , n307027 );
and ( n16601 , n307016 , n307022 );
or ( n307030 , n307028 , n16601 );
buf ( n307031 , n307030 );
nand ( n16604 , n307031 , n303515 );
or ( n307033 , n307015 , n16604 );
nand ( n307034 , n16586 , n12980 );
nand ( n16607 , n307033 , n307034 );
not ( n307036 , n16607 );
nor ( n307037 , n303477 , n13544 );
xor ( n16610 , n307000 , n307006 );
and ( n307039 , n16610 , n307011 );
and ( n307040 , n307000 , n307006 );
or ( n16613 , n307039 , n307040 );
buf ( n307042 , n16613 );
nor ( n16615 , n303511 , n307042 );
nor ( n16616 , n307037 , n16615 );
not ( n307045 , n16616 );
or ( n307046 , n307036 , n307045 );
or ( n307047 , n303477 , n13544 );
and ( n16620 , n303511 , n307042 );
and ( n307049 , n307047 , n16620 );
not ( n307050 , n303477 );
not ( n16623 , n13544 );
nor ( n307052 , n307050 , n16623 );
nor ( n307053 , n307049 , n307052 );
nand ( n16626 , n307046 , n307053 );
not ( n307055 , n16626 );
xor ( n307056 , n296370 , n296376 );
xor ( n16629 , n307056 , n296397 );
buf ( n307058 , n16629 );
nor ( n16631 , n307058 , n293580 );
xor ( n16632 , n292347 , n293267 );
xor ( n16633 , n16632 , n293576 );
buf ( n307062 , n16633 );
buf ( n307063 , n842 );
xor ( n16636 , n298346 , n298351 );
and ( n307065 , n16636 , n298356 );
and ( n307066 , n298346 , n298351 );
or ( n16639 , n307065 , n307066 );
buf ( n307068 , n16639 );
buf ( n307069 , n307068 );
xor ( n16642 , n307063 , n307069 );
buf ( n307071 , n304557 );
and ( n16644 , n16642 , n307071 );
and ( n16645 , n307063 , n307069 );
or ( n307074 , n16644 , n16645 );
buf ( n307075 , n307074 );
nor ( n16648 , n307062 , n307075 );
nor ( n307077 , n16631 , n16648 );
xor ( n307078 , n297878 , n298339 );
xor ( n16651 , n307078 , n298359 );
buf ( n307080 , n16651 );
xor ( n307081 , n303423 , n303469 );
and ( n16654 , n307081 , n303474 );
and ( n307083 , n303423 , n303469 );
or ( n16656 , n16654 , n307083 );
buf ( n307085 , n16656 );
nor ( n307086 , n307080 , n307085 );
xor ( n307087 , n307063 , n307069 );
xor ( n307088 , n307087 , n307071 );
buf ( n307089 , n307088 );
nor ( n307090 , n307089 , n298363 );
nor ( n307091 , n307086 , n307090 );
and ( n16664 , n307077 , n307091 );
not ( n307093 , n16664 );
or ( n307094 , n307055 , n307093 );
nand ( n16667 , n307085 , n307080 );
not ( n307096 , n16667 );
not ( n307097 , n307096 );
not ( n16670 , n307090 );
not ( n16671 , n16670 );
or ( n16672 , n307097 , n16671 );
buf ( n16673 , n307089 );
nand ( n16674 , n16673 , n298363 );
nand ( n307103 , n16672 , n16674 );
not ( n307104 , n307103 );
not ( n16677 , n307077 );
or ( n307106 , n307104 , n16677 );
nand ( n307107 , n307075 , n307062 );
not ( n16680 , n307107 );
not ( n16681 , n16631 );
and ( n16682 , n16680 , n16681 );
and ( n16683 , n307058 , n293580 );
nor ( n307112 , n16682 , n16683 );
nand ( n307113 , n307106 , n307112 );
not ( n16686 , n307113 );
nand ( n307115 , n307094 , n16686 );
nor ( n307116 , n12994 , n13539 );
nor ( n16689 , n16434 , n307116 );
and ( n307118 , n16463 , n16689 );
nand ( n307119 , n307115 , n306977 , n307118 );
xor ( n16692 , n307016 , n307022 );
xor ( n307121 , n16692 , n307027 );
buf ( n307122 , n307121 );
not ( n16695 , n307122 );
not ( n307124 , n292327 );
nand ( n307125 , n16695 , n307124 );
xor ( n16698 , n291648 , n292137 );
xor ( n307127 , n16698 , n292323 );
buf ( n307128 , n307127 );
not ( n16701 , n307128 );
xor ( n16702 , n303516 , n303551 );
and ( n307131 , n16702 , n303556 );
and ( n16704 , n303516 , n303551 );
or ( n307133 , n307131 , n16704 );
buf ( n307134 , n307133 );
not ( n16707 , n307134 );
nand ( n16708 , n16701 , n16707 );
nand ( n307137 , n307125 , n16708 );
not ( n16710 , n13131 );
buf ( n16711 , n851 );
xor ( n16712 , n1469 , n291911 );
xor ( n307141 , n16712 , n291954 );
buf ( n16714 , n307141 );
xor ( n307143 , n4581 , n295014 );
and ( n16716 , n307143 , n295049 );
and ( n16717 , n4581 , n295014 );
or ( n16718 , n16716 , n16717 );
buf ( n16719 , n16718 );
xor ( n16720 , n16714 , n16719 );
xor ( n307149 , n303526 , n303532 );
xor ( n307150 , n307149 , n13108 );
buf ( n307151 , n307150 );
buf ( n307152 , n307151 );
and ( n307153 , n16720 , n307152 );
and ( n16726 , n16714 , n16719 );
or ( n307155 , n307153 , n16726 );
buf ( n307156 , n307155 );
buf ( n307157 , n307156 );
xor ( n307158 , n16711 , n307157 );
xor ( n16731 , n303520 , n303541 );
xor ( n307160 , n16731 , n303546 );
buf ( n307161 , n307160 );
buf ( n307162 , n307161 );
and ( n16735 , n307158 , n307162 );
and ( n16736 , n16711 , n307157 );
or ( n307165 , n16735 , n16736 );
buf ( n307166 , n307165 );
not ( n16739 , n307166 );
nand ( n307168 , n16710 , n16739 );
xor ( n16741 , n16711 , n307157 );
xor ( n307170 , n16741 , n307162 );
buf ( n307171 , n307170 );
not ( n16744 , n307171 );
buf ( n307173 , n852 );
xor ( n307174 , n294997 , n4579 );
and ( n16747 , n307174 , n4622 );
and ( n307176 , n294997 , n4579 );
or ( n307177 , n16747 , n307176 );
buf ( n307178 , n307177 );
xor ( n307179 , n307173 , n307178 );
xor ( n307180 , n16714 , n16719 );
xor ( n16753 , n307180 , n307152 );
buf ( n307182 , n16753 );
buf ( n307183 , n307182 );
and ( n16756 , n307179 , n307183 );
and ( n307185 , n307173 , n307178 );
or ( n307186 , n16756 , n307185 );
buf ( n307187 , n307186 );
not ( n307188 , n307187 );
nand ( n307189 , n16744 , n307188 );
nand ( n16762 , n307168 , n307189 );
nor ( n307191 , n307137 , n16762 );
xor ( n307192 , n307173 , n307178 );
xor ( n16765 , n307192 , n307183 );
buf ( n307194 , n16765 );
not ( n307195 , n307194 );
not ( n16768 , n295056 );
nand ( n16769 , n307195 , n16768 );
not ( n307198 , n16769 );
nor ( n16771 , n13135 , n12779 );
nor ( n307200 , n307198 , n16771 );
not ( n307201 , n307200 );
nor ( n16774 , n303567 , n303280 );
buf ( n307203 , n856 );
buf ( n307204 , n303378 );
not ( n16777 , n307204 );
buf ( n307206 , n1453 );
not ( n307207 , n307206 );
or ( n16780 , n16777 , n307207 );
buf ( n307209 , n291886 );
buf ( n307210 , n295074 );
nand ( n16783 , n307209 , n307210 );
buf ( n307212 , n16783 );
buf ( n307213 , n307212 );
nand ( n16786 , n16780 , n307213 );
buf ( n307215 , n16786 );
buf ( n307216 , n307215 );
and ( n307217 , n12920 , n303361 );
buf ( n307218 , n307217 );
buf ( n307219 , n307218 );
xor ( n16792 , n307216 , n307219 );
xor ( n16793 , n303218 , n303235 );
xor ( n16794 , n16793 , n303253 );
buf ( n307223 , n16794 );
buf ( n307224 , n307223 );
and ( n16797 , n16792 , n307224 );
and ( n16798 , n307216 , n307219 );
or ( n16799 , n16797 , n16798 );
buf ( n307228 , n16799 );
buf ( n307229 , n307228 );
xor ( n307230 , n307203 , n307229 );
xor ( n16803 , n12784 , n303258 );
xnor ( n16804 , n16803 , n12782 );
buf ( n307233 , n16804 );
and ( n16806 , n307230 , n307233 );
and ( n307235 , n307203 , n307229 );
or ( n307236 , n16806 , n307235 );
buf ( n307237 , n307236 );
nand ( n307238 , n13143 , n307237 );
or ( n16811 , n16774 , n307238 );
nand ( n16812 , n303567 , n303280 );
nand ( n16813 , n16811 , n16812 );
not ( n307242 , n16813 );
or ( n307243 , n307201 , n307242 );
nand ( n16816 , n13135 , n12779 );
not ( n307245 , n16816 );
and ( n16818 , n307245 , n16769 );
not ( n307247 , n307194 );
nor ( n16820 , n307247 , n16768 );
nor ( n307249 , n16818 , n16820 );
nand ( n307250 , n307243 , n307249 );
nand ( n16823 , n307191 , n307250 );
nor ( n307252 , n13143 , n307237 );
nor ( n307253 , n16774 , n307252 );
not ( n16826 , n16771 );
nand ( n307255 , n16769 , n307253 , n16826 );
xor ( n16828 , n303281 , n303331 );
xor ( n16829 , n16828 , n303402 );
buf ( n307258 , n16829 );
buf ( n16831 , n859 );
buf ( n307260 , n797 );
buf ( n307261 , n830 );
xor ( n307262 , n307260 , n307261 );
buf ( n307263 , n307262 );
buf ( n307264 , n307263 );
not ( n16837 , n307264 );
buf ( n307266 , n1271 );
not ( n307267 , n307266 );
or ( n16840 , n16837 , n307267 );
buf ( n307269 , n303287 );
buf ( n307270 , n831 );
nand ( n16843 , n307269 , n307270 );
buf ( n307272 , n16843 );
buf ( n307273 , n307272 );
nand ( n307274 , n16840 , n307273 );
buf ( n307275 , n307274 );
buf ( n307276 , n307275 );
buf ( n307277 , n799 );
buf ( n307278 , n829 );
or ( n307279 , n307277 , n307278 );
buf ( n16852 , n830 );
nand ( n16853 , n307279 , n16852 );
buf ( n16854 , n16853 );
buf ( n16855 , n16854 );
buf ( n16856 , n799 );
buf ( n16857 , n829 );
nand ( n16858 , n16856 , n16857 );
buf ( n307287 , n16858 );
buf ( n16860 , n307287 );
buf ( n307289 , n828 );
nand ( n307290 , n16855 , n16860 , n307289 );
buf ( n307291 , n307290 );
buf ( n16864 , n307291 );
not ( n307293 , n16864 );
buf ( n307294 , n307293 );
buf ( n307295 , n307294 );
and ( n307296 , n307276 , n307295 );
buf ( n307297 , n307296 );
buf ( n307298 , n307297 );
xor ( n16871 , n16831 , n307298 );
xor ( n16872 , n303286 , n303304 );
xor ( n307301 , n16872 , n303326 );
buf ( n307302 , n307301 );
buf ( n307303 , n307302 );
and ( n16876 , n16871 , n307303 );
and ( n307305 , n16831 , n307298 );
or ( n307306 , n16876 , n307305 );
buf ( n307307 , n307306 );
nor ( n307308 , n307258 , n307307 );
not ( n307309 , n307308 );
buf ( n307310 , n861 );
buf ( n307311 , n291939 );
buf ( n307312 , n799 );
and ( n307313 , n307311 , n307312 );
buf ( n307314 , n307313 );
buf ( n307315 , n307314 );
xor ( n307316 , n307310 , n307315 );
buf ( n16889 , n291656 );
not ( n16890 , n16889 );
buf ( n307319 , n798 );
buf ( n307320 , n830 );
xor ( n16893 , n307319 , n307320 );
buf ( n307322 , n16893 );
buf ( n307323 , n307322 );
not ( n16896 , n307323 );
or ( n307325 , n16890 , n16896 );
buf ( n307326 , n307263 );
buf ( n307327 , n831 );
nand ( n307328 , n307326 , n307327 );
buf ( n307329 , n307328 );
buf ( n307330 , n307329 );
nand ( n307331 , n307325 , n307330 );
buf ( n307332 , n307331 );
buf ( n307333 , n307332 );
xor ( n307334 , n307316 , n307333 );
buf ( n307335 , n307334 );
buf ( n307336 , n862 );
buf ( n307337 , n799 );
buf ( n307338 , n831 );
nand ( n16911 , n307337 , n307338 );
buf ( n307340 , n16911 );
buf ( n16913 , n307340 );
buf ( n16914 , n830 );
and ( n16915 , n16913 , n16914 );
buf ( n307344 , n16915 );
buf ( n16917 , n307344 );
xor ( n16918 , n307336 , n16917 );
buf ( n307347 , n799 );
not ( n307348 , n307347 );
buf ( n307349 , n307348 );
buf ( n307350 , n307349 );
not ( n307351 , n307350 );
buf ( n307352 , n291656 );
not ( n307353 , n307352 );
or ( n16926 , n307351 , n307353 );
buf ( n307355 , n307322 );
buf ( n307356 , n831 );
nand ( n307357 , n307355 , n307356 );
buf ( n307358 , n307357 );
buf ( n307359 , n307358 );
nand ( n307360 , n16926 , n307359 );
buf ( n307361 , n307360 );
buf ( n307362 , n307361 );
and ( n16935 , n16918 , n307362 );
and ( n307364 , n307336 , n16917 );
or ( n307365 , n16935 , n307364 );
buf ( n307366 , n307365 );
or ( n307367 , n307335 , n307366 );
xor ( n307368 , n307336 , n16917 );
xor ( n16941 , n307368 , n307362 );
buf ( n307370 , n16941 );
buf ( n16943 , n863 );
buf ( n307372 , n307340 );
not ( n16945 , n307372 );
buf ( n16946 , n16945 );
buf ( n307375 , n16946 );
and ( n16948 , n16943 , n307375 );
buf ( n307377 , n16948 );
nand ( n16950 , n307367 , n307370 , n307377 );
not ( n307379 , n16950 );
xor ( n16952 , n307310 , n307315 );
and ( n16953 , n16952 , n307333 );
and ( n307382 , n307310 , n307315 );
or ( n307383 , n16953 , n307382 );
buf ( n307384 , n307383 );
buf ( n307385 , n860 );
buf ( n16958 , n799 );
buf ( n16959 , n828 );
xor ( n16960 , n16958 , n16959 );
buf ( n16961 , n16960 );
buf ( n16962 , n16961 );
not ( n16963 , n16962 );
buf ( n307392 , n291808 );
buf ( n307393 , n307392 );
not ( n16966 , n307393 );
or ( n307395 , n16963 , n16966 );
buf ( n307396 , n291939 );
buf ( n307397 , n303309 );
nand ( n307398 , n307396 , n307397 );
buf ( n307399 , n307398 );
buf ( n307400 , n307399 );
nand ( n307401 , n307395 , n307400 );
buf ( n307402 , n307401 );
buf ( n307403 , n307402 );
xor ( n307404 , n307385 , n307403 );
xnor ( n307405 , n307291 , n307275 );
buf ( n307406 , n307405 );
xor ( n16979 , n307404 , n307406 );
buf ( n307408 , n16979 );
or ( n16981 , n307384 , n307408 );
nand ( n307410 , n307379 , n16981 );
and ( n307411 , n307335 , n307366 );
nand ( n16984 , n16981 , n307411 );
nand ( n307413 , n307408 , n307384 );
nand ( n307414 , n307410 , n16984 , n307413 );
xor ( n16987 , n16831 , n307298 );
xor ( n307416 , n16987 , n307303 );
buf ( n307417 , n307416 );
xor ( n16990 , n307385 , n307403 );
and ( n16991 , n16990 , n307406 );
and ( n16992 , n307385 , n307403 );
or ( n307421 , n16991 , n16992 );
buf ( n307422 , n307421 );
or ( n16995 , n307417 , n307422 );
nand ( n307424 , n307309 , n307414 , n16995 );
not ( n307425 , n307424 );
xor ( n16998 , n307203 , n307229 );
xor ( n307427 , n16998 , n307233 );
buf ( n307428 , n307427 );
not ( n17001 , n307428 );
buf ( n307430 , n857 );
xor ( n17003 , n303364 , n303385 );
and ( n17004 , n17003 , n303399 );
and ( n307433 , n303364 , n303385 );
or ( n17006 , n17004 , n307433 );
buf ( n307435 , n17006 );
buf ( n307436 , n307435 );
xor ( n307437 , n307430 , n307436 );
xor ( n307438 , n307216 , n307219 );
xor ( n17011 , n307438 , n307224 );
buf ( n307440 , n17011 );
buf ( n307441 , n307440 );
and ( n17014 , n307437 , n307441 );
and ( n307443 , n307430 , n307436 );
or ( n17016 , n17014 , n307443 );
buf ( n307445 , n17016 );
not ( n307446 , n307445 );
nand ( n307447 , n17001 , n307446 );
xor ( n307448 , n307430 , n307436 );
xor ( n17021 , n307448 , n307441 );
buf ( n17022 , n17021 );
not ( n307451 , n17022 );
not ( n17024 , n303407 );
nand ( n307453 , n307451 , n17024 );
nand ( n307454 , n307425 , n307447 , n307453 );
nand ( n17027 , n307422 , n307417 );
or ( n307456 , n307308 , n17027 );
nand ( n17029 , n307258 , n307307 );
nand ( n307458 , n307456 , n17029 );
nand ( n307459 , n307447 , n307453 , n307458 );
nand ( n17032 , n17022 , n303407 );
not ( n17033 , n17032 );
and ( n307462 , n307447 , n17033 );
nor ( n17035 , n17001 , n307446 );
nor ( n17036 , n307462 , n17035 );
and ( n307465 , n307454 , n307459 , n17036 );
not ( n307466 , n307465 );
not ( n17039 , n307466 );
nor ( n307468 , n307255 , n17039 );
nand ( n307469 , n307191 , n307468 );
not ( n307470 , n307137 );
not ( n17043 , n307171 );
nor ( n307472 , n17043 , n307188 );
not ( n17045 , n307472 );
not ( n17046 , n307168 );
or ( n307475 , n17045 , n17046 );
nand ( n307476 , n13131 , n307166 );
nand ( n17049 , n307475 , n307476 );
and ( n307478 , n307470 , n17049 );
not ( n307479 , n307125 );
nand ( n17052 , n307128 , n307134 );
not ( n307481 , n17052 );
not ( n307482 , n307481 );
or ( n307483 , n307479 , n307482 );
nand ( n17056 , n292327 , n307122 );
nand ( n307485 , n307483 , n17056 );
nor ( n307486 , n307478 , n307485 );
nand ( n17059 , n16823 , n307469 , n307486 );
not ( n307488 , n17059 );
not ( n17061 , n307488 );
nand ( n17062 , n307050 , n16623 );
not ( n307491 , n16615 );
nor ( n307492 , n303515 , n307031 );
nor ( n17065 , n307015 , n307492 );
and ( n307494 , n17062 , n307491 , n17065 );
and ( n307495 , n16664 , n307494 );
not ( n17068 , n306947 );
nor ( n307497 , n17068 , n306976 );
nand ( n17070 , n17061 , n307495 , n307497 , n307118 );
nand ( n17071 , n306999 , n307119 , n17070 );
buf ( n307500 , n17071 );
not ( n307501 , n307500 );
or ( n17074 , n306859 , n307501 );
not ( n307503 , n16426 );
nand ( n307504 , n306847 , n16421 );
not ( n17077 , n307504 );
and ( n307506 , n307503 , n17077 );
nand ( n17079 , n306852 , n16425 );
not ( n17080 , n17079 );
nor ( n307509 , n307506 , n17080 );
nand ( n307510 , n306799 , n16359 );
or ( n17083 , n16405 , n307510 );
nand ( n307512 , n306827 , n306832 );
nand ( n307513 , n17083 , n307512 );
nand ( n17086 , n306855 , n307513 );
nand ( n307515 , n307509 , n17086 );
buf ( n17088 , n307515 );
not ( n17089 , n17088 );
nand ( n17090 , n17074 , n17089 );
not ( n17091 , n17090 );
or ( n307520 , n16261 , n17091 );
or ( n307521 , n17090 , n306688 );
nand ( n17094 , n307520 , n307521 );
xor ( n307523 , n300444 , n300840 );
nor ( n307524 , n303959 , n307523 );
nor ( n17097 , n307524 , n306685 );
buf ( n307526 , n17097 );
not ( n17099 , n307526 );
nor ( n17100 , n17099 , n16429 );
not ( n307529 , n17100 );
not ( n307530 , n307500 );
or ( n17103 , n307529 , n307530 );
not ( n307532 , n307509 );
not ( n307533 , n17086 );
or ( n17106 , n307532 , n307533 );
nand ( n307535 , n17106 , n17097 );
not ( n307536 , n307535 );
nor ( n307537 , n303959 , n307523 );
or ( n307538 , n307537 , n16259 );
nand ( n17111 , n303959 , n307523 );
nand ( n307540 , n307538 , n17111 );
nor ( n307541 , n307536 , n307540 );
nand ( n17114 , n17103 , n307541 );
xor ( n307543 , n300583 , n300591 );
and ( n17116 , n307543 , n300838 );
and ( n17117 , n300583 , n300591 );
or ( n307546 , n17116 , n17117 );
buf ( n307547 , n307546 );
not ( n17120 , n307547 );
not ( n307549 , n300457 );
not ( n307550 , n300462 );
or ( n17123 , n307549 , n307550 );
nor ( n307552 , n300462 , n300457 );
not ( n307553 , n300581 );
or ( n17126 , n307552 , n307553 );
nand ( n17127 , n17123 , n17126 );
buf ( n307556 , n17127 );
not ( n17129 , n300740 );
not ( n307558 , n300748 );
or ( n17131 , n17129 , n307558 );
not ( n17132 , n300740 );
nand ( n307561 , n10321 , n17132 );
nand ( n307562 , n300824 , n307561 );
nand ( n307563 , n17131 , n307562 );
xor ( n17136 , n300629 , n300682 );
and ( n307565 , n17136 , n300738 );
and ( n307566 , n300629 , n300682 );
or ( n17139 , n307565 , n307566 );
buf ( n307568 , n17139 );
buf ( n307569 , n307568 );
xor ( n17142 , n302994 , n302998 );
xor ( n307571 , n17142 , n303003 );
buf ( n307572 , n307571 );
buf ( n307573 , n307572 );
xor ( n17146 , n307569 , n307573 );
xor ( n17147 , n300757 , n300815 );
and ( n307576 , n17147 , n300822 );
and ( n17149 , n300757 , n300815 );
or ( n17150 , n307576 , n17149 );
buf ( n307579 , n17150 );
buf ( n307580 , n307579 );
xor ( n17153 , n17146 , n307580 );
buf ( n307582 , n17153 );
xor ( n307583 , n307563 , n307582 );
xor ( n307584 , n303047 , n303065 );
xor ( n307585 , n307584 , n303070 );
buf ( n307586 , n307585 );
buf ( n307587 , n307586 );
not ( n307588 , n300576 );
not ( n17161 , n300493 );
or ( n307590 , n307588 , n17161 );
or ( n17163 , n300493 , n300576 );
nand ( n17164 , n17163 , n300468 );
nand ( n307593 , n307590 , n17164 );
buf ( n17166 , n307593 );
xor ( n17167 , n307587 , n17166 );
xor ( n307596 , n303079 , n303084 );
xor ( n307597 , n307596 , n303088 );
buf ( n307598 , n307597 );
xor ( n307599 , n17167 , n307598 );
buf ( n307600 , n307599 );
xor ( n17173 , n307583 , n307600 );
buf ( n307602 , n17173 );
xor ( n307603 , n307556 , n307602 );
xor ( n17176 , n300597 , n10397 );
and ( n307605 , n17176 , n10408 );
and ( n17178 , n300597 , n10397 );
or ( n17179 , n307605 , n17178 );
buf ( n307608 , n17179 );
xor ( n307609 , n307603 , n307608 );
buf ( n307610 , n307609 );
not ( n17183 , n307610 );
not ( n307612 , n17183 );
or ( n307613 , n17120 , n307612 );
not ( n17186 , n307547 );
nand ( n307615 , n17186 , n307610 );
nand ( n307616 , n307613 , n307615 );
nor ( n17189 , n303572 , n307616 );
not ( n307618 , n17189 );
nand ( n307619 , n303572 , n307616 );
nand ( n17192 , n307618 , n307619 );
not ( n17193 , n17192 );
and ( n17194 , n17114 , n17193 );
not ( n307623 , n17114 );
and ( n17196 , n307623 , n17192 );
nor ( n17197 , n17194 , n17196 );
xor ( n17198 , n307556 , n307602 );
and ( n17199 , n17198 , n307608 );
and ( n17200 , n307556 , n307602 );
or ( n17201 , n17199 , n17200 );
buf ( n307630 , n17201 );
xor ( n307631 , n307587 , n17166 );
and ( n17204 , n307631 , n307598 );
and ( n17205 , n307587 , n17166 );
or ( n17206 , n17204 , n17205 );
buf ( n307635 , n17206 );
buf ( n307636 , n307635 );
xor ( n17209 , n307563 , n307582 );
and ( n17210 , n17209 , n307600 );
and ( n307639 , n307563 , n307582 );
or ( n307640 , n17210 , n307639 );
buf ( n307641 , n307640 );
xor ( n307642 , n307636 , n307641 );
xor ( n307643 , n307569 , n307573 );
and ( n307644 , n307643 , n307580 );
and ( n17217 , n307569 , n307573 );
or ( n307646 , n307644 , n17217 );
buf ( n307647 , n307646 );
buf ( n307648 , n307647 );
xor ( n307649 , n303007 , n12595 );
xor ( n307650 , n307649 , n303027 );
buf ( n17223 , n307650 );
xor ( n17224 , n307648 , n17223 );
xor ( n307653 , n303075 , n303092 );
xor ( n307654 , n307653 , n303097 );
buf ( n307655 , n307654 );
buf ( n307656 , n307655 );
xor ( n307657 , n17224 , n307656 );
buf ( n307658 , n307657 );
buf ( n307659 , n307658 );
xor ( n307660 , n307642 , n307659 );
buf ( n307661 , n307660 );
and ( n307662 , n307630 , n307661 );
xor ( n17235 , n307636 , n307641 );
and ( n307664 , n17235 , n307659 );
and ( n17237 , n307636 , n307641 );
or ( n17238 , n307664 , n17237 );
buf ( n307667 , n17238 );
buf ( n17240 , n307667 );
xor ( n307669 , n302874 , n302941 );
xor ( n17242 , n307669 , n302946 );
buf ( n307671 , n17242 );
buf ( n307672 , n307671 );
xor ( n17245 , n307648 , n17223 );
and ( n307674 , n17245 , n307656 );
and ( n307675 , n307648 , n17223 );
or ( n17248 , n307674 , n307675 );
buf ( n307677 , n17248 );
buf ( n307678 , n307677 );
xor ( n17251 , n307672 , n307678 );
xor ( n17252 , n303031 , n303035 );
xor ( n17253 , n17252 , n303102 );
buf ( n307682 , n17253 );
buf ( n307683 , n307682 );
xor ( n17256 , n17251 , n307683 );
buf ( n307685 , n17256 );
buf ( n307686 , n307685 );
xor ( n17259 , n17240 , n307686 );
buf ( n307688 , n17259 );
and ( n307689 , n307662 , n307688 );
not ( n307690 , n307689 );
or ( n17263 , n307688 , n307662 );
nand ( n307692 , n307690 , n17263 );
not ( n17265 , n307692 );
not ( n17266 , n307661 );
not ( n307695 , n17266 );
not ( n307696 , n307630 );
or ( n307697 , n307695 , n307696 );
not ( n17270 , n307630 );
nand ( n307699 , n17270 , n307661 );
nand ( n307700 , n307697 , n307699 );
buf ( n17273 , n307700 );
buf ( n307702 , n307610 );
buf ( n307703 , n307547 );
and ( n17276 , n307702 , n307703 );
buf ( n17277 , n17276 );
buf ( n307706 , n17277 );
nor ( n17279 , n17273 , n307706 );
nor ( n307708 , n17279 , n17189 );
nand ( n17281 , n307708 , n17097 );
nor ( n307710 , n306856 , n17281 );
buf ( n17283 , n307710 );
not ( n17284 , n17283 );
not ( n307713 , n307500 );
or ( n17286 , n17284 , n307713 );
not ( n307715 , n307515 );
and ( n17288 , n307708 , n17097 );
not ( n307717 , n17288 );
or ( n307718 , n307715 , n307717 );
not ( n17291 , n307540 );
not ( n307720 , n307708 );
or ( n307721 , n17291 , n307720 );
nor ( n17294 , n17273 , n307706 );
or ( n307723 , n17294 , n307619 );
nand ( n17296 , n307706 , n17273 );
nand ( n307725 , n307723 , n17296 );
not ( n17298 , n307725 );
nand ( n17299 , n307721 , n17298 );
not ( n17300 , n17299 );
nand ( n307729 , n307718 , n17300 );
not ( n307730 , n307729 );
nand ( n17303 , n17286 , n307730 );
not ( n17304 , n17303 );
or ( n307733 , n17265 , n17304 );
or ( n307734 , n17303 , n307692 );
nand ( n17307 , n307733 , n307734 );
buf ( n307736 , n16518 );
not ( n17309 , n307736 );
buf ( n307738 , n16473 );
not ( n17311 , n307738 );
or ( n17312 , n17309 , n17311 );
not ( n307741 , n306982 );
nand ( n17314 , n17312 , n307741 );
not ( n307743 , n17314 );
and ( n17316 , n307118 , n307736 );
buf ( n307745 , n307495 );
not ( n307746 , n307488 );
buf ( n17319 , n307746 );
nand ( n307748 , n17316 , n307745 , n17319 );
buf ( n307749 , n307115 );
nand ( n307750 , n17316 , n307749 );
nand ( n17323 , n307743 , n307748 , n307750 );
buf ( n307752 , n306940 );
nand ( n17325 , n307752 , n306988 );
not ( n17326 , n17325 );
and ( n307755 , n17323 , n17326 );
not ( n307756 , n17323 );
and ( n17329 , n307756 , n17325 );
nor ( n307758 , n307755 , n17329 );
not ( n307759 , n307738 );
buf ( n17332 , n307118 );
nand ( n307761 , n307749 , n17332 );
buf ( n307762 , n17059 );
buf ( n17335 , n307762 );
nand ( n17336 , n307745 , n17332 , n17335 );
nand ( n17337 , n307759 , n307761 , n17336 );
not ( n17338 , n306982 );
nand ( n17339 , n17338 , n307736 );
not ( n17340 , n17339 );
and ( n307769 , n17337 , n17340 );
not ( n17342 , n17337 );
and ( n17343 , n17342 , n17339 );
nor ( n307772 , n307769 , n17343 );
buf ( n307773 , n16689 );
not ( n17346 , n306890 );
and ( n307775 , n307773 , n17346 );
nand ( n17348 , n307745 , n17335 , n307775 );
nand ( n307777 , n307749 , n307775 );
not ( n17350 , n17346 );
not ( n17351 , n16438 );
or ( n307780 , n17350 , n17351 );
nand ( n307781 , n307780 , n306895 );
not ( n17354 , n307781 );
nand ( n307783 , n17348 , n307777 , n17354 );
not ( n307784 , n16470 );
nor ( n17357 , n307784 , n306886 );
and ( n307786 , n307783 , n17357 );
not ( n307787 , n307783 );
not ( n17360 , n17357 );
and ( n307789 , n307787 , n17360 );
nor ( n307790 , n307786 , n307789 );
or ( n17363 , n307037 , n307052 );
not ( n307792 , n17363 );
and ( n307793 , n307491 , n17065 );
not ( n17366 , n307793 );
not ( n307795 , n307762 );
or ( n307796 , n17366 , n307795 );
not ( n17369 , n16607 );
not ( n307798 , n307491 );
or ( n307799 , n17369 , n307798 );
not ( n307800 , n16620 );
nand ( n17373 , n307799 , n307800 );
not ( n307802 , n17373 );
nand ( n17375 , n307796 , n307802 );
not ( n17376 , n17375 );
or ( n307805 , n307792 , n17376 );
or ( n307806 , n17375 , n17363 );
nand ( n17379 , n307805 , n307806 );
not ( n307808 , n307116 );
buf ( n307809 , n16435 );
nand ( n17382 , n307808 , n307809 );
not ( n307811 , n17382 );
not ( n307812 , n307745 );
not ( n17385 , n307746 );
or ( n307814 , n307812 , n17385 );
not ( n17387 , n307749 );
nand ( n307816 , n307814 , n17387 );
not ( n17389 , n307816 );
or ( n17390 , n307811 , n17389 );
or ( n307819 , n307816 , n17382 );
nand ( n307820 , n17390 , n307819 );
nand ( n17393 , n16670 , n16674 );
not ( n307822 , n17393 );
not ( n307823 , n307494 );
nor ( n17396 , n307823 , n307086 );
not ( n307825 , n17396 );
not ( n307826 , n307488 );
not ( n17399 , n307826 );
or ( n17400 , n307825 , n17399 );
not ( n17401 , n307086 );
not ( n307830 , n17401 );
not ( n307831 , n16626 );
or ( n17404 , n307830 , n307831 );
buf ( n17405 , n16667 );
nand ( n17406 , n17404 , n17405 );
not ( n307835 , n17406 );
nand ( n307836 , n17400 , n307835 );
not ( n17409 , n307836 );
or ( n17410 , n307822 , n17409 );
or ( n17411 , n307836 , n17393 );
nand ( n307840 , n17410 , n17411 );
not ( n307841 , n307823 );
not ( n17414 , n307841 );
not ( n307843 , n307762 );
or ( n307844 , n17414 , n307843 );
not ( n17417 , n16626 );
nand ( n17418 , n307844 , n17417 );
nand ( n17419 , n17401 , n17405 );
not ( n307848 , n17419 );
and ( n307849 , n17418 , n307848 );
not ( n17422 , n17418 );
and ( n17423 , n17422 , n17419 );
nor ( n307852 , n307849 , n17423 );
buf ( n307853 , n307773 );
nand ( n17426 , n307749 , n307853 );
nand ( n17427 , n307745 , n307826 , n307853 );
not ( n307856 , n16438 );
nand ( n307857 , n17426 , n17427 , n307856 );
not ( n17430 , n17065 );
not ( n17431 , n17059 );
or ( n307860 , n17430 , n17431 );
not ( n17433 , n16607 );
nand ( n17434 , n307860 , n17433 );
not ( n307863 , n307762 );
not ( n307864 , n307492 );
nand ( n17437 , n307864 , n16604 );
not ( n17438 , n17437 );
or ( n17439 , n307863 , n17438 );
or ( n307868 , n307826 , n17437 );
nand ( n307869 , n17439 , n307868 );
nand ( n17442 , n307745 , n307826 , n307808 );
and ( n17443 , n306940 , n16518 );
buf ( n17444 , n17443 );
and ( n17445 , n17444 , n306975 );
and ( n17446 , n17332 , n17445 );
nand ( n17447 , n17446 , n307745 , n17319 );
buf ( n17448 , n307091 );
not ( n307877 , n16648 );
and ( n17450 , n17448 , n307877 );
nand ( n17451 , n307746 , n17450 , n307841 );
not ( n17452 , n307468 );
not ( n307881 , n307250 );
nand ( n307882 , n17452 , n307881 );
not ( n17455 , n307472 );
nand ( n17456 , n307189 , n17455 );
not ( n17457 , n17456 );
and ( n307886 , n307882 , n17457 );
not ( n307887 , n307882 );
and ( n17460 , n307887 , n17456 );
nor ( n307889 , n307886 , n17460 );
nand ( n307890 , n307125 , n17056 );
not ( n307891 , n307890 );
not ( n17464 , n16762 );
buf ( n307893 , n16708 );
and ( n17466 , n17464 , n307893 );
not ( n17467 , n307255 );
nand ( n307896 , n17466 , n17467 , n307466 );
nand ( n307897 , n17466 , n307250 );
and ( n17470 , n17049 , n307893 );
nor ( n307899 , n17470 , n307481 );
nand ( n307900 , n307896 , n307897 , n307899 );
not ( n17473 , n307900 );
or ( n307902 , n307891 , n17473 );
or ( n307903 , n307900 , n307890 );
nand ( n307904 , n307902 , n307903 );
nand ( n17477 , n307189 , n307250 );
nand ( n307906 , n17467 , n307466 , n307189 );
nand ( n17479 , n17477 , n307906 , n17455 );
nand ( n17480 , n307168 , n307476 );
not ( n307909 , n17480 );
and ( n307910 , n17479 , n307909 );
not ( n17483 , n17479 );
and ( n307912 , n17483 , n17480 );
nor ( n307913 , n307910 , n307912 );
xor ( n17486 , n297868 , n297528 );
buf ( n307915 , n17486 );
nor ( n307916 , n13584 , n307915 );
not ( n17489 , n307916 );
and ( n307918 , n17240 , n307686 );
buf ( n307919 , n307918 );
not ( n307920 , n307919 );
not ( n307921 , n307920 );
xor ( n17494 , n307672 , n307678 );
and ( n17495 , n17494 , n307683 );
and ( n17496 , n307672 , n307678 );
or ( n307925 , n17495 , n17496 );
buf ( n307926 , n307925 );
xor ( n17499 , n302984 , n302988 );
xor ( n17500 , n17499 , n303107 );
buf ( n17501 , n17500 );
xor ( n307930 , n307926 , n17501 );
not ( n17503 , n307930 );
not ( n17504 , n17503 );
or ( n17505 , n307921 , n17504 );
nand ( n17506 , n17505 , n17263 );
buf ( n307935 , n17501 );
buf ( n307936 , n307926 );
and ( n307937 , n307935 , n307936 );
buf ( n307938 , n307937 );
not ( n17511 , n307938 );
xor ( n17512 , n303112 , n303116 );
buf ( n307941 , n17512 );
not ( n307942 , n307941 );
nand ( n307943 , n17511 , n307942 );
not ( n17516 , n303118 );
buf ( n307945 , n302965 );
buf ( n307946 , n302754 );
and ( n17519 , n307945 , n307946 );
not ( n17520 , n307945 );
buf ( n307949 , n302754 );
not ( n307950 , n307949 );
buf ( n307951 , n307950 );
buf ( n307952 , n307951 );
and ( n17525 , n17520 , n307952 );
nor ( n307954 , n17519 , n17525 );
buf ( n307955 , n307954 );
not ( n17528 , n307955 );
nand ( n17529 , n17516 , n17528 );
nand ( n17530 , n307943 , n17529 );
nor ( n307959 , n17506 , n17530 );
xor ( n307960 , n302391 , n302747 );
and ( n17533 , n307960 , n302752 );
and ( n17534 , n302391 , n302747 );
or ( n307963 , n17533 , n17534 );
buf ( n307964 , n307963 );
xor ( n17537 , n10860 , n301832 );
xor ( n17538 , n17537 , n302112 );
buf ( n307967 , n17538 );
xor ( n307968 , n307964 , n307967 );
or ( n307969 , n307968 , n302968 );
xor ( n17542 , n302117 , n302163 );
buf ( n307971 , n17542 );
buf ( n307972 , n307971 );
not ( n17545 , n307972 );
nand ( n17546 , n307964 , n307967 );
buf ( n17547 , n17546 );
nand ( n307976 , n17545 , n17547 );
nand ( n307977 , n307969 , n307976 );
xor ( n17550 , n303989 , n303993 );
xor ( n17551 , n17550 , n304000 );
buf ( n307980 , n17551 );
xor ( n307981 , n302123 , n302129 );
and ( n307982 , n307981 , n302160 );
and ( n17555 , n302123 , n302129 );
or ( n17556 , n307982 , n17555 );
buf ( n307985 , n17556 );
xor ( n307986 , n307980 , n307985 );
or ( n17559 , n302165 , n307986 );
buf ( n307988 , n307985 );
buf ( n307989 , n307980 );
and ( n17562 , n307988 , n307989 );
buf ( n307991 , n17562 );
not ( n307992 , n307991 );
xor ( n307993 , n304005 , n304009 );
buf ( n307994 , n307993 );
not ( n17567 , n307994 );
nand ( n17568 , n307992 , n17567 );
nand ( n17569 , n17559 , n17568 );
nor ( n307998 , n307977 , n17569 );
nand ( n307999 , n307959 , n307998 );
not ( n17572 , n307999 );
nor ( n17573 , n307540 , n307725 );
nand ( n17574 , n307535 , n17573 );
not ( n308003 , n307708 );
nand ( n308004 , n308003 , n17298 );
nand ( n17577 , n17572 , n17574 , n308004 );
not ( n17578 , n307998 );
not ( n17579 , n17530 );
not ( n308008 , n17579 );
nand ( n308009 , n307920 , n17503 );
not ( n17582 , n308009 );
not ( n17583 , n307689 );
or ( n17584 , n17582 , n17583 );
not ( n308013 , n307920 );
nand ( n308014 , n308013 , n307930 );
nand ( n17587 , n17584 , n308014 );
not ( n17588 , n17587 );
or ( n17589 , n308008 , n17588 );
buf ( n308018 , n17529 );
and ( n308019 , n307941 , n307938 );
and ( n17592 , n308018 , n308019 );
not ( n308021 , n17528 );
not ( n308022 , n308021 );
nor ( n17595 , n308022 , n17516 );
nor ( n308024 , n17592 , n17595 );
nand ( n308025 , n17589 , n308024 );
not ( n17598 , n308025 );
or ( n17599 , n17578 , n17598 );
not ( n308028 , n17569 );
not ( n308029 , n308028 );
not ( n17602 , n17546 );
nor ( n17603 , n17602 , n307972 );
nand ( n308032 , n307968 , n302968 );
or ( n308033 , n17603 , n308032 );
nand ( n17606 , n307972 , n17602 );
nand ( n17607 , n308033 , n17606 );
not ( n17608 , n17607 );
or ( n17609 , n308029 , n17608 );
and ( n308038 , n307986 , n302165 );
and ( n308039 , n308038 , n17568 );
not ( n17612 , n307991 );
nor ( n17613 , n17612 , n17567 );
nor ( n308042 , n308039 , n17613 );
nand ( n308043 , n17609 , n308042 );
not ( n17616 , n308043 );
nand ( n17617 , n17599 , n17616 );
not ( n17618 , n17617 );
nand ( n17619 , n17577 , n17618 );
nand ( n17620 , n17489 , n17619 );
xor ( n308049 , n302184 , n11773 );
and ( n308050 , n308049 , n302208 );
and ( n17623 , n302184 , n11773 );
or ( n17624 , n308050 , n17623 );
buf ( n308053 , n17624 );
buf ( n308054 , n308053 );
xor ( n308055 , n302224 , n302361 );
and ( n17628 , n308055 , n302368 );
and ( n17629 , n302224 , n302361 );
or ( n17630 , n17628 , n17629 );
buf ( n308059 , n17630 );
buf ( n308060 , n308059 );
xor ( n17633 , n308054 , n308060 );
xor ( n17634 , n302227 , n302244 );
and ( n17635 , n17634 , n302259 );
and ( n308064 , n302227 , n302244 );
or ( n308065 , n17635 , n308064 );
buf ( n308066 , n308065 );
buf ( n308067 , n308066 );
xor ( n308068 , n302320 , n11909 );
and ( n17641 , n308068 , n302355 );
and ( n308070 , n302320 , n11909 );
or ( n308071 , n17641 , n308070 );
buf ( n308072 , n308071 );
buf ( n308073 , n308072 );
xor ( n308074 , n308067 , n308073 );
buf ( n308075 , n302313 );
not ( n17648 , n308075 );
buf ( n308077 , n296508 );
not ( n308078 , n308077 );
or ( n17651 , n17648 , n308078 );
buf ( n308080 , n296749 );
buf ( n308081 , n777 );
buf ( n308082 , n802 );
xor ( n17655 , n308081 , n308082 );
buf ( n308084 , n17655 );
buf ( n308085 , n308084 );
nand ( n308086 , n308080 , n308085 );
buf ( n308087 , n308086 );
buf ( n308088 , n308087 );
nand ( n17661 , n17651 , n308088 );
buf ( n308090 , n17661 );
buf ( n308091 , n308090 );
buf ( n308092 , n11841 );
not ( n308093 , n308092 );
buf ( n308094 , n296594 );
not ( n17667 , n308094 );
or ( n17668 , n308093 , n17667 );
buf ( n308097 , n294557 );
buf ( n308098 , n771 );
buf ( n308099 , n808 );
xor ( n308100 , n308098 , n308099 );
buf ( n308101 , n308100 );
buf ( n308102 , n308101 );
nand ( n17675 , n308097 , n308102 );
buf ( n308104 , n17675 );
buf ( n308105 , n308104 );
nand ( n17678 , n17668 , n308105 );
buf ( n17679 , n17678 );
buf ( n17680 , n17679 );
xor ( n17681 , n308091 , n17680 );
buf ( n308110 , n302350 );
not ( n308111 , n308110 );
buf ( n308112 , n308111 );
buf ( n308113 , n308112 );
not ( n308114 , n308113 );
buf ( n308115 , n296441 );
not ( n17688 , n308115 );
or ( n17689 , n308114 , n17688 );
buf ( n17690 , n6017 );
buf ( n308119 , n17690 );
buf ( n308120 , n804 );
buf ( n308121 , n775 );
xor ( n308122 , n308120 , n308121 );
buf ( n308123 , n308122 );
buf ( n308124 , n308123 );
nand ( n17697 , n308119 , n308124 );
buf ( n308126 , n17697 );
buf ( n308127 , n308126 );
nand ( n17700 , n17689 , n308127 );
buf ( n17701 , n17700 );
buf ( n308130 , n17701 );
xor ( n308131 , n17681 , n308130 );
buf ( n308132 , n308131 );
buf ( n308133 , n308132 );
xor ( n308134 , n308074 , n308133 );
buf ( n308135 , n308134 );
buf ( n308136 , n308135 );
xor ( n17709 , n302262 , n302302 );
and ( n308138 , n17709 , n302358 );
and ( n17711 , n302262 , n302302 );
or ( n308140 , n308138 , n17711 );
buf ( n308141 , n308140 );
buf ( n308142 , n308141 );
xor ( n17715 , n308136 , n308142 );
and ( n308144 , n6908 , n6909 );
buf ( n308145 , n308144 );
buf ( n308146 , n308145 );
buf ( n308147 , n302252 );
not ( n308148 , n308147 );
buf ( n308149 , n296617 );
not ( n17722 , n308149 );
or ( n308151 , n308148 , n17722 );
buf ( n308152 , n295437 );
xor ( n17725 , n806 , n773 );
buf ( n308154 , n17725 );
nand ( n308155 , n308152 , n308154 );
buf ( n308156 , n308155 );
buf ( n308157 , n308156 );
nand ( n308158 , n308151 , n308157 );
buf ( n308159 , n308158 );
buf ( n308160 , n308159 );
xor ( n308161 , n308146 , n308160 );
buf ( n308162 , n302330 );
not ( n308163 , n308162 );
buf ( n308164 , n297175 );
not ( n17737 , n308164 );
or ( n308166 , n308163 , n17737 );
buf ( n17739 , n292841 );
buf ( n308168 , n810 );
buf ( n308169 , n769 );
and ( n308170 , n308168 , n308169 );
not ( n17743 , n308168 );
buf ( n308172 , n299244 );
and ( n17745 , n17743 , n308172 );
nor ( n17746 , n308170 , n17745 );
buf ( n308175 , n17746 );
buf ( n308176 , n308175 );
nand ( n308177 , n17739 , n308176 );
buf ( n308178 , n308177 );
buf ( n308179 , n308178 );
nand ( n17752 , n308166 , n308179 );
buf ( n308181 , n17752 );
buf ( n308182 , n308181 );
xor ( n308183 , n308161 , n308182 );
buf ( n308184 , n308183 );
buf ( n308185 , n308184 );
buf ( n308186 , n11866 );
not ( n17759 , n308186 );
buf ( n308188 , n2376 );
not ( n308189 , n308188 );
or ( n17762 , n17759 , n308189 );
buf ( n308191 , n2383 );
buf ( n308192 , n812 );
nand ( n308193 , n308191 , n308192 );
buf ( n308194 , n308193 );
buf ( n308195 , n308194 );
nand ( n308196 , n17762 , n308195 );
buf ( n308197 , n308196 );
buf ( n308198 , n308197 );
not ( n308199 , n308198 );
buf ( n308200 , n308199 );
buf ( n308201 , n308200 );
buf ( n308202 , n302237 );
not ( n308203 , n308202 );
buf ( n308204 , n296480 );
not ( n308205 , n308204 );
or ( n308206 , n308203 , n308205 );
buf ( n308207 , n6057 );
buf ( n308208 , n800 );
buf ( n308209 , n779 );
xor ( n308210 , n308208 , n308209 );
buf ( n308211 , n308210 );
buf ( n308212 , n308211 );
nand ( n308213 , n308207 , n308212 );
buf ( n308214 , n308213 );
buf ( n308215 , n308214 );
nand ( n17788 , n308206 , n308215 );
buf ( n17789 , n17788 );
buf ( n17790 , n17789 );
xor ( n17791 , n308201 , n17790 );
buf ( n308220 , n302275 );
buf ( n308221 , n302300 );
or ( n17794 , n308220 , n308221 );
buf ( n308223 , n302286 );
nand ( n17796 , n17794 , n308223 );
buf ( n308225 , n17796 );
buf ( n308226 , n308225 );
buf ( n308227 , n297322 );
not ( n308228 , n308227 );
buf ( n308229 , n296594 );
not ( n308230 , n308229 );
or ( n308231 , n308228 , n308230 );
buf ( n308232 , n302272 );
nand ( n17805 , n308231 , n308232 );
buf ( n308234 , n17805 );
buf ( n308235 , n308234 );
buf ( n308236 , n302300 );
nand ( n17809 , n308235 , n308236 );
buf ( n308238 , n17809 );
buf ( n308239 , n308238 );
nand ( n308240 , n308226 , n308239 );
buf ( n308241 , n308240 );
buf ( n308242 , n308241 );
xor ( n308243 , n17791 , n308242 );
buf ( n308244 , n308243 );
buf ( n308245 , n308244 );
xor ( n308246 , n308185 , n308245 );
xor ( n308247 , n302185 , n302191 );
and ( n308248 , n308247 , n302198 );
and ( n17821 , n302185 , n302191 );
or ( n308250 , n308248 , n17821 );
buf ( n308251 , n308250 );
buf ( n308252 , n308251 );
xor ( n308253 , n308246 , n308252 );
buf ( n308254 , n308253 );
buf ( n308255 , n308254 );
xor ( n17828 , n17715 , n308255 );
buf ( n308257 , n17828 );
buf ( n308258 , n308257 );
xor ( n17831 , n17633 , n308258 );
buf ( n308260 , n17831 );
buf ( n17833 , n308260 );
xor ( n308262 , n302210 , n302215 );
and ( n17835 , n308262 , n302370 );
and ( n308264 , n302210 , n302215 );
or ( n308265 , n17835 , n308264 );
buf ( n308266 , n308265 );
xor ( n308267 , n17833 , n308266 );
buf ( n308268 , n308267 );
or ( n17841 , n11951 , n308268 );
and ( n308270 , n11806 , n302235 );
buf ( n308271 , n308270 );
buf ( n308272 , n308271 );
buf ( n308273 , n308101 );
not ( n308274 , n308273 );
buf ( n308275 , n296594 );
not ( n17848 , n308275 );
or ( n308277 , n308274 , n17848 );
buf ( n308278 , n294557 );
xor ( n308279 , n808 , n770 );
buf ( n308280 , n308279 );
nand ( n308281 , n308278 , n308280 );
buf ( n308282 , n308281 );
buf ( n308283 , n308282 );
nand ( n308284 , n308277 , n308283 );
buf ( n308285 , n308284 );
buf ( n308286 , n308285 );
xor ( n308287 , n308272 , n308286 );
buf ( n308288 , n308123 );
not ( n308289 , n308288 );
buf ( n308290 , n296441 );
not ( n17863 , n308290 );
or ( n308292 , n308289 , n17863 );
buf ( n17865 , n296446 );
buf ( n308294 , n774 );
buf ( n308295 , n804 );
xor ( n308296 , n308294 , n308295 );
buf ( n308297 , n308296 );
buf ( n308298 , n308297 );
nand ( n308299 , n17865 , n308298 );
buf ( n308300 , n308299 );
buf ( n308301 , n308300 );
nand ( n308302 , n308292 , n308301 );
buf ( n308303 , n308302 );
buf ( n308304 , n308303 );
xor ( n308305 , n308287 , n308304 );
buf ( n308306 , n308305 );
buf ( n308307 , n308306 );
buf ( n308308 , n308211 );
not ( n308309 , n308308 );
buf ( n308310 , n296480 );
not ( n17883 , n308310 );
or ( n308312 , n308309 , n17883 );
buf ( n308313 , n6057 );
buf ( n308314 , n800 );
buf ( n308315 , n778 );
xor ( n17888 , n308314 , n308315 );
buf ( n308317 , n17888 );
buf ( n308318 , n308317 );
nand ( n308319 , n308313 , n308318 );
buf ( n308320 , n308319 );
buf ( n308321 , n308320 );
nand ( n308322 , n308312 , n308321 );
buf ( n308323 , n308322 );
buf ( n17896 , n308084 );
not ( n17897 , n17896 );
buf ( n17898 , n296508 );
not ( n17899 , n17898 );
or ( n17900 , n17897 , n17899 );
buf ( n17901 , n296749 );
xor ( n308330 , n802 , n776 );
buf ( n17903 , n308330 );
nand ( n17904 , n17901 , n17903 );
buf ( n308333 , n17904 );
buf ( n308334 , n308333 );
nand ( n17907 , n17900 , n308334 );
buf ( n17908 , n17907 );
xor ( n308337 , n308323 , n17908 );
buf ( n308338 , n308337 );
buf ( n308339 , n308197 );
and ( n17912 , n308338 , n308339 );
not ( n308341 , n308338 );
buf ( n308342 , n308200 );
and ( n308343 , n308341 , n308342 );
nor ( n308344 , n17912 , n308343 );
buf ( n308345 , n308344 );
buf ( n308346 , n308345 );
xor ( n308347 , n308307 , n308346 );
xor ( n17920 , n308201 , n17790 );
and ( n308349 , n17920 , n308242 );
and ( n308350 , n308201 , n17790 );
or ( n17923 , n308349 , n308350 );
buf ( n308352 , n17923 );
buf ( n308353 , n308352 );
xor ( n17926 , n308347 , n308353 );
buf ( n308355 , n17926 );
buf ( n308356 , n308355 );
xor ( n17929 , n308067 , n308073 );
and ( n308358 , n17929 , n308133 );
and ( n308359 , n308067 , n308073 );
or ( n17932 , n308358 , n308359 );
buf ( n17933 , n17932 );
buf ( n308362 , n17933 );
xor ( n17935 , n308146 , n308160 );
and ( n17936 , n17935 , n308182 );
and ( n17937 , n308146 , n308160 );
or ( n308366 , n17936 , n17937 );
buf ( n308367 , n308366 );
buf ( n308368 , n308367 );
xor ( n308369 , n308091 , n17680 );
and ( n17942 , n308369 , n308130 );
and ( n17943 , n308091 , n17680 );
or ( n308372 , n17942 , n17943 );
buf ( n308373 , n308372 );
buf ( n17946 , n308373 );
xor ( n17947 , n308368 , n17946 );
not ( n308376 , n308175 );
not ( n308377 , n293058 );
or ( n17950 , n308376 , n308377 );
buf ( n308379 , n295259 );
buf ( n308380 , n768 );
buf ( n308381 , n810 );
xor ( n308382 , n308380 , n308381 );
buf ( n308383 , n308382 );
buf ( n308384 , n308383 );
nand ( n17957 , n308379 , n308384 );
buf ( n308386 , n17957 );
nand ( n17959 , n17950 , n308386 );
not ( n17960 , n17959 );
buf ( n308389 , n772 );
buf ( n308390 , n806 );
xor ( n308391 , n308389 , n308390 );
buf ( n308392 , n308391 );
not ( n17965 , n308392 );
not ( n308394 , n295437 );
or ( n17967 , n17965 , n308394 );
nand ( n308396 , n17725 , n296617 );
nand ( n17969 , n17967 , n308396 );
not ( n17970 , n17969 );
and ( n308399 , n17960 , n17970 );
not ( n308400 , n17960 );
and ( n308401 , n308400 , n17969 );
nor ( n17974 , n308399 , n308401 );
buf ( n308403 , n296700 );
not ( n308404 , n308403 );
buf ( n308405 , n6209 );
not ( n308406 , n308405 );
buf ( n308407 , n308406 );
buf ( n308408 , n308407 );
not ( n308409 , n308408 );
or ( n308410 , n308404 , n308409 );
buf ( n308411 , n812 );
nand ( n308412 , n308410 , n308411 );
buf ( n308413 , n308412 );
and ( n17986 , n17974 , n308413 );
not ( n308415 , n17974 );
not ( n17988 , n308413 );
and ( n308417 , n308415 , n17988 );
nor ( n17990 , n17986 , n308417 );
buf ( n308419 , n17990 );
xor ( n308420 , n17947 , n308419 );
buf ( n308421 , n308420 );
buf ( n17994 , n308421 );
xor ( n17995 , n308362 , n17994 );
xor ( n308424 , n308185 , n308245 );
and ( n308425 , n308424 , n308252 );
and ( n17998 , n308185 , n308245 );
or ( n308427 , n308425 , n17998 );
buf ( n308428 , n308427 );
buf ( n308429 , n308428 );
xor ( n308430 , n17995 , n308429 );
buf ( n308431 , n308430 );
buf ( n308432 , n308431 );
xor ( n18005 , n308356 , n308432 );
xor ( n308434 , n308136 , n308142 );
and ( n18007 , n308434 , n308255 );
and ( n18008 , n308136 , n308142 );
or ( n308437 , n18007 , n18008 );
buf ( n308438 , n308437 );
buf ( n308439 , n308438 );
xor ( n18012 , n18005 , n308439 );
buf ( n308441 , n18012 );
buf ( n308442 , n308441 );
xor ( n18015 , n308054 , n308060 );
and ( n308444 , n18015 , n308258 );
and ( n308445 , n308054 , n308060 );
or ( n18018 , n308444 , n308445 );
buf ( n308447 , n18018 );
buf ( n18020 , n308447 );
xor ( n18021 , n308442 , n18020 );
buf ( n308450 , n18021 );
and ( n18023 , n17833 , n308266 );
buf ( n308452 , n18023 );
or ( n18025 , n308450 , n308452 );
and ( n18026 , n17841 , n18025 );
not ( n308455 , n13584 );
not ( n308456 , n307915 );
and ( n308457 , n308455 , n308456 );
and ( n18030 , n302371 , n302377 );
not ( n308459 , n302371 );
and ( n308460 , n308459 , n302378 );
nor ( n18033 , n18030 , n308460 );
and ( n308462 , n297868 , n297528 );
or ( n308463 , n18033 , n308462 );
not ( n18036 , n308463 );
nor ( n308465 , n308457 , n18036 );
nand ( n308466 , n18026 , n308465 );
buf ( n18039 , n308466 );
and ( n308468 , n308442 , n18020 );
buf ( n308469 , n308468 );
buf ( n18042 , n308469 );
xor ( n308471 , n308356 , n308432 );
and ( n308472 , n308471 , n308439 );
and ( n18045 , n308356 , n308432 );
or ( n308474 , n308472 , n18045 );
buf ( n308475 , n308474 );
xor ( n308476 , n308307 , n308346 );
and ( n18049 , n308476 , n308353 );
and ( n18050 , n308307 , n308346 );
or ( n18051 , n18049 , n18050 );
buf ( n308480 , n18051 );
buf ( n308481 , n308480 );
xor ( n308482 , n308362 , n17994 );
and ( n308483 , n308482 , n308429 );
and ( n18056 , n308362 , n17994 );
or ( n308485 , n308483 , n18056 );
buf ( n308486 , n308485 );
buf ( n308487 , n308486 );
xor ( n18060 , n308481 , n308487 );
buf ( n308489 , n308383 );
not ( n18062 , n308489 );
buf ( n308491 , n293058 );
not ( n308492 , n308491 );
or ( n18065 , n18062 , n308492 );
buf ( n308494 , n295259 );
buf ( n308495 , n810 );
nand ( n18068 , n308494 , n308495 );
buf ( n308497 , n18068 );
buf ( n308498 , n308497 );
nand ( n308499 , n18065 , n308498 );
buf ( n308500 , n308499 );
buf ( n308501 , n308500 );
not ( n308502 , n308501 );
buf ( n308503 , n308502 );
buf ( n308504 , n308503 );
xor ( n18077 , n308272 , n308286 );
and ( n18078 , n18077 , n308304 );
and ( n18079 , n308272 , n308286 );
or ( n308508 , n18078 , n18079 );
buf ( n308509 , n308508 );
buf ( n308510 , n308509 );
xor ( n308511 , n308504 , n308510 );
nand ( n308512 , n17970 , n17960 );
not ( n18085 , n308512 );
not ( n18086 , n308413 );
or ( n18087 , n18085 , n18086 );
nand ( n18088 , n17969 , n17959 );
nand ( n308517 , n18087 , n18088 );
buf ( n308518 , n308517 );
xor ( n18091 , n308511 , n308518 );
buf ( n18092 , n18091 );
buf ( n308521 , n18092 );
xor ( n308522 , n308368 , n17946 );
and ( n18095 , n308522 , n308419 );
and ( n308524 , n308368 , n17946 );
or ( n308525 , n18095 , n308524 );
buf ( n308526 , n308525 );
buf ( n308527 , n308526 );
xor ( n308528 , n308521 , n308527 );
not ( n18101 , n308323 );
not ( n308530 , n17908 );
or ( n308531 , n18101 , n308530 );
buf ( n308532 , n308323 );
buf ( n308533 , n17908 );
nor ( n308534 , n308532 , n308533 );
buf ( n308535 , n308534 );
or ( n308536 , n308200 , n308535 );
nand ( n18109 , n308531 , n308536 );
buf ( n18110 , n18109 );
and ( n308539 , n308208 , n308209 );
buf ( n308540 , n308539 );
buf ( n308541 , n308540 );
buf ( n308542 , n308317 );
not ( n308543 , n308542 );
buf ( n308544 , n296480 );
not ( n308545 , n308544 );
or ( n18118 , n308543 , n308545 );
buf ( n308547 , n6057 );
buf ( n308548 , n800 );
buf ( n308549 , n777 );
xor ( n308550 , n308548 , n308549 );
buf ( n308551 , n308550 );
buf ( n308552 , n308551 );
nand ( n308553 , n308547 , n308552 );
buf ( n308554 , n308553 );
buf ( n308555 , n308554 );
nand ( n308556 , n18118 , n308555 );
buf ( n308557 , n308556 );
buf ( n308558 , n308557 );
xor ( n308559 , n308541 , n308558 );
buf ( n308560 , n308392 );
not ( n308561 , n308560 );
buf ( n308562 , n296617 );
not ( n18135 , n308562 );
or ( n308564 , n308561 , n18135 );
buf ( n18137 , n295437 );
buf ( n308566 , n806 );
buf ( n308567 , n771 );
xor ( n308568 , n308566 , n308567 );
buf ( n308569 , n308568 );
buf ( n308570 , n308569 );
nand ( n308571 , n18137 , n308570 );
buf ( n308572 , n308571 );
buf ( n308573 , n308572 );
nand ( n308574 , n308564 , n308573 );
buf ( n308575 , n308574 );
buf ( n308576 , n308575 );
xor ( n308577 , n308559 , n308576 );
buf ( n308578 , n308577 );
buf ( n308579 , n308578 );
xor ( n18152 , n18110 , n308579 );
buf ( n308581 , n308330 );
not ( n18154 , n308581 );
buf ( n308583 , n296508 );
not ( n18156 , n308583 );
or ( n18157 , n18154 , n18156 );
buf ( n308586 , n296749 );
xor ( n308587 , n802 , n775 );
buf ( n308588 , n308587 );
nand ( n18161 , n308586 , n308588 );
buf ( n308590 , n18161 );
buf ( n308591 , n308590 );
nand ( n308592 , n18157 , n308591 );
buf ( n308593 , n308592 );
buf ( n308594 , n308593 );
buf ( n308595 , n308279 );
not ( n18168 , n308595 );
buf ( n308597 , n296594 );
not ( n308598 , n308597 );
or ( n18171 , n18168 , n308598 );
buf ( n18172 , n294557 );
xor ( n308601 , n808 , n769 );
buf ( n308602 , n308601 );
nand ( n308603 , n18172 , n308602 );
buf ( n308604 , n308603 );
buf ( n308605 , n308604 );
nand ( n308606 , n18171 , n308605 );
buf ( n308607 , n308606 );
buf ( n308608 , n308607 );
xor ( n308609 , n308594 , n308608 );
buf ( n308610 , n308297 );
not ( n18183 , n308610 );
buf ( n308612 , n296441 );
not ( n308613 , n308612 );
or ( n18186 , n18183 , n308613 );
buf ( n308615 , n296446 );
buf ( n308616 , n773 );
buf ( n308617 , n804 );
xor ( n308618 , n308616 , n308617 );
buf ( n308619 , n308618 );
buf ( n308620 , n308619 );
nand ( n308621 , n308615 , n308620 );
buf ( n308622 , n308621 );
buf ( n308623 , n308622 );
nand ( n308624 , n18186 , n308623 );
buf ( n308625 , n308624 );
buf ( n308626 , n308625 );
xor ( n308627 , n308609 , n308626 );
buf ( n308628 , n308627 );
buf ( n308629 , n308628 );
xor ( n18202 , n18152 , n308629 );
buf ( n308631 , n18202 );
buf ( n308632 , n308631 );
xor ( n18205 , n308528 , n308632 );
buf ( n308634 , n18205 );
buf ( n308635 , n308634 );
xor ( n18208 , n18060 , n308635 );
buf ( n308637 , n18208 );
xor ( n308638 , n308475 , n308637 );
nor ( n18211 , n18042 , n308638 );
nor ( n308640 , n18039 , n18211 );
nand ( n308641 , n17619 , n308640 );
buf ( n18214 , n17619 );
not ( n308643 , n307253 );
not ( n308644 , n307465 );
not ( n18217 , n308644 );
or ( n308646 , n308643 , n18217 );
not ( n18219 , n16813 );
nand ( n18220 , n308646 , n18219 );
nor ( n308649 , n17530 , n17506 );
not ( n308650 , n17559 );
nor ( n18223 , n308650 , n307977 );
nand ( n18224 , n308649 , n18223 );
not ( n18225 , n18224 );
not ( n18226 , n18225 );
not ( n308655 , n307729 );
or ( n308656 , n18226 , n308655 );
buf ( n18229 , n308025 );
and ( n18230 , n18223 , n18229 );
not ( n18231 , n17559 );
not ( n18232 , n17607 );
or ( n308661 , n18231 , n18232 );
not ( n308662 , n308038 );
nand ( n18235 , n308661 , n308662 );
nor ( n308664 , n18230 , n18235 );
nand ( n18237 , n308656 , n308664 );
not ( n308666 , n18237 );
not ( n18239 , n308649 );
not ( n18240 , n307729 );
or ( n308669 , n18239 , n18240 );
not ( n308670 , n18229 );
nand ( n308671 , n308669 , n308670 );
not ( n18244 , n308671 );
nand ( n308673 , n307749 , n307808 );
nand ( n308674 , n17446 , n307749 );
not ( n18247 , n16995 );
not ( n308676 , n307414 );
or ( n308677 , n18247 , n308676 );
nand ( n18250 , n308677 , n17027 );
nand ( n308679 , n307309 , n17029 );
not ( n308680 , n308679 );
and ( n18253 , n18250 , n308680 );
not ( n308682 , n18250 );
and ( n18255 , n308682 , n308679 );
nor ( n18256 , n18253 , n18255 );
not ( n308685 , n308638 );
not ( n308686 , n308469 );
and ( n18259 , n308685 , n308686 );
xor ( n308688 , n308481 , n308487 );
and ( n308689 , n308688 , n308635 );
and ( n18262 , n308481 , n308487 );
or ( n308691 , n308689 , n18262 );
buf ( n308692 , n308691 );
xor ( n308693 , n308541 , n308558 );
and ( n18266 , n308693 , n308576 );
and ( n308695 , n308541 , n308558 );
or ( n18268 , n18266 , n308695 );
buf ( n308697 , n18268 );
buf ( n18270 , n308697 );
buf ( n308699 , n308569 );
not ( n308700 , n308699 );
buf ( n308701 , n296617 );
not ( n308702 , n308701 );
or ( n308703 , n308700 , n308702 );
buf ( n308704 , n295437 );
buf ( n308705 , n806 );
buf ( n308706 , n770 );
xor ( n18279 , n308705 , n308706 );
buf ( n18280 , n18279 );
buf ( n308709 , n18280 );
nand ( n308710 , n308704 , n308709 );
buf ( n308711 , n308710 );
buf ( n308712 , n308711 );
nand ( n308713 , n308703 , n308712 );
buf ( n308714 , n308713 );
buf ( n308715 , n308714 );
buf ( n308716 , n308587 );
not ( n308717 , n308716 );
buf ( n308718 , n296508 );
not ( n308719 , n308718 );
or ( n18292 , n308717 , n308719 );
buf ( n308721 , n296749 );
buf ( n18294 , n802 );
buf ( n308723 , n774 );
xor ( n308724 , n18294 , n308723 );
buf ( n308725 , n308724 );
buf ( n308726 , n308725 );
nand ( n308727 , n308721 , n308726 );
buf ( n308728 , n308727 );
buf ( n308729 , n308728 );
nand ( n308730 , n18292 , n308729 );
buf ( n308731 , n308730 );
buf ( n308732 , n308731 );
xor ( n308733 , n308715 , n308732 );
buf ( n308734 , n308551 );
not ( n308735 , n308734 );
buf ( n308736 , n296480 );
not ( n308737 , n308736 );
or ( n18310 , n308735 , n308737 );
buf ( n308739 , n6057 );
buf ( n18312 , n800 );
buf ( n308741 , n776 );
xor ( n308742 , n18312 , n308741 );
buf ( n308743 , n308742 );
buf ( n308744 , n308743 );
nand ( n308745 , n308739 , n308744 );
buf ( n308746 , n308745 );
buf ( n308747 , n308746 );
nand ( n308748 , n18310 , n308747 );
buf ( n308749 , n308748 );
buf ( n308750 , n308749 );
xor ( n308751 , n308733 , n308750 );
buf ( n308752 , n308751 );
buf ( n308753 , n308752 );
xor ( n308754 , n18270 , n308753 );
buf ( n308755 , n308601 );
not ( n18328 , n308755 );
buf ( n308757 , n296594 );
not ( n18330 , n308757 );
or ( n308759 , n18328 , n18330 );
buf ( n308760 , n294557 );
xor ( n18333 , n808 , n768 );
buf ( n308762 , n18333 );
nand ( n18335 , n308760 , n308762 );
buf ( n308764 , n18335 );
buf ( n308765 , n308764 );
nand ( n308766 , n308759 , n308765 );
buf ( n308767 , n308766 );
buf ( n308768 , n308767 );
buf ( n308769 , n295259 );
buf ( n308770 , n293058 );
or ( n18343 , n308769 , n308770 );
buf ( n308772 , n810 );
nand ( n18345 , n18343 , n308772 );
buf ( n308774 , n18345 );
buf ( n308775 , n308774 );
xor ( n308776 , n308768 , n308775 );
buf ( n308777 , n308619 );
not ( n18350 , n308777 );
buf ( n308779 , n296441 );
not ( n308780 , n308779 );
or ( n18353 , n18350 , n308780 );
not ( n18354 , n296664 );
not ( n18355 , n18354 );
buf ( n308784 , n18355 );
buf ( n308785 , n772 );
buf ( n18358 , n804 );
xor ( n18359 , n308785 , n18358 );
buf ( n308788 , n18359 );
buf ( n18361 , n308788 );
nand ( n18362 , n308784 , n18361 );
buf ( n18363 , n18362 );
buf ( n308792 , n18363 );
nand ( n18365 , n18353 , n308792 );
buf ( n18366 , n18365 );
buf ( n308795 , n18366 );
xor ( n308796 , n308776 , n308795 );
buf ( n308797 , n308796 );
buf ( n308798 , n308797 );
xor ( n18371 , n308754 , n308798 );
buf ( n308800 , n18371 );
buf ( n308801 , n308800 );
and ( n18374 , n308314 , n308315 );
buf ( n308803 , n18374 );
buf ( n308804 , n308803 );
buf ( n308805 , n308500 );
xor ( n308806 , n308804 , n308805 );
xor ( n308807 , n308594 , n308608 );
and ( n18380 , n308807 , n308626 );
and ( n308809 , n308594 , n308608 );
or ( n308810 , n18380 , n308809 );
buf ( n308811 , n308810 );
buf ( n308812 , n308811 );
xor ( n18385 , n308806 , n308812 );
buf ( n308814 , n18385 );
buf ( n18387 , n308814 );
xor ( n18388 , n308504 , n308510 );
and ( n308817 , n18388 , n308518 );
and ( n308818 , n308504 , n308510 );
or ( n18391 , n308817 , n308818 );
buf ( n308820 , n18391 );
buf ( n308821 , n308820 );
xor ( n18394 , n18387 , n308821 );
xor ( n308823 , n18110 , n308579 );
and ( n18396 , n308823 , n308629 );
and ( n308825 , n18110 , n308579 );
or ( n308826 , n18396 , n308825 );
buf ( n308827 , n308826 );
buf ( n308828 , n308827 );
xor ( n308829 , n18394 , n308828 );
buf ( n308830 , n308829 );
buf ( n308831 , n308830 );
xor ( n308832 , n308801 , n308831 );
xor ( n18405 , n308521 , n308527 );
and ( n308834 , n18405 , n308632 );
and ( n308835 , n308521 , n308527 );
or ( n308836 , n308834 , n308835 );
buf ( n308837 , n308836 );
buf ( n308838 , n308837 );
xor ( n308839 , n308832 , n308838 );
buf ( n308840 , n308839 );
xor ( n18413 , n308692 , n308840 );
and ( n308842 , n308637 , n308475 );
nor ( n308843 , n18413 , n308842 );
nor ( n18416 , n18259 , n308843 );
not ( n18417 , n18416 );
nand ( n308846 , n13584 , n307915 );
not ( n18419 , n308463 );
or ( n18420 , n308846 , n18419 );
nand ( n308849 , n18033 , n308462 );
nand ( n18422 , n18420 , n308849 );
not ( n308851 , n18422 );
and ( n18424 , n17841 , n18025 );
not ( n18425 , n18424 );
or ( n18426 , n308851 , n18425 );
nor ( n308855 , n308452 , n308450 );
not ( n18428 , n308855 );
nand ( n18429 , n308268 , n11951 );
not ( n18430 , n18429 );
and ( n18431 , n18428 , n18430 );
and ( n18432 , n308452 , n308450 );
nor ( n18433 , n18431 , n18432 );
nand ( n18434 , n18426 , n18433 );
buf ( n18435 , n18434 );
not ( n308864 , n18435 );
or ( n18437 , n18417 , n308864 );
and ( n308866 , n308638 , n308469 );
not ( n308867 , n308866 );
not ( n18440 , n308843 );
not ( n308869 , n18440 );
or ( n308870 , n308867 , n308869 );
nand ( n308871 , n308842 , n18413 );
nand ( n308872 , n308870 , n308871 );
buf ( n18445 , n308872 );
not ( n308874 , n18445 );
nand ( n308875 , n18437 , n308874 );
not ( n18448 , n308875 );
not ( n18449 , n18211 );
and ( n308878 , n18435 , n18449 );
nor ( n18451 , n308878 , n308866 );
buf ( n308880 , n18280 );
not ( n308881 , n308880 );
buf ( n308882 , n296617 );
not ( n18455 , n308882 );
or ( n308884 , n308881 , n18455 );
buf ( n308885 , n769 );
buf ( n308886 , n806 );
xnor ( n18459 , n308885 , n308886 );
buf ( n308888 , n18459 );
buf ( n308889 , n308888 );
not ( n18462 , n308889 );
buf ( n308891 , n295437 );
nand ( n18464 , n18462 , n308891 );
buf ( n18465 , n18464 );
buf ( n308894 , n18465 );
nand ( n18467 , n308884 , n308894 );
buf ( n308896 , n18467 );
buf ( n308897 , n308896 );
buf ( n308898 , n18333 );
not ( n308899 , n308898 );
buf ( n308900 , n296594 );
not ( n18473 , n308900 );
or ( n308902 , n308899 , n18473 );
buf ( n308903 , n6301 );
buf ( n308904 , n808 );
nand ( n308905 , n308903 , n308904 );
buf ( n308906 , n308905 );
buf ( n308907 , n308906 );
nand ( n18480 , n308902 , n308907 );
buf ( n18481 , n18480 );
buf ( n308910 , n18481 );
buf ( n308911 , n308725 );
not ( n308912 , n308911 );
buf ( n308913 , n296508 );
not ( n308914 , n308913 );
or ( n18487 , n308912 , n308914 );
buf ( n308916 , n296749 );
buf ( n18489 , n773 );
buf ( n308918 , n802 );
xor ( n18491 , n18489 , n308918 );
buf ( n18492 , n18491 );
buf ( n18493 , n18492 );
nand ( n18494 , n308916 , n18493 );
buf ( n18495 , n18494 );
buf ( n308924 , n18495 );
nand ( n18497 , n18487 , n308924 );
buf ( n18498 , n18497 );
buf ( n308927 , n18498 );
or ( n18500 , n308910 , n308927 );
buf ( n308929 , n308743 );
not ( n18502 , n308929 );
buf ( n308931 , n296480 );
not ( n18504 , n308931 );
or ( n308933 , n18502 , n18504 );
buf ( n308934 , n775 );
buf ( n308935 , n800 );
xnor ( n18508 , n308934 , n308935 );
buf ( n18509 , n18508 );
buf ( n308938 , n18509 );
not ( n18511 , n308938 );
buf ( n308940 , n6057 );
nand ( n308941 , n18511 , n308940 );
buf ( n308942 , n308941 );
buf ( n308943 , n308942 );
nand ( n18516 , n308933 , n308943 );
buf ( n18517 , n18516 );
buf ( n308946 , n18517 );
nand ( n18519 , n18500 , n308946 );
buf ( n308948 , n18519 );
buf ( n308949 , n308948 );
buf ( n308950 , n18481 );
buf ( n308951 , n18498 );
nand ( n308952 , n308950 , n308951 );
buf ( n308953 , n308952 );
buf ( n308954 , n308953 );
nand ( n308955 , n308949 , n308954 );
buf ( n308956 , n308955 );
buf ( n308957 , n308956 );
xor ( n18530 , n308897 , n308957 );
and ( n308959 , n18312 , n308741 );
buf ( n308960 , n308959 );
buf ( n308961 , n308960 );
buf ( n18534 , n804 );
buf ( n308963 , n771 );
xor ( n308964 , n18534 , n308963 );
buf ( n308965 , n308964 );
buf ( n308966 , n308965 );
not ( n18539 , n308966 );
buf ( n308968 , n296441 );
not ( n18541 , n308968 );
or ( n308970 , n18539 , n18541 );
buf ( n308971 , n297395 );
buf ( n308972 , n804 );
buf ( n308973 , n770 );
xor ( n308974 , n308972 , n308973 );
buf ( n308975 , n308974 );
buf ( n308976 , n308975 );
nand ( n18549 , n308971 , n308976 );
buf ( n308978 , n18549 );
buf ( n308979 , n308978 );
nand ( n18552 , n308970 , n308979 );
buf ( n308981 , n18552 );
buf ( n308982 , n308981 );
xor ( n18555 , n308961 , n308982 );
buf ( n18556 , n296480 );
not ( n18557 , n18556 );
buf ( n18558 , n18557 );
buf ( n308987 , n18558 );
buf ( n308988 , n18509 );
or ( n308989 , n308987 , n308988 );
buf ( n308990 , n6056 );
not ( n18563 , n308990 );
buf ( n308992 , n18563 );
buf ( n308993 , n308992 );
buf ( n308994 , n774 );
buf ( n308995 , n800 );
xnor ( n308996 , n308994 , n308995 );
buf ( n308997 , n308996 );
buf ( n308998 , n308997 );
or ( n308999 , n308993 , n308998 );
nand ( n309000 , n308989 , n308999 );
buf ( n309001 , n309000 );
buf ( n309002 , n309001 );
xor ( n18575 , n18555 , n309002 );
buf ( n309004 , n18575 );
buf ( n309005 , n309004 );
and ( n18578 , n18530 , n309005 );
and ( n309007 , n308897 , n308957 );
or ( n309008 , n18578 , n309007 );
buf ( n309009 , n309008 );
buf ( n309010 , n775 );
buf ( n309011 , n800 );
and ( n18584 , n309010 , n309011 );
buf ( n18585 , n18584 );
buf ( n18586 , n18585 );
buf ( n309015 , n806 );
buf ( n309016 , n768 );
xor ( n309017 , n309015 , n309016 );
buf ( n309018 , n309017 );
buf ( n309019 , n309018 );
not ( n309020 , n309019 );
buf ( n309021 , n296617 );
not ( n309022 , n309021 );
or ( n18595 , n309020 , n309022 );
buf ( n309024 , n295437 );
buf ( n18597 , n806 );
nand ( n18598 , n309024 , n18597 );
buf ( n309027 , n18598 );
buf ( n309028 , n309027 );
nand ( n18601 , n18595 , n309028 );
buf ( n18602 , n18601 );
buf ( n309031 , n18602 );
xor ( n18604 , n18586 , n309031 );
buf ( n309033 , n308997 );
not ( n309034 , n309033 );
buf ( n309035 , n309034 );
buf ( n309036 , n309035 );
not ( n18609 , n309036 );
buf ( n309038 , n296480 );
not ( n18611 , n309038 );
or ( n309040 , n18609 , n18611 );
buf ( n309041 , n800 );
buf ( n309042 , n773 );
xnor ( n309043 , n309041 , n309042 );
buf ( n309044 , n309043 );
buf ( n309045 , n309044 );
not ( n309046 , n309045 );
buf ( n309047 , n6057 );
nand ( n18620 , n309046 , n309047 );
buf ( n309049 , n18620 );
buf ( n309050 , n309049 );
nand ( n309051 , n309040 , n309050 );
buf ( n309052 , n309051 );
buf ( n309053 , n309052 );
xor ( n309054 , n18604 , n309053 );
buf ( n309055 , n309054 );
buf ( n18628 , n309055 );
buf ( n309057 , n11650 );
not ( n18630 , n309057 );
buf ( n309059 , n296594 );
not ( n309060 , n309059 );
buf ( n309061 , n309060 );
buf ( n309062 , n309061 );
not ( n309063 , n309062 );
or ( n18636 , n18630 , n309063 );
buf ( n309065 , n808 );
nand ( n309066 , n18636 , n309065 );
buf ( n309067 , n309066 );
buf ( n309068 , n309067 );
buf ( n309069 , n18492 );
not ( n18642 , n309069 );
buf ( n309071 , n296508 );
not ( n18644 , n309071 );
or ( n309073 , n18642 , n18644 );
buf ( n309074 , n296749 );
buf ( n309075 , n772 );
buf ( n309076 , n802 );
xor ( n18649 , n309075 , n309076 );
buf ( n18650 , n18649 );
buf ( n309079 , n18650 );
nand ( n18652 , n309074 , n309079 );
buf ( n18653 , n18652 );
buf ( n309082 , n18653 );
nand ( n18655 , n309073 , n309082 );
buf ( n309084 , n18655 );
buf ( n18657 , n309084 );
xor ( n18658 , n309068 , n18657 );
buf ( n309087 , n296617 );
not ( n309088 , n309087 );
buf ( n309089 , n309088 );
buf ( n309090 , n309089 );
buf ( n309091 , n308888 );
or ( n18664 , n309090 , n309091 );
not ( n18665 , n295437 );
buf ( n309094 , n18665 );
buf ( n309095 , n309018 );
not ( n18668 , n309095 );
buf ( n18669 , n18668 );
buf ( n309098 , n18669 );
or ( n309099 , n309094 , n309098 );
nand ( n18672 , n18664 , n309099 );
buf ( n18673 , n18672 );
buf ( n309102 , n18673 );
and ( n309103 , n18658 , n309102 );
and ( n18676 , n309068 , n18657 );
or ( n309105 , n309103 , n18676 );
buf ( n309106 , n309105 );
buf ( n309107 , n309106 );
xor ( n309108 , n18628 , n309107 );
buf ( n309109 , n308975 );
not ( n18682 , n309109 );
buf ( n309111 , n296441 );
not ( n18684 , n309111 );
or ( n18685 , n18682 , n18684 );
buf ( n309114 , n804 );
buf ( n309115 , n769 );
xnor ( n18688 , n309114 , n309115 );
buf ( n18689 , n18688 );
buf ( n309118 , n18689 );
not ( n18691 , n309118 );
buf ( n309120 , n296446 );
nand ( n18693 , n18691 , n309120 );
buf ( n309122 , n18693 );
buf ( n309123 , n309122 );
nand ( n18696 , n18685 , n309123 );
buf ( n309125 , n18696 );
buf ( n309126 , n309125 );
not ( n18699 , n309126 );
buf ( n309128 , n18699 );
buf ( n309129 , n309128 );
buf ( n309130 , n18650 );
not ( n309131 , n309130 );
buf ( n309132 , n296508 );
not ( n18705 , n309132 );
or ( n309134 , n309131 , n18705 );
buf ( n309135 , n296749 );
buf ( n309136 , n771 );
buf ( n309137 , n802 );
xor ( n309138 , n309136 , n309137 );
buf ( n309139 , n309138 );
buf ( n309140 , n309139 );
nand ( n309141 , n309135 , n309140 );
buf ( n309142 , n309141 );
buf ( n309143 , n309142 );
nand ( n309144 , n309134 , n309143 );
buf ( n309145 , n309144 );
buf ( n309146 , n309145 );
xor ( n309147 , n309129 , n309146 );
xor ( n18720 , n308961 , n308982 );
and ( n309149 , n18720 , n309002 );
and ( n309150 , n308961 , n308982 );
or ( n18723 , n309149 , n309150 );
buf ( n309152 , n18723 );
buf ( n309153 , n309152 );
xor ( n18726 , n309147 , n309153 );
buf ( n309155 , n18726 );
buf ( n309156 , n309155 );
xor ( n18729 , n309108 , n309156 );
buf ( n309158 , n18729 );
xor ( n18731 , n309009 , n309158 );
xor ( n309160 , n309068 , n18657 );
xor ( n309161 , n309160 , n309102 );
buf ( n309162 , n309161 );
not ( n309163 , n309162 );
and ( n309164 , n308548 , n308549 );
buf ( n309165 , n309164 );
buf ( n309166 , n309165 );
buf ( n309167 , n308788 );
not ( n18740 , n309167 );
buf ( n309169 , n296441 );
not ( n309170 , n309169 );
or ( n18743 , n18740 , n309170 );
buf ( n309172 , n6017 );
buf ( n309173 , n308965 );
nand ( n18746 , n309172 , n309173 );
buf ( n309175 , n18746 );
buf ( n309176 , n309175 );
nand ( n18749 , n18743 , n309176 );
buf ( n309178 , n18749 );
buf ( n309179 , n309178 );
xor ( n18752 , n309166 , n309179 );
buf ( n309181 , n308896 );
not ( n309182 , n309181 );
buf ( n309183 , n309182 );
buf ( n309184 , n309183 );
and ( n309185 , n18752 , n309184 );
and ( n18758 , n309166 , n309179 );
or ( n309187 , n309185 , n18758 );
buf ( n309188 , n309187 );
not ( n309189 , n309188 );
nand ( n18762 , n309163 , n309189 );
not ( n309191 , n18762 );
xor ( n18764 , n308897 , n308957 );
xor ( n309193 , n18764 , n309005 );
buf ( n309194 , n309193 );
buf ( n309195 , n309194 );
not ( n18768 , n309195 );
or ( n309197 , n309191 , n18768 );
nand ( n309198 , n309188 , n309162 );
nand ( n18771 , n309197 , n309198 );
and ( n309200 , n18731 , n18771 );
and ( n18773 , n309009 , n309158 );
or ( n18774 , n309200 , n18773 );
buf ( n309203 , n18774 );
xor ( n309204 , n309129 , n309146 );
and ( n18777 , n309204 , n309153 );
and ( n309206 , n309129 , n309146 );
or ( n18779 , n18777 , n309206 );
buf ( n309208 , n18779 );
buf ( n309209 , n309208 );
xor ( n18782 , n18586 , n309031 );
and ( n309211 , n18782 , n309053 );
and ( n309212 , n18586 , n309031 );
or ( n309213 , n309211 , n309212 );
buf ( n309214 , n309213 );
buf ( n309215 , n18558 );
buf ( n309216 , n309044 );
or ( n18789 , n309215 , n309216 );
buf ( n309218 , n308992 );
buf ( n18791 , n772 );
buf ( n18792 , n800 );
xnor ( n18793 , n18791 , n18792 );
buf ( n18794 , n18793 );
buf ( n309223 , n18794 );
or ( n18796 , n309218 , n309223 );
nand ( n18797 , n18789 , n18796 );
buf ( n309226 , n18797 );
buf ( n309227 , n302341 );
buf ( n309228 , n18689 );
or ( n18801 , n309227 , n309228 );
not ( n18802 , n17690 );
buf ( n309231 , n18802 );
buf ( n309232 , n768 );
buf ( n309233 , n804 );
not ( n18806 , n309233 );
buf ( n309235 , n18806 );
buf ( n309236 , n309235 );
and ( n18809 , n309232 , n309236 );
not ( n309238 , n309232 );
buf ( n309239 , n804 );
and ( n309240 , n309238 , n309239 );
nor ( n18813 , n18809 , n309240 );
buf ( n309242 , n18813 );
buf ( n309243 , n309242 );
or ( n309244 , n309231 , n309243 );
nand ( n18817 , n18801 , n309244 );
buf ( n309246 , n18817 );
xor ( n18819 , n309226 , n309246 );
buf ( n309248 , n18665 );
not ( n309249 , n309248 );
buf ( n309250 , n309089 );
not ( n309251 , n309250 );
or ( n309252 , n309249 , n309251 );
buf ( n309253 , n806 );
nand ( n309254 , n309252 , n309253 );
buf ( n309255 , n309254 );
xor ( n18828 , n18819 , n309255 );
xor ( n18829 , n309214 , n18828 );
buf ( n18830 , n774 );
buf ( n309259 , n800 );
and ( n18832 , n18830 , n309259 );
buf ( n18833 , n18832 );
buf ( n309262 , n18833 );
buf ( n309263 , n309139 );
not ( n309264 , n309263 );
buf ( n309265 , n296508 );
not ( n309266 , n309265 );
or ( n309267 , n309264 , n309266 );
buf ( n309268 , n802 );
buf ( n309269 , n770 );
not ( n18842 , n309269 );
buf ( n309271 , n18842 );
buf ( n309272 , n309271 );
and ( n18845 , n309268 , n309272 );
not ( n18846 , n309268 );
buf ( n309275 , n770 );
and ( n18848 , n18846 , n309275 );
nor ( n18849 , n18845 , n18848 );
buf ( n309278 , n18849 );
buf ( n309279 , n309278 );
not ( n18852 , n309279 );
buf ( n309281 , n296749 );
nand ( n18854 , n18852 , n309281 );
buf ( n309283 , n18854 );
buf ( n309284 , n309283 );
nand ( n18857 , n309267 , n309284 );
buf ( n309286 , n18857 );
buf ( n309287 , n309286 );
xor ( n18860 , n309262 , n309287 );
buf ( n309289 , n309125 );
xor ( n309290 , n18860 , n309289 );
buf ( n309291 , n309290 );
xor ( n309292 , n18829 , n309291 );
buf ( n309293 , n309292 );
xor ( n18866 , n309209 , n309293 );
xor ( n309295 , n18628 , n309107 );
and ( n309296 , n309295 , n309156 );
and ( n309297 , n18628 , n309107 );
or ( n309298 , n309296 , n309297 );
buf ( n309299 , n309298 );
buf ( n309300 , n309299 );
xor ( n309301 , n18866 , n309300 );
buf ( n309302 , n309301 );
buf ( n309303 , n309302 );
and ( n18876 , n309203 , n309303 );
buf ( n309305 , n18876 );
xor ( n309306 , n309262 , n309287 );
and ( n309307 , n309306 , n309289 );
and ( n18880 , n309262 , n309287 );
or ( n309309 , n309307 , n18880 );
buf ( n309310 , n309309 );
or ( n18883 , n309242 , n302341 );
or ( n309312 , n18354 , n309235 );
nand ( n309313 , n18883 , n309312 );
not ( n18886 , n309313 );
buf ( n309315 , n773 );
buf ( n309316 , n800 );
and ( n18889 , n309315 , n309316 );
buf ( n309318 , n18889 );
buf ( n309319 , n18794 );
not ( n18892 , n309319 );
buf ( n309321 , n18892 );
buf ( n309322 , n309321 );
not ( n309323 , n309322 );
buf ( n309324 , n296480 );
not ( n18897 , n309324 );
or ( n309326 , n309323 , n18897 );
buf ( n18899 , n771 );
buf ( n309328 , n800 );
xnor ( n309329 , n18899 , n309328 );
buf ( n309330 , n309329 );
buf ( n309331 , n309330 );
not ( n309332 , n309331 );
buf ( n309333 , n6057 );
nand ( n309334 , n309332 , n309333 );
buf ( n309335 , n309334 );
buf ( n309336 , n309335 );
nand ( n309337 , n309326 , n309336 );
buf ( n309338 , n309337 );
xor ( n18911 , n309318 , n309338 );
buf ( n18912 , n296508 );
not ( n309341 , n18912 );
buf ( n309342 , n309341 );
buf ( n309343 , n309342 );
buf ( n309344 , n309278 );
or ( n18917 , n309343 , n309344 );
buf ( n309346 , n296749 );
not ( n18919 , n309346 );
buf ( n309348 , n18919 );
buf ( n309349 , n309348 );
buf ( n309350 , n802 );
not ( n18923 , n309350 );
buf ( n309352 , n18923 );
buf ( n309353 , n309352 );
buf ( n309354 , n769 );
and ( n309355 , n309353 , n309354 );
buf ( n309356 , n299244 );
buf ( n309357 , n802 );
and ( n18930 , n309356 , n309357 );
nor ( n309359 , n309355 , n18930 );
buf ( n309360 , n309359 );
buf ( n309361 , n309360 );
or ( n18934 , n309349 , n309361 );
nand ( n309363 , n18917 , n18934 );
buf ( n309364 , n309363 );
xor ( n18937 , n18911 , n309364 );
xor ( n309366 , n18886 , n18937 );
xor ( n309367 , n309226 , n309246 );
and ( n18940 , n309367 , n309255 );
and ( n309369 , n309226 , n309246 );
or ( n309370 , n18940 , n309369 );
xor ( n18943 , n309366 , n309370 );
xor ( n309372 , n309310 , n18943 );
xor ( n309373 , n309214 , n18828 );
and ( n309374 , n309373 , n309291 );
and ( n309375 , n309214 , n18828 );
or ( n18948 , n309374 , n309375 );
xor ( n309377 , n309372 , n18948 );
buf ( n309378 , n309377 );
xor ( n18951 , n309209 , n309293 );
and ( n309380 , n18951 , n309300 );
and ( n309381 , n309209 , n309293 );
or ( n18954 , n309380 , n309381 );
buf ( n309383 , n18954 );
buf ( n309384 , n309383 );
xor ( n309385 , n309378 , n309384 );
buf ( n309386 , n309385 );
nor ( n18959 , n309305 , n309386 );
and ( n309388 , n309378 , n309384 );
buf ( n309389 , n309388 );
buf ( n309390 , n296441 );
buf ( n309391 , n18355 );
or ( n18964 , n309390 , n309391 );
buf ( n309393 , n804 );
nand ( n18966 , n18964 , n309393 );
buf ( n18967 , n18966 );
buf ( n309396 , n18967 );
buf ( n309397 , n772 );
buf ( n18970 , n800 );
and ( n18971 , n309397 , n18970 );
buf ( n18972 , n18971 );
buf ( n309401 , n18972 );
xor ( n18974 , n309396 , n309401 );
buf ( n309403 , n309342 );
buf ( n309404 , n309360 );
or ( n309405 , n309403 , n309404 );
buf ( n309406 , n309348 );
buf ( n309407 , n768 );
buf ( n309408 , n309352 );
and ( n18981 , n309407 , n309408 );
not ( n309410 , n309407 );
buf ( n309411 , n802 );
and ( n309412 , n309410 , n309411 );
nor ( n309413 , n18981 , n309412 );
buf ( n309414 , n309413 );
buf ( n309415 , n309414 );
or ( n309416 , n309406 , n309415 );
nand ( n309417 , n309405 , n309416 );
buf ( n309418 , n309417 );
buf ( n309419 , n309418 );
xor ( n309420 , n18974 , n309419 );
buf ( n309421 , n309420 );
xor ( n18994 , n309318 , n309338 );
and ( n309423 , n18994 , n309364 );
and ( n309424 , n309318 , n309338 );
nor ( n18997 , n309423 , n309424 );
buf ( n309426 , n18558 );
buf ( n309427 , n309330 );
or ( n19000 , n309426 , n309427 );
buf ( n309429 , n308992 );
buf ( n309430 , n298423 );
buf ( n309431 , n770 );
and ( n19004 , n309430 , n309431 );
buf ( n309433 , n309271 );
buf ( n309434 , n800 );
and ( n19007 , n309433 , n309434 );
nor ( n19008 , n19004 , n19007 );
buf ( n309437 , n19008 );
buf ( n309438 , n309437 );
or ( n19011 , n309429 , n309438 );
nand ( n19012 , n19000 , n19011 );
buf ( n309441 , n19012 );
not ( n309442 , n309441 );
and ( n19015 , n309313 , n309442 );
not ( n309444 , n309313 );
and ( n309445 , n309444 , n309441 );
nor ( n309446 , n19015 , n309445 );
xor ( n309447 , n18997 , n309446 );
xor ( n19020 , n309421 , n309447 );
xor ( n309449 , n18886 , n18937 );
and ( n309450 , n309449 , n309370 );
and ( n19023 , n18886 , n18937 );
or ( n309452 , n309450 , n19023 );
xor ( n309453 , n19020 , n309452 );
buf ( n309454 , n309453 );
xor ( n309455 , n309310 , n18943 );
and ( n309456 , n309455 , n18948 );
and ( n19029 , n309310 , n18943 );
or ( n309458 , n309456 , n19029 );
buf ( n309459 , n309458 );
xor ( n19032 , n309454 , n309459 );
buf ( n309461 , n19032 );
nor ( n309462 , n309389 , n309461 );
nor ( n309463 , n18959 , n309462 );
xor ( n309464 , n308768 , n308775 );
and ( n19037 , n309464 , n308795 );
and ( n309466 , n308768 , n308775 );
or ( n309467 , n19037 , n309466 );
buf ( n309468 , n309467 );
buf ( n309469 , n309468 );
xor ( n309470 , n308715 , n308732 );
and ( n19043 , n309470 , n308750 );
and ( n19044 , n308715 , n308732 );
or ( n309473 , n19043 , n19044 );
buf ( n309474 , n309473 );
buf ( n309475 , n309474 );
xor ( n19048 , n309469 , n309475 );
buf ( n309477 , n18498 );
buf ( n309478 , n18481 );
xor ( n309479 , n309477 , n309478 );
buf ( n309480 , n309479 );
buf ( n309481 , n309480 );
buf ( n309482 , n18517 );
xor ( n309483 , n309481 , n309482 );
buf ( n309484 , n309483 );
buf ( n309485 , n309484 );
and ( n309486 , n19048 , n309485 );
and ( n19059 , n309469 , n309475 );
or ( n309488 , n309486 , n19059 );
buf ( n309489 , n309488 );
not ( n309490 , n309489 );
xor ( n309491 , n309166 , n309179 );
xor ( n19064 , n309491 , n309184 );
buf ( n309493 , n19064 );
buf ( n309494 , n309493 );
xor ( n19067 , n308804 , n308805 );
and ( n19068 , n19067 , n308812 );
and ( n19069 , n308804 , n308805 );
or ( n19070 , n19068 , n19069 );
buf ( n309499 , n19070 );
buf ( n309500 , n309499 );
xor ( n19073 , n309494 , n309500 );
xor ( n19074 , n18270 , n308753 );
and ( n19075 , n19074 , n308798 );
and ( n19076 , n18270 , n308753 );
or ( n19077 , n19075 , n19076 );
buf ( n309506 , n19077 );
buf ( n309507 , n309506 );
and ( n19080 , n19073 , n309507 );
and ( n19081 , n309494 , n309500 );
or ( n19082 , n19080 , n19081 );
buf ( n309511 , n19082 );
not ( n19084 , n309511 );
nand ( n309513 , n309490 , n19084 );
not ( n309514 , n309513 );
and ( n309515 , n309162 , n309189 );
not ( n309516 , n309162 );
and ( n19089 , n309516 , n309188 );
nor ( n309518 , n309515 , n19089 );
and ( n309519 , n309518 , n309195 );
not ( n19092 , n309518 );
not ( n309521 , n309195 );
and ( n309522 , n19092 , n309521 );
or ( n19095 , n309519 , n309522 );
not ( n309524 , n19095 );
or ( n19097 , n309514 , n309524 );
not ( n19098 , n19084 );
nand ( n309527 , n19098 , n309489 );
nand ( n309528 , n19097 , n309527 );
xor ( n19101 , n309009 , n309158 );
xor ( n309530 , n19101 , n18771 );
and ( n309531 , n309528 , n309530 );
xor ( n19104 , n309203 , n309303 );
buf ( n309533 , n19104 );
nor ( n19106 , n309531 , n309533 );
xor ( n19107 , n309489 , n19095 );
xor ( n19108 , n19107 , n309511 );
xor ( n309537 , n309469 , n309475 );
xor ( n19110 , n309537 , n309485 );
buf ( n309539 , n19110 );
buf ( n309540 , n309539 );
xor ( n309541 , n18387 , n308821 );
and ( n19114 , n309541 , n308828 );
and ( n309543 , n18387 , n308821 );
or ( n19116 , n19114 , n309543 );
buf ( n309545 , n19116 );
buf ( n309546 , n309545 );
xor ( n309547 , n309540 , n309546 );
xor ( n309548 , n309494 , n309500 );
xor ( n19121 , n309548 , n309507 );
buf ( n309550 , n19121 );
buf ( n309551 , n309550 );
and ( n19124 , n309547 , n309551 );
and ( n309553 , n309540 , n309546 );
or ( n309554 , n19124 , n309553 );
buf ( n309555 , n309554 );
and ( n19128 , n19108 , n309555 );
not ( n309557 , n309530 );
not ( n19130 , n309557 );
not ( n309559 , n309528 );
or ( n309560 , n19130 , n309559 );
or ( n19133 , n309528 , n309557 );
nand ( n309562 , n309560 , n19133 );
nand ( n309563 , n19128 , n309562 );
or ( n309564 , n19106 , n309563 );
nand ( n309565 , n309531 , n309533 );
nand ( n19138 , n309564 , n309565 );
and ( n309567 , n309463 , n19138 );
nand ( n309568 , n309305 , n309386 );
or ( n19141 , n309462 , n309568 );
nand ( n309570 , n309389 , n309461 );
nand ( n309571 , n19141 , n309570 );
nor ( n19144 , n309567 , n309571 );
not ( n309573 , n19144 );
and ( n19146 , n309454 , n309459 );
buf ( n309575 , n19146 );
xor ( n309576 , n309396 , n309401 );
and ( n19149 , n309576 , n309419 );
and ( n309578 , n309396 , n309401 );
or ( n309579 , n19149 , n309578 );
buf ( n309580 , n309579 );
buf ( n309581 , n309580 );
buf ( n309582 , n18558 );
buf ( n309583 , n309437 );
or ( n19156 , n309582 , n309583 );
buf ( n309585 , n308992 );
buf ( n309586 , n298423 );
buf ( n309587 , n769 );
and ( n309588 , n309586 , n309587 );
buf ( n19161 , n299244 );
buf ( n309590 , n800 );
and ( n309591 , n19161 , n309590 );
nor ( n19164 , n309588 , n309591 );
buf ( n309593 , n19164 );
buf ( n309594 , n309593 );
or ( n19167 , n309585 , n309594 );
nand ( n309596 , n19156 , n19167 );
buf ( n309597 , n309596 );
buf ( n309598 , n309597 );
buf ( n309599 , n771 );
buf ( n309600 , n800 );
and ( n19173 , n309599 , n309600 );
buf ( n309602 , n19173 );
buf ( n309603 , n309602 );
xor ( n309604 , n309598 , n309603 );
buf ( n309605 , n309342 );
buf ( n309606 , n309414 );
or ( n309607 , n309605 , n309606 );
buf ( n309608 , n309348 );
buf ( n309609 , n309352 );
or ( n309610 , n309608 , n309609 );
nand ( n19183 , n309607 , n309610 );
buf ( n19184 , n19183 );
buf ( n309613 , n19184 );
not ( n19186 , n309613 );
buf ( n309615 , n19186 );
buf ( n309616 , n309615 );
xor ( n19189 , n309604 , n309616 );
buf ( n309618 , n19189 );
buf ( n309619 , n309618 );
xor ( n19192 , n309581 , n309619 );
not ( n309621 , n309313 );
not ( n19194 , n309441 );
or ( n19195 , n309621 , n19194 );
not ( n309624 , n18886 );
not ( n309625 , n309442 );
or ( n19198 , n309624 , n309625 );
not ( n309627 , n18997 );
nand ( n309628 , n19198 , n309627 );
nand ( n19201 , n19195 , n309628 );
buf ( n309630 , n19201 );
xor ( n19203 , n19192 , n309630 );
buf ( n309632 , n19203 );
buf ( n19205 , n309632 );
xor ( n309634 , n309421 , n309447 );
and ( n19207 , n309634 , n309452 );
and ( n309636 , n309421 , n309447 );
or ( n19209 , n19207 , n309636 );
buf ( n309638 , n19209 );
xor ( n309639 , n19205 , n309638 );
buf ( n309640 , n309639 );
nor ( n19213 , n309575 , n309640 );
and ( n309642 , n19205 , n309638 );
buf ( n309643 , n309642 );
buf ( n309644 , n19184 );
xor ( n19217 , n309598 , n309603 );
and ( n309646 , n19217 , n309616 );
and ( n309647 , n309598 , n309603 );
or ( n19220 , n309646 , n309647 );
buf ( n309649 , n19220 );
buf ( n309650 , n309649 );
xor ( n19223 , n309644 , n309650 );
buf ( n309652 , n296508 );
buf ( n309653 , n296749 );
or ( n309654 , n309652 , n309653 );
buf ( n309655 , n802 );
nand ( n309656 , n309654 , n309655 );
buf ( n309657 , n309656 );
buf ( n309658 , n309657 );
buf ( n309659 , n770 );
buf ( n309660 , n800 );
and ( n19233 , n309659 , n309660 );
buf ( n309662 , n19233 );
buf ( n309663 , n309662 );
xor ( n309664 , n309658 , n309663 );
buf ( n309665 , n18558 );
buf ( n309666 , n309593 );
or ( n19239 , n309665 , n309666 );
buf ( n309668 , n308992 );
buf ( n309669 , n768 );
buf ( n309670 , n298423 );
and ( n309671 , n309669 , n309670 );
not ( n309672 , n309669 );
buf ( n309673 , n800 );
and ( n309674 , n309672 , n309673 );
nor ( n19247 , n309671 , n309674 );
buf ( n309676 , n19247 );
buf ( n309677 , n309676 );
or ( n19250 , n309668 , n309677 );
nand ( n309679 , n19239 , n19250 );
buf ( n309680 , n309679 );
buf ( n309681 , n309680 );
xor ( n19254 , n309664 , n309681 );
buf ( n309683 , n19254 );
buf ( n309684 , n309683 );
xor ( n309685 , n19223 , n309684 );
buf ( n309686 , n309685 );
buf ( n309687 , n309686 );
xor ( n309688 , n309581 , n309619 );
and ( n19261 , n309688 , n309630 );
and ( n19262 , n309581 , n309619 );
or ( n309691 , n19261 , n19262 );
buf ( n309692 , n309691 );
buf ( n309693 , n309692 );
xor ( n309694 , n309687 , n309693 );
buf ( n309695 , n309694 );
nor ( n309696 , n309643 , n309695 );
nor ( n19269 , n19213 , n309696 );
and ( n309698 , n309573 , n19269 );
nand ( n309699 , n309575 , n309640 );
or ( n19272 , n309699 , n309696 );
nand ( n309701 , n309643 , n309695 );
nand ( n309702 , n19272 , n309701 );
nor ( n19275 , n309698 , n309702 );
or ( n309704 , n19144 , n19213 );
nand ( n19277 , n309704 , n309699 );
buf ( n309706 , n308692 );
buf ( n309707 , n308840 );
and ( n19280 , n309706 , n309707 );
buf ( n309709 , n19280 );
xor ( n19282 , n309540 , n309546 );
xor ( n309711 , n19282 , n309551 );
buf ( n309712 , n309711 );
buf ( n309713 , n309712 );
xor ( n19286 , n308801 , n308831 );
and ( n309715 , n19286 , n308838 );
and ( n19288 , n308801 , n308831 );
or ( n19289 , n309715 , n19288 );
buf ( n309718 , n19289 );
buf ( n309719 , n309718 );
xor ( n19292 , n309713 , n309719 );
buf ( n309721 , n19292 );
or ( n19294 , n309709 , n309721 );
and ( n309723 , n18416 , n19294 );
not ( n309724 , n309723 );
not ( n19297 , n18435 );
or ( n309726 , n309724 , n19297 );
and ( n309727 , n18445 , n19294 );
and ( n309728 , n309709 , n309721 );
nor ( n19301 , n309727 , n309728 );
nand ( n309730 , n309726 , n19301 );
not ( n19303 , n309730 );
and ( n19304 , n309687 , n309693 );
buf ( n309733 , n19304 );
buf ( n19306 , n769 );
buf ( n19307 , n800 );
nand ( n19308 , n19306 , n19307 );
buf ( n19309 , n19308 );
buf ( n309738 , n19309 );
buf ( n309739 , n18558 );
buf ( n309740 , n309676 );
or ( n309741 , n309739 , n309740 );
buf ( n309742 , n308992 );
buf ( n309743 , n298423 );
or ( n309744 , n309742 , n309743 );
nand ( n19317 , n309741 , n309744 );
buf ( n309746 , n19317 );
buf ( n19319 , n309746 );
xor ( n19320 , n309738 , n19319 );
xor ( n309749 , n309658 , n309663 );
and ( n19322 , n309749 , n309681 );
and ( n19323 , n309658 , n309663 );
or ( n19324 , n19322 , n19323 );
buf ( n309753 , n19324 );
buf ( n309754 , n309753 );
xor ( n19327 , n19320 , n309754 );
buf ( n309756 , n19327 );
buf ( n309757 , n309756 );
xor ( n19330 , n309644 , n309650 );
and ( n309759 , n19330 , n309684 );
and ( n19332 , n309644 , n309650 );
or ( n19333 , n309759 , n19332 );
buf ( n309762 , n19333 );
buf ( n309763 , n309762 );
xor ( n309764 , n309757 , n309763 );
buf ( n309765 , n309764 );
or ( n309766 , n309733 , n309765 );
and ( n309767 , n19269 , n309766 );
not ( n19340 , n309767 );
not ( n309769 , n309573 );
or ( n309770 , n19340 , n309769 );
and ( n19343 , n309702 , n309766 );
and ( n19344 , n309733 , n309765 );
nor ( n19345 , n19343 , n19344 );
nand ( n309774 , n309770 , n19345 );
nand ( n309775 , n307526 , n307618 );
not ( n19348 , n309775 );
and ( n309777 , n17088 , n19348 );
not ( n19350 , n307618 );
not ( n309779 , n307540 );
or ( n19352 , n19350 , n309779 );
nand ( n19353 , n19352 , n307619 );
nor ( n309782 , n309777 , n19353 );
not ( n309783 , n307453 );
nor ( n309784 , n309783 , n307424 );
not ( n19357 , n307453 );
not ( n309786 , n307458 );
or ( n309787 , n19357 , n309786 );
nand ( n19360 , n309787 , n17032 );
nor ( n309789 , n309784 , n19360 );
not ( n309790 , n307999 );
nand ( n19363 , n309790 , n307710 );
not ( n309792 , n19363 );
xor ( n309793 , n19108 , n309555 );
and ( n309794 , n309713 , n309719 );
buf ( n309795 , n309794 );
or ( n19368 , n309793 , n309795 );
and ( n309797 , n19368 , n19294 );
nand ( n19370 , n18416 , n309797 );
nor ( n309799 , n308466 , n19370 );
or ( n309800 , n19128 , n309562 );
not ( n19373 , n19106 );
and ( n309802 , n309800 , n19373 );
and ( n19375 , n309799 , n309802 );
and ( n309804 , n309792 , n19375 );
not ( n19377 , n309792 );
nor ( n19378 , n19377 , n307916 );
buf ( n309807 , n309799 );
nand ( n309808 , n309802 , n309463 );
not ( n309809 , n309808 );
and ( n19382 , n309809 , n309767 );
nand ( n309811 , n309807 , n19382 );
nor ( n309812 , n19377 , n309811 );
not ( n19385 , n307458 );
nand ( n309814 , n19385 , n307424 );
not ( n309815 , n309792 );
not ( n19388 , n308466 );
nand ( n309817 , n19388 , n309723 );
nor ( n309818 , n309815 , n309817 );
nand ( n19391 , n19388 , n18416 );
nor ( n19392 , n19377 , n19391 );
nor ( n19393 , n309815 , n18039 );
buf ( n309822 , n19363 );
not ( n309823 , n18959 );
and ( n19396 , n309802 , n309823 );
nand ( n309825 , n309807 , n19396 );
nor ( n309826 , n309822 , n309825 );
not ( n19399 , n309799 );
nor ( n309828 , n309815 , n19399 );
and ( n309829 , n309809 , n19269 );
nand ( n309830 , n309807 , n309829 );
nor ( n309831 , n309822 , n309830 );
not ( n19404 , n19399 );
nand ( n309833 , n19404 , n309809 );
nor ( n309834 , n19377 , n309833 );
not ( n309835 , n307977 );
nand ( n19408 , n308649 , n309835 );
not ( n309837 , n306856 );
not ( n19410 , n17281 );
nand ( n19411 , n309837 , n19410 );
nor ( n309840 , n19408 , n19411 );
not ( n19413 , n308649 );
nor ( n309842 , n19411 , n19413 );
not ( n19415 , n16826 );
not ( n309844 , n16813 );
or ( n309845 , n19415 , n309844 );
nand ( n19418 , n309845 , n16816 );
not ( n309847 , n19418 );
not ( n309848 , n306850 );
not ( n19421 , n309848 );
buf ( n309850 , n307513 );
not ( n19423 , n309850 );
or ( n309852 , n19421 , n19423 );
not ( n19425 , n17077 );
nand ( n19426 , n309852 , n19425 );
not ( n309855 , n19426 );
not ( n19428 , n18435 );
not ( n309857 , n309823 );
not ( n19430 , n19138 );
or ( n309859 , n309857 , n19430 );
nand ( n309860 , n309859 , n309568 );
not ( n19433 , n307943 );
buf ( n309862 , n17587 );
not ( n309863 , n309862 );
or ( n19436 , n19433 , n309863 );
not ( n309865 , n308019 );
nand ( n309866 , n19436 , n309865 );
not ( n309867 , n306975 );
not ( n19440 , n306989 );
or ( n309869 , n309867 , n19440 );
nand ( n19442 , n309869 , n16565 );
nor ( n19443 , n16429 , n309775 );
buf ( n309872 , n306834 );
and ( n309873 , n309872 , n309848 );
and ( n309874 , n307253 , n16826 );
and ( n19447 , n308465 , n17841 );
not ( n309876 , n309850 );
not ( n309877 , n307103 );
and ( n19450 , n309728 , n19368 );
and ( n309879 , n309795 , n309793 );
nor ( n309880 , n19450 , n309879 );
nand ( n19453 , n307893 , n17052 );
not ( n309882 , n19453 );
nand ( n309883 , n17346 , n306895 );
not ( n309884 , n309883 );
not ( n19457 , n19213 );
nand ( n309886 , n19457 , n309699 );
not ( n19459 , n309886 );
nand ( n19460 , n16826 , n16816 );
not ( n19461 , n309696 );
nand ( n309890 , n19461 , n309701 );
not ( n309891 , n309462 );
nand ( n309892 , n309891 , n309570 );
nand ( n19465 , n307453 , n17032 );
not ( n309894 , n17294 );
nand ( n309895 , n309894 , n17296 );
nand ( n19468 , n309848 , n19425 );
not ( n309897 , n19468 );
buf ( n309898 , n307510 );
nand ( n19471 , n306801 , n309898 );
nand ( n309900 , n307943 , n309865 );
nand ( n309901 , n18440 , n308871 );
nand ( n19474 , n307800 , n307491 );
nand ( n309903 , n17559 , n308662 );
nand ( n19476 , n309823 , n309568 );
not ( n309905 , n19106 );
nand ( n19478 , n309905 , n309565 );
not ( n309907 , n307252 );
not ( n309908 , n307969 );
and ( n19481 , n17445 , n307738 );
nor ( n19482 , n19481 , n19442 );
not ( n309911 , n309809 );
not ( n309912 , n19370 );
not ( n19485 , n309912 );
not ( n309914 , n18434 );
or ( n309915 , n19485 , n309914 );
not ( n19488 , n309797 );
not ( n309917 , n308872 );
or ( n309918 , n19488 , n309917 );
nand ( n19491 , n309918 , n309880 );
not ( n309920 , n19491 );
nand ( n309921 , n309915 , n309920 );
not ( n19494 , n309921 );
not ( n309923 , n19494 );
not ( n309924 , n309923 );
or ( n19497 , n309911 , n309924 );
nand ( n309926 , n19497 , n19144 );
not ( n19499 , n309926 );
buf ( n309928 , n307500 );
nand ( n19501 , n309834 , n309928 );
not ( n19502 , n309833 );
nand ( n309931 , n19502 , n18214 );
nand ( n19504 , n19499 , n19501 , n309931 );
not ( n309933 , n309825 );
nand ( n19506 , n309933 , n18214 );
not ( n309935 , n309811 );
nand ( n309936 , n309935 , n18214 );
not ( n19509 , n17283 );
nor ( n309938 , n19509 , n18224 );
buf ( n309939 , n17506 );
not ( n309940 , n309939 );
and ( n19513 , n307943 , n309940 );
not ( n309942 , n19513 );
nor ( n19515 , n309942 , n19411 );
not ( n19516 , n17613 );
nand ( n309945 , n19516 , n17568 );
not ( n19518 , n17035 );
nand ( n309947 , n19518 , n307447 );
not ( n19520 , n17595 );
nand ( n309949 , n19520 , n308018 );
buf ( n309950 , n831 );
buf ( n309951 , n307166 );
buf ( n309952 , n883 );
buf ( n19525 , n307156 );
xor ( n19526 , n309952 , n19525 );
buf ( n309955 , n307161 );
and ( n19528 , n19526 , n309955 );
and ( n309957 , n309952 , n19525 );
or ( n19530 , n19528 , n309957 );
buf ( n309959 , n19530 );
buf ( n19532 , n309959 );
buf ( n309961 , n5980 );
nand ( n309962 , n19532 , n309961 );
buf ( n309963 , n309962 );
buf ( n309964 , n309963 );
not ( n309965 , n309950 );
not ( n19538 , n309951 );
or ( n309967 , n309965 , n19538 );
nand ( n309968 , n309967 , n309964 );
buf ( n309969 , n309968 );
buf ( n309970 , n831 );
buf ( n309971 , n308452 );
buf ( n309972 , n831 );
not ( n309973 , n309972 );
buf ( n19546 , n308260 );
buf ( n309975 , n308265 );
and ( n19548 , n19546 , n309975 );
buf ( n309977 , n19548 );
buf ( n309978 , n309977 );
nand ( n19551 , n309973 , n309978 );
buf ( n309980 , n19551 );
buf ( n309981 , n309980 );
not ( n309982 , n309970 );
not ( n19555 , n309971 );
or ( n19556 , n309982 , n19555 );
nand ( n19557 , n19556 , n309981 );
buf ( n309986 , n19557 );
buf ( n309987 , n768 );
not ( n19560 , n309987 );
buf ( n309989 , n298423 );
nor ( n19562 , n19560 , n309989 );
buf ( n309991 , n19562 );
buf ( n309992 , n309991 );
buf ( n309993 , n19309 );
not ( n309994 , n309993 );
buf ( n309995 , n309994 );
buf ( n309996 , n309995 );
xor ( n19569 , n309992 , n309996 );
buf ( n19570 , n308992 );
not ( n19571 , n19570 );
buf ( n310000 , n18558 );
not ( n19573 , n310000 );
or ( n19574 , n19571 , n19573 );
buf ( n310003 , n800 );
nand ( n19576 , n19574 , n310003 );
buf ( n310005 , n19576 );
buf ( n310006 , n310005 );
xor ( n19579 , n19569 , n310006 );
buf ( n310008 , n19579 );
buf ( n19581 , n310008 );
xor ( n19582 , n309738 , n19319 );
and ( n310011 , n19582 , n309754 );
and ( n310012 , n309738 , n19319 );
or ( n19585 , n310011 , n310012 );
buf ( n310014 , n19585 );
buf ( n310015 , n310014 );
and ( n19588 , n19581 , n310015 );
buf ( n310017 , n19588 );
buf ( n19590 , n310017 );
buf ( n19591 , n310008 );
buf ( n19592 , n310014 );
and ( n19593 , n19591 , n19592 );
buf ( n310022 , n19593 );
buf ( n310023 , n310022 );
buf ( n310024 , n831 );
and ( n310025 , n310024 , n310023 );
not ( n19598 , n310024 );
and ( n19599 , n19598 , n19590 );
or ( n310028 , n310025 , n19599 );
buf ( n310029 , n310028 );
buf ( n310030 , n304008 );
buf ( n310031 , n304004 );
and ( n310032 , n310030 , n310031 );
buf ( n310033 , n310032 );
buf ( n310034 , n310033 );
buf ( n19607 , n296412 );
nand ( n19608 , n310034 , n19607 );
buf ( n310037 , n19608 );
and ( n310038 , n307926 , n17501 );
buf ( n310039 , n310038 );
buf ( n310040 , n296412 );
nand ( n19613 , n310039 , n310040 );
buf ( n19614 , n19613 );
buf ( n310043 , n831 );
buf ( n310044 , n877 );
buf ( n310045 , n303509 );
xor ( n310046 , n310044 , n310045 );
buf ( n310047 , n303505 );
and ( n19620 , n310046 , n310047 );
and ( n310049 , n310044 , n310045 );
or ( n310050 , n19620 , n310049 );
buf ( n310051 , n310050 );
buf ( n310052 , n310051 );
not ( n310053 , n310043 );
nand ( n19626 , n310053 , n310052 );
buf ( n310055 , n19626 );
buf ( n310056 , n831 );
buf ( n310057 , n869 );
buf ( n310058 , n306875 );
xor ( n19631 , n310057 , n310058 );
buf ( n310060 , n306880 );
and ( n310061 , n19631 , n310060 );
and ( n19634 , n310057 , n310058 );
or ( n19635 , n310061 , n19634 );
buf ( n310064 , n19635 );
buf ( n310065 , n310064 );
not ( n19638 , n310056 );
nand ( n310067 , n19638 , n310065 );
buf ( n310068 , n310067 );
xor ( n19641 , n303192 , n303193 );
xor ( n310070 , n19641 , n303195 );
buf ( n310071 , n310070 );
buf ( n310072 , n880 );
buf ( n310073 , n307021 );
buf ( n310074 , n307026 );
xor ( n19647 , n310072 , n310073 );
xor ( n310076 , n19647 , n310074 );
buf ( n310077 , n310076 );
xor ( n19650 , n310072 , n310073 );
and ( n310079 , n19650 , n310074 );
and ( n310080 , n310072 , n310073 );
or ( n19653 , n310079 , n310080 );
buf ( n310082 , n19653 );
xor ( n310083 , n292332 , n292333 );
xor ( n19656 , n310083 , n292335 );
buf ( n310085 , n19656 );
xor ( n19658 , n3158 , n293587 );
xor ( n19659 , n19658 , n293589 );
buf ( n310088 , n19659 );
buf ( n310089 , n882 );
buf ( n310090 , n303550 );
buf ( n310091 , n303555 );
xor ( n310092 , n310089 , n310090 );
xor ( n19665 , n310092 , n310091 );
buf ( n310094 , n19665 );
xor ( n310095 , n310089 , n310090 );
and ( n19668 , n310095 , n310091 );
and ( n19669 , n310089 , n310090 );
or ( n310098 , n19668 , n19669 );
buf ( n310099 , n310098 );
xor ( n310100 , n309952 , n19525 );
xor ( n310101 , n310100 , n309955 );
buf ( n310102 , n310101 );
buf ( n19675 , n884 );
buf ( n310104 , n307177 );
buf ( n310105 , n307182 );
xor ( n310106 , n19675 , n310104 );
xor ( n19679 , n310106 , n310105 );
buf ( n310108 , n19679 );
xor ( n310109 , n19675 , n310104 );
and ( n310110 , n310109 , n310105 );
and ( n19683 , n19675 , n310104 );
or ( n310112 , n310110 , n19683 );
buf ( n310113 , n310112 );
xor ( n19686 , n298368 , n298369 );
xor ( n310115 , n19686 , n298371 );
buf ( n310116 , n310115 );
xor ( n19689 , n295139 , n295140 );
xor ( n310118 , n19689 , n295142 );
buf ( n310119 , n310118 );
buf ( n310120 , n887 );
buf ( n310121 , n303263 );
buf ( n310122 , n303274 );
xor ( n19695 , n310120 , n310121 );
xor ( n310124 , n19695 , n310122 );
buf ( n310125 , n310124 );
xor ( n19698 , n310120 , n310121 );
and ( n310127 , n19698 , n310122 );
and ( n310128 , n310120 , n310121 );
or ( n19701 , n310127 , n310128 );
buf ( n310130 , n19701 );
xor ( n310131 , n296353 , n296354 );
xor ( n19704 , n310131 , n296356 );
buf ( n310133 , n19704 );
buf ( n19706 , n876 );
buf ( n310135 , n303468 );
buf ( n310136 , n303473 );
xor ( n310137 , n19706 , n310135 );
xor ( n19710 , n310137 , n310136 );
buf ( n310139 , n19710 );
xor ( n310140 , n19706 , n310135 );
and ( n19713 , n310140 , n310136 );
and ( n310142 , n19706 , n310135 );
or ( n310143 , n19713 , n310142 );
buf ( n310144 , n310143 );
buf ( n310145 , n888 );
buf ( n310146 , n307228 );
buf ( n310147 , n16804 );
xor ( n19720 , n310145 , n310146 );
xor ( n19721 , n19720 , n310147 );
buf ( n19722 , n19721 );
xor ( n19723 , n310145 , n310146 );
and ( n19724 , n19723 , n310147 );
and ( n19725 , n310145 , n310146 );
or ( n19726 , n19724 , n19725 );
buf ( n310155 , n19726 );
xor ( n310156 , n310044 , n310045 );
xor ( n19729 , n310156 , n310047 );
buf ( n310158 , n19729 );
buf ( n310159 , n890 );
buf ( n310160 , n303330 );
buf ( n310161 , n303401 );
xor ( n310162 , n310159 , n310160 );
xor ( n19735 , n310162 , n310161 );
buf ( n310164 , n19735 );
xor ( n19737 , n310159 , n310160 );
and ( n310166 , n19737 , n310161 );
and ( n19739 , n310159 , n310160 );
or ( n19740 , n310166 , n19739 );
buf ( n310169 , n19740 );
buf ( n19742 , n871 );
buf ( n19743 , n303414 );
buf ( n310172 , n12990 );
xor ( n310173 , n19742 , n19743 );
xor ( n19746 , n310173 , n310172 );
buf ( n310175 , n19746 );
xor ( n310176 , n19742 , n19743 );
and ( n310177 , n310176 , n310172 );
and ( n19750 , n19742 , n19743 );
or ( n310179 , n310177 , n19750 );
buf ( n310180 , n310179 );
buf ( n310181 , n878 );
buf ( n310182 , n307005 );
buf ( n310183 , n307010 );
xor ( n19756 , n310181 , n310182 );
xor ( n19757 , n19756 , n310183 );
buf ( n310186 , n19757 );
xor ( n19759 , n310181 , n310182 );
and ( n310188 , n19759 , n310183 );
and ( n19761 , n310181 , n310182 );
or ( n19762 , n310188 , n19761 );
buf ( n310191 , n19762 );
buf ( n310192 , n892 );
buf ( n310193 , n307402 );
buf ( n310194 , n307405 );
xor ( n19767 , n310192 , n310193 );
xor ( n19768 , n19767 , n310194 );
buf ( n310197 , n19768 );
xor ( n19770 , n310192 , n310193 );
and ( n19771 , n19770 , n310194 );
and ( n310200 , n310192 , n310193 );
or ( n19773 , n19771 , n310200 );
buf ( n310202 , n19773 );
buf ( n310203 , n893 );
buf ( n310204 , n307314 );
buf ( n19777 , n307332 );
xor ( n19778 , n310203 , n310204 );
xor ( n310207 , n19778 , n19777 );
buf ( n310208 , n310207 );
xor ( n19781 , n310203 , n310204 );
and ( n19782 , n19781 , n19777 );
and ( n19783 , n310203 , n310204 );
or ( n310212 , n19782 , n19783 );
buf ( n310213 , n310212 );
xor ( n310214 , n301133 , n301134 );
xor ( n310215 , n310214 , n301136 );
buf ( n310216 , n310215 );
buf ( n310217 , n894 );
buf ( n310218 , n307344 );
buf ( n310219 , n307361 );
xor ( n19792 , n310217 , n310218 );
xor ( n310221 , n19792 , n310219 );
buf ( n310222 , n310221 );
xor ( n19795 , n310217 , n310218 );
and ( n19796 , n19795 , n310219 );
and ( n310225 , n310217 , n310218 );
or ( n310226 , n19796 , n310225 );
buf ( n310227 , n310226 );
buf ( n310228 , n309686 );
buf ( n310229 , n309692 );
xor ( n19802 , n310228 , n310229 );
buf ( n310231 , n19802 );
and ( n19804 , n310228 , n310229 );
buf ( n310233 , n19804 );
buf ( n310234 , n309756 );
buf ( n310235 , n309762 );
xor ( n310236 , n310234 , n310235 );
buf ( n310237 , n310236 );
and ( n19810 , n310234 , n310235 );
buf ( n310239 , n19810 );
xor ( n310240 , n19581 , n310015 );
buf ( n310241 , n310240 );
buf ( n310242 , n18774 );
buf ( n19815 , n309302 );
xor ( n19816 , n310242 , n19815 );
buf ( n310245 , n19816 );
and ( n310246 , n310242 , n19815 );
buf ( n310247 , n310246 );
buf ( n310248 , n309712 );
buf ( n310249 , n309718 );
xor ( n19822 , n310248 , n310249 );
buf ( n310251 , n19822 );
and ( n19824 , n310248 , n310249 );
buf ( n310253 , n19824 );
buf ( n19826 , n308840 );
buf ( n19827 , n308692 );
xor ( n19828 , n19826 , n19827 );
buf ( n310257 , n19828 );
and ( n310258 , n19826 , n19827 );
buf ( n310259 , n310258 );
xor ( n310260 , n19546 , n309975 );
buf ( n310261 , n310260 );
xor ( n19834 , n302382 , n302383 );
buf ( n310263 , n19834 );
xor ( n19836 , n310030 , n310031 );
buf ( n310265 , n19836 );
buf ( n19838 , n307985 );
buf ( n310267 , n307980 );
xor ( n19840 , n19838 , n310267 );
buf ( n310269 , n19840 );
and ( n19842 , n19838 , n310267 );
buf ( n310271 , n19842 );
xor ( n310272 , n303121 , n303122 );
buf ( n310273 , n310272 );
buf ( n310274 , n307630 );
buf ( n310275 , n307661 );
xor ( n19848 , n310274 , n310275 );
buf ( n310277 , n19848 );
and ( n19850 , n310274 , n310275 );
buf ( n310279 , n19850 );
buf ( n19852 , n16946 );
buf ( n19853 , n895 );
xor ( n19854 , n19852 , n19853 );
buf ( n310283 , n19854 );
buf ( n310284 , n309377 );
buf ( n310285 , n309383 );
xor ( n19860 , n310284 , n310285 );
buf ( n310287 , n19860 );
and ( n19862 , n310284 , n310285 );
buf ( n310289 , n19862 );
buf ( n310290 , n308447 );
buf ( n310291 , n308441 );
xor ( n310292 , n310290 , n310291 );
buf ( n310293 , n310292 );
and ( n19868 , n310290 , n310291 );
buf ( n310295 , n19868 );
xor ( n310296 , n7101 , n297869 );
buf ( n310297 , n310296 );
xor ( n310298 , n302972 , n302973 );
buf ( n310299 , n310298 );
buf ( n310300 , n303951 );
buf ( n310301 , n303955 );
xor ( n310302 , n310300 , n310301 );
buf ( n310303 , n310302 );
and ( n310304 , n310300 , n310301 );
buf ( n310305 , n310304 );
buf ( n310306 , n309453 );
buf ( n310307 , n309458 );
xor ( n310308 , n310306 , n310307 );
buf ( n310309 , n310308 );
and ( n310310 , n310306 , n310307 );
buf ( n310311 , n310310 );
buf ( n310312 , n309632 );
buf ( n310313 , n19209 );
xor ( n310314 , n310312 , n310313 );
buf ( n310315 , n310314 );
and ( n19890 , n310312 , n310313 );
buf ( n310317 , n19890 );
xor ( n310318 , n302170 , n302171 );
buf ( n310319 , n310318 );
and ( n310320 , n309757 , n309763 );
buf ( n310321 , n310320 );
xor ( n19896 , n309992 , n309996 );
and ( n310323 , n19896 , n310006 );
and ( n310324 , n309992 , n309996 );
or ( n19899 , n310323 , n310324 );
buf ( n310326 , n19899 );
xor ( n19901 , n870 , n847 );
buf ( n310328 , n19901 );
not ( n19903 , n310328 );
buf ( n310330 , n14323 );
not ( n19905 , n310330 );
or ( n19906 , n19903 , n19905 );
buf ( n310333 , n304763 );
xor ( n19908 , n870 , n846 );
buf ( n310335 , n19908 );
nand ( n19910 , n310333 , n310335 );
buf ( n310337 , n19910 );
buf ( n310338 , n310337 );
nand ( n19913 , n19906 , n310338 );
buf ( n19914 , n19913 );
buf ( n310341 , n19914 );
xor ( n19916 , n872 , n845 );
buf ( n310343 , n19916 );
not ( n310344 , n310343 );
buf ( n310345 , n304851 );
not ( n310346 , n310345 );
or ( n19921 , n310344 , n310346 );
buf ( n310348 , n304845 );
buf ( n310349 , n844 );
buf ( n310350 , n872 );
xor ( n310351 , n310349 , n310350 );
buf ( n310352 , n310351 );
buf ( n310353 , n310352 );
nand ( n310354 , n310348 , n310353 );
buf ( n310355 , n310354 );
buf ( n310356 , n310355 );
nand ( n310357 , n19921 , n310356 );
buf ( n310358 , n310357 );
buf ( n310359 , n310358 );
xor ( n310360 , n310341 , n310359 );
buf ( n310361 , n304941 );
buf ( n310362 , n839 );
buf ( n310363 , n878 );
xnor ( n310364 , n310362 , n310363 );
buf ( n310365 , n310364 );
buf ( n310366 , n310365 );
or ( n310367 , n310361 , n310366 );
buf ( n310368 , n14523 );
buf ( n310369 , n878 );
not ( n19944 , n310369 );
buf ( n310371 , n19944 );
buf ( n310372 , n310371 );
buf ( n310373 , n838 );
and ( n19948 , n310372 , n310373 );
buf ( n310375 , n838 );
not ( n310376 , n310375 );
buf ( n310377 , n310376 );
buf ( n310378 , n310377 );
buf ( n310379 , n878 );
and ( n19954 , n310378 , n310379 );
nor ( n19955 , n19948 , n19954 );
buf ( n310382 , n19955 );
buf ( n310383 , n310382 );
or ( n310384 , n310368 , n310383 );
nand ( n19959 , n310367 , n310384 );
buf ( n310386 , n19959 );
buf ( n310387 , n310386 );
xor ( n19962 , n310360 , n310387 );
buf ( n310389 , n19962 );
buf ( n310390 , n310389 );
not ( n310391 , n310390 );
buf ( n310392 , n884 );
buf ( n310393 , n833 );
xor ( n310394 , n310392 , n310393 );
buf ( n310395 , n310394 );
buf ( n310396 , n310395 );
not ( n310397 , n310396 );
buf ( n310398 , n304802 );
buf ( n310399 , n304807 );
nor ( n310400 , n310398 , n310399 );
buf ( n310401 , n310400 );
buf ( n310402 , n310401 );
not ( n310403 , n310402 );
or ( n310404 , n310397 , n310403 );
buf ( n310405 , n304807 );
buf ( n310406 , n884 );
buf ( n19981 , n832 );
xor ( n19982 , n310406 , n19981 );
buf ( n310409 , n19982 );
buf ( n19984 , n310409 );
nand ( n19985 , n310405 , n19984 );
buf ( n19986 , n19985 );
buf ( n310413 , n19986 );
nand ( n19988 , n310404 , n310413 );
buf ( n310415 , n19988 );
buf ( n310416 , n310415 );
buf ( n310417 , n305363 );
not ( n310418 , n310417 );
buf ( n310419 , n305356 );
not ( n19994 , n310419 );
or ( n310421 , n310418 , n19994 );
buf ( n19996 , n886 );
nand ( n19997 , n310421 , n19996 );
buf ( n19998 , n19997 );
buf ( n310425 , n19998 );
xor ( n20000 , n310416 , n310425 );
buf ( n310427 , n304987 );
buf ( n310428 , n880 );
not ( n310429 , n310428 );
buf ( n310430 , n837 );
nor ( n20005 , n310429 , n310430 );
buf ( n310432 , n20005 );
buf ( n310433 , n310432 );
buf ( n310434 , n837 );
not ( n310435 , n310434 );
buf ( n310436 , n880 );
nor ( n20011 , n310435 , n310436 );
buf ( n310438 , n20011 );
buf ( n310439 , n310438 );
nor ( n310440 , n310433 , n310439 );
buf ( n310441 , n310440 );
buf ( n310442 , n310441 );
or ( n20017 , n310427 , n310442 );
buf ( n310444 , n836 );
buf ( n310445 , n880 );
xor ( n310446 , n310444 , n310445 );
buf ( n310447 , n310446 );
buf ( n310448 , n310447 );
not ( n20023 , n310448 );
buf ( n310450 , n20023 );
buf ( n310451 , n310450 );
buf ( n310452 , n304976 );
or ( n20027 , n310451 , n310452 );
nand ( n20028 , n20017 , n20027 );
buf ( n310455 , n20028 );
buf ( n310456 , n310455 );
xor ( n20031 , n20000 , n310456 );
buf ( n310458 , n20031 );
buf ( n310459 , n310458 );
buf ( n310460 , n851 );
buf ( n310461 , n866 );
xor ( n20036 , n310460 , n310461 );
buf ( n310463 , n20036 );
buf ( n310464 , n310463 );
not ( n20039 , n310464 );
buf ( n310466 , n867 );
buf ( n310467 , n868 );
xor ( n20042 , n310466 , n310467 );
buf ( n310469 , n20042 );
buf ( n310470 , n310469 );
not ( n310471 , n310470 );
buf ( n310472 , n310471 );
buf ( n310473 , n310472 );
xor ( n20048 , n866 , n867 );
buf ( n310475 , n20048 );
and ( n20050 , n310473 , n310475 );
buf ( n310477 , n20050 );
buf ( n310478 , n310477 );
not ( n20053 , n310478 );
or ( n310480 , n20039 , n20053 );
buf ( n310481 , n310469 );
buf ( n310482 , n310481 );
buf ( n310483 , n310482 );
buf ( n310484 , n310483 );
buf ( n310485 , n850 );
buf ( n310486 , n866 );
xor ( n310487 , n310485 , n310486 );
buf ( n310488 , n310487 );
buf ( n310489 , n310488 );
nand ( n20064 , n310484 , n310489 );
buf ( n20065 , n20064 );
buf ( n310492 , n20065 );
nand ( n310493 , n310480 , n310492 );
buf ( n310494 , n310493 );
buf ( n310495 , n310494 );
xor ( n310496 , n882 , n835 );
buf ( n310497 , n310496 );
not ( n20072 , n310497 );
buf ( n310499 , n304584 );
not ( n310500 , n310499 );
or ( n20075 , n20072 , n310500 );
buf ( n310502 , n304596 );
buf ( n310503 , n882 );
buf ( n310504 , n834 );
xor ( n310505 , n310503 , n310504 );
buf ( n310506 , n310505 );
buf ( n310507 , n310506 );
nand ( n310508 , n310502 , n310507 );
buf ( n310509 , n310508 );
buf ( n310510 , n310509 );
nand ( n310511 , n20075 , n310510 );
buf ( n310512 , n310511 );
buf ( n310513 , n310512 );
xor ( n310514 , n310495 , n310513 );
buf ( n310515 , n849 );
buf ( n310516 , n868 );
and ( n20091 , n310515 , n310516 );
not ( n310518 , n310515 );
buf ( n310519 , n868 );
not ( n20094 , n310519 );
buf ( n310521 , n20094 );
buf ( n310522 , n310521 );
and ( n310523 , n310518 , n310522 );
nor ( n310524 , n20091 , n310523 );
buf ( n310525 , n310524 );
buf ( n310526 , n310525 );
not ( n310527 , n310526 );
buf ( n310528 , n305213 );
not ( n20103 , n310528 );
or ( n310530 , n310527 , n20103 );
buf ( n310531 , n305202 );
buf ( n310532 , n848 );
buf ( n310533 , n868 );
xor ( n310534 , n310532 , n310533 );
buf ( n310535 , n310534 );
buf ( n310536 , n310535 );
nand ( n310537 , n310531 , n310536 );
buf ( n310538 , n310537 );
buf ( n310539 , n310538 );
nand ( n310540 , n310530 , n310539 );
buf ( n310541 , n310540 );
buf ( n310542 , n310541 );
xor ( n310543 , n310514 , n310542 );
buf ( n310544 , n310543 );
buf ( n310545 , n310544 );
xnor ( n310546 , n310459 , n310545 );
buf ( n310547 , n310546 );
buf ( n310548 , n310547 );
not ( n310549 , n310548 );
or ( n310550 , n310391 , n310549 );
buf ( n310551 , n310547 );
buf ( n310552 , n310389 );
or ( n20127 , n310551 , n310552 );
nand ( n20128 , n310550 , n20127 );
buf ( n310555 , n20128 );
buf ( n310556 , n310555 );
buf ( n310557 , n864 );
buf ( n310558 , n854 );
and ( n20133 , n310557 , n310558 );
buf ( n310560 , n20133 );
buf ( n310561 , n310560 );
buf ( n310562 , n864 );
buf ( n20137 , n853 );
xor ( n20138 , n310562 , n20137 );
buf ( n310565 , n20138 );
buf ( n310566 , n310565 );
not ( n20141 , n310566 );
xnor ( n310568 , n864 , n865 );
buf ( n310569 , n310568 );
buf ( n310570 , n865 );
buf ( n310571 , n866 );
xor ( n20146 , n310570 , n310571 );
buf ( n310573 , n20146 );
buf ( n310574 , n310573 );
nor ( n20149 , n310569 , n310574 );
buf ( n310576 , n20149 );
buf ( n310577 , n310576 );
not ( n20152 , n310577 );
or ( n20153 , n20141 , n20152 );
buf ( n310580 , n310573 );
buf ( n20155 , n310580 );
buf ( n310582 , n20155 );
buf ( n20157 , n310582 );
buf ( n310584 , n864 );
buf ( n310585 , n852 );
xor ( n310586 , n310584 , n310585 );
buf ( n310587 , n310586 );
buf ( n310588 , n310587 );
nand ( n20163 , n20157 , n310588 );
buf ( n310590 , n20163 );
buf ( n310591 , n310590 );
nand ( n20166 , n20153 , n310591 );
buf ( n20167 , n20166 );
buf ( n310594 , n20167 );
xor ( n20169 , n310561 , n310594 );
buf ( n310596 , n305650 );
buf ( n310597 , n876 );
buf ( n310598 , n841 );
not ( n310599 , n310598 );
buf ( n310600 , n310599 );
buf ( n310601 , n310600 );
and ( n310602 , n310597 , n310601 );
not ( n20177 , n310597 );
buf ( n310604 , n841 );
and ( n20179 , n20177 , n310604 );
nor ( n310606 , n310602 , n20179 );
buf ( n310607 , n310606 );
buf ( n310608 , n310607 );
or ( n20183 , n310596 , n310608 );
buf ( n310610 , n305664 );
buf ( n310611 , n876 );
buf ( n310612 , n305261 );
and ( n20187 , n310611 , n310612 );
not ( n20188 , n310611 );
buf ( n310615 , n840 );
and ( n310616 , n20188 , n310615 );
nor ( n310617 , n20187 , n310616 );
buf ( n310618 , n310617 );
buf ( n310619 , n310618 );
or ( n310620 , n310610 , n310619 );
nand ( n310621 , n20183 , n310620 );
buf ( n310622 , n310621 );
buf ( n310623 , n310622 );
xor ( n20198 , n20169 , n310623 );
buf ( n310625 , n20198 );
buf ( n20200 , n310625 );
buf ( n310627 , n305627 );
not ( n310628 , n310627 );
buf ( n310629 , n310628 );
buf ( n310630 , n310629 );
buf ( n310631 , n874 );
buf ( n310632 , n843 );
xnor ( n20207 , n310631 , n310632 );
buf ( n310634 , n20207 );
buf ( n310635 , n310634 );
or ( n20210 , n310630 , n310635 );
buf ( n310637 , n306346 );
buf ( n310638 , n874 );
buf ( n310639 , n842 );
and ( n310640 , n310638 , n310639 );
not ( n20215 , n310638 );
buf ( n310642 , n304610 );
and ( n20217 , n20215 , n310642 );
nor ( n310644 , n310640 , n20217 );
buf ( n310645 , n310644 );
buf ( n310646 , n310645 );
not ( n20221 , n310646 );
buf ( n310648 , n20221 );
buf ( n310649 , n310648 );
or ( n20224 , n310637 , n310649 );
nand ( n20225 , n20210 , n20224 );
buf ( n310652 , n20225 );
buf ( n310653 , n310652 );
buf ( n310654 , n15804 );
buf ( n310655 , n884 );
buf ( n310656 , n834 );
not ( n310657 , n310656 );
buf ( n310658 , n310657 );
buf ( n310659 , n310658 );
and ( n20234 , n310655 , n310659 );
not ( n20235 , n310655 );
buf ( n310662 , n834 );
and ( n20237 , n20235 , n310662 );
nor ( n20238 , n20234 , n20237 );
buf ( n310665 , n20238 );
buf ( n310666 , n310665 );
or ( n20241 , n310654 , n310666 );
buf ( n310668 , n306238 );
buf ( n310669 , n310395 );
not ( n20244 , n310669 );
buf ( n310671 , n20244 );
buf ( n310672 , n310671 );
or ( n310673 , n310668 , n310672 );
nand ( n20248 , n20241 , n310673 );
buf ( n310675 , n20248 );
buf ( n310676 , n310675 );
xor ( n310677 , n310653 , n310676 );
buf ( n310678 , n866 );
buf ( n310679 , n852 );
and ( n20254 , n310678 , n310679 );
not ( n20255 , n310678 );
buf ( n310682 , n305168 );
and ( n20257 , n20255 , n310682 );
nor ( n20258 , n20254 , n20257 );
buf ( n310685 , n20258 );
buf ( n310686 , n310685 );
not ( n20261 , n310686 );
buf ( n310688 , n310472 );
buf ( n310689 , n20048 );
nand ( n20264 , n310688 , n310689 );
buf ( n310691 , n20264 );
buf ( n310692 , n310691 );
not ( n20267 , n310692 );
buf ( n310694 , n20267 );
buf ( n310695 , n310694 );
not ( n310696 , n310695 );
or ( n20271 , n20261 , n310696 );
buf ( n310698 , n310483 );
buf ( n310699 , n310463 );
nand ( n310700 , n310698 , n310699 );
buf ( n310701 , n310700 );
buf ( n310702 , n310701 );
nand ( n310703 , n20271 , n310702 );
buf ( n310704 , n310703 );
buf ( n310705 , n310704 );
buf ( n310706 , n304941 );
buf ( n310707 , n878 );
buf ( n310708 , n305261 );
and ( n310709 , n310707 , n310708 );
not ( n310710 , n310707 );
buf ( n310711 , n840 );
and ( n310712 , n310710 , n310711 );
nor ( n20287 , n310709 , n310712 );
buf ( n310714 , n20287 );
buf ( n310715 , n310714 );
or ( n20290 , n310706 , n310715 );
buf ( n310717 , n14523 );
buf ( n310718 , n310365 );
or ( n20293 , n310717 , n310718 );
nand ( n310720 , n20290 , n20293 );
buf ( n310721 , n310720 );
buf ( n310722 , n310721 );
xor ( n310723 , n310705 , n310722 );
buf ( n310724 , n305213 );
not ( n310725 , n310724 );
buf ( n310726 , n310725 );
buf ( n310727 , n310726 );
buf ( n310728 , n868 );
buf ( n310729 , n850 );
xnor ( n20304 , n310728 , n310729 );
buf ( n310731 , n20304 );
buf ( n310732 , n310731 );
or ( n20307 , n310727 , n310732 );
buf ( n20308 , n305205 );
buf ( n310735 , n310525 );
not ( n310736 , n310735 );
buf ( n310737 , n310736 );
buf ( n310738 , n310737 );
or ( n310739 , n20308 , n310738 );
nand ( n310740 , n20307 , n310739 );
buf ( n310741 , n310740 );
buf ( n310742 , n310741 );
and ( n310743 , n310723 , n310742 );
and ( n20318 , n310705 , n310722 );
or ( n310745 , n310743 , n20318 );
buf ( n310746 , n310745 );
buf ( n310747 , n310746 );
xor ( n310748 , n310677 , n310747 );
buf ( n310749 , n310748 );
buf ( n310750 , n310749 );
xor ( n20325 , n20200 , n310750 );
buf ( n20326 , n310675 );
not ( n310753 , n20326 );
buf ( n310754 , n310753 );
buf ( n310755 , n310754 );
xor ( n310756 , n872 , n847 );
buf ( n310757 , n310756 );
not ( n20332 , n310757 );
buf ( n310759 , n304851 );
not ( n310760 , n310759 );
or ( n20335 , n20332 , n310760 );
buf ( n310762 , n304864 );
buf ( n20337 , n872 );
buf ( n310764 , n846 );
xor ( n310765 , n20337 , n310764 );
buf ( n310766 , n310765 );
buf ( n310767 , n310766 );
nand ( n20342 , n310762 , n310767 );
buf ( n310769 , n20342 );
buf ( n310770 , n310769 );
nand ( n20345 , n20335 , n310770 );
buf ( n20346 , n20345 );
buf ( n310773 , n20346 );
buf ( n310774 , n874 );
buf ( n310775 , n845 );
not ( n20350 , n310775 );
buf ( n310777 , n20350 );
buf ( n310778 , n310777 );
and ( n20353 , n310774 , n310778 );
not ( n20354 , n310774 );
buf ( n310781 , n845 );
and ( n20356 , n20354 , n310781 );
nor ( n20357 , n20353 , n20356 );
buf ( n310784 , n20357 );
buf ( n310785 , n310784 );
not ( n20360 , n310785 );
buf ( n310787 , n20360 );
buf ( n310788 , n310787 );
not ( n20363 , n310788 );
buf ( n310790 , n305627 );
not ( n20365 , n310790 );
or ( n310792 , n20363 , n20365 );
buf ( n310793 , n874 );
buf ( n310794 , n844 );
and ( n310795 , n310793 , n310794 );
not ( n20370 , n310793 );
buf ( n310797 , n305458 );
and ( n310798 , n20370 , n310797 );
nor ( n20373 , n310795 , n310798 );
buf ( n20374 , n20373 );
buf ( n20375 , n20374 );
buf ( n310802 , n305289 );
nand ( n310803 , n20375 , n310802 );
buf ( n310804 , n310803 );
buf ( n310805 , n310804 );
nand ( n310806 , n310792 , n310805 );
buf ( n310807 , n310806 );
buf ( n310808 , n310807 );
xor ( n20383 , n310773 , n310808 );
buf ( n310810 , n304987 );
buf ( n310811 , n880 );
not ( n20386 , n310811 );
buf ( n310813 , n839 );
nor ( n310814 , n20386 , n310813 );
buf ( n310815 , n310814 );
buf ( n310816 , n310815 );
buf ( n310817 , n839 );
not ( n20392 , n310817 );
buf ( n310819 , n880 );
nor ( n310820 , n20392 , n310819 );
buf ( n310821 , n310820 );
buf ( n310822 , n310821 );
nor ( n20397 , n310816 , n310822 );
buf ( n310824 , n20397 );
buf ( n310825 , n310824 );
or ( n310826 , n310810 , n310825 );
buf ( n310827 , n304976 );
buf ( n310828 , n838 );
buf ( n310829 , n880 );
xor ( n20404 , n310828 , n310829 );
buf ( n310831 , n20404 );
buf ( n310832 , n310831 );
not ( n20407 , n310832 );
buf ( n310834 , n20407 );
buf ( n310835 , n310834 );
or ( n310836 , n310827 , n310835 );
nand ( n20411 , n310826 , n310836 );
buf ( n20412 , n20411 );
buf ( n310839 , n20412 );
and ( n20414 , n20383 , n310839 );
and ( n310841 , n310773 , n310808 );
or ( n310842 , n20414 , n310841 );
buf ( n310843 , n310842 );
buf ( n310844 , n310843 );
xor ( n20419 , n310755 , n310844 );
buf ( n20420 , n849 );
buf ( n20421 , n870 );
xor ( n20422 , n20420 , n20421 );
buf ( n310849 , n20422 );
buf ( n310850 , n310849 );
not ( n20425 , n310850 );
buf ( n310852 , n14323 );
not ( n20427 , n310852 );
or ( n20428 , n20425 , n20427 );
buf ( n310855 , n304763 );
buf ( n310856 , n870 );
buf ( n310857 , n848 );
xor ( n20432 , n310856 , n310857 );
buf ( n310859 , n20432 );
buf ( n310860 , n310859 );
nand ( n20435 , n310855 , n310860 );
buf ( n310862 , n20435 );
buf ( n310863 , n310862 );
nand ( n310864 , n20428 , n310863 );
buf ( n310865 , n310864 );
buf ( n310866 , n310865 );
buf ( n310867 , n851 );
buf ( n310868 , n310521 );
and ( n20443 , n310867 , n310868 );
not ( n310870 , n310867 );
buf ( n310871 , n868 );
and ( n310872 , n310870 , n310871 );
nor ( n20447 , n20443 , n310872 );
buf ( n310874 , n20447 );
buf ( n20449 , n310874 );
not ( n310876 , n20449 );
buf ( n310877 , n310876 );
buf ( n310878 , n310877 );
not ( n310879 , n310878 );
buf ( n310880 , n305213 );
not ( n20455 , n310880 );
or ( n310882 , n310879 , n20455 );
buf ( n310883 , n310731 );
not ( n20458 , n310883 );
buf ( n310885 , n305219 );
nand ( n310886 , n20458 , n310885 );
buf ( n310887 , n310886 );
buf ( n310888 , n310887 );
nand ( n310889 , n310882 , n310888 );
buf ( n310890 , n310889 );
buf ( n20465 , n310890 );
xor ( n20466 , n310866 , n20465 );
buf ( n310893 , n15804 );
buf ( n310894 , n835 );
buf ( n310895 , n884 );
and ( n310896 , n310894 , n310895 );
not ( n310897 , n310894 );
buf ( n310898 , n304827 );
and ( n20473 , n310897 , n310898 );
nor ( n310900 , n310896 , n20473 );
buf ( n310901 , n310900 );
buf ( n310902 , n310901 );
not ( n310903 , n310902 );
buf ( n310904 , n310903 );
buf ( n310905 , n310904 );
or ( n20480 , n310893 , n310905 );
buf ( n310907 , n304807 );
not ( n310908 , n310907 );
buf ( n310909 , n310908 );
buf ( n310910 , n310909 );
buf ( n310911 , n310665 );
or ( n20486 , n310910 , n310911 );
nand ( n310913 , n20480 , n20486 );
buf ( n310914 , n310913 );
buf ( n310915 , n310914 );
and ( n310916 , n20466 , n310915 );
and ( n310917 , n310866 , n20465 );
or ( n310918 , n310916 , n310917 );
buf ( n310919 , n310918 );
buf ( n310920 , n310919 );
and ( n310921 , n20419 , n310920 );
and ( n20496 , n310755 , n310844 );
or ( n310923 , n310921 , n20496 );
buf ( n310924 , n310923 );
buf ( n310925 , n310924 );
xor ( n310926 , n20325 , n310925 );
buf ( n310927 , n310926 );
buf ( n310928 , n310927 );
xor ( n20503 , n310556 , n310928 );
buf ( n310930 , n856 );
buf ( n310931 , n864 );
and ( n20506 , n310930 , n310931 );
buf ( n310933 , n20506 );
buf ( n310934 , n310933 );
and ( n20509 , n876 , n843 );
not ( n310936 , n876 );
and ( n20511 , n310936 , n305117 );
nor ( n310938 , n20509 , n20511 );
not ( n20513 , n310938 );
not ( n20514 , n305338 );
or ( n20515 , n20513 , n20514 );
buf ( n310942 , n842 );
buf ( n310943 , n876 );
xnor ( n310944 , n310942 , n310943 );
buf ( n310945 , n310944 );
not ( n20520 , n310945 );
nand ( n20521 , n20520 , n305344 );
nand ( n310948 , n20515 , n20521 );
buf ( n310949 , n310948 );
xor ( n20524 , n310934 , n310949 );
xor ( n20525 , n886 , n834 );
buf ( n310952 , n20525 );
not ( n310953 , n310952 );
buf ( n310954 , n304912 );
not ( n20529 , n310954 );
or ( n310956 , n310953 , n20529 );
buf ( n310957 , n304901 );
buf ( n310958 , n886 );
buf ( n310959 , n833 );
and ( n310960 , n310958 , n310959 );
not ( n20535 , n310958 );
buf ( n310962 , n833 );
not ( n20537 , n310962 );
buf ( n310964 , n20537 );
buf ( n310965 , n310964 );
and ( n20540 , n20535 , n310965 );
nor ( n310967 , n310960 , n20540 );
buf ( n310968 , n310967 );
buf ( n310969 , n310968 );
nand ( n310970 , n310957 , n310969 );
buf ( n310971 , n310970 );
buf ( n310972 , n310971 );
nand ( n20547 , n310956 , n310972 );
buf ( n20548 , n20547 );
buf ( n310975 , n20548 );
and ( n310976 , n20524 , n310975 );
and ( n20551 , n310934 , n310949 );
or ( n20552 , n310976 , n20551 );
buf ( n310979 , n20552 );
buf ( n310980 , n310979 );
buf ( n310981 , n838 );
buf ( n310982 , n882 );
xor ( n20557 , n310981 , n310982 );
buf ( n310984 , n20557 );
buf ( n310985 , n310984 );
not ( n310986 , n310985 );
buf ( n310987 , n304584 );
not ( n20562 , n310987 );
or ( n310989 , n310986 , n20562 );
buf ( n310990 , n304596 );
buf ( n310991 , n837 );
buf ( n310992 , n882 );
xor ( n310993 , n310991 , n310992 );
buf ( n310994 , n310993 );
buf ( n310995 , n310994 );
nand ( n310996 , n310990 , n310995 );
buf ( n310997 , n310996 );
buf ( n310998 , n310997 );
nand ( n20573 , n310989 , n310998 );
buf ( n20574 , n20573 );
buf ( n311001 , n20574 );
buf ( n311002 , n872 );
buf ( n311003 , n848 );
xor ( n20578 , n311002 , n311003 );
buf ( n311005 , n20578 );
buf ( n311006 , n311005 );
not ( n20581 , n311006 );
buf ( n311008 , n306132 );
not ( n20583 , n311008 );
or ( n311010 , n20581 , n20583 );
buf ( n311011 , n304845 );
buf ( n311012 , n310756 );
nand ( n311013 , n311011 , n311012 );
buf ( n311014 , n311013 );
buf ( n311015 , n311014 );
nand ( n311016 , n311010 , n311015 );
buf ( n311017 , n311016 );
buf ( n311018 , n311017 );
xor ( n311019 , n311001 , n311018 );
buf ( n311020 , n310629 );
buf ( n311021 , n874 );
buf ( n311022 , n846 );
not ( n311023 , n311022 );
buf ( n311024 , n311023 );
buf ( n311025 , n311024 );
and ( n20600 , n311021 , n311025 );
not ( n20601 , n311021 );
buf ( n311028 , n846 );
and ( n311029 , n20601 , n311028 );
nor ( n311030 , n20600 , n311029 );
buf ( n311031 , n311030 );
buf ( n311032 , n311031 );
or ( n20607 , n311020 , n311032 );
buf ( n311034 , n305298 );
buf ( n311035 , n310784 );
or ( n20610 , n311034 , n311035 );
nand ( n311037 , n20607 , n20610 );
buf ( n311038 , n311037 );
buf ( n311039 , n311038 );
and ( n311040 , n311019 , n311039 );
and ( n311041 , n311001 , n311018 );
or ( n20616 , n311040 , n311041 );
buf ( n311043 , n20616 );
buf ( n311044 , n311043 );
xor ( n20619 , n870 , n850 );
buf ( n20620 , n20619 );
not ( n20621 , n20620 );
buf ( n311048 , n14320 );
not ( n20623 , n311048 );
buf ( n311050 , n14318 );
not ( n311051 , n311050 );
buf ( n311052 , n311051 );
buf ( n20627 , n311052 );
nor ( n20628 , n20623 , n20627 );
buf ( n20629 , n20628 );
buf ( n311056 , n20629 );
not ( n20631 , n311056 );
or ( n311058 , n20621 , n20631 );
buf ( n311059 , n311052 );
buf ( n311060 , n310849 );
nand ( n20635 , n311059 , n311060 );
buf ( n311062 , n20635 );
buf ( n311063 , n311062 );
nand ( n20638 , n311058 , n311063 );
buf ( n311065 , n20638 );
buf ( n311066 , n880 );
buf ( n311067 , n840 );
xor ( n20642 , n311066 , n311067 );
buf ( n311069 , n20642 );
not ( n20644 , n311069 );
not ( n20645 , n304984 );
or ( n20646 , n20644 , n20645 );
buf ( n311073 , n304973 );
not ( n20648 , n311073 );
buf ( n311075 , n20648 );
or ( n20650 , n311075 , n310824 );
nand ( n311077 , n20646 , n20650 );
xor ( n20652 , n311065 , n311077 );
buf ( n311079 , n310726 );
buf ( n20654 , n852 );
buf ( n311081 , n868 );
xnor ( n311082 , n20654 , n311081 );
buf ( n311083 , n311082 );
buf ( n311084 , n311083 );
or ( n311085 , n311079 , n311084 );
buf ( n311086 , n305449 );
buf ( n311087 , n310874 );
or ( n20662 , n311086 , n311087 );
nand ( n311089 , n311085 , n20662 );
buf ( n311090 , n311089 );
and ( n20665 , n20652 , n311090 );
and ( n311092 , n311065 , n311077 );
or ( n311093 , n20665 , n311092 );
buf ( n311094 , n311093 );
xor ( n311095 , n311044 , n311094 );
buf ( n311096 , n854 );
buf ( n311097 , n866 );
xor ( n311098 , n311096 , n311097 );
buf ( n311099 , n311098 );
buf ( n20674 , n311099 );
not ( n20675 , n20674 );
buf ( n311102 , n310694 );
not ( n311103 , n311102 );
or ( n20678 , n20675 , n311103 );
buf ( n311105 , n310472 );
not ( n20680 , n311105 );
buf ( n311107 , n20680 );
buf ( n20682 , n311107 );
buf ( n311109 , n866 );
buf ( n311110 , n853 );
xor ( n20685 , n311109 , n311110 );
buf ( n311112 , n20685 );
buf ( n20687 , n311112 );
nand ( n20688 , n20682 , n20687 );
buf ( n20689 , n20688 );
buf ( n311116 , n20689 );
nand ( n20691 , n20678 , n311116 );
buf ( n311118 , n20691 );
buf ( n311119 , n311118 );
buf ( n311120 , n888 );
buf ( n311121 , n832 );
and ( n20696 , n311120 , n311121 );
not ( n20697 , n311120 );
buf ( n20698 , n832 );
not ( n20699 , n20698 );
buf ( n20700 , n20699 );
buf ( n20701 , n20700 );
and ( n311128 , n20697 , n20701 );
nor ( n20703 , n20696 , n311128 );
buf ( n20704 , n20703 );
buf ( n311131 , n20704 );
not ( n20706 , n311131 );
buf ( n311133 , n305138 );
not ( n20708 , n311133 );
or ( n311135 , n20706 , n20708 );
buf ( n311136 , n305127 );
buf ( n311137 , n888 );
nand ( n311138 , n311136 , n311137 );
buf ( n311139 , n311138 );
buf ( n311140 , n311139 );
nand ( n311141 , n311135 , n311140 );
buf ( n311142 , n311141 );
buf ( n311143 , n311142 );
xor ( n311144 , n311119 , n311143 );
buf ( n311145 , n304941 );
buf ( n311146 , n310371 );
buf ( n311147 , n842 );
and ( n311148 , n311146 , n311147 );
buf ( n311149 , n304610 );
buf ( n311150 , n878 );
and ( n311151 , n311149 , n311150 );
nor ( n20726 , n311148 , n311151 );
buf ( n20727 , n20726 );
buf ( n311154 , n20727 );
or ( n20729 , n311145 , n311154 );
buf ( n311156 , n14523 );
buf ( n311157 , n310371 );
buf ( n311158 , n841 );
and ( n311159 , n311157 , n311158 );
buf ( n311160 , n310600 );
buf ( n311161 , n878 );
and ( n20736 , n311160 , n311161 );
nor ( n311163 , n311159 , n20736 );
buf ( n311164 , n311163 );
buf ( n311165 , n311164 );
or ( n311166 , n311156 , n311165 );
nand ( n311167 , n20729 , n311166 );
buf ( n311168 , n311167 );
buf ( n311169 , n311168 );
and ( n311170 , n311144 , n311169 );
and ( n20745 , n311119 , n311143 );
or ( n311172 , n311170 , n20745 );
buf ( n311173 , n311172 );
buf ( n311174 , n311173 );
and ( n311175 , n311095 , n311174 );
and ( n311176 , n311044 , n311094 );
or ( n20751 , n311175 , n311176 );
buf ( n311178 , n20751 );
buf ( n311179 , n311178 );
xor ( n20754 , n310980 , n311179 );
xor ( n20755 , n310755 , n310844 );
xor ( n20756 , n20755 , n310920 );
buf ( n311183 , n20756 );
buf ( n311184 , n311183 );
and ( n311185 , n20754 , n311184 );
and ( n20760 , n310980 , n311179 );
or ( n20761 , n311185 , n20760 );
buf ( n311188 , n20761 );
buf ( n311189 , n311188 );
xor ( n20764 , n20503 , n311189 );
buf ( n311191 , n20764 );
buf ( n311192 , n311191 );
buf ( n311193 , n857 );
buf ( n311194 , n864 );
and ( n311195 , n311193 , n311194 );
buf ( n311196 , n311195 );
buf ( n311197 , n311196 );
buf ( n311198 , n884 );
buf ( n20773 , n836 );
and ( n20774 , n311198 , n20773 );
not ( n311201 , n311198 );
buf ( n311202 , n836 );
not ( n20777 , n311202 );
buf ( n311204 , n20777 );
buf ( n311205 , n311204 );
and ( n311206 , n311201 , n311205 );
nor ( n311207 , n20774 , n311206 );
buf ( n311208 , n311207 );
buf ( n311209 , n311208 );
not ( n20784 , n311209 );
buf ( n311211 , n304813 );
not ( n20786 , n311211 );
or ( n311213 , n20784 , n20786 );
buf ( n20788 , n304819 );
buf ( n20789 , n310901 );
nand ( n20790 , n20788 , n20789 );
buf ( n20791 , n20790 );
buf ( n311218 , n20791 );
nand ( n20793 , n311213 , n311218 );
buf ( n20794 , n20793 );
buf ( n311221 , n20794 );
xor ( n20796 , n311197 , n311221 );
buf ( n20797 , n310573 );
buf ( n311224 , n310568 );
nor ( n311225 , n20797 , n311224 );
buf ( n311226 , n311225 );
buf ( n311227 , n311226 );
not ( n311228 , n311227 );
buf ( n311229 , n311228 );
buf ( n311230 , n311229 );
buf ( n311231 , n856 );
buf ( n311232 , n864 );
not ( n20807 , n311232 );
buf ( n311234 , n20807 );
buf ( n311235 , n311234 );
and ( n20810 , n311231 , n311235 );
not ( n311237 , n311231 );
buf ( n311238 , n864 );
and ( n20813 , n311237 , n311238 );
nor ( n20814 , n20810 , n20813 );
buf ( n311241 , n20814 );
buf ( n311242 , n311241 );
or ( n20817 , n311230 , n311242 );
buf ( n311244 , n310582 );
not ( n20819 , n311244 );
buf ( n311246 , n20819 );
buf ( n311247 , n311246 );
buf ( n311248 , n311234 );
buf ( n311249 , n855 );
and ( n20824 , n311248 , n311249 );
buf ( n311251 , n305319 );
buf ( n311252 , n864 );
and ( n20827 , n311251 , n311252 );
nor ( n20828 , n20824 , n20827 );
buf ( n311255 , n20828 );
buf ( n311256 , n311255 );
or ( n311257 , n311247 , n311256 );
nand ( n20832 , n20817 , n311257 );
buf ( n20833 , n20832 );
buf ( n311260 , n20833 );
and ( n20835 , n20796 , n311260 );
and ( n311262 , n311197 , n311221 );
or ( n311263 , n20835 , n311262 );
buf ( n311264 , n311263 );
buf ( n311265 , n311264 );
xor ( n20840 , n310773 , n310808 );
xor ( n311267 , n20840 , n310839 );
buf ( n311268 , n311267 );
buf ( n311269 , n311268 );
xor ( n20844 , n311265 , n311269 );
buf ( n311271 , n305130 );
not ( n20846 , n311271 );
buf ( n311273 , n305138 );
not ( n311274 , n311273 );
buf ( n311275 , n311274 );
buf ( n311276 , n311275 );
not ( n20851 , n311276 );
or ( n311278 , n20846 , n20851 );
buf ( n311279 , n888 );
nand ( n20854 , n311278 , n311279 );
buf ( n20855 , n20854 );
buf ( n311282 , n20855 );
buf ( n311283 , n310968 );
not ( n311284 , n311283 );
buf ( n311285 , n304912 );
not ( n311286 , n311285 );
or ( n20861 , n311284 , n311286 );
buf ( n311288 , n304901 );
buf ( n311289 , n886 );
buf ( n311290 , n832 );
and ( n311291 , n311289 , n311290 );
not ( n311292 , n311289 );
buf ( n311293 , n20700 );
and ( n311294 , n311292 , n311293 );
nor ( n20869 , n311291 , n311294 );
buf ( n311296 , n20869 );
buf ( n311297 , n311296 );
nand ( n20872 , n311288 , n311297 );
buf ( n20873 , n20872 );
buf ( n311300 , n20873 );
nand ( n311301 , n20861 , n311300 );
buf ( n311302 , n311301 );
buf ( n311303 , n311302 );
xor ( n20878 , n311282 , n311303 );
buf ( n311305 , n304581 );
buf ( n20880 , n310994 );
not ( n311307 , n20880 );
buf ( n311308 , n311307 );
buf ( n311309 , n311308 );
or ( n311310 , n311305 , n311309 );
buf ( n311311 , n14959 );
buf ( n311312 , n882 );
buf ( n311313 , n836 );
xor ( n20888 , n311312 , n311313 );
buf ( n311315 , n20888 );
buf ( n311316 , n311315 );
not ( n20891 , n311316 );
buf ( n311318 , n20891 );
buf ( n311319 , n311318 );
or ( n20894 , n311311 , n311319 );
nand ( n20895 , n311310 , n20894 );
buf ( n311322 , n20895 );
buf ( n311323 , n311322 );
xor ( n20898 , n20878 , n311323 );
buf ( n311325 , n20898 );
buf ( n311326 , n311325 );
and ( n311327 , n20844 , n311326 );
and ( n20902 , n311265 , n311269 );
or ( n311329 , n311327 , n20902 );
buf ( n311330 , n311329 );
buf ( n311331 , n311330 );
xor ( n311332 , n310934 , n310949 );
xor ( n311333 , n311332 , n310975 );
buf ( n311334 , n311333 );
buf ( n311335 , n311334 );
buf ( n20910 , n311255 );
not ( n311337 , n20910 );
buf ( n311338 , n311337 );
buf ( n311339 , n311338 );
not ( n311340 , n311339 );
buf ( n311341 , n310576 );
not ( n20916 , n311341 );
or ( n311343 , n311340 , n20916 );
buf ( n311344 , n310582 );
xor ( n20919 , n310557 , n310558 );
buf ( n311346 , n20919 );
buf ( n311347 , n311346 );
nand ( n311348 , n311344 , n311347 );
buf ( n311349 , n311348 );
buf ( n311350 , n311349 );
nand ( n20925 , n311343 , n311350 );
buf ( n311352 , n20925 );
buf ( n311353 , n311352 );
buf ( n311354 , n311112 );
not ( n311355 , n311354 );
buf ( n311356 , n310694 );
not ( n20931 , n311356 );
or ( n311358 , n311355 , n20931 );
buf ( n20933 , n311107 );
buf ( n20934 , n310685 );
nand ( n20935 , n20933 , n20934 );
buf ( n20936 , n20935 );
buf ( n311363 , n20936 );
nand ( n20938 , n311358 , n311363 );
buf ( n311365 , n20938 );
buf ( n311366 , n311365 );
xor ( n20941 , n311353 , n311366 );
buf ( n311368 , n304941 );
buf ( n311369 , n311164 );
or ( n20944 , n311368 , n311369 );
buf ( n311371 , n14523 );
buf ( n311372 , n310714 );
or ( n311373 , n311371 , n311372 );
nand ( n311374 , n20944 , n311373 );
buf ( n311375 , n311374 );
buf ( n311376 , n311375 );
xor ( n311377 , n20941 , n311376 );
buf ( n311378 , n311377 );
buf ( n311379 , n311378 );
xor ( n311380 , n311335 , n311379 );
xor ( n20955 , n310866 , n20465 );
xor ( n20956 , n20955 , n310915 );
buf ( n311383 , n20956 );
buf ( n311384 , n311383 );
and ( n20959 , n311380 , n311384 );
and ( n20960 , n311335 , n311379 );
or ( n20961 , n20959 , n20960 );
buf ( n311388 , n20961 );
buf ( n311389 , n311388 );
xor ( n20964 , n311331 , n311389 );
buf ( n311391 , n855 );
buf ( n311392 , n864 );
and ( n311393 , n311391 , n311392 );
buf ( n311394 , n311393 );
buf ( n311395 , n311394 );
buf ( n311396 , n311315 );
not ( n311397 , n311396 );
buf ( n311398 , n304584 );
not ( n20973 , n311398 );
or ( n311400 , n311397 , n20973 );
buf ( n311401 , n304596 );
buf ( n311402 , n310496 );
nand ( n20977 , n311401 , n311402 );
buf ( n311404 , n20977 );
buf ( n311405 , n311404 );
nand ( n311406 , n311400 , n311405 );
buf ( n311407 , n311406 );
buf ( n20982 , n311407 );
xor ( n20983 , n311395 , n20982 );
buf ( n311410 , n20374 );
not ( n311411 , n311410 );
buf ( n311412 , n305627 );
not ( n311413 , n311412 );
or ( n20988 , n311411 , n311413 );
buf ( n311415 , n310634 );
not ( n311416 , n311415 );
buf ( n311417 , n305301 );
nand ( n311418 , n311416 , n311417 );
buf ( n311419 , n311418 );
buf ( n311420 , n311419 );
nand ( n311421 , n20988 , n311420 );
buf ( n311422 , n311421 );
buf ( n311423 , n311422 );
xor ( n20998 , n20983 , n311423 );
buf ( n311425 , n20998 );
buf ( n311426 , n311425 );
xor ( n21001 , n311282 , n311303 );
and ( n311428 , n21001 , n311323 );
and ( n21003 , n311282 , n311303 );
or ( n21004 , n311428 , n21003 );
buf ( n311431 , n21004 );
buf ( n311432 , n311431 );
xor ( n21007 , n311426 , n311432 );
xor ( n21008 , n311353 , n311366 );
and ( n21009 , n21008 , n311376 );
and ( n21010 , n311353 , n311366 );
or ( n21011 , n21009 , n21010 );
buf ( n311438 , n21011 );
buf ( n311439 , n311438 );
xor ( n21014 , n21007 , n311439 );
buf ( n311441 , n21014 );
buf ( n311442 , n311441 );
and ( n21017 , n20964 , n311442 );
and ( n21018 , n311331 , n311389 );
or ( n21019 , n21017 , n21018 );
buf ( n311446 , n21019 );
buf ( n311447 , n311446 );
xor ( n21022 , n311426 , n311432 );
and ( n311449 , n21022 , n311439 );
and ( n21024 , n311426 , n311432 );
or ( n311451 , n311449 , n21024 );
buf ( n311452 , n311451 );
buf ( n311453 , n311452 );
buf ( n311454 , n310859 );
not ( n21029 , n311454 );
buf ( n311456 , n20629 );
not ( n21031 , n311456 );
or ( n311458 , n21029 , n21031 );
buf ( n311459 , n304763 );
buf ( n311460 , n19901 );
nand ( n311461 , n311459 , n311460 );
buf ( n311462 , n311461 );
buf ( n311463 , n311462 );
nand ( n21038 , n311458 , n311463 );
buf ( n311465 , n21038 );
buf ( n311466 , n311465 );
buf ( n311467 , n310766 );
not ( n21042 , n311467 );
buf ( n311469 , n306132 );
not ( n311470 , n311469 );
or ( n21045 , n21042 , n311470 );
buf ( n311472 , n304864 );
buf ( n311473 , n19916 );
nand ( n311474 , n311472 , n311473 );
buf ( n311475 , n311474 );
buf ( n311476 , n311475 );
nand ( n21051 , n21045 , n311476 );
buf ( n311478 , n21051 );
buf ( n311479 , n311478 );
or ( n21054 , n311466 , n311479 );
buf ( n311481 , n310831 );
not ( n21056 , n311481 );
buf ( n311483 , n305098 );
not ( n311484 , n311483 );
or ( n21059 , n21056 , n311484 );
buf ( n311486 , n310441 );
not ( n21061 , n311486 );
buf ( n311488 , n304997 );
nand ( n21063 , n21061 , n311488 );
buf ( n311490 , n21063 );
buf ( n311491 , n311490 );
nand ( n311492 , n21059 , n311491 );
buf ( n311493 , n311492 );
buf ( n311494 , n311493 );
nand ( n311495 , n21054 , n311494 );
buf ( n311496 , n311495 );
buf ( n311497 , n311496 );
buf ( n311498 , n311465 );
buf ( n311499 , n311478 );
nand ( n311500 , n311498 , n311499 );
buf ( n311501 , n311500 );
buf ( n311502 , n311501 );
nand ( n311503 , n311497 , n311502 );
buf ( n311504 , n311503 );
buf ( n311505 , n311504 );
xor ( n311506 , n311395 , n20982 );
and ( n21081 , n311506 , n311423 );
and ( n21082 , n311395 , n20982 );
or ( n21083 , n21081 , n21082 );
buf ( n311510 , n21083 );
buf ( n311511 , n311510 );
xor ( n21086 , n311505 , n311511 );
buf ( n311513 , n311346 );
not ( n21088 , n311513 );
buf ( n311515 , n311226 );
not ( n311516 , n311515 );
or ( n311517 , n21088 , n311516 );
buf ( n311518 , n310582 );
buf ( n311519 , n310565 );
nand ( n311520 , n311518 , n311519 );
buf ( n311521 , n311520 );
buf ( n311522 , n311521 );
nand ( n21097 , n311517 , n311522 );
buf ( n311524 , n21097 );
buf ( n311525 , n311524 );
buf ( n311526 , n311296 );
not ( n311527 , n311526 );
buf ( n311528 , n304912 );
not ( n311529 , n311528 );
or ( n21104 , n311527 , n311529 );
buf ( n311531 , n304901 );
buf ( n21106 , n886 );
nand ( n21107 , n311531 , n21106 );
buf ( n21108 , n21107 );
buf ( n21109 , n21108 );
nand ( n21110 , n21104 , n21109 );
buf ( n21111 , n21110 );
buf ( n311538 , n21111 );
xor ( n21113 , n311525 , n311538 );
buf ( n311540 , n305650 );
buf ( n311541 , n310945 );
or ( n21116 , n311540 , n311541 );
buf ( n311543 , n305664 );
buf ( n311544 , n310607 );
or ( n21119 , n311543 , n311544 );
nand ( n21120 , n21116 , n21119 );
buf ( n21121 , n21120 );
buf ( n311548 , n21121 );
and ( n21123 , n21113 , n311548 );
and ( n311550 , n311525 , n311538 );
or ( n21125 , n21123 , n311550 );
buf ( n311552 , n21125 );
buf ( n311553 , n311552 );
xor ( n21128 , n21086 , n311553 );
buf ( n311555 , n21128 );
buf ( n311556 , n311555 );
xor ( n21131 , n311453 , n311556 );
buf ( n311558 , n311493 );
buf ( n311559 , n311478 );
xor ( n311560 , n311558 , n311559 );
buf ( n311561 , n311560 );
buf ( n311562 , n311561 );
buf ( n311563 , n311465 );
xor ( n21138 , n311562 , n311563 );
buf ( n21139 , n21138 );
buf ( n21140 , n21139 );
xor ( n311567 , n311525 , n311538 );
xor ( n311568 , n311567 , n311548 );
buf ( n311569 , n311568 );
buf ( n311570 , n311569 );
xor ( n311571 , n21140 , n311570 );
xor ( n21146 , n310705 , n310722 );
xor ( n311573 , n21146 , n310742 );
buf ( n311574 , n311573 );
buf ( n311575 , n311574 );
and ( n21150 , n311571 , n311575 );
and ( n21151 , n21140 , n311570 );
or ( n21152 , n21150 , n21151 );
buf ( n311579 , n21152 );
buf ( n311580 , n311579 );
xor ( n21155 , n21131 , n311580 );
buf ( n311582 , n21155 );
buf ( n311583 , n311582 );
xor ( n311584 , n311447 , n311583 );
xor ( n21159 , n21140 , n311570 );
xor ( n21160 , n21159 , n311575 );
buf ( n311587 , n21160 );
buf ( n311588 , n311587 );
xor ( n21163 , n876 , n844 );
buf ( n311590 , n21163 );
not ( n21165 , n311590 );
buf ( n311592 , n305338 );
not ( n21167 , n311592 );
or ( n21168 , n21165 , n21167 );
buf ( n311595 , n305344 );
buf ( n311596 , n310938 );
nand ( n21171 , n311595 , n311596 );
buf ( n311598 , n21171 );
buf ( n311599 , n311598 );
nand ( n21174 , n21168 , n311599 );
buf ( n21175 , n21174 );
buf ( n311602 , n21175 );
buf ( n311603 , n20548 );
not ( n311604 , n311603 );
buf ( n311605 , n311604 );
buf ( n311606 , n311605 );
xor ( n311607 , n311602 , n311606 );
xor ( n21182 , n866 , n855 );
buf ( n311609 , n21182 );
not ( n311610 , n311609 );
buf ( n311611 , n310477 );
not ( n21186 , n311611 );
or ( n311613 , n311610 , n21186 );
buf ( n21188 , n311107 );
buf ( n311615 , n311099 );
nand ( n311616 , n21188 , n311615 );
buf ( n311617 , n311616 );
buf ( n311618 , n311617 );
nand ( n21193 , n311613 , n311618 );
buf ( n311620 , n21193 );
buf ( n311621 , n311620 );
buf ( n311622 , n880 );
buf ( n311623 , n841 );
and ( n311624 , n311622 , n311623 );
not ( n21199 , n311622 );
buf ( n311626 , n310600 );
and ( n311627 , n21199 , n311626 );
nor ( n311628 , n311624 , n311627 );
buf ( n311629 , n311628 );
buf ( n311630 , n311629 );
not ( n311631 , n311630 );
buf ( n311632 , n304984 );
not ( n311633 , n311632 );
or ( n311634 , n311631 , n311633 );
buf ( n21209 , n311069 );
buf ( n311636 , n304973 );
nand ( n311637 , n21209 , n311636 );
buf ( n311638 , n311637 );
buf ( n311639 , n311638 );
nand ( n21214 , n311634 , n311639 );
buf ( n311641 , n21214 );
buf ( n311642 , n311641 );
xor ( n21217 , n311621 , n311642 );
buf ( n311644 , n305210 );
xor ( n311645 , n868 , n853 );
buf ( n311646 , n311645 );
not ( n311647 , n311646 );
buf ( n311648 , n311647 );
buf ( n311649 , n311648 );
or ( n21224 , n311644 , n311649 );
buf ( n311651 , n305205 );
buf ( n311652 , n311083 );
or ( n21227 , n311651 , n311652 );
nand ( n21228 , n21224 , n21227 );
buf ( n311655 , n21228 );
buf ( n311656 , n311655 );
and ( n21231 , n21217 , n311656 );
and ( n21232 , n311621 , n311642 );
or ( n311659 , n21231 , n21232 );
buf ( n311660 , n311659 );
buf ( n311661 , n311660 );
and ( n311662 , n311607 , n311661 );
and ( n311663 , n311602 , n311606 );
or ( n311664 , n311662 , n311663 );
buf ( n311665 , n311664 );
buf ( n311666 , n311665 );
xor ( n311667 , n870 , n851 );
buf ( n21242 , n311667 );
not ( n21243 , n21242 );
buf ( n21244 , n14323 );
not ( n21245 , n21244 );
or ( n21246 , n21243 , n21245 );
buf ( n21247 , n304763 );
buf ( n311674 , n20619 );
nand ( n311675 , n21247 , n311674 );
buf ( n311676 , n311675 );
buf ( n311677 , n311676 );
nand ( n21252 , n21246 , n311677 );
buf ( n21253 , n21252 );
buf ( n311680 , n21253 );
buf ( n311681 , n886 );
buf ( n311682 , n835 );
and ( n311683 , n311681 , n311682 );
not ( n311684 , n311681 );
buf ( n311685 , n835 );
not ( n21260 , n311685 );
buf ( n21261 , n21260 );
buf ( n311688 , n21261 );
and ( n21263 , n311684 , n311688 );
nor ( n311690 , n311683 , n21263 );
buf ( n311691 , n311690 );
buf ( n311692 , n311691 );
not ( n311693 , n311692 );
buf ( n311694 , n304906 );
buf ( n311695 , n304901 );
nor ( n311696 , n311694 , n311695 );
buf ( n311697 , n311696 );
buf ( n311698 , n311697 );
not ( n311699 , n311698 );
or ( n311700 , n311693 , n311699 );
buf ( n311701 , n304901 );
buf ( n311702 , n20525 );
nand ( n311703 , n311701 , n311702 );
buf ( n311704 , n311703 );
buf ( n21279 , n311704 );
nand ( n21280 , n311700 , n21279 );
buf ( n21281 , n21280 );
buf ( n311708 , n21281 );
or ( n311709 , n311680 , n311708 );
buf ( n311710 , n872 );
buf ( n311711 , n849 );
and ( n311712 , n311710 , n311711 );
not ( n311713 , n311710 );
buf ( n311714 , n305596 );
and ( n21289 , n311713 , n311714 );
nor ( n311716 , n311712 , n21289 );
buf ( n311717 , n311716 );
buf ( n311718 , n311717 );
not ( n311719 , n311718 );
buf ( n311720 , n304851 );
not ( n21295 , n311720 );
or ( n21296 , n311719 , n21295 );
buf ( n311723 , n304845 );
buf ( n311724 , n311005 );
nand ( n21299 , n311723 , n311724 );
buf ( n311726 , n21299 );
buf ( n311727 , n311726 );
nand ( n311728 , n21296 , n311727 );
buf ( n311729 , n311728 );
buf ( n311730 , n311729 );
nand ( n311731 , n311709 , n311730 );
buf ( n311732 , n311731 );
buf ( n311733 , n311732 );
buf ( n311734 , n21253 );
buf ( n311735 , n21281 );
nand ( n311736 , n311734 , n311735 );
buf ( n311737 , n311736 );
buf ( n311738 , n311737 );
nand ( n311739 , n311733 , n311738 );
buf ( n311740 , n311739 );
buf ( n311741 , n311740 );
xor ( n311742 , n882 , n839 );
buf ( n311743 , n311742 );
not ( n21318 , n311743 );
buf ( n311745 , n304584 );
not ( n311746 , n311745 );
or ( n21321 , n21318 , n311746 );
buf ( n311748 , n304596 );
buf ( n311749 , n310984 );
nand ( n21324 , n311748 , n311749 );
buf ( n311751 , n21324 );
buf ( n311752 , n311751 );
nand ( n311753 , n21321 , n311752 );
buf ( n311754 , n311753 );
buf ( n311755 , n311754 );
buf ( n311756 , n845 );
buf ( n311757 , n876 );
xor ( n311758 , n311756 , n311757 );
buf ( n311759 , n311758 );
buf ( n311760 , n311759 );
not ( n311761 , n311760 );
buf ( n311762 , n305338 );
not ( n21337 , n311762 );
or ( n311764 , n311761 , n21337 );
buf ( n311765 , n305344 );
buf ( n311766 , n21163 );
nand ( n311767 , n311765 , n311766 );
buf ( n311768 , n311767 );
buf ( n311769 , n311768 );
nand ( n311770 , n311764 , n311769 );
buf ( n311771 , n311770 );
buf ( n311772 , n311771 );
xor ( n311773 , n311755 , n311772 );
buf ( n311774 , n305627 );
not ( n21349 , n311774 );
buf ( n21350 , n874 );
buf ( n311777 , n847 );
xor ( n311778 , n21350 , n311777 );
buf ( n311779 , n311778 );
buf ( n311780 , n311779 );
not ( n311781 , n311780 );
or ( n21356 , n21349 , n311781 );
buf ( n311783 , n305298 );
buf ( n311784 , n311031 );
or ( n21359 , n311783 , n311784 );
nand ( n311786 , n21356 , n21359 );
buf ( n311787 , n311786 );
buf ( n311788 , n311787 );
and ( n311789 , n311773 , n311788 );
and ( n311790 , n311755 , n311772 );
or ( n21365 , n311789 , n311790 );
buf ( n311792 , n21365 );
buf ( n311793 , n311792 );
xor ( n311794 , n311741 , n311793 );
xor ( n21369 , n888 , n833 );
buf ( n311796 , n21369 );
not ( n21371 , n311796 );
buf ( n311798 , n305138 );
not ( n311799 , n311798 );
or ( n311800 , n21371 , n311799 );
buf ( n311801 , n305144 );
buf ( n311802 , n20704 );
nand ( n311803 , n311801 , n311802 );
buf ( n311804 , n311803 );
buf ( n311805 , n311804 );
nand ( n311806 , n311800 , n311805 );
buf ( n311807 , n311806 );
buf ( n311808 , n311807 );
buf ( n311809 , n304655 );
not ( n311810 , n311809 );
buf ( n311811 , n306152 );
not ( n311812 , n311811 );
buf ( n311813 , n311812 );
buf ( n311814 , n311813 );
not ( n311815 , n311814 );
or ( n21390 , n311810 , n311815 );
buf ( n311817 , n890 );
nand ( n311818 , n21390 , n311817 );
buf ( n311819 , n311818 );
buf ( n311820 , n311819 );
xor ( n311821 , n311808 , n311820 );
buf ( n311822 , n15804 );
buf ( n311823 , n837 );
buf ( n311824 , n884 );
xnor ( n311825 , n311823 , n311824 );
buf ( n311826 , n311825 );
buf ( n311827 , n311826 );
or ( n21402 , n311822 , n311827 );
buf ( n311829 , n306238 );
buf ( n21404 , n311208 );
not ( n311831 , n21404 );
buf ( n311832 , n311831 );
buf ( n311833 , n311832 );
or ( n311834 , n311829 , n311833 );
nand ( n21409 , n21402 , n311834 );
buf ( n21410 , n21409 );
buf ( n311837 , n21410 );
and ( n311838 , n311821 , n311837 );
and ( n311839 , n311808 , n311820 );
or ( n21414 , n311838 , n311839 );
buf ( n311841 , n21414 );
buf ( n311842 , n311841 );
and ( n21417 , n311794 , n311842 );
and ( n21418 , n311741 , n311793 );
or ( n311845 , n21417 , n21418 );
buf ( n311846 , n311845 );
buf ( n21421 , n311846 );
xor ( n21422 , n311666 , n21421 );
xor ( n311849 , n311044 , n311094 );
xor ( n311850 , n311849 , n311174 );
buf ( n311851 , n311850 );
buf ( n311852 , n311851 );
and ( n21427 , n21422 , n311852 );
and ( n21428 , n311666 , n21421 );
or ( n311855 , n21427 , n21428 );
buf ( n311856 , n311855 );
buf ( n311857 , n311856 );
xor ( n311858 , n311588 , n311857 );
xor ( n21433 , n310980 , n311179 );
xor ( n21434 , n21433 , n311184 );
buf ( n311861 , n21434 );
buf ( n311862 , n311861 );
and ( n21437 , n311858 , n311862 );
and ( n21438 , n311588 , n311857 );
or ( n311865 , n21437 , n21438 );
buf ( n311866 , n311865 );
buf ( n311867 , n311866 );
xor ( n21442 , n311584 , n311867 );
buf ( n311869 , n21442 );
buf ( n311870 , n311869 );
xor ( n311871 , n311197 , n311221 );
xor ( n311872 , n311871 , n311260 );
buf ( n311873 , n311872 );
buf ( n311874 , n311873 );
xor ( n311875 , n311001 , n311018 );
xor ( n21450 , n311875 , n311039 );
buf ( n311877 , n21450 );
buf ( n311878 , n311877 );
xor ( n21453 , n311874 , n311878 );
buf ( n311880 , n864 );
buf ( n311881 , n858 );
and ( n311882 , n311880 , n311881 );
buf ( n311883 , n311882 );
buf ( n21458 , n311883 );
buf ( n311885 , n310568 );
buf ( n311886 , n310573 );
nor ( n311887 , n311885 , n311886 );
buf ( n311888 , n311887 );
buf ( n311889 , n311888 );
not ( n311890 , n311889 );
buf ( n311891 , n311890 );
buf ( n311892 , n311891 );
buf ( n21467 , n864 );
buf ( n311894 , n857 );
xnor ( n311895 , n21467 , n311894 );
buf ( n311896 , n311895 );
buf ( n311897 , n311896 );
or ( n311898 , n311892 , n311897 );
buf ( n311899 , n311246 );
buf ( n311900 , n311241 );
or ( n311901 , n311899 , n311900 );
nand ( n21476 , n311898 , n311901 );
buf ( n21477 , n21476 );
buf ( n311904 , n21477 );
xor ( n21479 , n21458 , n311904 );
buf ( n311906 , n304941 );
buf ( n311907 , n878 );
buf ( n311908 , n843 );
and ( n311909 , n311907 , n311908 );
not ( n21484 , n311907 );
buf ( n311911 , n305117 );
and ( n21486 , n21484 , n311911 );
nor ( n21487 , n311909 , n21486 );
buf ( n311914 , n21487 );
buf ( n311915 , n311914 );
not ( n21490 , n311915 );
buf ( n311917 , n21490 );
buf ( n311918 , n311917 );
or ( n21493 , n311906 , n311918 );
buf ( n311920 , n14523 );
buf ( n311921 , n20727 );
or ( n21496 , n311920 , n311921 );
nand ( n311923 , n21493 , n21496 );
buf ( n311924 , n311923 );
buf ( n311925 , n311924 );
and ( n21500 , n21479 , n311925 );
and ( n21501 , n21458 , n311904 );
or ( n311928 , n21500 , n21501 );
buf ( n311929 , n311928 );
buf ( n311930 , n311929 );
and ( n311931 , n21453 , n311930 );
and ( n311932 , n311874 , n311878 );
or ( n21507 , n311931 , n311932 );
buf ( n311934 , n21507 );
buf ( n311935 , n311934 );
xor ( n21510 , n311265 , n311269 );
xor ( n311937 , n21510 , n311326 );
buf ( n311938 , n311937 );
buf ( n311939 , n311938 );
xor ( n311940 , n311935 , n311939 );
xor ( n311941 , n311335 , n311379 );
xor ( n311942 , n311941 , n311384 );
buf ( n311943 , n311942 );
buf ( n311944 , n311943 );
and ( n311945 , n311940 , n311944 );
and ( n21520 , n311935 , n311939 );
or ( n311947 , n311945 , n21520 );
buf ( n311948 , n311947 );
buf ( n311949 , n311948 );
xor ( n311950 , n311331 , n311389 );
xor ( n21525 , n311950 , n311442 );
buf ( n311952 , n21525 );
buf ( n311953 , n311952 );
xor ( n21528 , n311949 , n311953 );
xor ( n311955 , n311119 , n311143 );
xor ( n311956 , n311955 , n311169 );
buf ( n311957 , n311956 );
xor ( n311958 , n311065 , n311077 );
xor ( n21533 , n311958 , n311090 );
and ( n311960 , n311957 , n21533 );
xor ( n311961 , n311602 , n311606 );
xor ( n21536 , n311961 , n311661 );
buf ( n311963 , n21536 );
xor ( n311964 , n311065 , n311077 );
xor ( n21539 , n311964 , n311090 );
and ( n21540 , n311963 , n21539 );
and ( n21541 , n311957 , n311963 );
or ( n311968 , n311960 , n21540 , n21541 );
buf ( n311969 , n311968 );
xor ( n21544 , n311666 , n21421 );
xor ( n21545 , n21544 , n311852 );
buf ( n311972 , n21545 );
buf ( n311973 , n311972 );
xor ( n21548 , n311969 , n311973 );
buf ( n311975 , n890 );
buf ( n311976 , n832 );
xor ( n21551 , n311975 , n311976 );
buf ( n311978 , n21551 );
buf ( n311979 , n311978 );
not ( n21554 , n311979 );
buf ( n311981 , n306152 );
not ( n311982 , n311981 );
or ( n21557 , n21554 , n311982 );
buf ( n311984 , n304658 );
buf ( n311985 , n890 );
nand ( n311986 , n311984 , n311985 );
buf ( n311987 , n311986 );
buf ( n311988 , n311987 );
nand ( n311989 , n21557 , n311988 );
buf ( n311990 , n311989 );
buf ( n311991 , n311990 );
xor ( n21566 , n888 , n834 );
buf ( n311993 , n21566 );
not ( n21568 , n311993 );
buf ( n311995 , n305130 );
buf ( n311996 , n305132 );
and ( n311997 , n311995 , n311996 );
buf ( n311998 , n311997 );
buf ( n311999 , n311998 );
not ( n312000 , n311999 );
or ( n21575 , n21568 , n312000 );
buf ( n312002 , n305127 );
buf ( n312003 , n21369 );
nand ( n21578 , n312002 , n312003 );
buf ( n312005 , n21578 );
buf ( n312006 , n312005 );
nand ( n21581 , n21575 , n312006 );
buf ( n312008 , n21581 );
buf ( n312009 , n312008 );
xor ( n312010 , n876 , n846 );
buf ( n312011 , n312010 );
not ( n21586 , n312011 );
buf ( n312013 , n305338 );
not ( n21588 , n312013 );
or ( n21589 , n21586 , n21588 );
buf ( n21590 , n305344 );
buf ( n312017 , n311759 );
nand ( n312018 , n21590 , n312017 );
buf ( n312019 , n312018 );
buf ( n312020 , n312019 );
nand ( n21595 , n21589 , n312020 );
buf ( n21596 , n21595 );
buf ( n312023 , n21596 );
xor ( n21598 , n312009 , n312023 );
buf ( n312025 , n884 );
buf ( n312026 , n838 );
and ( n21601 , n312025 , n312026 );
not ( n21602 , n312025 );
buf ( n312029 , n310377 );
and ( n21604 , n21602 , n312029 );
nor ( n21605 , n21601 , n21604 );
buf ( n312032 , n21605 );
buf ( n312033 , n312032 );
not ( n21608 , n312033 );
buf ( n312035 , n310401 );
not ( n21610 , n312035 );
or ( n21611 , n21608 , n21610 );
buf ( n312038 , n311826 );
not ( n21613 , n312038 );
buf ( n312040 , n304807 );
nand ( n21615 , n21613 , n312040 );
buf ( n312042 , n21615 );
buf ( n312043 , n312042 );
nand ( n21618 , n21611 , n312043 );
buf ( n312045 , n21618 );
buf ( n312046 , n312045 );
and ( n21621 , n21598 , n312046 );
and ( n21622 , n312009 , n312023 );
or ( n21623 , n21621 , n21622 );
buf ( n312050 , n21623 );
buf ( n312051 , n312050 );
xor ( n21626 , n311991 , n312051 );
buf ( n312053 , n848 );
buf ( n312054 , n874 );
xor ( n312055 , n312053 , n312054 );
buf ( n312056 , n312055 );
buf ( n312057 , n312056 );
not ( n312058 , n312057 );
buf ( n312059 , n305624 );
not ( n21634 , n312059 );
or ( n21635 , n312058 , n21634 );
buf ( n312062 , n311779 );
buf ( n312063 , n305289 );
nand ( n312064 , n312062 , n312063 );
buf ( n312065 , n312064 );
buf ( n312066 , n312065 );
nand ( n312067 , n21635 , n312066 );
buf ( n312068 , n312067 );
buf ( n312069 , n312068 );
buf ( n312070 , n882 );
buf ( n312071 , n840 );
and ( n21646 , n312070 , n312071 );
not ( n21647 , n312070 );
buf ( n21648 , n305261 );
and ( n312075 , n21647 , n21648 );
nor ( n21650 , n21646 , n312075 );
buf ( n21651 , n21650 );
buf ( n312078 , n21651 );
not ( n21653 , n312078 );
buf ( n312080 , n304584 );
not ( n312081 , n312080 );
or ( n21656 , n21653 , n312081 );
buf ( n312083 , n304596 );
buf ( n312084 , n311742 );
nand ( n312085 , n312083 , n312084 );
buf ( n312086 , n312085 );
buf ( n312087 , n312086 );
nand ( n312088 , n21656 , n312087 );
buf ( n312089 , n312088 );
buf ( n312090 , n312089 );
xor ( n312091 , n312069 , n312090 );
buf ( n312092 , n304854 );
buf ( n312093 , n872 );
buf ( n312094 , n304565 );
and ( n312095 , n312093 , n312094 );
not ( n21670 , n312093 );
buf ( n312097 , n850 );
and ( n312098 , n21670 , n312097 );
nor ( n21673 , n312095 , n312098 );
buf ( n21674 , n21673 );
buf ( n312101 , n21674 );
or ( n21676 , n312092 , n312101 );
buf ( n312103 , n14439 );
buf ( n312104 , n311717 );
not ( n21679 , n312104 );
buf ( n312106 , n21679 );
buf ( n312107 , n312106 );
or ( n312108 , n312103 , n312107 );
nand ( n21683 , n21676 , n312108 );
buf ( n21684 , n21683 );
buf ( n312111 , n21684 );
and ( n21686 , n312091 , n312111 );
and ( n312113 , n312069 , n312090 );
or ( n21688 , n21686 , n312113 );
buf ( n312115 , n21688 );
buf ( n312116 , n312115 );
and ( n312117 , n21626 , n312116 );
and ( n21692 , n311991 , n312051 );
or ( n312119 , n312117 , n21692 );
buf ( n312120 , n312119 );
buf ( n312121 , n312120 );
xor ( n312122 , n868 , n854 );
buf ( n312123 , n312122 );
not ( n21698 , n312123 );
buf ( n312125 , n305205 );
buf ( n312126 , n305207 );
and ( n21701 , n312125 , n312126 );
buf ( n21702 , n21701 );
buf ( n312129 , n21702 );
not ( n21704 , n312129 );
or ( n21705 , n21698 , n21704 );
buf ( n312132 , n305219 );
buf ( n312133 , n311645 );
nand ( n312134 , n312132 , n312133 );
buf ( n312135 , n312134 );
buf ( n312136 , n312135 );
nand ( n312137 , n21705 , n312136 );
buf ( n312138 , n312137 );
xor ( n21713 , n866 , n856 );
buf ( n312140 , n21713 );
not ( n21715 , n312140 );
buf ( n312142 , n310477 );
not ( n312143 , n312142 );
or ( n21718 , n21715 , n312143 );
buf ( n312145 , n310472 );
not ( n21720 , n312145 );
buf ( n312147 , n21182 );
nand ( n312148 , n21720 , n312147 );
buf ( n312149 , n312148 );
buf ( n312150 , n312149 );
nand ( n312151 , n21718 , n312150 );
buf ( n312152 , n312151 );
or ( n312153 , n312138 , n312152 );
not ( n312154 , n312153 );
buf ( n312155 , n878 );
buf ( n312156 , n844 );
and ( n312157 , n312155 , n312156 );
not ( n21732 , n312155 );
buf ( n312159 , n305458 );
and ( n21734 , n21732 , n312159 );
nor ( n21735 , n312157 , n21734 );
buf ( n312162 , n21735 );
buf ( n312163 , n312162 );
not ( n21738 , n312163 );
buf ( n312165 , n15836 );
not ( n21740 , n312165 );
or ( n312167 , n21738 , n21740 );
buf ( n312168 , n306272 );
buf ( n312169 , n311914 );
nand ( n312170 , n312168 , n312169 );
buf ( n312171 , n312170 );
buf ( n312172 , n312171 );
nand ( n21747 , n312167 , n312172 );
buf ( n312174 , n21747 );
not ( n21749 , n312174 );
or ( n312176 , n312154 , n21749 );
nand ( n312177 , n312138 , n312152 );
nand ( n21752 , n312176 , n312177 );
xor ( n312179 , n311755 , n311772 );
xor ( n21754 , n312179 , n311788 );
buf ( n312181 , n21754 );
xor ( n21756 , n21752 , n312181 );
buf ( n312183 , n870 );
buf ( n21758 , n852 );
and ( n21759 , n312183 , n21758 );
not ( n312186 , n312183 );
buf ( n312187 , n305168 );
and ( n21762 , n312186 , n312187 );
nor ( n21763 , n21759 , n21762 );
buf ( n312190 , n21763 );
buf ( n312191 , n312190 );
not ( n312192 , n312191 );
buf ( n312193 , n14323 );
not ( n21768 , n312193 );
or ( n312195 , n312192 , n21768 );
buf ( n312196 , n311052 );
buf ( n312197 , n311667 );
nand ( n21772 , n312196 , n312197 );
buf ( n312199 , n21772 );
buf ( n312200 , n312199 );
nand ( n312201 , n312195 , n312200 );
buf ( n312202 , n312201 );
buf ( n312203 , n312202 );
buf ( n312204 , n886 );
buf ( n312205 , n836 );
xor ( n312206 , n312204 , n312205 );
buf ( n312207 , n312206 );
buf ( n312208 , n312207 );
not ( n312209 , n312208 );
buf ( n312210 , n304912 );
not ( n21785 , n312210 );
or ( n312212 , n312209 , n21785 );
buf ( n312213 , n304901 );
buf ( n312214 , n311691 );
nand ( n312215 , n312213 , n312214 );
buf ( n312216 , n312215 );
buf ( n312217 , n312216 );
nand ( n21792 , n312212 , n312217 );
buf ( n312219 , n21792 );
buf ( n312220 , n312219 );
xor ( n312221 , n312203 , n312220 );
buf ( n21796 , n304987 );
buf ( n312223 , n842 );
buf ( n312224 , n880 );
not ( n21799 , n312224 );
buf ( n21800 , n21799 );
buf ( n312227 , n21800 );
and ( n21802 , n312223 , n312227 );
not ( n312229 , n312223 );
buf ( n312230 , n880 );
and ( n21805 , n312229 , n312230 );
nor ( n312232 , n21802 , n21805 );
buf ( n312233 , n312232 );
buf ( n312234 , n312233 );
or ( n312235 , n21796 , n312234 );
buf ( n21810 , n311075 );
buf ( n312237 , n311629 );
not ( n312238 , n312237 );
buf ( n312239 , n312238 );
buf ( n312240 , n312239 );
or ( n312241 , n21810 , n312240 );
nand ( n21816 , n312235 , n312241 );
buf ( n312243 , n21816 );
buf ( n312244 , n312243 );
and ( n21819 , n312221 , n312244 );
and ( n21820 , n312203 , n312220 );
or ( n312247 , n21819 , n21820 );
buf ( n312248 , n312247 );
and ( n21823 , n21756 , n312248 );
and ( n312250 , n21752 , n312181 );
or ( n312251 , n21823 , n312250 );
buf ( n312252 , n312251 );
xor ( n312253 , n312121 , n312252 );
xor ( n312254 , n311741 , n311793 );
xor ( n21829 , n312254 , n311842 );
buf ( n312256 , n21829 );
buf ( n312257 , n312256 );
and ( n312258 , n312253 , n312257 );
and ( n21833 , n312121 , n312252 );
or ( n312260 , n312258 , n21833 );
buf ( n312261 , n312260 );
buf ( n312262 , n312261 );
and ( n312263 , n21548 , n312262 );
and ( n312264 , n311969 , n311973 );
or ( n21839 , n312263 , n312264 );
buf ( n312266 , n21839 );
buf ( n312267 , n312266 );
and ( n21842 , n21528 , n312267 );
and ( n312269 , n311949 , n311953 );
or ( n312270 , n21842 , n312269 );
buf ( n312271 , n312270 );
buf ( n312272 , n312271 );
xor ( n312273 , n311192 , n311870 );
xor ( n21848 , n312273 , n312272 );
buf ( n312275 , n21848 );
xor ( n312276 , n311192 , n311870 );
and ( n21851 , n312276 , n312272 );
and ( n312278 , n311192 , n311870 );
or ( n312279 , n21851 , n312278 );
buf ( n312280 , n312279 );
buf ( n312281 , n310582 );
buf ( n312282 , n863 );
and ( n21857 , n312281 , n312282 );
buf ( n312284 , n21857 );
buf ( n312285 , n312284 );
buf ( n312286 , n834 );
buf ( n312287 , n894 );
xor ( n21862 , n312286 , n312287 );
buf ( n312289 , n21862 );
buf ( n312290 , n312289 );
not ( n21865 , n312290 );
buf ( n312292 , n305032 );
not ( n312293 , n312292 );
or ( n21868 , n21865 , n312293 );
buf ( n312295 , n833 );
buf ( n312296 , n894 );
xor ( n21871 , n312295 , n312296 );
buf ( n312298 , n21871 );
buf ( n312299 , n312298 );
buf ( n312300 , n895 );
nand ( n21875 , n312299 , n312300 );
buf ( n312302 , n21875 );
buf ( n312303 , n312302 );
nand ( n312304 , n21868 , n312303 );
buf ( n312305 , n312304 );
buf ( n312306 , n312305 );
xor ( n312307 , n312285 , n312306 );
buf ( n312308 , n836 );
buf ( n312309 , n892 );
xor ( n312310 , n312308 , n312309 );
buf ( n312311 , n312310 );
buf ( n312312 , n312311 );
not ( n21887 , n312312 );
buf ( n312314 , n14272 );
not ( n21889 , n312314 );
or ( n312316 , n21887 , n21889 );
buf ( n312317 , n892 );
buf ( n312318 , n835 );
xor ( n312319 , n312317 , n312318 );
buf ( n312320 , n312319 );
buf ( n312321 , n312320 );
buf ( n312322 , n304694 );
nand ( n312323 , n312321 , n312322 );
buf ( n312324 , n312323 );
buf ( n312325 , n312324 );
nand ( n21900 , n312316 , n312325 );
buf ( n312327 , n21900 );
buf ( n312328 , n312327 );
xor ( n312329 , n312307 , n312328 );
buf ( n312330 , n312329 );
buf ( n312331 , n312330 );
buf ( n312332 , n858 );
buf ( n312333 , n870 );
xor ( n312334 , n312332 , n312333 );
buf ( n312335 , n312334 );
buf ( n312336 , n312335 );
not ( n312337 , n312336 );
buf ( n312338 , n20629 );
not ( n21913 , n312338 );
or ( n312340 , n312337 , n21913 );
buf ( n312341 , n311052 );
buf ( n312342 , n857 );
buf ( n312343 , n870 );
xor ( n312344 , n312342 , n312343 );
buf ( n312345 , n312344 );
buf ( n312346 , n312345 );
nand ( n21921 , n312341 , n312346 );
buf ( n312348 , n21921 );
buf ( n312349 , n312348 );
nand ( n21924 , n312340 , n312349 );
buf ( n312351 , n21924 );
buf ( n312352 , n312351 );
xor ( n312353 , n868 , n860 );
buf ( n312354 , n312353 );
not ( n312355 , n312354 );
buf ( n312356 , n21702 );
not ( n312357 , n312356 );
or ( n312358 , n312355 , n312357 );
buf ( n312359 , n305219 );
xor ( n312360 , n868 , n859 );
buf ( n312361 , n312360 );
nand ( n21936 , n312359 , n312361 );
buf ( n312363 , n21936 );
buf ( n312364 , n312363 );
nand ( n312365 , n312358 , n312364 );
buf ( n312366 , n312365 );
buf ( n312367 , n312366 );
xor ( n312368 , n312352 , n312367 );
xor ( n21943 , n882 , n846 );
buf ( n312370 , n21943 );
not ( n312371 , n312370 );
buf ( n312372 , n304584 );
not ( n312373 , n312372 );
or ( n312374 , n312371 , n312373 );
buf ( n312375 , n304596 );
buf ( n312376 , n845 );
buf ( n312377 , n882 );
and ( n21952 , n312376 , n312377 );
not ( n312379 , n312376 );
buf ( n312380 , n305526 );
and ( n21955 , n312379 , n312380 );
nor ( n312382 , n21952 , n21955 );
buf ( n312383 , n312382 );
buf ( n312384 , n312383 );
nand ( n312385 , n312375 , n312384 );
buf ( n312386 , n312385 );
buf ( n312387 , n312386 );
nand ( n21962 , n312374 , n312387 );
buf ( n312389 , n21962 );
buf ( n312390 , n312389 );
xor ( n312391 , n312368 , n312390 );
buf ( n312392 , n312391 );
buf ( n312393 , n312392 );
xor ( n312394 , n312331 , n312393 );
buf ( n312395 , n872 );
buf ( n312396 , n856 );
and ( n312397 , n312395 , n312396 );
not ( n21972 , n312395 );
buf ( n312399 , n15582 );
and ( n21974 , n21972 , n312399 );
nor ( n21975 , n312397 , n21974 );
buf ( n312402 , n21975 );
buf ( n312403 , n312402 );
not ( n312404 , n312403 );
buf ( n312405 , n14420 );
not ( n312406 , n312405 );
or ( n312407 , n312404 , n312406 );
buf ( n312408 , n304864 );
xor ( n312409 , n872 , n855 );
buf ( n312410 , n312409 );
nand ( n21985 , n312408 , n312410 );
buf ( n312412 , n21985 );
buf ( n312413 , n312412 );
nand ( n21988 , n312407 , n312413 );
buf ( n312415 , n21988 );
buf ( n312416 , n312415 );
buf ( n312417 , n884 );
buf ( n312418 , n844 );
and ( n21993 , n312417 , n312418 );
not ( n21994 , n312417 );
buf ( n21995 , n305458 );
and ( n312422 , n21994 , n21995 );
nor ( n21997 , n21993 , n312422 );
buf ( n21998 , n21997 );
buf ( n312425 , n21998 );
not ( n22000 , n312425 );
buf ( n312427 , n304810 );
not ( n312428 , n312427 );
or ( n22003 , n22000 , n312428 );
buf ( n312430 , n304807 );
buf ( n312431 , n884 );
buf ( n312432 , n843 );
and ( n312433 , n312431 , n312432 );
not ( n312434 , n312431 );
buf ( n312435 , n305117 );
and ( n312436 , n312434 , n312435 );
nor ( n22011 , n312433 , n312436 );
buf ( n22012 , n22011 );
buf ( n312439 , n22012 );
nand ( n22014 , n312430 , n312439 );
buf ( n312441 , n22014 );
buf ( n312442 , n312441 );
nand ( n312443 , n22003 , n312442 );
buf ( n312444 , n312443 );
buf ( n312445 , n312444 );
xor ( n312446 , n312416 , n312445 );
buf ( n312447 , n304630 );
buf ( n312448 , n890 );
not ( n22023 , n312448 );
buf ( n312450 , n838 );
nor ( n312451 , n22023 , n312450 );
buf ( n312452 , n312451 );
buf ( n312453 , n312452 );
buf ( n312454 , n838 );
not ( n312455 , n312454 );
buf ( n312456 , n890 );
nor ( n312457 , n312455 , n312456 );
buf ( n312458 , n312457 );
buf ( n312459 , n312458 );
nor ( n312460 , n312453 , n312459 );
buf ( n312461 , n312460 );
buf ( n312462 , n312461 );
or ( n312463 , n312447 , n312462 );
buf ( n312464 , n837 );
buf ( n312465 , n890 );
not ( n22040 , n312465 );
buf ( n312467 , n22040 );
buf ( n312468 , n312467 );
and ( n22043 , n312464 , n312468 );
not ( n22044 , n312464 );
buf ( n312471 , n890 );
and ( n312472 , n22044 , n312471 );
nor ( n22047 , n22043 , n312472 );
buf ( n312474 , n22047 );
buf ( n312475 , n312474 );
buf ( n312476 , n304655 );
or ( n22051 , n312475 , n312476 );
nand ( n22052 , n312463 , n22051 );
buf ( n312479 , n22052 );
buf ( n312480 , n312479 );
xor ( n22055 , n312446 , n312480 );
buf ( n312482 , n22055 );
buf ( n312483 , n312482 );
xor ( n22058 , n312394 , n312483 );
buf ( n312485 , n22058 );
buf ( n312486 , n312485 );
buf ( n312487 , n866 );
buf ( n312488 , n863 );
and ( n22063 , n312487 , n312488 );
not ( n312490 , n312487 );
buf ( n312491 , n305192 );
and ( n22066 , n312490 , n312491 );
nor ( n22067 , n22063 , n22066 );
buf ( n312494 , n22067 );
buf ( n312495 , n312494 );
not ( n22070 , n312495 );
buf ( n312497 , n310694 );
not ( n22072 , n312497 );
or ( n22073 , n22070 , n22072 );
buf ( n312500 , n310483 );
buf ( n312501 , n866 );
buf ( n312502 , n862 );
xor ( n312503 , n312501 , n312502 );
buf ( n312504 , n312503 );
buf ( n312505 , n312504 );
nand ( n22080 , n312500 , n312505 );
buf ( n312507 , n22080 );
buf ( n22082 , n312507 );
nand ( n22083 , n22073 , n22082 );
buf ( n22084 , n22083 );
buf ( n22085 , n22084 );
buf ( n312512 , n867 );
buf ( n312513 , n863 );
or ( n22088 , n312512 , n312513 );
buf ( n312515 , n868 );
nand ( n22090 , n22088 , n312515 );
buf ( n22091 , n22090 );
buf ( n312518 , n22091 );
buf ( n312519 , n863 );
buf ( n312520 , n867 );
nand ( n22095 , n312519 , n312520 );
buf ( n312522 , n22095 );
buf ( n312523 , n312522 );
buf ( n312524 , n866 );
and ( n22099 , n312518 , n312523 , n312524 );
buf ( n312526 , n22099 );
buf ( n312527 , n312526 );
buf ( n312528 , n835 );
buf ( n312529 , n894 );
xor ( n312530 , n312528 , n312529 );
buf ( n312531 , n312530 );
buf ( n312532 , n312531 );
not ( n312533 , n312532 );
buf ( n312534 , n305032 );
not ( n312535 , n312534 );
or ( n312536 , n312533 , n312535 );
buf ( n312537 , n312289 );
buf ( n312538 , n895 );
nand ( n312539 , n312537 , n312538 );
buf ( n312540 , n312539 );
buf ( n312541 , n312540 );
nand ( n22116 , n312536 , n312541 );
buf ( n312543 , n22116 );
buf ( n312544 , n312543 );
xor ( n22119 , n312527 , n312544 );
buf ( n312546 , n22119 );
buf ( n312547 , n312546 );
xor ( n22122 , n22085 , n312547 );
buf ( n312549 , n310726 );
buf ( n312550 , n861 );
buf ( n312551 , n868 );
xor ( n22126 , n312550 , n312551 );
buf ( n312553 , n22126 );
buf ( n312554 , n312553 );
not ( n312555 , n312554 );
buf ( n312556 , n312555 );
buf ( n312557 , n312556 );
or ( n22132 , n312549 , n312557 );
buf ( n312559 , n305449 );
buf ( n22134 , n312353 );
not ( n312561 , n22134 );
buf ( n312562 , n312561 );
buf ( n312563 , n312562 );
or ( n22138 , n312559 , n312563 );
nand ( n22139 , n22132 , n22138 );
buf ( n312566 , n22139 );
buf ( n312567 , n312566 );
xor ( n312568 , n22122 , n312567 );
buf ( n312569 , n312568 );
buf ( n312570 , n312569 );
buf ( n312571 , n14918 );
not ( n22146 , n312571 );
buf ( n312573 , n305338 );
not ( n312574 , n312573 );
or ( n22149 , n22146 , n312574 );
buf ( n312576 , n305344 );
buf ( n312577 , n876 );
buf ( n312578 , n853 );
xor ( n22153 , n312577 , n312578 );
buf ( n312580 , n22153 );
buf ( n312581 , n312580 );
nand ( n312582 , n312576 , n312581 );
buf ( n312583 , n312582 );
buf ( n312584 , n312583 );
nand ( n312585 , n22149 , n312584 );
buf ( n312586 , n312585 );
buf ( n312587 , n305039 );
not ( n22162 , n312587 );
buf ( n312589 , n305032 );
not ( n22164 , n312589 );
or ( n312591 , n22162 , n22164 );
buf ( n22166 , n312531 );
buf ( n312593 , n895 );
nand ( n22168 , n22166 , n312593 );
buf ( n312595 , n22168 );
buf ( n312596 , n312595 );
nand ( n22171 , n312591 , n312596 );
buf ( n312598 , n22171 );
xor ( n22173 , n312586 , n312598 );
buf ( n312600 , n305306 );
not ( n312601 , n312600 );
buf ( n312602 , n305627 );
not ( n22177 , n312602 );
or ( n312604 , n312601 , n22177 );
buf ( n312605 , n305289 );
buf ( n312606 , n874 );
buf ( n312607 , n855 );
xor ( n312608 , n312606 , n312607 );
buf ( n312609 , n312608 );
buf ( n312610 , n312609 );
nand ( n312611 , n312605 , n312610 );
buf ( n312612 , n312611 );
buf ( n312613 , n312612 );
nand ( n312614 , n312604 , n312613 );
buf ( n312615 , n312614 );
xnor ( n22190 , n22173 , n312615 );
buf ( n312617 , n22190 );
not ( n312618 , n312617 );
buf ( n312619 , n312618 );
buf ( n22194 , n312619 );
not ( n22195 , n22194 );
buf ( n312622 , n311107 );
buf ( n312623 , n863 );
and ( n22198 , n312622 , n312623 );
buf ( n312625 , n22198 );
buf ( n22200 , n312625 );
buf ( n312627 , n305435 );
not ( n22202 , n312627 );
buf ( n312629 , n14272 );
not ( n312630 , n312629 );
or ( n22205 , n22202 , n312630 );
buf ( n312632 , n892 );
buf ( n312633 , n837 );
xor ( n22208 , n312632 , n312633 );
buf ( n22209 , n22208 );
buf ( n312636 , n22209 );
buf ( n312637 , n304694 );
nand ( n312638 , n312636 , n312637 );
buf ( n312639 , n312638 );
buf ( n312640 , n312639 );
nand ( n22215 , n22205 , n312640 );
buf ( n312642 , n22215 );
buf ( n312643 , n312642 );
xor ( n312644 , n22200 , n312643 );
buf ( n312645 , n305149 );
not ( n22220 , n312645 );
buf ( n312647 , n305138 );
not ( n22222 , n312647 );
or ( n312649 , n22220 , n22222 );
buf ( n22224 , n305144 );
buf ( n312651 , n841 );
buf ( n312652 , n888 );
xor ( n312653 , n312651 , n312652 );
buf ( n312654 , n312653 );
buf ( n312655 , n312654 );
nand ( n312656 , n22224 , n312655 );
buf ( n312657 , n312656 );
buf ( n312658 , n312657 );
nand ( n312659 , n312649 , n312658 );
buf ( n312660 , n312659 );
buf ( n312661 , n312660 );
xnor ( n312662 , n312644 , n312661 );
buf ( n312663 , n312662 );
buf ( n312664 , n312663 );
not ( n312665 , n312664 );
buf ( n312666 , n312665 );
buf ( n312667 , n312666 );
not ( n22242 , n312667 );
or ( n312669 , n22195 , n22242 );
not ( n312670 , n312663 );
not ( n312671 , n22190 );
or ( n22246 , n312670 , n312671 );
buf ( n312673 , n14793 );
not ( n312674 , n312673 );
buf ( n312675 , n21702 );
not ( n312676 , n312675 );
or ( n312677 , n312674 , n312676 );
buf ( n312678 , n305202 );
buf ( n312679 , n312553 );
nand ( n312680 , n312678 , n312679 );
buf ( n312681 , n312680 );
buf ( n312682 , n312681 );
nand ( n22257 , n312677 , n312682 );
buf ( n312684 , n22257 );
buf ( n312685 , n312684 );
buf ( n312686 , n14961 );
not ( n22261 , n312686 );
buf ( n312688 , n304584 );
not ( n22263 , n312688 );
or ( n312690 , n22261 , n22263 );
buf ( n312691 , n304596 );
buf ( n312692 , n882 );
buf ( n312693 , n847 );
xor ( n312694 , n312692 , n312693 );
buf ( n312695 , n312694 );
buf ( n312696 , n312695 );
nand ( n22271 , n312691 , n312696 );
buf ( n312698 , n22271 );
buf ( n312699 , n312698 );
nand ( n312700 , n312690 , n312699 );
buf ( n312701 , n312700 );
buf ( n312702 , n312701 );
xor ( n312703 , n312685 , n312702 );
buf ( n312704 , n311813 );
buf ( n312705 , n305268 );
or ( n312706 , n312704 , n312705 );
buf ( n312707 , n304655 );
buf ( n312708 , n890 );
buf ( n312709 , n839 );
xor ( n22284 , n312708 , n312709 );
buf ( n312711 , n22284 );
buf ( n312712 , n312711 );
not ( n22287 , n312712 );
buf ( n312714 , n22287 );
buf ( n312715 , n312714 );
or ( n312716 , n312707 , n312715 );
nand ( n22291 , n312706 , n312716 );
buf ( n22292 , n22291 );
buf ( n312719 , n22292 );
xor ( n22294 , n312703 , n312719 );
buf ( n312721 , n22294 );
nand ( n22296 , n22246 , n312721 );
buf ( n312723 , n22296 );
nand ( n22298 , n312669 , n312723 );
buf ( n312725 , n22298 );
buf ( n312726 , n312725 );
xor ( n22301 , n312570 , n312726 );
and ( n22302 , n305413 , n305442 );
buf ( n312729 , n22302 );
buf ( n312730 , n312729 );
xor ( n22305 , n305110 , n305156 );
and ( n312732 , n22305 , n305180 );
and ( n312733 , n305110 , n305156 );
or ( n312734 , n312732 , n312733 );
buf ( n312735 , n312734 );
buf ( n312736 , n312735 );
xor ( n312737 , n312730 , n312736 );
xor ( n22312 , n305312 , n305352 );
and ( n312739 , n22312 , n14944 );
and ( n22314 , n305312 , n305352 );
or ( n22315 , n312739 , n22314 );
buf ( n312742 , n22315 );
and ( n312743 , n312737 , n312742 );
and ( n22318 , n312730 , n312736 );
or ( n312745 , n312743 , n22318 );
buf ( n312746 , n312745 );
buf ( n312747 , n312746 );
and ( n312748 , n22301 , n312747 );
and ( n22323 , n312570 , n312726 );
or ( n312750 , n312748 , n22323 );
buf ( n312751 , n312750 );
buf ( n312752 , n312751 );
xor ( n312753 , n312486 , n312752 );
buf ( n312754 , n305245 );
not ( n312755 , n312754 );
buf ( n312756 , n14323 );
not ( n312757 , n312756 );
or ( n22332 , n312755 , n312757 );
buf ( n312759 , n304763 );
xor ( n312760 , n870 , n859 );
buf ( n312761 , n312760 );
nand ( n22336 , n312759 , n312761 );
buf ( n312763 , n22336 );
buf ( n312764 , n312763 );
nand ( n312765 , n22332 , n312764 );
buf ( n312766 , n312765 );
buf ( n312767 , n305082 );
not ( n22342 , n312767 );
buf ( n312769 , n304813 );
not ( n312770 , n312769 );
or ( n312771 , n22342 , n312770 );
buf ( n312772 , n304819 );
buf ( n312773 , n884 );
buf ( n22348 , n845 );
xor ( n22349 , n312773 , n22348 );
buf ( n22350 , n22349 );
buf ( n312777 , n22350 );
nand ( n312778 , n312772 , n312777 );
buf ( n312779 , n312778 );
buf ( n312780 , n312779 );
nand ( n22355 , n312771 , n312780 );
buf ( n312782 , n22355 );
xor ( n22357 , n312766 , n312782 );
buf ( n312784 , n305064 );
not ( n312785 , n312784 );
buf ( n312786 , n306132 );
not ( n312787 , n312786 );
or ( n22362 , n312785 , n312787 );
buf ( n312789 , n304864 );
buf ( n312790 , n872 );
buf ( n312791 , n857 );
and ( n312792 , n312790 , n312791 );
not ( n312793 , n312790 );
buf ( n312794 , n305939 );
and ( n312795 , n312793 , n312794 );
nor ( n312796 , n312792 , n312795 );
buf ( n312797 , n312796 );
buf ( n312798 , n312797 );
nand ( n312799 , n312789 , n312798 );
buf ( n312800 , n312799 );
buf ( n312801 , n312800 );
nand ( n312802 , n22362 , n312801 );
buf ( n312803 , n312802 );
and ( n312804 , n22357 , n312803 );
and ( n22379 , n312766 , n312782 );
or ( n312806 , n312804 , n22379 );
buf ( n312807 , n312806 );
xor ( n22382 , n312685 , n312702 );
and ( n312809 , n22382 , n312719 );
and ( n312810 , n312685 , n312702 );
or ( n312811 , n312809 , n312810 );
buf ( n312812 , n312811 );
buf ( n312813 , n312812 );
xor ( n22388 , n312807 , n312813 );
buf ( n312815 , n22209 );
not ( n312816 , n312815 );
buf ( n312817 , n304697 );
not ( n22392 , n312817 );
or ( n312819 , n312816 , n22392 );
buf ( n22394 , n312311 );
buf ( n22395 , n304694 );
nand ( n22396 , n22394 , n22395 );
buf ( n22397 , n22396 );
buf ( n22398 , n22397 );
nand ( n22399 , n312819 , n22398 );
buf ( n22400 , n22399 );
buf ( n22401 , n22400 );
buf ( n312828 , n312654 );
not ( n312829 , n312828 );
buf ( n312830 , n311998 );
not ( n22405 , n312830 );
or ( n22406 , n312829 , n22405 );
buf ( n22407 , n305144 );
buf ( n312834 , n888 );
buf ( n312835 , n840 );
xor ( n312836 , n312834 , n312835 );
buf ( n312837 , n312836 );
buf ( n312838 , n312837 );
nand ( n22413 , n22407 , n312838 );
buf ( n312840 , n22413 );
buf ( n312841 , n312840 );
nand ( n312842 , n22406 , n312841 );
buf ( n312843 , n312842 );
buf ( n312844 , n312843 );
xor ( n22419 , n22401 , n312844 );
buf ( n312846 , n880 );
buf ( n22421 , n849 );
and ( n22422 , n312846 , n22421 );
not ( n22423 , n312846 );
buf ( n312850 , n305596 );
and ( n22425 , n22423 , n312850 );
nor ( n22426 , n22422 , n22425 );
buf ( n312853 , n22426 );
buf ( n312854 , n312853 );
not ( n312855 , n312854 );
buf ( n312856 , n304984 );
not ( n22431 , n312856 );
or ( n312858 , n312855 , n22431 );
buf ( n312859 , n304997 );
xor ( n22434 , n880 , n848 );
buf ( n312861 , n22434 );
nand ( n312862 , n312859 , n312861 );
buf ( n312863 , n312862 );
buf ( n312864 , n312863 );
nand ( n312865 , n312858 , n312864 );
buf ( n312866 , n312865 );
buf ( n312867 , n312866 );
xor ( n312868 , n22419 , n312867 );
buf ( n312869 , n312868 );
buf ( n312870 , n312869 );
xor ( n312871 , n22388 , n312870 );
buf ( n312872 , n312871 );
buf ( n312873 , n312872 );
buf ( n312874 , n312615 );
buf ( n312875 , n312598 );
or ( n22450 , n312874 , n312875 );
buf ( n312877 , n312586 );
nand ( n312878 , n22450 , n312877 );
buf ( n312879 , n312878 );
buf ( n312880 , n312879 );
buf ( n312881 , n312615 );
buf ( n312882 , n312598 );
nand ( n22457 , n312881 , n312882 );
buf ( n312884 , n22457 );
buf ( n312885 , n312884 );
nand ( n22460 , n312880 , n312885 );
buf ( n312887 , n22460 );
buf ( n312888 , n312887 );
buf ( n312889 , n305172 );
not ( n312890 , n312889 );
buf ( n312891 , n15836 );
not ( n22466 , n312891 );
or ( n312893 , n312890 , n22466 );
buf ( n312894 , n306272 );
buf ( n312895 , n878 );
buf ( n312896 , n851 );
and ( n312897 , n312895 , n312896 );
not ( n22472 , n312895 );
buf ( n312899 , n305532 );
and ( n312900 , n22472 , n312899 );
nor ( n22475 , n312897 , n312900 );
buf ( n312902 , n22475 );
buf ( n312903 , n312902 );
nand ( n312904 , n312894 , n312903 );
buf ( n312905 , n312904 );
buf ( n312906 , n312905 );
nand ( n22481 , n312893 , n312906 );
buf ( n312908 , n22481 );
buf ( n22483 , n312908 );
buf ( n312910 , n305368 );
not ( n22485 , n312910 );
buf ( n22486 , n22485 );
buf ( n312913 , n22486 );
not ( n22488 , n312913 );
buf ( n312915 , n304912 );
not ( n22490 , n312915 );
or ( n312917 , n22488 , n22490 );
buf ( n312918 , n304901 );
and ( n22493 , n886 , n305117 );
not ( n312920 , n886 );
and ( n22495 , n312920 , n843 );
or ( n312922 , n22493 , n22495 );
buf ( n312923 , n312922 );
nand ( n22498 , n312918 , n312923 );
buf ( n22499 , n22498 );
buf ( n312926 , n22499 );
nand ( n22501 , n312917 , n312926 );
buf ( n312928 , n22501 );
buf ( n312929 , n312928 );
xor ( n22504 , n22483 , n312929 );
buf ( n312931 , n305103 );
not ( n22506 , n312931 );
buf ( n312933 , n304984 );
not ( n22508 , n312933 );
or ( n22509 , n22506 , n22508 );
buf ( n312936 , n304997 );
buf ( n312937 , n312853 );
nand ( n22512 , n312936 , n312937 );
buf ( n312939 , n22512 );
buf ( n22514 , n312939 );
nand ( n22515 , n22509 , n22514 );
buf ( n22516 , n22515 );
buf ( n312943 , n22516 );
and ( n312944 , n22504 , n312943 );
and ( n22519 , n22483 , n312929 );
or ( n312946 , n312944 , n22519 );
buf ( n312947 , n312946 );
buf ( n312948 , n312947 );
xor ( n312949 , n312888 , n312948 );
buf ( n312950 , n312625 );
not ( n312951 , n312950 );
buf ( n312952 , n312660 );
not ( n312953 , n312952 );
or ( n22528 , n312951 , n312953 );
buf ( n312955 , n312660 );
buf ( n312956 , n312625 );
or ( n312957 , n312955 , n312956 );
buf ( n312958 , n312642 );
nand ( n312959 , n312957 , n312958 );
buf ( n312960 , n312959 );
buf ( n312961 , n312960 );
nand ( n312962 , n22528 , n312961 );
buf ( n312963 , n312962 );
buf ( n312964 , n312963 );
xor ( n22539 , n312949 , n312964 );
buf ( n312966 , n22539 );
buf ( n22541 , n312966 );
xor ( n22542 , n312873 , n22541 );
xor ( n312969 , n305047 , n305071 );
and ( n312970 , n312969 , n305089 );
and ( n22545 , n305047 , n305071 );
or ( n22546 , n312970 , n22545 );
buf ( n312973 , n22546 );
buf ( n312974 , n312973 );
xor ( n22549 , n305228 , n305252 );
and ( n22550 , n22549 , n305273 );
and ( n22551 , n305228 , n305252 );
or ( n22552 , n22550 , n22551 );
buf ( n312979 , n22552 );
buf ( n312980 , n312979 );
xor ( n312981 , n312974 , n312980 );
xor ( n22556 , n22483 , n312929 );
xor ( n22557 , n22556 , n312943 );
buf ( n312984 , n22557 );
buf ( n312985 , n312984 );
and ( n22560 , n312981 , n312985 );
and ( n22561 , n312974 , n312980 );
or ( n22562 , n22560 , n22561 );
buf ( n312989 , n22562 );
buf ( n312990 , n312989 );
and ( n22565 , n22542 , n312990 );
and ( n22566 , n312873 , n22541 );
or ( n22567 , n22565 , n22566 );
buf ( n312994 , n22567 );
buf ( n312995 , n312994 );
xor ( n22570 , n312753 , n312995 );
buf ( n312997 , n22570 );
buf ( n312998 , n312997 );
xor ( n22573 , n312570 , n312726 );
xor ( n313000 , n22573 , n312747 );
buf ( n313001 , n313000 );
buf ( n313002 , n313001 );
xor ( n22577 , n312873 , n22541 );
xor ( n22578 , n22577 , n312990 );
buf ( n313005 , n22578 );
buf ( n22580 , n313005 );
xor ( n22581 , n313002 , n22580 );
buf ( n313008 , n312922 );
not ( n313009 , n313008 );
buf ( n313010 , n311697 );
not ( n313011 , n313010 );
or ( n22586 , n313009 , n313011 );
buf ( n22587 , n304901 );
buf ( n313014 , n842 );
buf ( n313015 , n886 );
xor ( n313016 , n313014 , n313015 );
buf ( n313017 , n313016 );
buf ( n313018 , n313017 );
nand ( n313019 , n22587 , n313018 );
buf ( n313020 , n313019 );
buf ( n313021 , n313020 );
nand ( n313022 , n22586 , n313021 );
buf ( n313023 , n313022 );
buf ( n313024 , n313023 );
buf ( n313025 , n312902 );
not ( n313026 , n313025 );
buf ( n313027 , n304938 );
not ( n313028 , n313027 );
buf ( n313029 , n313028 );
buf ( n313030 , n313029 );
not ( n313031 , n313030 );
or ( n313032 , n313026 , n313031 );
buf ( n313033 , n850 );
buf ( n313034 , n878 );
xor ( n313035 , n313033 , n313034 );
buf ( n313036 , n313035 );
buf ( n313037 , n313036 );
buf ( n313038 , n304932 );
nand ( n22613 , n313037 , n313038 );
buf ( n313040 , n22613 );
buf ( n313041 , n313040 );
nand ( n22616 , n313032 , n313041 );
buf ( n313043 , n22616 );
buf ( n22618 , n313043 );
xor ( n22619 , n313024 , n22618 );
buf ( n313046 , n312580 );
not ( n313047 , n313046 );
buf ( n313048 , n305338 );
not ( n313049 , n313048 );
or ( n313050 , n313047 , n313049 );
buf ( n313051 , n305344 );
buf ( n313052 , n876 );
buf ( n313053 , n852 );
xor ( n313054 , n313052 , n313053 );
buf ( n313055 , n313054 );
buf ( n313056 , n313055 );
nand ( n313057 , n313051 , n313056 );
buf ( n313058 , n313057 );
buf ( n313059 , n313058 );
nand ( n313060 , n313050 , n313059 );
buf ( n313061 , n313060 );
buf ( n313062 , n313061 );
xor ( n313063 , n22619 , n313062 );
buf ( n313064 , n313063 );
buf ( n313065 , n313064 );
buf ( n313066 , n312609 );
not ( n313067 , n313066 );
buf ( n313068 , n305292 );
not ( n313069 , n313068 );
or ( n22644 , n313067 , n313069 );
buf ( n22645 , n305301 );
buf ( n313072 , n854 );
buf ( n313073 , n874 );
xor ( n313074 , n313072 , n313073 );
buf ( n313075 , n313074 );
buf ( n313076 , n313075 );
nand ( n313077 , n22645 , n313076 );
buf ( n313078 , n313077 );
buf ( n313079 , n313078 );
nand ( n313080 , n22644 , n313079 );
buf ( n313081 , n313080 );
buf ( n313082 , n313081 );
buf ( n313083 , n312711 );
not ( n313084 , n313083 );
buf ( n313085 , n306152 );
not ( n22660 , n313085 );
or ( n22661 , n313084 , n22660 );
buf ( n313088 , n312461 );
not ( n22663 , n313088 );
buf ( n313090 , n304658 );
nand ( n22665 , n22663 , n313090 );
buf ( n313092 , n22665 );
buf ( n313093 , n313092 );
nand ( n22668 , n22661 , n313093 );
buf ( n313095 , n22668 );
buf ( n22670 , n313095 );
xor ( n22671 , n313082 , n22670 );
buf ( n313098 , n22350 );
not ( n313099 , n313098 );
buf ( n313100 , n304813 );
not ( n313101 , n313100 );
or ( n22676 , n313099 , n313101 );
buf ( n313103 , n304819 );
buf ( n313104 , n21998 );
nand ( n313105 , n313103 , n313104 );
buf ( n313106 , n313105 );
buf ( n313107 , n313106 );
nand ( n313108 , n22676 , n313107 );
buf ( n313109 , n313108 );
buf ( n313110 , n313109 );
xor ( n22685 , n22671 , n313110 );
buf ( n313112 , n22685 );
buf ( n22687 , n313112 );
xor ( n22688 , n313065 , n22687 );
buf ( n313115 , n312695 );
not ( n313116 , n313115 );
buf ( n313117 , n304584 );
not ( n313118 , n313117 );
or ( n22693 , n313116 , n313118 );
buf ( n313120 , n304596 );
buf ( n313121 , n21943 );
nand ( n313122 , n313120 , n313121 );
buf ( n313123 , n313122 );
buf ( n313124 , n313123 );
nand ( n313125 , n22693 , n313124 );
buf ( n313126 , n313125 );
buf ( n313127 , n313126 );
buf ( n313128 , n312335 );
not ( n22703 , n313128 );
buf ( n313130 , n304763 );
not ( n313131 , n313130 );
or ( n22706 , n22703 , n313131 );
buf ( n22707 , n14323 );
buf ( n22708 , n312760 );
nand ( n22709 , n22707 , n22708 );
buf ( n22710 , n22709 );
buf ( n313137 , n22710 );
nand ( n22712 , n22706 , n313137 );
buf ( n313139 , n22712 );
buf ( n313140 , n313139 );
xor ( n22715 , n313127 , n313140 );
buf ( n313142 , n304854 );
buf ( n313143 , n312797 );
not ( n22718 , n313143 );
buf ( n22719 , n22718 );
buf ( n313146 , n22719 );
or ( n22721 , n313142 , n313146 );
buf ( n313148 , n14439 );
buf ( n313149 , n312402 );
not ( n22724 , n313149 );
buf ( n22725 , n22724 );
buf ( n313152 , n22725 );
or ( n22727 , n313148 , n313152 );
nand ( n22728 , n22721 , n22727 );
buf ( n313155 , n22728 );
buf ( n313156 , n313155 );
xor ( n22731 , n22715 , n313156 );
buf ( n313158 , n22731 );
buf ( n313159 , n313158 );
xor ( n22734 , n22688 , n313159 );
buf ( n313161 , n22734 );
buf ( n313162 , n313161 );
xor ( n22737 , n312766 , n312782 );
xor ( n22738 , n22737 , n312803 );
buf ( n313165 , n22738 );
xor ( n313166 , n14969 , n305445 );
and ( n22741 , n313166 , n305503 );
and ( n22742 , n14969 , n305445 );
or ( n22743 , n22741 , n22742 );
buf ( n22744 , n22743 );
buf ( n313171 , n22744 );
xor ( n22746 , n313165 , n313171 );
xor ( n22747 , n306493 , n306499 );
and ( n313174 , n22747 , n306506 );
and ( n22749 , n306493 , n306499 );
or ( n22750 , n313174 , n22749 );
buf ( n313177 , n22750 );
buf ( n313178 , n313177 );
and ( n313179 , n22746 , n313178 );
and ( n313180 , n313165 , n313171 );
or ( n313181 , n313179 , n313180 );
buf ( n313182 , n313181 );
buf ( n313183 , n313182 );
xor ( n22758 , n313162 , n313183 );
xor ( n313185 , n312730 , n312736 );
xor ( n313186 , n313185 , n312742 );
buf ( n313187 , n313186 );
buf ( n313188 , n313187 );
xor ( n22763 , n312974 , n312980 );
xor ( n313190 , n22763 , n312985 );
buf ( n313191 , n313190 );
buf ( n313192 , n313191 );
xor ( n22767 , n313188 , n313192 );
xor ( n313194 , n305092 , n305183 );
and ( n313195 , n313194 , n305276 );
and ( n313196 , n305092 , n305183 );
or ( n313197 , n313195 , n313196 );
buf ( n313198 , n313197 );
buf ( n313199 , n313198 );
and ( n313200 , n22767 , n313199 );
and ( n22775 , n313188 , n313192 );
or ( n22776 , n313200 , n22775 );
buf ( n313203 , n22776 );
buf ( n313204 , n313203 );
xor ( n22779 , n22758 , n313204 );
buf ( n313206 , n22779 );
buf ( n313207 , n313206 );
and ( n22782 , n22581 , n313207 );
and ( n313209 , n313002 , n22580 );
or ( n313210 , n22782 , n313209 );
buf ( n313211 , n313210 );
buf ( n313212 , n313211 );
buf ( n313213 , n310694 );
not ( n22788 , n313213 );
buf ( n313215 , n22788 );
buf ( n313216 , n313215 );
buf ( n22791 , n312504 );
not ( n313218 , n22791 );
buf ( n313219 , n313218 );
buf ( n313220 , n313219 );
or ( n313221 , n313216 , n313220 );
buf ( n313222 , n310483 );
not ( n313223 , n313222 );
buf ( n313224 , n313223 );
buf ( n313225 , n313224 );
buf ( n22800 , n866 );
buf ( n22801 , n861 );
xor ( n22802 , n22800 , n22801 );
buf ( n22803 , n22802 );
buf ( n313230 , n22803 );
not ( n22805 , n313230 );
buf ( n22806 , n22805 );
buf ( n313233 , n22806 );
or ( n22808 , n313225 , n313233 );
nand ( n313235 , n313221 , n22808 );
buf ( n313236 , n313235 );
buf ( n313237 , n313236 );
and ( n313238 , n312527 , n312544 );
buf ( n313239 , n313238 );
buf ( n313240 , n313239 );
xor ( n22815 , n313237 , n313240 );
xor ( n313242 , n22401 , n312844 );
and ( n22817 , n313242 , n312867 );
and ( n313244 , n22401 , n312844 );
or ( n313245 , n22817 , n313244 );
buf ( n313246 , n313245 );
buf ( n313247 , n313246 );
xor ( n313248 , n22815 , n313247 );
buf ( n313249 , n313248 );
buf ( n313250 , n313249 );
xor ( n22825 , n313065 , n22687 );
and ( n22826 , n22825 , n313159 );
and ( n22827 , n313065 , n22687 );
or ( n22828 , n22826 , n22827 );
buf ( n313255 , n22828 );
buf ( n313256 , n313255 );
xor ( n22831 , n313250 , n313256 );
xor ( n22832 , n312888 , n312948 );
and ( n22833 , n22832 , n312964 );
and ( n22834 , n312888 , n312948 );
or ( n22835 , n22833 , n22834 );
buf ( n313262 , n22835 );
buf ( n313263 , n313262 );
xor ( n22838 , n22831 , n313263 );
buf ( n313265 , n22838 );
buf ( n313266 , n313265 );
xor ( n22841 , n313024 , n22618 );
and ( n313268 , n22841 , n313062 );
and ( n313269 , n313024 , n22618 );
or ( n313270 , n313268 , n313269 );
buf ( n313271 , n313270 );
buf ( n313272 , n313271 );
xor ( n22847 , n313127 , n313140 );
and ( n22848 , n22847 , n313156 );
and ( n22849 , n313127 , n313140 );
or ( n22850 , n22848 , n22849 );
buf ( n313277 , n22850 );
buf ( n313278 , n313277 );
xor ( n22853 , n313272 , n313278 );
xor ( n22854 , n313082 , n22670 );
and ( n313281 , n22854 , n313110 );
and ( n313282 , n313082 , n22670 );
or ( n22857 , n313281 , n313282 );
buf ( n313284 , n22857 );
buf ( n313285 , n313284 );
xor ( n313286 , n22853 , n313285 );
buf ( n313287 , n313286 );
buf ( n22862 , n313287 );
xor ( n313289 , n312807 , n312813 );
and ( n22864 , n313289 , n312870 );
and ( n313291 , n312807 , n312813 );
or ( n313292 , n22864 , n313291 );
buf ( n313293 , n313292 );
buf ( n313294 , n313293 );
xor ( n313295 , n22862 , n313294 );
xor ( n313296 , n22085 , n312547 );
and ( n22871 , n313296 , n312567 );
and ( n22872 , n22085 , n312547 );
or ( n22873 , n22871 , n22872 );
buf ( n22874 , n22873 );
buf ( n313301 , n22874 );
buf ( n313302 , n22434 );
not ( n22877 , n313302 );
buf ( n313304 , n305098 );
not ( n22879 , n313304 );
or ( n22880 , n22877 , n22879 );
buf ( n313307 , n880 );
buf ( n313308 , n847 );
xor ( n22883 , n313307 , n313308 );
buf ( n313310 , n22883 );
buf ( n313311 , n313310 );
buf ( n313312 , n304973 );
nand ( n313313 , n313311 , n313312 );
buf ( n313314 , n313313 );
buf ( n313315 , n313314 );
nand ( n313316 , n22880 , n313315 );
buf ( n313317 , n313316 );
buf ( n313318 , n313317 );
buf ( n313319 , n313036 );
not ( n313320 , n313319 );
buf ( n313321 , n15836 );
not ( n22896 , n313321 );
or ( n313323 , n313320 , n22896 );
buf ( n313324 , n849 );
buf ( n313325 , n878 );
xnor ( n22900 , n313324 , n313325 );
buf ( n313327 , n22900 );
buf ( n313328 , n313327 );
not ( n22903 , n313328 );
buf ( n313330 , n306272 );
nand ( n22905 , n22903 , n313330 );
buf ( n313332 , n22905 );
buf ( n313333 , n313332 );
nand ( n313334 , n313323 , n313333 );
buf ( n313335 , n313334 );
buf ( n313336 , n313335 );
xor ( n313337 , n313318 , n313336 );
buf ( n313338 , n306283 );
buf ( n313339 , n312837 );
not ( n22914 , n313339 );
buf ( n313341 , n22914 );
buf ( n313342 , n313341 );
or ( n313343 , n313338 , n313342 );
buf ( n313344 , n15861 );
buf ( n313345 , n888 );
buf ( n313346 , n14992 );
and ( n313347 , n313345 , n313346 );
not ( n22922 , n313345 );
buf ( n313349 , n839 );
and ( n313350 , n22922 , n313349 );
nor ( n22925 , n313347 , n313350 );
buf ( n313352 , n22925 );
buf ( n313353 , n313352 );
or ( n313354 , n313344 , n313353 );
nand ( n22929 , n313343 , n313354 );
buf ( n313356 , n22929 );
buf ( n313357 , n313356 );
xor ( n22932 , n313337 , n313357 );
buf ( n313359 , n22932 );
buf ( n313360 , n313359 );
xor ( n22935 , n313301 , n313360 );
buf ( n313362 , n313055 );
not ( n22937 , n313362 );
buf ( n313364 , n305338 );
not ( n313365 , n313364 );
or ( n313366 , n22937 , n313365 );
buf ( n313367 , n305344 );
buf ( n22942 , n851 );
buf ( n22943 , n876 );
xor ( n22944 , n22942 , n22943 );
buf ( n22945 , n22944 );
buf ( n313372 , n22945 );
nand ( n22947 , n313367 , n313372 );
buf ( n313374 , n22947 );
buf ( n313375 , n313374 );
nand ( n313376 , n313366 , n313375 );
buf ( n313377 , n313376 );
buf ( n313378 , n313377 );
buf ( n313379 , n313075 );
not ( n313380 , n313379 );
buf ( n313381 , n305627 );
not ( n313382 , n313381 );
or ( n313383 , n313380 , n313382 );
buf ( n313384 , n305301 );
buf ( n313385 , n874 );
buf ( n313386 , n853 );
and ( n22961 , n313385 , n313386 );
not ( n22962 , n313385 );
buf ( n313389 , n304956 );
and ( n22964 , n22962 , n313389 );
nor ( n313391 , n22961 , n22964 );
buf ( n313392 , n313391 );
buf ( n313393 , n313392 );
nand ( n313394 , n313384 , n313393 );
buf ( n313395 , n313394 );
buf ( n313396 , n313395 );
nand ( n22971 , n313383 , n313396 );
buf ( n22972 , n22971 );
buf ( n313399 , n22972 );
xor ( n22974 , n313378 , n313399 );
buf ( n22975 , n304912 );
not ( n22976 , n22975 );
buf ( n313403 , n22976 );
buf ( n313404 , n313403 );
buf ( n313405 , n313017 );
not ( n313406 , n313405 );
buf ( n313407 , n313406 );
buf ( n313408 , n313407 );
or ( n313409 , n313404 , n313408 );
buf ( n313410 , n305363 );
xor ( n22985 , n886 , n841 );
buf ( n313412 , n22985 );
not ( n22987 , n313412 );
buf ( n313414 , n22987 );
buf ( n313415 , n313414 );
or ( n313416 , n313410 , n313415 );
nand ( n22991 , n313409 , n313416 );
buf ( n313418 , n22991 );
buf ( n313419 , n313418 );
xor ( n313420 , n22974 , n313419 );
buf ( n313421 , n313420 );
buf ( n313422 , n313421 );
xor ( n313423 , n22935 , n313422 );
buf ( n313424 , n313423 );
buf ( n313425 , n313424 );
xor ( n23000 , n313295 , n313425 );
buf ( n313427 , n23000 );
buf ( n313428 , n313427 );
xor ( n23003 , n313266 , n313428 );
xor ( n23004 , n313162 , n313183 );
and ( n23005 , n23004 , n313204 );
and ( n313432 , n313162 , n313183 );
or ( n313433 , n23005 , n313432 );
buf ( n313434 , n313433 );
buf ( n313435 , n313434 );
xor ( n23010 , n23003 , n313435 );
buf ( n313437 , n23010 );
buf ( n23012 , n313437 );
xor ( n23013 , n312998 , n313212 );
xor ( n313440 , n23013 , n23012 );
buf ( n313441 , n313440 );
xor ( n313442 , n312998 , n313212 );
and ( n313443 , n313442 , n23012 );
and ( n23018 , n312998 , n313212 );
or ( n313445 , n313443 , n23018 );
buf ( n313446 , n313445 );
buf ( n313447 , n310488 );
not ( n313448 , n313447 );
buf ( n313449 , n310694 );
not ( n313450 , n313449 );
or ( n313451 , n313448 , n313450 );
buf ( n313452 , n311107 );
buf ( n313453 , n866 );
buf ( n313454 , n849 );
xor ( n23029 , n313453 , n313454 );
buf ( n313456 , n23029 );
buf ( n313457 , n313456 );
nand ( n313458 , n313452 , n313457 );
buf ( n313459 , n313458 );
buf ( n313460 , n313459 );
nand ( n313461 , n313451 , n313460 );
buf ( n313462 , n313461 );
buf ( n313463 , n313462 );
buf ( n313464 , n310587 );
not ( n313465 , n313464 );
buf ( n313466 , n310576 );
not ( n313467 , n313466 );
or ( n313468 , n313465 , n313467 );
buf ( n313469 , n310582 );
buf ( n313470 , n864 );
buf ( n313471 , n851 );
xor ( n313472 , n313470 , n313471 );
buf ( n313473 , n313472 );
buf ( n313474 , n313473 );
nand ( n23049 , n313469 , n313474 );
buf ( n313476 , n23049 );
buf ( n313477 , n313476 );
nand ( n313478 , n313468 , n313477 );
buf ( n313479 , n313478 );
buf ( n313480 , n313479 );
xor ( n313481 , n313463 , n313480 );
buf ( n313482 , n305650 );
buf ( n313483 , n310618 );
or ( n313484 , n313482 , n313483 );
buf ( n313485 , n839 );
buf ( n313486 , n876 );
xnor ( n313487 , n313485 , n313486 );
buf ( n313488 , n313487 );
buf ( n313489 , n313488 );
buf ( n313490 , n305664 );
or ( n23065 , n313489 , n313490 );
nand ( n313492 , n313484 , n23065 );
buf ( n313493 , n313492 );
buf ( n313494 , n313493 );
and ( n313495 , n313481 , n313494 );
and ( n23070 , n313463 , n313480 );
or ( n23071 , n313495 , n23070 );
buf ( n313498 , n23071 );
buf ( n23073 , n313498 );
and ( n313500 , n310584 , n310585 );
buf ( n313501 , n313500 );
buf ( n313502 , n313501 );
buf ( n313503 , n872 );
buf ( n313504 , n843 );
and ( n313505 , n313503 , n313504 );
not ( n313506 , n313503 );
buf ( n313507 , n305117 );
and ( n313508 , n313506 , n313507 );
nor ( n23083 , n313505 , n313508 );
buf ( n313510 , n23083 );
buf ( n313511 , n313510 );
not ( n313512 , n313511 );
buf ( n313513 , n304851 );
not ( n313514 , n313513 );
or ( n313515 , n313512 , n313514 );
buf ( n313516 , n304864 );
buf ( n313517 , n872 );
buf ( n313518 , n842 );
and ( n23093 , n313517 , n313518 );
not ( n23094 , n313517 );
buf ( n23095 , n304610 );
and ( n313522 , n23094 , n23095 );
nor ( n23097 , n23093 , n313522 );
buf ( n23098 , n23097 );
buf ( n313525 , n23098 );
nand ( n23100 , n313516 , n313525 );
buf ( n23101 , n23100 );
buf ( n313528 , n23101 );
nand ( n313529 , n313515 , n313528 );
buf ( n313530 , n313529 );
buf ( n313531 , n313530 );
xor ( n313532 , n313502 , n313531 );
buf ( n313533 , n310629 );
buf ( n313534 , n874 );
buf ( n313535 , n841 );
xnor ( n313536 , n313534 , n313535 );
buf ( n313537 , n313536 );
buf ( n313538 , n313537 );
or ( n313539 , n313533 , n313538 );
buf ( n313540 , n306346 );
buf ( n313541 , n874 );
buf ( n313542 , n840 );
and ( n313543 , n313541 , n313542 );
not ( n23118 , n313541 );
buf ( n313545 , n305261 );
and ( n23120 , n23118 , n313545 );
nor ( n23121 , n313543 , n23120 );
buf ( n313548 , n23121 );
buf ( n313549 , n313548 );
not ( n23124 , n313549 );
buf ( n313551 , n23124 );
buf ( n313552 , n313551 );
or ( n313553 , n313540 , n313552 );
nand ( n313554 , n313539 , n313553 );
buf ( n313555 , n313554 );
buf ( n313556 , n313555 );
xor ( n313557 , n313532 , n313556 );
buf ( n313558 , n313557 );
buf ( n313559 , n313558 );
xor ( n23134 , n23073 , n313559 );
buf ( n313561 , n313473 );
not ( n313562 , n313561 );
buf ( n313563 , n311888 );
not ( n23138 , n313563 );
or ( n313565 , n313562 , n23138 );
buf ( n313566 , n310582 );
buf ( n313567 , n864 );
buf ( n313568 , n850 );
xor ( n23143 , n313567 , n313568 );
buf ( n313570 , n23143 );
buf ( n313571 , n313570 );
nand ( n23146 , n313566 , n313571 );
buf ( n313573 , n23146 );
buf ( n313574 , n313573 );
nand ( n313575 , n313565 , n313574 );
buf ( n313576 , n313575 );
buf ( n313577 , n313576 );
buf ( n313578 , n313456 );
not ( n313579 , n313578 );
buf ( n313580 , n310694 );
not ( n313581 , n313580 );
or ( n313582 , n313579 , n313581 );
buf ( n313583 , n866 );
buf ( n313584 , n848 );
xnor ( n313585 , n313583 , n313584 );
buf ( n313586 , n313585 );
buf ( n313587 , n313586 );
not ( n313588 , n313587 );
buf ( n313589 , n310483 );
nand ( n313590 , n313588 , n313589 );
buf ( n313591 , n313590 );
buf ( n313592 , n313591 );
nand ( n313593 , n313582 , n313592 );
buf ( n313594 , n313593 );
buf ( n313595 , n313594 );
xor ( n313596 , n313577 , n313595 );
buf ( n313597 , n304987 );
buf ( n313598 , n880 );
buf ( n313599 , n835 );
xnor ( n23174 , n313598 , n313599 );
buf ( n23175 , n23174 );
buf ( n313602 , n23175 );
or ( n23177 , n313597 , n313602 );
buf ( n313604 , n311075 );
buf ( n313605 , n880 );
buf ( n313606 , n310658 );
and ( n313607 , n313605 , n313606 );
not ( n313608 , n313605 );
buf ( n23183 , n834 );
and ( n313610 , n313608 , n23183 );
nor ( n23185 , n313607 , n313610 );
buf ( n23186 , n23185 );
buf ( n313613 , n23186 );
or ( n23188 , n313604 , n313613 );
nand ( n313615 , n23177 , n23188 );
buf ( n313616 , n313615 );
buf ( n313617 , n313616 );
xor ( n313618 , n313596 , n313617 );
buf ( n313619 , n313618 );
buf ( n313620 , n313619 );
and ( n313621 , n23134 , n313620 );
and ( n313622 , n23073 , n313559 );
or ( n23197 , n313621 , n313622 );
buf ( n313624 , n23197 );
buf ( n313625 , n313624 );
buf ( n313626 , n310352 );
not ( n313627 , n313626 );
buf ( n313628 , n304851 );
not ( n313629 , n313628 );
or ( n23204 , n313627 , n313629 );
buf ( n313631 , n304864 );
buf ( n23206 , n313510 );
nand ( n313633 , n313631 , n23206 );
buf ( n313634 , n313633 );
buf ( n313635 , n313634 );
nand ( n313636 , n23204 , n313635 );
buf ( n313637 , n313636 );
buf ( n313638 , n313637 );
buf ( n313639 , n310645 );
not ( n313640 , n313639 );
buf ( n313641 , n305627 );
not ( n23216 , n313641 );
or ( n313643 , n313640 , n23216 );
buf ( n313644 , n313537 );
not ( n23219 , n313644 );
buf ( n313646 , n305289 );
nand ( n23221 , n23219 , n313646 );
buf ( n313648 , n23221 );
buf ( n313649 , n313648 );
nand ( n23224 , n313643 , n313649 );
buf ( n313651 , n23224 );
buf ( n313652 , n313651 );
xor ( n313653 , n313638 , n313652 );
buf ( n313654 , n304584 );
not ( n313655 , n313654 );
buf ( n313656 , n310506 );
not ( n313657 , n313656 );
or ( n23232 , n313655 , n313657 );
buf ( n313659 , n14959 );
buf ( n313660 , n882 );
buf ( n313661 , n310964 );
and ( n313662 , n313660 , n313661 );
not ( n23237 , n313660 );
buf ( n313664 , n833 );
and ( n313665 , n23237 , n313664 );
nor ( n23240 , n313662 , n313665 );
buf ( n23241 , n23240 );
buf ( n313668 , n23241 );
or ( n313669 , n313659 , n313668 );
nand ( n313670 , n23232 , n313669 );
buf ( n313671 , n313670 );
buf ( n313672 , n313671 );
not ( n313673 , n313672 );
buf ( n313674 , n313673 );
buf ( n313675 , n313674 );
and ( n23250 , n313653 , n313675 );
and ( n23251 , n313638 , n313652 );
or ( n313678 , n23250 , n23251 );
buf ( n313679 , n313678 );
buf ( n313680 , n313679 );
buf ( n313681 , n305650 );
buf ( n313682 , n313488 );
or ( n313683 , n313681 , n313682 );
buf ( n313684 , n305664 );
buf ( n313685 , n876 );
buf ( n313686 , n838 );
xnor ( n23261 , n313685 , n313686 );
buf ( n23262 , n23261 );
buf ( n313689 , n23262 );
or ( n23264 , n313684 , n313689 );
nand ( n313691 , n313683 , n23264 );
buf ( n313692 , n313691 );
buf ( n313693 , n847 );
buf ( n313694 , n868 );
and ( n23269 , n313693 , n313694 );
not ( n313696 , n313693 );
buf ( n23271 , n310521 );
and ( n313698 , n313696 , n23271 );
nor ( n23273 , n23269 , n313698 );
buf ( n23274 , n23273 );
buf ( n313701 , n23274 );
not ( n23276 , n313701 );
buf ( n313703 , n305213 );
not ( n313704 , n313703 );
or ( n23279 , n23276 , n313704 );
buf ( n313706 , n868 );
buf ( n313707 , n846 );
xnor ( n23282 , n313706 , n313707 );
buf ( n313709 , n23282 );
buf ( n313710 , n313709 );
not ( n23285 , n313710 );
buf ( n313712 , n305219 );
nand ( n23287 , n23285 , n313712 );
buf ( n313714 , n23287 );
buf ( n313715 , n313714 );
nand ( n23290 , n23279 , n313715 );
buf ( n313717 , n23290 );
xor ( n313718 , n313692 , n313717 );
buf ( n313719 , n845 );
buf ( n313720 , n870 );
xor ( n313721 , n313719 , n313720 );
buf ( n313722 , n313721 );
buf ( n313723 , n313722 );
not ( n313724 , n313723 );
buf ( n313725 , n14323 );
not ( n313726 , n313725 );
or ( n23301 , n313724 , n313726 );
buf ( n313728 , n870 );
not ( n23303 , n313728 );
buf ( n313730 , n844 );
nor ( n313731 , n23303 , n313730 );
buf ( n313732 , n313731 );
buf ( n313733 , n313732 );
buf ( n313734 , n844 );
not ( n313735 , n313734 );
buf ( n313736 , n870 );
nor ( n313737 , n313735 , n313736 );
buf ( n313738 , n313737 );
buf ( n313739 , n313738 );
nor ( n23314 , n313733 , n313739 );
buf ( n313741 , n23314 );
buf ( n313742 , n313741 );
not ( n313743 , n313742 );
buf ( n313744 , n304763 );
nand ( n23319 , n313743 , n313744 );
buf ( n313746 , n23319 );
buf ( n313747 , n313746 );
nand ( n313748 , n23301 , n313747 );
buf ( n313749 , n313748 );
xor ( n313750 , n313718 , n313749 );
buf ( n313751 , n313750 );
xor ( n23326 , n313680 , n313751 );
buf ( n313753 , n304941 );
buf ( n313754 , n878 );
buf ( n313755 , n837 );
not ( n23330 , n313755 );
buf ( n313757 , n23330 );
buf ( n313758 , n313757 );
and ( n313759 , n313754 , n313758 );
not ( n23334 , n313754 );
buf ( n313761 , n837 );
and ( n313762 , n23334 , n313761 );
nor ( n23337 , n313759 , n313762 );
buf ( n313764 , n23337 );
buf ( n313765 , n313764 );
or ( n313766 , n313753 , n313765 );
buf ( n313767 , n14523 );
buf ( n313768 , n878 );
buf ( n313769 , n311204 );
and ( n313770 , n313768 , n313769 );
not ( n313771 , n313768 );
buf ( n313772 , n836 );
and ( n313773 , n313771 , n313772 );
nor ( n23348 , n313770 , n313773 );
buf ( n313775 , n23348 );
buf ( n313776 , n313775 );
or ( n313777 , n313767 , n313776 );
nand ( n313778 , n313766 , n313777 );
buf ( n313779 , n313778 );
buf ( n313780 , n23241 );
not ( n313781 , n313780 );
buf ( n313782 , n313781 );
buf ( n313783 , n313782 );
not ( n313784 , n313783 );
buf ( n313785 , n304584 );
not ( n313786 , n313785 );
or ( n313787 , n313784 , n313786 );
buf ( n313788 , n304596 );
buf ( n313789 , n882 );
buf ( n313790 , n832 );
and ( n313791 , n313789 , n313790 );
not ( n23366 , n313789 );
buf ( n313793 , n20700 );
and ( n313794 , n23366 , n313793 );
nor ( n313795 , n313791 , n313794 );
buf ( n313796 , n313795 );
buf ( n313797 , n313796 );
nand ( n313798 , n313788 , n313797 );
buf ( n313799 , n313798 );
buf ( n313800 , n313799 );
nand ( n313801 , n313787 , n313800 );
buf ( n313802 , n313801 );
xor ( n313803 , n313779 , n313802 );
buf ( n313804 , n310909 );
not ( n23379 , n313804 );
buf ( n313806 , n15804 );
not ( n313807 , n313806 );
or ( n23382 , n23379 , n313807 );
buf ( n313809 , n884 );
nand ( n23384 , n23382 , n313809 );
buf ( n313811 , n23384 );
xor ( n313812 , n313803 , n313811 );
buf ( n313813 , n313812 );
and ( n23388 , n23326 , n313813 );
and ( n23389 , n313680 , n313751 );
or ( n23390 , n23388 , n23389 );
buf ( n313817 , n23390 );
buf ( n313818 , n313817 );
xor ( n23393 , n313625 , n313818 );
and ( n23394 , n313470 , n313471 );
buf ( n313821 , n23394 );
buf ( n313822 , n313821 );
buf ( n313823 , n313570 );
not ( n23398 , n313823 );
buf ( n313825 , n311888 );
not ( n23400 , n313825 );
or ( n313827 , n23398 , n23400 );
buf ( n313828 , n310582 );
buf ( n313829 , n864 );
buf ( n313830 , n849 );
xor ( n23405 , n313829 , n313830 );
buf ( n313832 , n23405 );
buf ( n313833 , n313832 );
nand ( n23408 , n313828 , n313833 );
buf ( n313835 , n23408 );
buf ( n313836 , n313835 );
nand ( n23411 , n313827 , n313836 );
buf ( n313838 , n23411 );
buf ( n313839 , n313838 );
xor ( n23414 , n313822 , n313839 );
buf ( n313841 , n313548 );
not ( n23416 , n313841 );
buf ( n313843 , n305627 );
not ( n23418 , n313843 );
or ( n313845 , n23416 , n23418 );
buf ( n313846 , n305301 );
buf ( n313847 , n874 );
buf ( n313848 , n839 );
and ( n313849 , n313847 , n313848 );
not ( n313850 , n313847 );
buf ( n313851 , n14992 );
and ( n313852 , n313850 , n313851 );
nor ( n313853 , n313849 , n313852 );
buf ( n313854 , n313853 );
buf ( n313855 , n313854 );
nand ( n313856 , n313846 , n313855 );
buf ( n313857 , n313856 );
buf ( n313858 , n313857 );
nand ( n313859 , n313845 , n313858 );
buf ( n313860 , n313859 );
buf ( n313861 , n313860 );
xor ( n313862 , n23414 , n313861 );
buf ( n313863 , n313862 );
buf ( n313864 , n313863 );
buf ( n313865 , n847 );
buf ( n23440 , n866 );
and ( n23441 , n313865 , n23440 );
not ( n313868 , n313865 );
buf ( n23443 , n866 );
not ( n313870 , n23443 );
buf ( n313871 , n313870 );
buf ( n313872 , n313871 );
and ( n313873 , n313868 , n313872 );
nor ( n23448 , n23441 , n313873 );
buf ( n23449 , n23448 );
buf ( n313876 , n23449 );
not ( n313877 , n313876 );
buf ( n313878 , n311107 );
not ( n313879 , n313878 );
or ( n23454 , n313877 , n313879 );
buf ( n313881 , n313586 );
not ( n23456 , n313881 );
buf ( n313883 , n310694 );
nand ( n23458 , n23456 , n313883 );
buf ( n313885 , n23458 );
buf ( n313886 , n313885 );
nand ( n313887 , n23454 , n313886 );
buf ( n313888 , n313887 );
buf ( n313889 , n313888 );
buf ( n313890 , n876 );
buf ( n313891 , n313757 );
and ( n23466 , n313890 , n313891 );
not ( n313893 , n313890 );
buf ( n313894 , n837 );
and ( n313895 , n313893 , n313894 );
nor ( n313896 , n23466 , n313895 );
buf ( n313897 , n313896 );
buf ( n313898 , n313897 );
not ( n313899 , n313898 );
buf ( n313900 , n313899 );
buf ( n313901 , n313900 );
not ( n313902 , n313901 );
buf ( n313903 , n305344 );
not ( n313904 , n313903 );
or ( n313905 , n313902 , n313904 );
buf ( n313906 , n23262 );
not ( n313907 , n313906 );
buf ( n313908 , n305338 );
nand ( n313909 , n313907 , n313908 );
buf ( n313910 , n313909 );
buf ( n313911 , n313910 );
nand ( n313912 , n313905 , n313911 );
buf ( n313913 , n313912 );
buf ( n313914 , n313913 );
xor ( n313915 , n313889 , n313914 );
buf ( n313916 , n305210 );
buf ( n313917 , n313709 );
or ( n313918 , n313916 , n313917 );
buf ( n313919 , n305205 );
buf ( n313920 , n310521 );
buf ( n313921 , n845 );
and ( n23496 , n313920 , n313921 );
buf ( n313923 , n310777 );
buf ( n313924 , n868 );
and ( n23499 , n313923 , n313924 );
nor ( n23500 , n23496 , n23499 );
buf ( n313927 , n23500 );
buf ( n313928 , n313927 );
or ( n23503 , n313919 , n313928 );
nand ( n23504 , n313918 , n23503 );
buf ( n313931 , n23504 );
buf ( n313932 , n313931 );
xor ( n23507 , n313915 , n313932 );
buf ( n313934 , n23507 );
buf ( n313935 , n313934 );
xor ( n313936 , n313864 , n313935 );
buf ( n313937 , n23098 );
not ( n313938 , n313937 );
buf ( n313939 , n304851 );
not ( n313940 , n313939 );
or ( n313941 , n313938 , n313940 );
buf ( n313942 , n872 );
buf ( n313943 , n841 );
xnor ( n23518 , n313942 , n313943 );
buf ( n313945 , n23518 );
buf ( n313946 , n313945 );
not ( n313947 , n313946 );
buf ( n313948 , n304864 );
nand ( n313949 , n313947 , n313948 );
buf ( n313950 , n313949 );
buf ( n313951 , n313950 );
nand ( n313952 , n313941 , n313951 );
buf ( n313953 , n313952 );
buf ( n313954 , n313953 );
buf ( n313955 , n313796 );
not ( n313956 , n313955 );
buf ( n313957 , n304584 );
not ( n23532 , n313957 );
or ( n313959 , n313956 , n23532 );
buf ( n313960 , n304596 );
buf ( n313961 , n882 );
nand ( n313962 , n313960 , n313961 );
buf ( n313963 , n313962 );
buf ( n313964 , n313963 );
nand ( n23539 , n313959 , n313964 );
buf ( n313966 , n23539 );
buf ( n313967 , n313966 );
xor ( n313968 , n313954 , n313967 );
buf ( n313969 , n304941 );
buf ( n313970 , n313775 );
or ( n23545 , n313969 , n313970 );
buf ( n313972 , n878 );
buf ( n313973 , n835 );
and ( n23548 , n313972 , n313973 );
not ( n313975 , n313972 );
buf ( n313976 , n21261 );
and ( n313977 , n313975 , n313976 );
nor ( n23552 , n23548 , n313977 );
buf ( n23553 , n23552 );
buf ( n313980 , n23553 );
not ( n23555 , n313980 );
buf ( n313982 , n23555 );
buf ( n313983 , n313982 );
buf ( n313984 , n14523 );
or ( n23559 , n313983 , n313984 );
nand ( n313986 , n23545 , n23559 );
buf ( n313987 , n313986 );
buf ( n313988 , n313987 );
xor ( n23563 , n313968 , n313988 );
buf ( n313990 , n23563 );
buf ( n313991 , n313990 );
xor ( n313992 , n313936 , n313991 );
buf ( n313993 , n313992 );
buf ( n313994 , n313993 );
xor ( n313995 , n23393 , n313994 );
buf ( n313996 , n313995 );
buf ( n313997 , n313996 );
xor ( n313998 , n310495 , n310513 );
and ( n313999 , n313998 , n310542 );
and ( n23574 , n310495 , n310513 );
or ( n314001 , n313999 , n23574 );
buf ( n314002 , n314001 );
buf ( n314003 , n314002 );
xor ( n23578 , n310416 , n310425 );
and ( n23579 , n23578 , n310456 );
and ( n23580 , n310416 , n310425 );
or ( n23581 , n23579 , n23580 );
buf ( n314008 , n23581 );
buf ( n314009 , n314008 );
xor ( n314010 , n314003 , n314009 );
xor ( n23585 , n310561 , n310594 );
and ( n23586 , n23585 , n310623 );
and ( n23587 , n310561 , n310594 );
or ( n23588 , n23586 , n23587 );
buf ( n314015 , n23588 );
buf ( n314016 , n314015 );
and ( n314017 , n314010 , n314016 );
and ( n314018 , n314003 , n314009 );
or ( n314019 , n314017 , n314018 );
buf ( n314020 , n314019 );
buf ( n314021 , n314020 );
buf ( n314022 , n313671 );
and ( n23597 , n310562 , n20137 );
buf ( n314024 , n23597 );
buf ( n314025 , n314024 );
buf ( n314026 , n310447 );
not ( n23601 , n314026 );
buf ( n314028 , n304984 );
not ( n314029 , n314028 );
or ( n23604 , n23601 , n314029 );
buf ( n314031 , n23175 );
not ( n23606 , n314031 );
buf ( n314033 , n304973 );
nand ( n23608 , n23606 , n314033 );
buf ( n314035 , n23608 );
buf ( n314036 , n314035 );
nand ( n23611 , n23604 , n314036 );
buf ( n314038 , n23611 );
buf ( n314039 , n314038 );
xor ( n314040 , n314025 , n314039 );
buf ( n314041 , n15804 );
buf ( n314042 , n310409 );
not ( n314043 , n314042 );
buf ( n314044 , n314043 );
buf ( n314045 , n314044 );
or ( n23620 , n314041 , n314045 );
buf ( n314047 , n306238 );
buf ( n314048 , n304827 );
or ( n23623 , n314047 , n314048 );
nand ( n23624 , n23620 , n23623 );
buf ( n314051 , n23624 );
buf ( n314052 , n314051 );
and ( n23627 , n314040 , n314052 );
and ( n23628 , n314025 , n314039 );
or ( n314055 , n23627 , n23628 );
buf ( n314056 , n314055 );
buf ( n314057 , n314056 );
xor ( n23632 , n314022 , n314057 );
buf ( n314059 , n19908 );
not ( n314060 , n314059 );
buf ( n314061 , n304754 );
not ( n314062 , n314061 );
or ( n23637 , n314060 , n314062 );
buf ( n314064 , n311052 );
buf ( n23639 , n313722 );
nand ( n23640 , n314064 , n23639 );
buf ( n23641 , n23640 );
buf ( n23642 , n23641 );
nand ( n23643 , n23637 , n23642 );
buf ( n23644 , n23643 );
buf ( n314071 , n23644 );
buf ( n314072 , n310535 );
not ( n314073 , n314072 );
buf ( n314074 , n305213 );
not ( n23649 , n314074 );
or ( n314076 , n314073 , n23649 );
buf ( n23651 , n305219 );
buf ( n23652 , n23274 );
nand ( n23653 , n23651 , n23652 );
buf ( n23654 , n23653 );
buf ( n314081 , n23654 );
nand ( n23656 , n314076 , n314081 );
buf ( n23657 , n23656 );
buf ( n314084 , n23657 );
xor ( n23659 , n314071 , n314084 );
buf ( n314086 , n304941 );
buf ( n314087 , n310382 );
or ( n23662 , n314086 , n314087 );
buf ( n314089 , n14523 );
buf ( n314090 , n313764 );
or ( n23665 , n314089 , n314090 );
nand ( n314092 , n23662 , n23665 );
buf ( n314093 , n314092 );
buf ( n314094 , n314093 );
and ( n23669 , n23659 , n314094 );
and ( n314096 , n314071 , n314084 );
or ( n314097 , n23669 , n314096 );
buf ( n314098 , n314097 );
buf ( n314099 , n314098 );
xor ( n23674 , n23632 , n314099 );
buf ( n314101 , n23674 );
buf ( n314102 , n314101 );
xor ( n23677 , n314021 , n314102 );
xor ( n23678 , n310341 , n310359 );
and ( n23679 , n23678 , n310387 );
and ( n23680 , n310341 , n310359 );
or ( n23681 , n23679 , n23680 );
buf ( n314108 , n23681 );
buf ( n314109 , n314108 );
xor ( n23684 , n314025 , n314039 );
xor ( n23685 , n23684 , n314052 );
buf ( n314112 , n23685 );
buf ( n314113 , n314112 );
xor ( n23688 , n314109 , n314113 );
xor ( n314115 , n314071 , n314084 );
xor ( n314116 , n314115 , n314094 );
buf ( n314117 , n314116 );
buf ( n314118 , n314117 );
and ( n23693 , n23688 , n314118 );
and ( n23694 , n314109 , n314113 );
or ( n314121 , n23693 , n23694 );
buf ( n314122 , n314121 );
buf ( n314123 , n314122 );
xor ( n314124 , n23677 , n314123 );
buf ( n314125 , n314124 );
buf ( n314126 , n314125 );
xor ( n23701 , n310653 , n310676 );
and ( n23702 , n23701 , n310747 );
and ( n314129 , n310653 , n310676 );
or ( n23704 , n23702 , n314129 );
buf ( n314131 , n23704 );
buf ( n23706 , n314131 );
buf ( n314133 , n310544 );
not ( n314134 , n314133 );
buf ( n314135 , n310389 );
not ( n314136 , n314135 );
or ( n314137 , n314134 , n314136 );
buf ( n314138 , n310389 );
buf ( n314139 , n310544 );
or ( n314140 , n314138 , n314139 );
buf ( n314141 , n310458 );
nand ( n314142 , n314140 , n314141 );
buf ( n314143 , n314142 );
buf ( n314144 , n314143 );
nand ( n23719 , n314137 , n314144 );
buf ( n314146 , n23719 );
buf ( n314147 , n314146 );
xor ( n314148 , n23706 , n314147 );
xor ( n314149 , n314003 , n314009 );
xor ( n23724 , n314149 , n314016 );
buf ( n314151 , n23724 );
buf ( n314152 , n314151 );
and ( n314153 , n314148 , n314152 );
and ( n23728 , n23706 , n314147 );
or ( n23729 , n314153 , n23728 );
buf ( n314156 , n23729 );
buf ( n314157 , n314156 );
xor ( n314158 , n314126 , n314157 );
xor ( n314159 , n314109 , n314113 );
xor ( n23734 , n314159 , n314118 );
buf ( n314161 , n23734 );
buf ( n314162 , n314161 );
xor ( n314163 , n313463 , n313480 );
xor ( n23738 , n314163 , n313494 );
buf ( n314165 , n23738 );
buf ( n314166 , n314165 );
xor ( n314167 , n313638 , n313652 );
xor ( n23742 , n314167 , n313675 );
buf ( n314169 , n23742 );
buf ( n314170 , n314169 );
xor ( n314171 , n314166 , n314170 );
xor ( n23746 , n311505 , n311511 );
and ( n314173 , n23746 , n311553 );
and ( n23748 , n311505 , n311511 );
or ( n23749 , n314173 , n23748 );
buf ( n314176 , n23749 );
buf ( n314177 , n314176 );
xor ( n314178 , n314171 , n314177 );
buf ( n314179 , n314178 );
buf ( n314180 , n314179 );
xor ( n23755 , n314162 , n314180 );
xor ( n314182 , n20200 , n310750 );
and ( n23757 , n314182 , n310925 );
and ( n314184 , n20200 , n310750 );
or ( n314185 , n23757 , n314184 );
buf ( n314186 , n314185 );
buf ( n314187 , n314186 );
and ( n314188 , n23755 , n314187 );
and ( n23763 , n314162 , n314180 );
or ( n23764 , n314188 , n23763 );
buf ( n314191 , n23764 );
buf ( n314192 , n314191 );
and ( n23767 , n314158 , n314192 );
and ( n314194 , n314126 , n314157 );
or ( n314195 , n23767 , n314194 );
buf ( n314196 , n314195 );
buf ( n314197 , n314196 );
buf ( n314198 , n304987 );
buf ( n314199 , n23186 );
or ( n314200 , n314198 , n314199 );
buf ( n314201 , n311075 );
buf ( n314202 , n880 );
buf ( n23777 , n310964 );
and ( n23778 , n314202 , n23777 );
not ( n23779 , n314202 );
buf ( n314206 , n833 );
and ( n23781 , n23779 , n314206 );
nor ( n23782 , n23778 , n23781 );
buf ( n314209 , n23782 );
buf ( n314210 , n314209 );
or ( n23785 , n314201 , n314210 );
nand ( n23786 , n314200 , n23785 );
buf ( n314213 , n23786 );
buf ( n314214 , n314213 );
not ( n23789 , n314214 );
buf ( n314216 , n23789 );
buf ( n314217 , n14323 );
not ( n23792 , n314217 );
buf ( n314219 , n23792 );
buf ( n314220 , n314219 );
buf ( n314221 , n313741 );
or ( n314222 , n314220 , n314221 );
buf ( n314223 , n311052 );
not ( n314224 , n314223 );
buf ( n314225 , n314224 );
buf ( n314226 , n314225 );
buf ( n314227 , n870 );
buf ( n314228 , n305117 );
and ( n23803 , n314227 , n314228 );
not ( n23804 , n314227 );
buf ( n23805 , n843 );
and ( n314232 , n23804 , n23805 );
nor ( n314233 , n23803 , n314232 );
buf ( n314234 , n314233 );
buf ( n314235 , n314234 );
or ( n314236 , n314226 , n314235 );
nand ( n23811 , n314222 , n314236 );
buf ( n23812 , n23811 );
xor ( n314239 , n314216 , n23812 );
xor ( n23814 , n313577 , n313595 );
and ( n314241 , n23814 , n313617 );
and ( n314242 , n313577 , n313595 );
or ( n23817 , n314241 , n314242 );
buf ( n314244 , n23817 );
xor ( n23819 , n314239 , n314244 );
xor ( n314246 , n314022 , n314057 );
and ( n23821 , n314246 , n314099 );
and ( n23822 , n314022 , n314057 );
or ( n314249 , n23821 , n23822 );
buf ( n314250 , n314249 );
buf ( n314251 , n313749 );
not ( n23826 , n314251 );
buf ( n314253 , n313692 );
not ( n314254 , n314253 );
or ( n23829 , n23826 , n314254 );
buf ( n314256 , n313749 );
buf ( n314257 , n313692 );
or ( n23832 , n314256 , n314257 );
buf ( n314259 , n313717 );
nand ( n314260 , n23832 , n314259 );
buf ( n314261 , n314260 );
buf ( n314262 , n314261 );
nand ( n314263 , n23829 , n314262 );
buf ( n314264 , n314263 );
buf ( n314265 , n314264 );
xor ( n23840 , n313779 , n313802 );
and ( n23841 , n23840 , n313811 );
and ( n23842 , n313779 , n313802 );
or ( n23843 , n23841 , n23842 );
buf ( n314270 , n23843 );
xor ( n314271 , n314265 , n314270 );
xor ( n314272 , n313502 , n313531 );
and ( n23847 , n314272 , n313556 );
and ( n314274 , n313502 , n313531 );
or ( n314275 , n23847 , n314274 );
buf ( n314276 , n314275 );
buf ( n314277 , n314276 );
xor ( n23852 , n314271 , n314277 );
buf ( n314279 , n23852 );
xor ( n23854 , n314250 , n314279 );
xor ( n23855 , n23819 , n23854 );
buf ( n314282 , n23855 );
xor ( n23857 , n314021 , n314102 );
and ( n23858 , n23857 , n314123 );
and ( n23859 , n314021 , n314102 );
or ( n23860 , n23858 , n23859 );
buf ( n314287 , n23860 );
buf ( n314288 , n314287 );
xor ( n314289 , n314282 , n314288 );
xor ( n23864 , n314166 , n314170 );
and ( n314291 , n23864 , n314177 );
and ( n314292 , n314166 , n314170 );
or ( n23867 , n314291 , n314292 );
buf ( n314294 , n23867 );
buf ( n314295 , n314294 );
xor ( n23870 , n313680 , n313751 );
xor ( n23871 , n23870 , n313813 );
buf ( n314298 , n23871 );
buf ( n314299 , n314298 );
xor ( n314300 , n314295 , n314299 );
xor ( n23875 , n23073 , n313559 );
xor ( n23876 , n23875 , n313620 );
buf ( n314303 , n23876 );
buf ( n314304 , n314303 );
and ( n314305 , n314300 , n314304 );
and ( n23880 , n314295 , n314299 );
or ( n314307 , n314305 , n23880 );
buf ( n314308 , n314307 );
buf ( n314309 , n314308 );
xor ( n314310 , n314289 , n314309 );
buf ( n314311 , n314310 );
buf ( n314312 , n314311 );
xor ( n314313 , n313997 , n314197 );
xor ( n314314 , n314313 , n314312 );
buf ( n314315 , n314314 );
xor ( n314316 , n313997 , n314197 );
and ( n314317 , n314316 , n314312 );
and ( n23892 , n313997 , n314197 );
or ( n314319 , n314317 , n23892 );
buf ( n314320 , n314319 );
xor ( n23895 , n314162 , n314180 );
xor ( n23896 , n23895 , n314187 );
buf ( n314323 , n23896 );
buf ( n23898 , n314323 );
xor ( n314325 , n311447 , n311583 );
and ( n23900 , n314325 , n311867 );
and ( n314327 , n311447 , n311583 );
or ( n314328 , n23900 , n314327 );
buf ( n314329 , n314328 );
buf ( n314330 , n314329 );
xor ( n314331 , n23706 , n314147 );
xor ( n23906 , n314331 , n314152 );
buf ( n314333 , n23906 );
buf ( n314334 , n314333 );
xor ( n314335 , n311453 , n311556 );
and ( n314336 , n314335 , n311580 );
and ( n23911 , n311453 , n311556 );
or ( n314338 , n314336 , n23911 );
buf ( n314339 , n314338 );
buf ( n314340 , n314339 );
xor ( n314341 , n314334 , n314340 );
xor ( n23916 , n310556 , n310928 );
and ( n314343 , n23916 , n311189 );
and ( n314344 , n310556 , n310928 );
or ( n314345 , n314343 , n314344 );
buf ( n314346 , n314345 );
buf ( n314347 , n314346 );
xor ( n314348 , n314341 , n314347 );
buf ( n314349 , n314348 );
buf ( n314350 , n314349 );
xor ( n314351 , n23898 , n314330 );
xor ( n314352 , n314351 , n314350 );
buf ( n314353 , n314352 );
xor ( n314354 , n23898 , n314330 );
and ( n314355 , n314354 , n314350 );
and ( n23930 , n23898 , n314330 );
or ( n314357 , n314355 , n23930 );
buf ( n314358 , n314357 );
xor ( n314359 , n314295 , n314299 );
xor ( n23934 , n314359 , n314304 );
buf ( n314361 , n23934 );
buf ( n314362 , n314361 );
xor ( n23937 , n314126 , n314157 );
xor ( n23938 , n23937 , n314192 );
buf ( n314365 , n23938 );
buf ( n314366 , n314365 );
xor ( n314367 , n314334 , n314340 );
and ( n23942 , n314367 , n314347 );
and ( n314369 , n314334 , n314340 );
or ( n23944 , n23942 , n314369 );
buf ( n314371 , n23944 );
buf ( n314372 , n314371 );
xor ( n314373 , n314362 , n314366 );
xor ( n314374 , n314373 , n314372 );
buf ( n314375 , n314374 );
xor ( n314376 , n314362 , n314366 );
and ( n314377 , n314376 , n314372 );
and ( n23952 , n314362 , n314366 );
or ( n314379 , n314377 , n23952 );
buf ( n314380 , n314379 );
xor ( n23955 , n305312 , n305352 );
xor ( n314382 , n23955 , n14944 );
and ( n314383 , n305378 , n314382 );
xor ( n23958 , n305312 , n305352 );
xor ( n314385 , n23958 , n14944 );
and ( n23960 , n305505 , n314385 );
and ( n23961 , n305378 , n305505 );
or ( n314388 , n314383 , n23960 , n23961 );
buf ( n23963 , n314388 );
buf ( n314390 , n312666 );
not ( n23965 , n314390 );
buf ( n314392 , n312721 );
buf ( n23967 , n22190 );
and ( n23968 , n314392 , n23967 );
not ( n314395 , n314392 );
buf ( n314396 , n312619 );
and ( n23971 , n314395 , n314396 );
nor ( n314398 , n23968 , n23971 );
buf ( n314399 , n314398 );
buf ( n314400 , n314399 );
not ( n23975 , n314400 );
or ( n314402 , n23965 , n23975 );
buf ( n314403 , n314399 );
buf ( n314404 , n312666 );
or ( n314405 , n314403 , n314404 );
nand ( n314406 , n314402 , n314405 );
buf ( n314407 , n314406 );
buf ( n314408 , n314407 );
xor ( n314409 , n23963 , n314408 );
xor ( n314410 , n306427 , n306486 );
and ( n23985 , n314410 , n306509 );
and ( n314412 , n306427 , n306486 );
or ( n314413 , n23985 , n314412 );
buf ( n314414 , n314413 );
buf ( n314415 , n314414 );
and ( n23990 , n314409 , n314415 );
and ( n314417 , n23963 , n314408 );
or ( n23992 , n23990 , n314417 );
buf ( n314419 , n23992 );
buf ( n314420 , n314419 );
xor ( n23995 , n313165 , n313171 );
xor ( n23996 , n23995 , n313178 );
buf ( n314423 , n23996 );
buf ( n314424 , n314423 );
xor ( n23999 , n313188 , n313192 );
xor ( n314426 , n23999 , n313199 );
buf ( n314427 , n314426 );
buf ( n314428 , n314427 );
xor ( n314429 , n314424 , n314428 );
xor ( n24004 , n305021 , n305279 );
and ( n24005 , n24004 , n305508 );
and ( n24006 , n305021 , n305279 );
or ( n314433 , n24005 , n24006 );
buf ( n314434 , n314433 );
buf ( n314435 , n314434 );
and ( n24010 , n314429 , n314435 );
and ( n24011 , n314424 , n314428 );
or ( n24012 , n24010 , n24011 );
buf ( n314439 , n24012 );
buf ( n314440 , n314439 );
xor ( n24015 , n313002 , n22580 );
xor ( n24016 , n24015 , n313207 );
buf ( n314443 , n24016 );
buf ( n314444 , n314443 );
xor ( n24019 , n314420 , n314440 );
xor ( n24020 , n24019 , n314444 );
buf ( n24021 , n24020 );
xor ( n314448 , n314420 , n314440 );
and ( n24023 , n314448 , n314444 );
and ( n24024 , n314420 , n314440 );
or ( n24025 , n24023 , n24024 );
buf ( n24026 , n24025 );
xor ( n24027 , n23963 , n314408 );
xor ( n24028 , n24027 , n314415 );
buf ( n314455 , n24028 );
buf ( n314456 , n314455 );
xor ( n24031 , n306512 , n306518 );
and ( n24032 , n24031 , n306537 );
and ( n314459 , n306512 , n306518 );
or ( n24034 , n24032 , n314459 );
buf ( n314461 , n24034 );
buf ( n314462 , n314461 );
xor ( n24037 , n314424 , n314428 );
xor ( n24038 , n24037 , n314435 );
buf ( n314465 , n24038 );
buf ( n314466 , n314465 );
xor ( n24041 , n314456 , n314462 );
xor ( n24042 , n24041 , n314466 );
buf ( n314469 , n24042 );
xor ( n24044 , n314456 , n314462 );
and ( n24045 , n24044 , n314466 );
and ( n24046 , n314456 , n314462 );
or ( n314473 , n24045 , n24046 );
buf ( n314474 , n314473 );
xor ( n24049 , n306523 , n306527 );
xor ( n314476 , n24049 , n306532 );
buf ( n314477 , n314476 );
buf ( n314478 , n314477 );
buf ( n314479 , n304581 );
buf ( n314480 , n882 );
not ( n314481 , n314480 );
buf ( n314482 , n853 );
nor ( n314483 , n314481 , n314482 );
buf ( n314484 , n314483 );
buf ( n314485 , n314484 );
buf ( n314486 , n853 );
not ( n24061 , n314486 );
buf ( n314488 , n882 );
nor ( n314489 , n24061 , n314488 );
buf ( n314490 , n314489 );
buf ( n314491 , n314490 );
nor ( n314492 , n314485 , n314491 );
buf ( n314493 , n314492 );
buf ( n314494 , n314493 );
or ( n24069 , n314479 , n314494 );
buf ( n314496 , n14959 );
buf ( n314497 , n305520 );
or ( n24072 , n314496 , n314497 );
nand ( n24073 , n24069 , n24072 );
buf ( n314500 , n24073 );
buf ( n314501 , n314500 );
buf ( n314502 , n15804 );
buf ( n314503 , n884 );
buf ( n314504 , n851 );
xnor ( n24079 , n314503 , n314504 );
buf ( n314506 , n24079 );
buf ( n314507 , n314506 );
or ( n24082 , n314502 , n314507 );
buf ( n314509 , n306238 );
buf ( n314510 , n305760 );
not ( n24085 , n314510 );
buf ( n314512 , n24085 );
buf ( n24087 , n314512 );
or ( n24088 , n314509 , n24087 );
nand ( n24089 , n24082 , n24088 );
buf ( n24090 , n24089 );
buf ( n314517 , n24090 );
xor ( n24092 , n314501 , n314517 );
xor ( n24093 , n305558 , n15157 );
buf ( n24094 , n24093 );
buf ( n314521 , n24094 );
and ( n314522 , n24092 , n314521 );
and ( n314523 , n314501 , n314517 );
or ( n24098 , n314522 , n314523 );
buf ( n314525 , n24098 );
buf ( n314526 , n314525 );
buf ( n314527 , n842 );
buf ( n314528 , n894 );
xor ( n24103 , n314527 , n314528 );
buf ( n314530 , n24103 );
buf ( n314531 , n314530 );
not ( n314532 , n314531 );
buf ( n314533 , n305032 );
not ( n314534 , n314533 );
or ( n314535 , n314532 , n314534 );
buf ( n314536 , n306106 );
buf ( n314537 , n895 );
nand ( n24112 , n314536 , n314537 );
buf ( n314539 , n24112 );
buf ( n314540 , n314539 );
nand ( n24115 , n314535 , n314540 );
buf ( n24116 , n24115 );
buf ( n314543 , n24116 );
buf ( n314544 , n874 );
buf ( n314545 , n862 );
and ( n314546 , n314544 , n314545 );
not ( n24121 , n314544 );
buf ( n314548 , n304739 );
and ( n314549 , n24121 , n314548 );
nor ( n314550 , n314546 , n314549 );
buf ( n314551 , n314550 );
buf ( n314552 , n314551 );
not ( n314553 , n314552 );
buf ( n314554 , n305627 );
not ( n314555 , n314554 );
or ( n24130 , n314553 , n314555 );
buf ( n314557 , n305289 );
buf ( n314558 , n305618 );
nand ( n314559 , n314557 , n314558 );
buf ( n314560 , n314559 );
buf ( n314561 , n314560 );
nand ( n314562 , n24130 , n314561 );
buf ( n314563 , n314562 );
buf ( n314564 , n314563 );
xor ( n314565 , n314543 , n314564 );
buf ( n314566 , n305650 );
buf ( n314567 , n860 );
buf ( n314568 , n876 );
xnor ( n24143 , n314567 , n314568 );
buf ( n314570 , n24143 );
buf ( n314571 , n314570 );
or ( n24146 , n314566 , n314571 );
buf ( n314573 , n305664 );
buf ( n314574 , n305659 );
or ( n24149 , n314573 , n314574 );
nand ( n314576 , n24146 , n24149 );
buf ( n314577 , n314576 );
buf ( n314578 , n314577 );
and ( n314579 , n314565 , n314578 );
and ( n24154 , n314543 , n314564 );
or ( n24155 , n314579 , n24154 );
buf ( n314582 , n24155 );
buf ( n314583 , n314582 );
buf ( n314584 , n304864 );
buf ( n314585 , n863 );
and ( n314586 , n314584 , n314585 );
buf ( n314587 , n314586 );
buf ( n314588 , n314587 );
xor ( n24163 , n888 , n848 );
buf ( n314590 , n24163 );
not ( n314591 , n314590 );
buf ( n314592 , n305138 );
not ( n314593 , n314592 );
or ( n24168 , n314591 , n314593 );
buf ( n314595 , n305144 );
buf ( n314596 , n306070 );
nand ( n314597 , n314595 , n314596 );
buf ( n314598 , n314597 );
buf ( n314599 , n314598 );
nand ( n314600 , n24168 , n314599 );
buf ( n314601 , n314600 );
buf ( n314602 , n314601 );
xor ( n314603 , n314588 , n314602 );
buf ( n314604 , n305561 );
buf ( n24179 , n844 );
buf ( n24180 , n892 );
xnor ( n24181 , n24179 , n24180 );
buf ( n24182 , n24181 );
buf ( n314609 , n24182 );
or ( n24184 , n314604 , n314609 );
buf ( n314611 , n305489 );
buf ( n314612 , n15145 );
or ( n24187 , n314611 , n314612 );
nand ( n314614 , n24184 , n24187 );
buf ( n314615 , n314614 );
buf ( n314616 , n314615 );
and ( n314617 , n314603 , n314616 );
and ( n314618 , n314588 , n314602 );
or ( n24193 , n314617 , n314618 );
buf ( n314620 , n24193 );
buf ( n314621 , n314620 );
xor ( n24196 , n314583 , n314621 );
buf ( n314623 , n854 );
buf ( n314624 , n882 );
xor ( n314625 , n314623 , n314624 );
buf ( n314626 , n314625 );
buf ( n314627 , n314626 );
not ( n314628 , n314627 );
buf ( n24203 , n304584 );
not ( n24204 , n24203 );
or ( n24205 , n314628 , n24204 );
buf ( n314632 , n314493 );
not ( n314633 , n314632 );
buf ( n314634 , n304596 );
nand ( n314635 , n314633 , n314634 );
buf ( n314636 , n314635 );
buf ( n314637 , n314636 );
nand ( n314638 , n24205 , n314637 );
buf ( n314639 , n314638 );
buf ( n314640 , n314639 );
buf ( n314641 , n884 );
buf ( n24216 , n852 );
and ( n24217 , n314641 , n24216 );
not ( n314644 , n314641 );
buf ( n314645 , n305168 );
and ( n24220 , n314644 , n314645 );
nor ( n314647 , n24217 , n24220 );
buf ( n314648 , n314647 );
buf ( n314649 , n314648 );
not ( n314650 , n314649 );
buf ( n314651 , n304813 );
not ( n314652 , n314651 );
or ( n24227 , n314650 , n314652 );
buf ( n314654 , n314506 );
not ( n24229 , n314654 );
buf ( n314656 , n304819 );
nand ( n314657 , n24229 , n314656 );
buf ( n314658 , n314657 );
buf ( n314659 , n314658 );
nand ( n24234 , n24227 , n314659 );
buf ( n314661 , n24234 );
buf ( n314662 , n314661 );
xor ( n314663 , n314640 , n314662 );
buf ( n314664 , n304630 );
buf ( n314665 , n890 );
buf ( n314666 , n846 );
xnor ( n314667 , n314665 , n314666 );
buf ( n314668 , n314667 );
buf ( n314669 , n314668 );
or ( n24244 , n314664 , n314669 );
buf ( n314671 , n304655 );
buf ( n314672 , n306147 );
not ( n24247 , n314672 );
buf ( n314674 , n24247 );
buf ( n24249 , n314674 );
or ( n24250 , n314671 , n24249 );
nand ( n24251 , n24244 , n24250 );
buf ( n24252 , n24251 );
buf ( n314679 , n24252 );
and ( n24254 , n314663 , n314679 );
and ( n24255 , n314640 , n314662 );
or ( n314682 , n24254 , n24255 );
buf ( n314683 , n314682 );
buf ( n314684 , n314683 );
and ( n314685 , n24196 , n314684 );
and ( n314686 , n314583 , n314621 );
or ( n314687 , n314685 , n314686 );
buf ( n314688 , n314687 );
buf ( n314689 , n314688 );
xor ( n314690 , n314526 , n314689 );
xor ( n24265 , n305542 , n15160 );
xor ( n314692 , n24265 , n305683 );
buf ( n314693 , n314692 );
buf ( n314694 , n314693 );
and ( n24269 , n314690 , n314694 );
and ( n24270 , n314526 , n314689 );
or ( n24271 , n24269 , n24270 );
buf ( n314698 , n24271 );
buf ( n314699 , n314698 );
xor ( n24274 , n305688 , n305874 );
xor ( n24275 , n24274 , n306044 );
buf ( n314702 , n24275 );
buf ( n314703 , n314702 );
xor ( n24278 , n314699 , n314703 );
buf ( n314705 , n880 );
buf ( n314706 , n856 );
and ( n24281 , n314705 , n314706 );
not ( n24282 , n314705 );
buf ( n314709 , n15582 );
and ( n24284 , n24282 , n314709 );
nor ( n24285 , n24281 , n24284 );
buf ( n314712 , n24285 );
buf ( n314713 , n314712 );
not ( n314714 , n314713 );
buf ( n314715 , n304984 );
not ( n314716 , n314715 );
or ( n24291 , n314714 , n314716 );
buf ( n24292 , n304997 );
buf ( n24293 , n15625 );
nand ( n24294 , n24292 , n24293 );
buf ( n24295 , n24294 );
buf ( n314722 , n24295 );
nand ( n314723 , n24291 , n314722 );
buf ( n314724 , n314723 );
buf ( n314725 , n314724 );
buf ( n314726 , n313029 );
buf ( n314727 , n858 );
buf ( n314728 , n878 );
xor ( n314729 , n314727 , n314728 );
buf ( n314730 , n314729 );
buf ( n314731 , n314730 );
nand ( n24306 , n314726 , n314731 );
buf ( n314733 , n24306 );
buf ( n314734 , n314733 );
buf ( n314735 , n306089 );
not ( n24310 , n314735 );
buf ( n314737 , n306272 );
nand ( n24312 , n24310 , n314737 );
buf ( n314739 , n24312 );
buf ( n314740 , n314739 );
nand ( n24315 , n314734 , n314740 );
buf ( n314742 , n24315 );
buf ( n314743 , n314742 );
xor ( n24318 , n314725 , n314743 );
buf ( n314745 , n304912 );
not ( n24320 , n314745 );
buf ( n314747 , n24320 );
buf ( n314748 , n314747 );
buf ( n314749 , n305993 );
buf ( n314750 , n850 );
and ( n24325 , n314749 , n314750 );
buf ( n314752 , n304565 );
buf ( n314753 , n886 );
and ( n24328 , n314752 , n314753 );
nor ( n24329 , n24325 , n24328 );
buf ( n314756 , n24329 );
buf ( n314757 , n314756 );
or ( n24332 , n314748 , n314757 );
buf ( n314759 , n305363 );
buf ( n314760 , n305600 );
not ( n24335 , n314760 );
buf ( n314762 , n24335 );
buf ( n314763 , n314762 );
or ( n24338 , n314759 , n314763 );
nand ( n314765 , n24332 , n24338 );
buf ( n314766 , n314765 );
buf ( n314767 , n314766 );
and ( n314768 , n24318 , n314767 );
and ( n24343 , n314725 , n314743 );
or ( n24344 , n314768 , n24343 );
buf ( n314771 , n24344 );
xor ( n314772 , n306118 , n306142 );
xor ( n24347 , n314772 , n306163 );
and ( n314774 , n314771 , n24347 );
xor ( n314775 , n305617 , n305646 );
xor ( n24350 , n314775 , n305678 );
buf ( n314777 , n24350 );
xor ( n24352 , n306118 , n306142 );
xor ( n24353 , n24352 , n306163 );
and ( n24354 , n314777 , n24353 );
and ( n314781 , n314771 , n314777 );
or ( n314782 , n314774 , n24354 , n314781 );
buf ( n314783 , n314782 );
xor ( n314784 , n306102 , n306167 );
xor ( n314785 , n314784 , n306172 );
buf ( n314786 , n314785 );
buf ( n314787 , n314786 );
xor ( n24362 , n314783 , n314787 );
xor ( n24363 , n305879 , n305954 );
xor ( n314790 , n24363 , n306039 );
buf ( n314791 , n314790 );
buf ( n314792 , n314791 );
and ( n314793 , n24362 , n314792 );
and ( n314794 , n314783 , n314787 );
or ( n24369 , n314793 , n314794 );
buf ( n314796 , n24369 );
buf ( n314797 , n314796 );
and ( n24372 , n24278 , n314797 );
and ( n314799 , n314699 , n314703 );
or ( n314800 , n24372 , n314799 );
buf ( n314801 , n314800 );
buf ( n314802 , n314801 );
xor ( n314803 , n306049 , n306374 );
xor ( n24378 , n314803 , n306397 );
buf ( n314805 , n24378 );
buf ( n314806 , n314805 );
xor ( n24381 , n314478 , n314802 );
xor ( n314808 , n24381 , n314806 );
buf ( n314809 , n314808 );
xor ( n24384 , n314478 , n314802 );
and ( n314811 , n24384 , n314806 );
and ( n314812 , n314478 , n314802 );
or ( n24387 , n314811 , n314812 );
buf ( n314814 , n24387 );
and ( n314815 , n313567 , n313568 );
buf ( n314816 , n314815 );
buf ( n24391 , n314816 );
buf ( n314818 , n23553 );
not ( n24393 , n314818 );
buf ( n314820 , n15836 );
not ( n314821 , n314820 );
or ( n24396 , n24393 , n314821 );
xnor ( n314823 , n878 , n834 );
buf ( n314824 , n314823 );
not ( n24399 , n314824 );
buf ( n314826 , n304932 );
nand ( n314827 , n24399 , n314826 );
buf ( n314828 , n314827 );
buf ( n314829 , n314828 );
nand ( n314830 , n24396 , n314829 );
buf ( n314831 , n314830 );
buf ( n314832 , n314831 );
xor ( n314833 , n24391 , n314832 );
buf ( n314834 , n313832 );
not ( n24409 , n314834 );
buf ( n314836 , n310576 );
not ( n314837 , n314836 );
or ( n314838 , n24409 , n314837 );
buf ( n314839 , n310582 );
buf ( n314840 , n864 );
buf ( n314841 , n848 );
xor ( n24416 , n314840 , n314841 );
buf ( n314843 , n24416 );
buf ( n314844 , n314843 );
nand ( n314845 , n314839 , n314844 );
buf ( n314846 , n314845 );
buf ( n314847 , n314846 );
nand ( n24422 , n314838 , n314847 );
buf ( n314849 , n24422 );
buf ( n314850 , n314849 );
xor ( n24425 , n314833 , n314850 );
buf ( n314852 , n24425 );
buf ( n314853 , n314852 );
buf ( n314854 , n14959 );
not ( n24429 , n314854 );
buf ( n314856 , n305381 );
not ( n24431 , n314856 );
or ( n24432 , n24429 , n24431 );
buf ( n314859 , n882 );
nand ( n24434 , n24432 , n314859 );
buf ( n314861 , n24434 );
buf ( n314862 , n314861 );
buf ( n314863 , n305650 );
buf ( n314864 , n313897 );
or ( n314865 , n314863 , n314864 );
buf ( n314866 , n876 );
buf ( n314867 , n311204 );
and ( n24442 , n314866 , n314867 );
not ( n314869 , n314866 );
buf ( n314870 , n836 );
and ( n24445 , n314869 , n314870 );
nor ( n24446 , n24442 , n24445 );
buf ( n314873 , n24446 );
buf ( n314874 , n314873 );
buf ( n314875 , n305664 );
or ( n24450 , n314874 , n314875 );
nand ( n24451 , n314865 , n24450 );
buf ( n314878 , n24451 );
buf ( n314879 , n314878 );
xor ( n24454 , n314862 , n314879 );
buf ( n314881 , n304987 );
buf ( n314882 , n314209 );
or ( n314883 , n314881 , n314882 );
buf ( n314884 , n304976 );
buf ( n314885 , n21800 );
buf ( n314886 , n832 );
and ( n314887 , n314885 , n314886 );
buf ( n314888 , n20700 );
buf ( n314889 , n880 );
and ( n314890 , n314888 , n314889 );
nor ( n314891 , n314887 , n314890 );
buf ( n314892 , n314891 );
buf ( n314893 , n314892 );
or ( n314894 , n314884 , n314893 );
nand ( n24469 , n314883 , n314894 );
buf ( n314896 , n24469 );
buf ( n314897 , n314896 );
xor ( n314898 , n24454 , n314897 );
buf ( n314899 , n314898 );
buf ( n314900 , n314899 );
xor ( n314901 , n314853 , n314900 );
buf ( n314902 , n23449 );
not ( n314903 , n314902 );
buf ( n314904 , n310694 );
not ( n314905 , n314904 );
or ( n24480 , n314903 , n314905 );
buf ( n314907 , n866 );
buf ( n314908 , n846 );
xnor ( n314909 , n314907 , n314908 );
buf ( n314910 , n314909 );
buf ( n314911 , n314910 );
not ( n24486 , n314911 );
buf ( n314913 , n311107 );
nand ( n24488 , n24486 , n314913 );
buf ( n314915 , n24488 );
buf ( n314916 , n314915 );
nand ( n314917 , n24480 , n314916 );
buf ( n314918 , n314917 );
buf ( n314919 , n314918 );
buf ( n314920 , n313854 );
not ( n24495 , n314920 );
buf ( n314922 , n305627 );
not ( n314923 , n314922 );
or ( n24498 , n24495 , n314923 );
buf ( n314925 , n874 );
buf ( n314926 , n310377 );
and ( n24501 , n314925 , n314926 );
not ( n314928 , n314925 );
buf ( n314929 , n838 );
and ( n314930 , n314928 , n314929 );
nor ( n24505 , n24501 , n314930 );
buf ( n314932 , n24505 );
buf ( n314933 , n314932 );
not ( n24508 , n314933 );
buf ( n314935 , n305301 );
nand ( n314936 , n24508 , n314935 );
buf ( n314937 , n314936 );
buf ( n314938 , n314937 );
nand ( n24513 , n24498 , n314938 );
buf ( n314940 , n24513 );
buf ( n314941 , n314940 );
xor ( n314942 , n314919 , n314941 );
buf ( n314943 , n310726 );
buf ( n314944 , n313927 );
or ( n314945 , n314943 , n314944 );
buf ( n314946 , n305449 );
buf ( n314947 , n868 );
buf ( n314948 , n844 );
and ( n24523 , n314947 , n314948 );
not ( n314950 , n314947 );
buf ( n314951 , n305458 );
and ( n24526 , n314950 , n314951 );
nor ( n314953 , n24523 , n24526 );
buf ( n314954 , n314953 );
buf ( n314955 , n314954 );
not ( n314956 , n314955 );
buf ( n314957 , n314956 );
buf ( n314958 , n314957 );
or ( n314959 , n314946 , n314958 );
nand ( n24534 , n314945 , n314959 );
buf ( n314961 , n24534 );
buf ( n314962 , n314961 );
xor ( n314963 , n314942 , n314962 );
buf ( n314964 , n314963 );
buf ( n314965 , n314964 );
and ( n314966 , n314901 , n314965 );
and ( n24541 , n314853 , n314900 );
or ( n314968 , n314966 , n24541 );
buf ( n314969 , n314968 );
buf ( n24544 , n314969 );
buf ( n314971 , n304981 );
buf ( n314972 , n314892 );
or ( n314973 , n314971 , n314972 );
buf ( n314974 , n311075 );
buf ( n314975 , n21800 );
or ( n314976 , n314974 , n314975 );
nand ( n314977 , n314973 , n314976 );
buf ( n314978 , n314977 );
buf ( n314979 , n314978 );
not ( n314980 , n314979 );
buf ( n314981 , n314980 );
buf ( n314982 , n314981 );
xor ( n24557 , n314862 , n314879 );
and ( n24558 , n24557 , n314897 );
and ( n314985 , n314862 , n314879 );
or ( n314986 , n24558 , n314985 );
buf ( n314987 , n314986 );
buf ( n314988 , n314987 );
xor ( n314989 , n314982 , n314988 );
xor ( n24564 , n314919 , n314941 );
and ( n314991 , n24564 , n314962 );
and ( n24566 , n314919 , n314941 );
or ( n314993 , n314991 , n24566 );
buf ( n314994 , n314993 );
buf ( n314995 , n314994 );
xor ( n314996 , n314989 , n314995 );
buf ( n314997 , n314996 );
buf ( n314998 , n314997 );
xor ( n314999 , n24544 , n314998 );
xor ( n24574 , n24391 , n314832 );
and ( n24575 , n24574 , n314850 );
and ( n315002 , n24391 , n314832 );
or ( n315003 , n24575 , n315002 );
buf ( n315004 , n315003 );
buf ( n315005 , n315004 );
and ( n315006 , n313829 , n313830 );
buf ( n315007 , n315006 );
buf ( n315008 , n315007 );
buf ( n315009 , n306132 );
buf ( n315010 , n872 );
buf ( n315011 , n840 );
xor ( n315012 , n315010 , n315011 );
buf ( n315013 , n315012 );
buf ( n315014 , n315013 );
nand ( n315015 , n315009 , n315014 );
buf ( n315016 , n315015 );
buf ( n315017 , n315016 );
buf ( n315018 , n304845 );
buf ( n315019 , n839 );
buf ( n315020 , n872 );
xor ( n24595 , n315019 , n315020 );
buf ( n315022 , n24595 );
buf ( n315023 , n315022 );
nand ( n24598 , n315018 , n315023 );
buf ( n315025 , n24598 );
buf ( n315026 , n315025 );
nand ( n24601 , n315017 , n315026 );
buf ( n315028 , n24601 );
buf ( n315029 , n315028 );
xor ( n24604 , n315008 , n315029 );
buf ( n315031 , n304941 );
buf ( n315032 , n314823 );
or ( n24607 , n315031 , n315032 );
buf ( n315034 , n14523 );
buf ( n315035 , n878 );
buf ( n315036 , n310964 );
and ( n315037 , n315035 , n315036 );
not ( n315038 , n315035 );
buf ( n315039 , n833 );
and ( n24614 , n315038 , n315039 );
nor ( n315041 , n315037 , n24614 );
buf ( n315042 , n315041 );
buf ( n315043 , n315042 );
or ( n315044 , n315034 , n315043 );
nand ( n24619 , n24607 , n315044 );
buf ( n315046 , n24619 );
buf ( n315047 , n315046 );
xor ( n24622 , n24604 , n315047 );
buf ( n315049 , n24622 );
buf ( n315050 , n315049 );
xor ( n24625 , n315005 , n315050 );
buf ( n315052 , n314843 );
not ( n24627 , n315052 );
buf ( n315054 , n310576 );
not ( n24629 , n315054 );
or ( n315056 , n24627 , n24629 );
buf ( n315057 , n864 );
buf ( n315058 , n847 );
xnor ( n315059 , n315057 , n315058 );
buf ( n315060 , n315059 );
buf ( n315061 , n315060 );
not ( n315062 , n315061 );
buf ( n315063 , n310582 );
nand ( n315064 , n315062 , n315063 );
buf ( n315065 , n315064 );
buf ( n315066 , n315065 );
nand ( n315067 , n315056 , n315066 );
buf ( n315068 , n315067 );
buf ( n315069 , n315068 );
buf ( n315070 , n313215 );
buf ( n315071 , n314910 );
or ( n24646 , n315070 , n315071 );
buf ( n315073 , n313224 );
buf ( n315074 , n845 );
buf ( n315075 , n866 );
xnor ( n315076 , n315074 , n315075 );
buf ( n315077 , n315076 );
buf ( n315078 , n315077 );
or ( n315079 , n315073 , n315078 );
nand ( n315080 , n24646 , n315079 );
buf ( n315081 , n315080 );
buf ( n315082 , n315081 );
xor ( n24657 , n315069 , n315082 );
buf ( n315084 , n306340 );
buf ( n315085 , n314932 );
or ( n24660 , n315084 , n315085 );
buf ( n315087 , n306346 );
buf ( n315088 , n874 );
not ( n24663 , n315088 );
buf ( n315090 , n24663 );
buf ( n315091 , n315090 );
buf ( n315092 , n837 );
and ( n24667 , n315091 , n315092 );
buf ( n315094 , n313757 );
buf ( n315095 , n874 );
and ( n24670 , n315094 , n315095 );
nor ( n24671 , n24667 , n24670 );
buf ( n315098 , n24671 );
buf ( n315099 , n315098 );
or ( n315100 , n315087 , n315099 );
nand ( n24675 , n24660 , n315100 );
buf ( n315102 , n24675 );
buf ( n315103 , n315102 );
xor ( n24678 , n24657 , n315103 );
buf ( n315105 , n24678 );
buf ( n315106 , n315105 );
xor ( n315107 , n24625 , n315106 );
buf ( n315108 , n315107 );
buf ( n315109 , n315108 );
xor ( n24684 , n314999 , n315109 );
buf ( n315111 , n24684 );
buf ( n315112 , n315111 );
xor ( n24687 , n314216 , n23812 );
and ( n315114 , n24687 , n314244 );
and ( n315115 , n314216 , n23812 );
or ( n24690 , n315114 , n315115 );
buf ( n315117 , n24690 );
buf ( n315118 , n304754 );
not ( n24693 , n315118 );
buf ( n315120 , n24693 );
buf ( n315121 , n315120 );
buf ( n315122 , n314234 );
or ( n315123 , n315121 , n315122 );
buf ( n24698 , n314225 );
buf ( n315125 , n842 );
buf ( n315126 , n870 );
xnor ( n315127 , n315125 , n315126 );
buf ( n315128 , n315127 );
buf ( n315129 , n315128 );
or ( n24704 , n24698 , n315129 );
nand ( n315131 , n315123 , n24704 );
buf ( n315132 , n315131 );
buf ( n315133 , n315132 );
buf ( n315134 , n304854 );
buf ( n315135 , n313945 );
or ( n24710 , n315134 , n315135 );
buf ( n315137 , n14439 );
buf ( n315138 , n315013 );
not ( n24713 , n315138 );
buf ( n24714 , n24713 );
buf ( n315141 , n24714 );
or ( n24716 , n315137 , n315141 );
nand ( n315143 , n24710 , n24716 );
buf ( n315144 , n315143 );
buf ( n315145 , n315144 );
xor ( n24720 , n315133 , n315145 );
buf ( n315147 , n314213 );
xor ( n24722 , n24720 , n315147 );
buf ( n315149 , n24722 );
buf ( n315150 , n315149 );
xor ( n24725 , n315117 , n315150 );
xor ( n315152 , n314265 , n314270 );
and ( n315153 , n315152 , n314277 );
and ( n24728 , n314265 , n314270 );
or ( n315155 , n315153 , n24728 );
buf ( n315156 , n315155 );
buf ( n315157 , n315156 );
and ( n315158 , n24725 , n315157 );
and ( n315159 , n315117 , n315150 );
or ( n24734 , n315158 , n315159 );
buf ( n315161 , n24734 );
buf ( n315162 , n315161 );
buf ( n315163 , n314219 );
buf ( n315164 , n315128 );
or ( n315165 , n315163 , n315164 );
buf ( n315166 , n304760 );
buf ( n315167 , n841 );
buf ( n315168 , n870 );
xnor ( n315169 , n315167 , n315168 );
buf ( n315170 , n315169 );
buf ( n315171 , n315170 );
or ( n24746 , n315166 , n315171 );
nand ( n24747 , n315165 , n24746 );
buf ( n315174 , n24747 );
buf ( n315175 , n314954 );
not ( n24750 , n315175 );
buf ( n315177 , n305213 );
not ( n315178 , n315177 );
or ( n24753 , n24750 , n315178 );
buf ( n315180 , n843 );
buf ( n315181 , n868 );
xnor ( n24756 , n315180 , n315181 );
buf ( n315183 , n24756 );
buf ( n315184 , n315183 );
not ( n24759 , n315184 );
buf ( n315186 , n305202 );
nand ( n315187 , n24759 , n315186 );
buf ( n315188 , n315187 );
buf ( n315189 , n315188 );
nand ( n24764 , n24753 , n315189 );
buf ( n315191 , n24764 );
xor ( n315192 , n315174 , n315191 );
buf ( n315193 , n305650 );
buf ( n315194 , n314873 );
or ( n315195 , n315193 , n315194 );
buf ( n24770 , n305664 );
buf ( n315197 , n876 );
buf ( n315198 , n21261 );
and ( n315199 , n315197 , n315198 );
not ( n24774 , n315197 );
buf ( n315201 , n835 );
and ( n315202 , n24774 , n315201 );
nor ( n315203 , n315199 , n315202 );
buf ( n315204 , n315203 );
buf ( n315205 , n315204 );
or ( n315206 , n24770 , n315205 );
nand ( n24781 , n315195 , n315206 );
buf ( n24782 , n24781 );
xor ( n315209 , n315192 , n24782 );
xor ( n24784 , n315133 , n315145 );
and ( n315211 , n24784 , n315147 );
and ( n24786 , n315133 , n315145 );
or ( n24787 , n315211 , n24786 );
buf ( n315214 , n24787 );
xor ( n315215 , n313822 , n313839 );
and ( n24790 , n315215 , n313861 );
and ( n315217 , n313822 , n313839 );
or ( n315218 , n24790 , n315217 );
buf ( n315219 , n315218 );
buf ( n315220 , n315219 );
xor ( n315221 , n313954 , n313967 );
and ( n24796 , n315221 , n313988 );
and ( n315223 , n313954 , n313967 );
or ( n315224 , n24796 , n315223 );
buf ( n315225 , n315224 );
buf ( n315226 , n315225 );
xor ( n315227 , n315220 , n315226 );
xor ( n24802 , n313889 , n313914 );
and ( n24803 , n24802 , n313932 );
and ( n24804 , n313889 , n313914 );
or ( n315231 , n24803 , n24804 );
buf ( n315232 , n315231 );
buf ( n315233 , n315232 );
and ( n24808 , n315227 , n315233 );
and ( n24809 , n315220 , n315226 );
or ( n315236 , n24808 , n24809 );
buf ( n315237 , n315236 );
xor ( n24812 , n315214 , n315237 );
xor ( n315239 , n315209 , n24812 );
buf ( n315240 , n315239 );
xor ( n315241 , n315162 , n315240 );
xor ( n24816 , n313864 , n313935 );
and ( n315243 , n24816 , n313991 );
and ( n24818 , n313864 , n313935 );
or ( n315245 , n315243 , n24818 );
buf ( n315246 , n315245 );
buf ( n315247 , n315246 );
xor ( n315248 , n315220 , n315226 );
xor ( n315249 , n315248 , n315233 );
buf ( n315250 , n315249 );
buf ( n315251 , n315250 );
xor ( n315252 , n315247 , n315251 );
xor ( n24827 , n314853 , n314900 );
xor ( n24828 , n24827 , n314965 );
buf ( n315255 , n24828 );
buf ( n315256 , n315255 );
and ( n315257 , n315252 , n315256 );
and ( n24832 , n315247 , n315251 );
or ( n24833 , n315257 , n24832 );
buf ( n315260 , n24833 );
buf ( n315261 , n315260 );
xor ( n315262 , n315241 , n315261 );
buf ( n315263 , n315262 );
buf ( n315264 , n315263 );
xor ( n24839 , n314216 , n23812 );
xor ( n315266 , n24839 , n314244 );
and ( n24841 , n314250 , n315266 );
xor ( n24842 , n314216 , n23812 );
xor ( n315269 , n24842 , n314244 );
and ( n315270 , n314279 , n315269 );
and ( n24845 , n314250 , n314279 );
or ( n24846 , n24841 , n315270 , n24845 );
buf ( n315273 , n24846 );
xor ( n315274 , n315117 , n315150 );
xor ( n315275 , n315274 , n315157 );
buf ( n315276 , n315275 );
buf ( n315277 , n315276 );
xor ( n315278 , n315273 , n315277 );
xor ( n24853 , n315247 , n315251 );
xor ( n315280 , n24853 , n315256 );
buf ( n315281 , n315280 );
buf ( n315282 , n315281 );
and ( n315283 , n315278 , n315282 );
and ( n24858 , n315273 , n315277 );
or ( n315285 , n315283 , n24858 );
buf ( n315286 , n315285 );
buf ( n315287 , n315286 );
xor ( n315288 , n315112 , n315264 );
xor ( n24863 , n315288 , n315287 );
buf ( n315290 , n24863 );
xor ( n315291 , n315112 , n315264 );
and ( n315292 , n315291 , n315287 );
and ( n315293 , n315112 , n315264 );
or ( n24868 , n315292 , n315293 );
buf ( n315295 , n24868 );
xor ( n315296 , n314783 , n314787 );
xor ( n24871 , n315296 , n314792 );
buf ( n315298 , n24871 );
buf ( n315299 , n315298 );
xor ( n24874 , n306066 , n306083 );
xor ( n315301 , n24874 , n306097 );
buf ( n315302 , n315301 );
xor ( n315303 , n314501 , n314517 );
xor ( n24878 , n315303 , n314521 );
buf ( n315305 , n24878 );
xor ( n315306 , n315302 , n315305 );
buf ( n315307 , n863 );
buf ( n315308 , n875 );
or ( n24883 , n315307 , n315308 );
buf ( n315310 , n876 );
nand ( n315311 , n24883 , n315310 );
buf ( n315312 , n315311 );
buf ( n315313 , n315312 );
buf ( n315314 , n863 );
buf ( n315315 , n875 );
nand ( n315316 , n315314 , n315315 );
buf ( n315317 , n315316 );
buf ( n315318 , n315317 );
buf ( n315319 , n874 );
and ( n24894 , n315313 , n315318 , n315319 );
buf ( n24895 , n24894 );
buf ( n315322 , n24895 );
buf ( n24897 , n892 );
buf ( n24898 , n845 );
xor ( n24899 , n24897 , n24898 );
buf ( n24900 , n24899 );
buf ( n24901 , n24900 );
not ( n24902 , n24901 );
buf ( n24903 , n14272 );
not ( n24904 , n24903 );
or ( n24905 , n24902 , n24904 );
buf ( n315332 , n24182 );
not ( n315333 , n315332 );
buf ( n24908 , n304694 );
nand ( n24909 , n315333 , n24908 );
buf ( n24910 , n24909 );
buf ( n315337 , n24910 );
nand ( n24912 , n24905 , n315337 );
buf ( n24913 , n24912 );
buf ( n315340 , n24913 );
and ( n24915 , n315322 , n315340 );
buf ( n315342 , n24915 );
buf ( n315343 , n315342 );
buf ( n315344 , n876 );
buf ( n315345 , n861 );
xor ( n24920 , n315344 , n315345 );
buf ( n315347 , n24920 );
buf ( n315348 , n315347 );
not ( n315349 , n315348 );
buf ( n315350 , n305338 );
not ( n315351 , n315350 );
or ( n315352 , n315349 , n315351 );
buf ( n315353 , n314570 );
not ( n315354 , n315353 );
buf ( n315355 , n305344 );
nand ( n24930 , n315354 , n315355 );
buf ( n315357 , n24930 );
buf ( n315358 , n315357 );
nand ( n315359 , n315352 , n315358 );
buf ( n315360 , n315359 );
buf ( n315361 , n315360 );
buf ( n315362 , n305192 );
buf ( n315363 , n874 );
or ( n315364 , n315362 , n315363 );
buf ( n24939 , n315090 );
buf ( n315366 , n863 );
or ( n315367 , n24939 , n315366 );
nand ( n315368 , n315364 , n315367 );
buf ( n315369 , n315368 );
buf ( n315370 , n315369 );
not ( n24945 , n315370 );
buf ( n315372 , n305627 );
not ( n315373 , n315372 );
or ( n24948 , n24945 , n315373 );
buf ( n315375 , n305301 );
buf ( n315376 , n314551 );
nand ( n24951 , n315375 , n315376 );
buf ( n315378 , n24951 );
buf ( n315379 , n315378 );
nand ( n315380 , n24948 , n315379 );
buf ( n315381 , n315380 );
buf ( n315382 , n315381 );
xor ( n315383 , n315361 , n315382 );
buf ( n315384 , n314747 );
buf ( n315385 , n886 );
buf ( n315386 , n305532 );
and ( n24961 , n315385 , n315386 );
not ( n315388 , n315385 );
buf ( n315389 , n851 );
and ( n24964 , n315388 , n315389 );
nor ( n315391 , n24961 , n24964 );
buf ( n315392 , n315391 );
buf ( n315393 , n315392 );
or ( n315394 , n315384 , n315393 );
buf ( n315395 , n305363 );
buf ( n315396 , n314756 );
or ( n315397 , n315395 , n315396 );
nand ( n24972 , n315394 , n315397 );
buf ( n315399 , n24972 );
buf ( n315400 , n315399 );
and ( n315401 , n315383 , n315400 );
and ( n315402 , n315361 , n315382 );
or ( n24977 , n315401 , n315402 );
buf ( n315404 , n24977 );
buf ( n24979 , n315404 );
xor ( n24980 , n315343 , n24979 );
buf ( n315407 , n305881 );
buf ( n315408 , n843 );
buf ( n315409 , n894 );
xor ( n315410 , n315408 , n315409 );
buf ( n315411 , n315410 );
buf ( n315412 , n315411 );
not ( n315413 , n315412 );
buf ( n315414 , n315413 );
buf ( n315415 , n315414 );
or ( n24990 , n315407 , n315415 );
buf ( n315417 , n314530 );
not ( n315418 , n315417 );
buf ( n315419 , n315418 );
buf ( n315420 , n315419 );
buf ( n315421 , n15469 );
or ( n24996 , n315420 , n315421 );
nand ( n24997 , n24990 , n24996 );
buf ( n315424 , n24997 );
buf ( n315425 , n315424 );
buf ( n315426 , n884 );
buf ( n315427 , n853 );
and ( n25002 , n315426 , n315427 );
not ( n25003 , n315426 );
buf ( n315430 , n304956 );
and ( n315431 , n25003 , n315430 );
nor ( n315432 , n25002 , n315431 );
buf ( n315433 , n315432 );
buf ( n315434 , n315433 );
not ( n315435 , n315434 );
buf ( n315436 , n304813 );
not ( n25011 , n315436 );
or ( n315438 , n315435 , n25011 );
buf ( n315439 , n304807 );
buf ( n315440 , n314648 );
nand ( n315441 , n315439 , n315440 );
buf ( n315442 , n315441 );
buf ( n315443 , n315442 );
nand ( n315444 , n315438 , n315443 );
buf ( n315445 , n315444 );
buf ( n315446 , n315445 );
xor ( n25021 , n315425 , n315446 );
buf ( n315448 , n847 );
buf ( n315449 , n890 );
and ( n25024 , n315448 , n315449 );
not ( n315451 , n315448 );
buf ( n25026 , n312467 );
and ( n315453 , n315451 , n25026 );
nor ( n25028 , n25024 , n315453 );
buf ( n25029 , n25028 );
buf ( n315456 , n25029 );
not ( n25031 , n315456 );
buf ( n315458 , n304633 );
not ( n25033 , n315458 );
or ( n25034 , n25031 , n25033 );
buf ( n315461 , n314668 );
not ( n315462 , n315461 );
buf ( n25037 , n304658 );
nand ( n25038 , n315462 , n25037 );
buf ( n25039 , n25038 );
buf ( n315466 , n25039 );
nand ( n315467 , n25034 , n315466 );
buf ( n315468 , n315467 );
buf ( n315469 , n315468 );
and ( n315470 , n25021 , n315469 );
and ( n315471 , n315425 , n315446 );
or ( n25046 , n315470 , n315471 );
buf ( n315473 , n25046 );
buf ( n315474 , n315473 );
and ( n25049 , n24980 , n315474 );
and ( n315476 , n315343 , n24979 );
or ( n315477 , n25049 , n315476 );
buf ( n315478 , n315477 );
and ( n25053 , n315306 , n315478 );
and ( n315480 , n315302 , n315305 );
or ( n315481 , n25053 , n315480 );
buf ( n315482 , n315481 );
xor ( n315483 , n314526 , n314689 );
xor ( n315484 , n315483 , n314694 );
buf ( n315485 , n315484 );
buf ( n315486 , n315485 );
xor ( n315487 , n315482 , n315486 );
xor ( n25062 , n314583 , n314621 );
xor ( n315489 , n25062 , n314684 );
buf ( n315490 , n315489 );
buf ( n315491 , n315490 );
buf ( n315492 , n849 );
buf ( n315493 , n888 );
xor ( n25068 , n315492 , n315493 );
buf ( n315495 , n25068 );
buf ( n315496 , n315495 );
not ( n25071 , n315496 );
buf ( n315498 , n305138 );
not ( n315499 , n315498 );
or ( n315500 , n25071 , n315499 );
buf ( n315501 , n305144 );
buf ( n315502 , n24163 );
nand ( n315503 , n315501 , n315502 );
buf ( n315504 , n315503 );
buf ( n315505 , n315504 );
nand ( n315506 , n315500 , n315505 );
buf ( n315507 , n315506 );
buf ( n315508 , n315507 );
buf ( n315509 , n859 );
buf ( n315510 , n878 );
xor ( n315511 , n315509 , n315510 );
buf ( n315512 , n315511 );
buf ( n315513 , n315512 );
not ( n315514 , n315513 );
buf ( n315515 , n15836 );
not ( n315516 , n315515 );
or ( n25091 , n315514 , n315516 );
buf ( n315518 , n304932 );
buf ( n315519 , n314730 );
nand ( n315520 , n315518 , n315519 );
buf ( n315521 , n315520 );
buf ( n315522 , n315521 );
nand ( n315523 , n25091 , n315522 );
buf ( n315524 , n315523 );
buf ( n315525 , n315524 );
xor ( n315526 , n315508 , n315525 );
buf ( n315527 , n304987 );
buf ( n315528 , n21800 );
buf ( n315529 , n857 );
and ( n315530 , n315528 , n315529 );
buf ( n315531 , n305939 );
buf ( n315532 , n880 );
and ( n25107 , n315531 , n315532 );
nor ( n315534 , n315530 , n25107 );
buf ( n315535 , n315534 );
buf ( n315536 , n315535 );
or ( n315537 , n315527 , n315536 );
buf ( n315538 , n311075 );
buf ( n315539 , n314712 );
not ( n315540 , n315539 );
buf ( n315541 , n315540 );
buf ( n315542 , n315541 );
or ( n315543 , n315538 , n315542 );
nand ( n315544 , n315537 , n315543 );
buf ( n315545 , n315544 );
buf ( n315546 , n315545 );
and ( n315547 , n315526 , n315546 );
and ( n25122 , n315508 , n315525 );
or ( n315549 , n315547 , n25122 );
buf ( n315550 , n315549 );
buf ( n315551 , n315550 );
xor ( n315552 , n314640 , n314662 );
xor ( n315553 , n315552 , n314679 );
buf ( n315554 , n315553 );
buf ( n315555 , n315554 );
xor ( n25130 , n315551 , n315555 );
xor ( n25131 , n314725 , n314743 );
xor ( n315558 , n25131 , n314767 );
buf ( n315559 , n315558 );
buf ( n315560 , n315559 );
and ( n315561 , n25130 , n315560 );
and ( n315562 , n315551 , n315555 );
or ( n25137 , n315561 , n315562 );
buf ( n315564 , n25137 );
buf ( n315565 , n315564 );
xor ( n315566 , n315491 , n315565 );
xor ( n315567 , n306118 , n306142 );
xor ( n25142 , n315567 , n306163 );
xor ( n315569 , n314771 , n314777 );
xor ( n315570 , n25142 , n315569 );
buf ( n315571 , n315570 );
and ( n315572 , n315566 , n315571 );
and ( n25147 , n315491 , n315565 );
or ( n25148 , n315572 , n25147 );
buf ( n315575 , n25148 );
buf ( n315576 , n315575 );
xor ( n25151 , n315487 , n315576 );
buf ( n315578 , n25151 );
buf ( n315579 , n315578 );
xor ( n25154 , n314588 , n314602 );
xor ( n315581 , n25154 , n314616 );
buf ( n315582 , n315581 );
buf ( n315583 , n315582 );
xor ( n315584 , n314543 , n314564 );
xor ( n315585 , n315584 , n314578 );
buf ( n315586 , n315585 );
buf ( n315587 , n315586 );
xor ( n315588 , n315583 , n315587 );
buf ( n315589 , n305381 );
buf ( n315590 , n882 );
buf ( n315591 , n855 );
xnor ( n315592 , n315590 , n315591 );
buf ( n315593 , n315592 );
buf ( n315594 , n315593 );
or ( n25169 , n315589 , n315594 );
buf ( n315596 , n14959 );
buf ( n25171 , n314626 );
not ( n315598 , n25171 );
buf ( n315599 , n315598 );
buf ( n315600 , n315599 );
or ( n315601 , n315596 , n315600 );
nand ( n25176 , n25169 , n315601 );
buf ( n25177 , n25176 );
buf ( n25178 , n25177 );
xor ( n25179 , n315322 , n315340 );
buf ( n315606 , n25179 );
buf ( n315607 , n315606 );
xor ( n25182 , n25178 , n315607 );
xor ( n315609 , n892 , n846 );
buf ( n315610 , n315609 );
not ( n315611 , n315610 );
buf ( n315612 , n304697 );
not ( n25187 , n315612 );
or ( n315614 , n315611 , n25187 );
buf ( n315615 , n24900 );
buf ( n315616 , n304694 );
nand ( n25191 , n315615 , n315616 );
buf ( n315618 , n25191 );
buf ( n25193 , n315618 );
nand ( n25194 , n315614 , n25193 );
buf ( n25195 , n25194 );
buf ( n25196 , n25195 );
buf ( n315623 , n860 );
buf ( n315624 , n878 );
xnor ( n315625 , n315623 , n315624 );
buf ( n315626 , n315625 );
buf ( n315627 , n315626 );
not ( n25202 , n315627 );
buf ( n25203 , n25202 );
buf ( n25204 , n25203 );
not ( n25205 , n25204 );
buf ( n25206 , n313029 );
not ( n25207 , n25206 );
or ( n25208 , n25205 , n25207 );
buf ( n25209 , n315512 );
buf ( n25210 , n306272 );
nand ( n25211 , n25209 , n25210 );
buf ( n25212 , n25211 );
buf ( n25213 , n25212 );
nand ( n25214 , n25208 , n25213 );
buf ( n25215 , n25214 );
buf ( n315642 , n25215 );
xor ( n25217 , n25196 , n315642 );
buf ( n315644 , n304981 );
buf ( n315645 , n880 );
buf ( n315646 , n858 );
xnor ( n315647 , n315645 , n315646 );
buf ( n315648 , n315647 );
buf ( n315649 , n315648 );
or ( n315650 , n315644 , n315649 );
buf ( n315651 , n311075 );
buf ( n315652 , n315535 );
or ( n315653 , n315651 , n315652 );
nand ( n315654 , n315650 , n315653 );
buf ( n315655 , n315654 );
buf ( n315656 , n315655 );
and ( n315657 , n25217 , n315656 );
and ( n315658 , n25196 , n315642 );
or ( n25233 , n315657 , n315658 );
buf ( n315660 , n25233 );
buf ( n315661 , n315660 );
and ( n25236 , n25182 , n315661 );
and ( n315663 , n25178 , n315607 );
or ( n315664 , n25236 , n315663 );
buf ( n315665 , n315664 );
buf ( n315666 , n315665 );
and ( n315667 , n315588 , n315666 );
and ( n25242 , n315583 , n315587 );
or ( n315669 , n315667 , n25242 );
buf ( n315670 , n315669 );
xor ( n25245 , n315302 , n315305 );
xor ( n315672 , n25245 , n315478 );
and ( n25247 , n315670 , n315672 );
xor ( n315674 , n315491 , n315565 );
xor ( n315675 , n315674 , n315571 );
buf ( n315676 , n315675 );
xor ( n25251 , n315302 , n315305 );
xor ( n315678 , n25251 , n315478 );
and ( n315679 , n315676 , n315678 );
and ( n25254 , n315670 , n315676 );
or ( n315681 , n25247 , n315679 , n25254 );
buf ( n315682 , n315681 );
xor ( n25257 , n315299 , n315579 );
xor ( n315684 , n25257 , n315682 );
buf ( n315685 , n315684 );
xor ( n25260 , n315299 , n315579 );
and ( n315687 , n25260 , n315682 );
and ( n25262 , n315299 , n315579 );
or ( n315689 , n315687 , n25262 );
buf ( n315690 , n315689 );
xor ( n315691 , n313625 , n313818 );
and ( n25266 , n315691 , n313994 );
and ( n315693 , n313625 , n313818 );
or ( n315694 , n25266 , n315693 );
buf ( n315695 , n315694 );
buf ( n315696 , n315695 );
xor ( n315697 , n314282 , n314288 );
and ( n25272 , n315697 , n314309 );
and ( n315699 , n314282 , n314288 );
or ( n315700 , n25272 , n315699 );
buf ( n315701 , n315700 );
buf ( n315702 , n315701 );
xor ( n315703 , n315273 , n315277 );
xor ( n25278 , n315703 , n315282 );
buf ( n315705 , n25278 );
buf ( n315706 , n315705 );
xor ( n25281 , n315696 , n315702 );
xor ( n315708 , n25281 , n315706 );
buf ( n315709 , n315708 );
xor ( n25284 , n315696 , n315702 );
and ( n25285 , n25284 , n315706 );
and ( n315712 , n315696 , n315702 );
or ( n25287 , n25285 , n315712 );
buf ( n315714 , n25287 );
buf ( n25289 , n864 );
buf ( n315716 , n862 );
and ( n315717 , n25289 , n315716 );
buf ( n315718 , n315717 );
buf ( n315719 , n315718 );
buf ( n315720 , n864 );
buf ( n315721 , n861 );
xor ( n315722 , n315720 , n315721 );
buf ( n315723 , n315722 );
buf ( n315724 , n315723 );
not ( n315725 , n315724 );
buf ( n315726 , n311226 );
not ( n315727 , n315726 );
or ( n315728 , n315725 , n315727 );
buf ( n315729 , n310582 );
buf ( n315730 , n864 );
buf ( n315731 , n860 );
xor ( n25306 , n315730 , n315731 );
buf ( n315733 , n25306 );
buf ( n315734 , n315733 );
nand ( n25309 , n315729 , n315734 );
buf ( n315736 , n25309 );
buf ( n315737 , n315736 );
nand ( n315738 , n315728 , n315737 );
buf ( n315739 , n315738 );
buf ( n315740 , n315739 );
xor ( n315741 , n315719 , n315740 );
xor ( n25316 , n880 , n845 );
buf ( n315743 , n25316 );
not ( n315744 , n315743 );
buf ( n315745 , n305098 );
not ( n315746 , n315745 );
or ( n315747 , n315744 , n315746 );
buf ( n315748 , n304973 );
buf ( n315749 , n880 );
buf ( n315750 , n844 );
and ( n25325 , n315749 , n315750 );
not ( n315752 , n315749 );
buf ( n315753 , n305458 );
and ( n25328 , n315752 , n315753 );
nor ( n315755 , n25325 , n25328 );
buf ( n315756 , n315755 );
buf ( n25331 , n315756 );
nand ( n25332 , n315748 , n25331 );
buf ( n25333 , n25332 );
buf ( n315760 , n25333 );
nand ( n25335 , n315747 , n315760 );
buf ( n25336 , n25335 );
buf ( n315763 , n25336 );
xor ( n25338 , n315741 , n315763 );
buf ( n315765 , n25338 );
buf ( n315766 , n315765 );
xor ( n25341 , n874 , n852 );
buf ( n315768 , n25341 );
not ( n25343 , n315768 );
buf ( n315770 , n305624 );
not ( n315771 , n315770 );
or ( n25346 , n25343 , n315771 );
buf ( n315773 , n305301 );
buf ( n315774 , n851 );
buf ( n315775 , n874 );
xor ( n315776 , n315774 , n315775 );
buf ( n315777 , n315776 );
buf ( n315778 , n315777 );
nand ( n25353 , n315773 , n315778 );
buf ( n315780 , n25353 );
buf ( n315781 , n315780 );
nand ( n25356 , n25346 , n315781 );
buf ( n25357 , n25356 );
buf ( n25358 , n25357 );
buf ( n315785 , n890 );
buf ( n25360 , n836 );
and ( n25361 , n315785 , n25360 );
not ( n315788 , n315785 );
buf ( n315789 , n311204 );
and ( n25364 , n315788 , n315789 );
nor ( n315791 , n25361 , n25364 );
buf ( n315792 , n315791 );
buf ( n315793 , n315792 );
not ( n315794 , n315793 );
buf ( n315795 , n306152 );
not ( n315796 , n315795 );
or ( n25371 , n315794 , n315796 );
buf ( n315798 , n890 );
buf ( n25373 , n835 );
xor ( n25374 , n315798 , n25373 );
buf ( n25375 , n25374 );
buf ( n315802 , n25375 );
buf ( n315803 , n304658 );
nand ( n315804 , n315802 , n315803 );
buf ( n315805 , n315804 );
buf ( n315806 , n315805 );
nand ( n315807 , n25371 , n315806 );
buf ( n315808 , n315807 );
buf ( n315809 , n315808 );
xor ( n25384 , n25358 , n315809 );
buf ( n315811 , n884 );
buf ( n315812 , n842 );
and ( n315813 , n315811 , n315812 );
not ( n315814 , n315811 );
buf ( n315815 , n304610 );
and ( n315816 , n315814 , n315815 );
nor ( n315817 , n315813 , n315816 );
buf ( n315818 , n315817 );
buf ( n315819 , n315818 );
not ( n315820 , n315819 );
buf ( n315821 , n304813 );
not ( n315822 , n315821 );
or ( n315823 , n315820 , n315822 );
buf ( n315824 , n304819 );
and ( n25399 , n884 , n310600 );
not ( n25400 , n884 );
and ( n315827 , n25400 , n841 );
or ( n315828 , n25399 , n315827 );
buf ( n315829 , n315828 );
nand ( n25404 , n315824 , n315829 );
buf ( n315831 , n25404 );
buf ( n315832 , n315831 );
nand ( n25407 , n315823 , n315832 );
buf ( n315834 , n25407 );
buf ( n315835 , n315834 );
and ( n25410 , n25384 , n315835 );
and ( n315837 , n25358 , n315809 );
or ( n315838 , n25410 , n315837 );
buf ( n315839 , n315838 );
buf ( n315840 , n315839 );
xor ( n315841 , n315766 , n315840 );
buf ( n315842 , n855 );
buf ( n315843 , n870 );
xor ( n315844 , n315842 , n315843 );
buf ( n315845 , n315844 );
buf ( n315846 , n315845 );
not ( n315847 , n315846 );
buf ( n315848 , n20629 );
not ( n25423 , n315848 );
or ( n315850 , n315847 , n25423 );
buf ( n315851 , n311052 );
buf ( n315852 , n854 );
buf ( n315853 , n870 );
xor ( n315854 , n315852 , n315853 );
buf ( n315855 , n315854 );
buf ( n315856 , n315855 );
nand ( n25431 , n315851 , n315856 );
buf ( n315858 , n25431 );
buf ( n315859 , n315858 );
nand ( n25434 , n315850 , n315859 );
buf ( n315861 , n25434 );
buf ( n315862 , n315861 );
xor ( n25437 , n868 , n857 );
buf ( n315864 , n25437 );
not ( n315865 , n315864 );
buf ( n315866 , n305213 );
not ( n315867 , n315866 );
or ( n315868 , n315865 , n315867 );
buf ( n315869 , n305202 );
xor ( n315870 , n868 , n856 );
buf ( n315871 , n315870 );
nand ( n315872 , n315869 , n315871 );
buf ( n315873 , n315872 );
buf ( n315874 , n315873 );
nand ( n315875 , n315868 , n315874 );
buf ( n315876 , n315875 );
buf ( n315877 , n315876 );
xor ( n315878 , n315862 , n315877 );
buf ( n25453 , n882 );
buf ( n315880 , n843 );
xor ( n315881 , n25453 , n315880 );
buf ( n315882 , n315881 );
buf ( n315883 , n315882 );
not ( n315884 , n315883 );
buf ( n315885 , n304584 );
not ( n25460 , n315885 );
or ( n315887 , n315884 , n25460 );
buf ( n25462 , n304596 );
buf ( n315889 , n882 );
buf ( n315890 , n842 );
and ( n315891 , n315889 , n315890 );
not ( n25466 , n315889 );
buf ( n315893 , n304610 );
and ( n25468 , n25466 , n315893 );
nor ( n315895 , n315891 , n25468 );
buf ( n315896 , n315895 );
buf ( n315897 , n315896 );
nand ( n315898 , n25462 , n315897 );
buf ( n315899 , n315898 );
buf ( n315900 , n315899 );
nand ( n315901 , n315887 , n315900 );
buf ( n315902 , n315901 );
buf ( n315903 , n315902 );
xor ( n25478 , n315878 , n315903 );
buf ( n315905 , n25478 );
buf ( n315906 , n315905 );
xor ( n25481 , n315841 , n315906 );
buf ( n315908 , n25481 );
buf ( n315909 , n315908 );
buf ( n315910 , n315828 );
not ( n25485 , n315910 );
buf ( n315912 , n310401 );
not ( n315913 , n315912 );
or ( n25488 , n25485 , n315913 );
buf ( n315915 , n304807 );
buf ( n315916 , n840 );
buf ( n315917 , n884 );
xor ( n315918 , n315916 , n315917 );
buf ( n315919 , n315918 );
buf ( n315920 , n315919 );
nand ( n25495 , n315915 , n315920 );
buf ( n315922 , n25495 );
buf ( n315923 , n315922 );
nand ( n315924 , n25488 , n315923 );
buf ( n315925 , n315924 );
buf ( n315926 , n315925 );
buf ( n315927 , n25375 );
not ( n25502 , n315927 );
buf ( n315929 , n304633 );
not ( n315930 , n315929 );
or ( n25505 , n25502 , n315930 );
xor ( n315932 , n890 , n834 );
buf ( n315933 , n315932 );
buf ( n315934 , n304658 );
nand ( n315935 , n315933 , n315934 );
buf ( n315936 , n315935 );
buf ( n315937 , n315936 );
nand ( n25512 , n25505 , n315937 );
buf ( n315939 , n25512 );
buf ( n315940 , n315939 );
xor ( n25515 , n315926 , n315940 );
buf ( n315942 , n853 );
buf ( n315943 , n872 );
xor ( n25518 , n315942 , n315943 );
buf ( n25519 , n25518 );
buf ( n25520 , n25519 );
not ( n25521 , n25520 );
buf ( n315948 , n14420 );
not ( n25523 , n315948 );
or ( n315950 , n25521 , n25523 );
buf ( n315951 , n304845 );
buf ( n315952 , n872 );
buf ( n315953 , n852 );
xor ( n315954 , n315952 , n315953 );
buf ( n315955 , n315954 );
buf ( n315956 , n315955 );
nand ( n315957 , n315951 , n315956 );
buf ( n315958 , n315957 );
buf ( n315959 , n315958 );
nand ( n315960 , n315950 , n315959 );
buf ( n315961 , n315960 );
buf ( n315962 , n315961 );
xor ( n315963 , n25515 , n315962 );
buf ( n315964 , n315963 );
buf ( n315965 , n315964 );
buf ( n315966 , n878 );
buf ( n315967 , n847 );
and ( n25542 , n315966 , n315967 );
not ( n25543 , n315966 );
buf ( n315970 , n847 );
not ( n25545 , n315970 );
buf ( n315972 , n25545 );
buf ( n315973 , n315972 );
and ( n25548 , n25543 , n315973 );
nor ( n315975 , n25542 , n25548 );
buf ( n315976 , n315975 );
buf ( n315977 , n315976 );
not ( n25552 , n315977 );
buf ( n315979 , n15836 );
not ( n315980 , n315979 );
or ( n25555 , n25552 , n315980 );
buf ( n315982 , n306272 );
buf ( n315983 , n846 );
buf ( n315984 , n878 );
xor ( n315985 , n315983 , n315984 );
buf ( n315986 , n315985 );
buf ( n315987 , n315986 );
nand ( n315988 , n315982 , n315987 );
buf ( n315989 , n315988 );
buf ( n315990 , n315989 );
nand ( n315991 , n25555 , n315990 );
buf ( n315992 , n315991 );
buf ( n315993 , n315992 );
buf ( n315994 , n892 );
buf ( n315995 , n833 );
and ( n315996 , n315994 , n315995 );
not ( n315997 , n315994 );
buf ( n315998 , n310964 );
and ( n25573 , n315997 , n315998 );
nor ( n25574 , n315996 , n25573 );
buf ( n316001 , n25574 );
buf ( n316002 , n316001 );
not ( n25577 , n316002 );
buf ( n316004 , n14272 );
not ( n25579 , n316004 );
or ( n316006 , n25577 , n25579 );
buf ( n316007 , n304694 );
buf ( n316008 , n892 );
buf ( n316009 , n832 );
and ( n25584 , n316008 , n316009 );
not ( n316011 , n316008 );
buf ( n316012 , n20700 );
and ( n316013 , n316011 , n316012 );
nor ( n316014 , n25584 , n316013 );
buf ( n316015 , n316014 );
buf ( n316016 , n316015 );
nand ( n25591 , n316007 , n316016 );
buf ( n316018 , n25591 );
buf ( n316019 , n316018 );
nand ( n316020 , n316006 , n316019 );
buf ( n316021 , n316020 );
buf ( n316022 , n316021 );
xor ( n316023 , n315993 , n316022 );
and ( n25598 , n888 , n313757 );
not ( n316025 , n888 );
and ( n316026 , n316025 , n837 );
or ( n25601 , n25598 , n316026 );
buf ( n25602 , n25601 );
not ( n25603 , n25602 );
buf ( n25604 , n305138 );
not ( n25605 , n25604 );
or ( n25606 , n25603 , n25605 );
buf ( n25607 , n305144 );
buf ( n316034 , n888 );
buf ( n316035 , n836 );
and ( n316036 , n316034 , n316035 );
not ( n316037 , n316034 );
buf ( n316038 , n311204 );
and ( n316039 , n316037 , n316038 );
nor ( n316040 , n316036 , n316039 );
buf ( n316041 , n316040 );
buf ( n316042 , n316041 );
nand ( n316043 , n25607 , n316042 );
buf ( n316044 , n316043 );
buf ( n316045 , n316044 );
nand ( n316046 , n25606 , n316045 );
buf ( n316047 , n316046 );
buf ( n316048 , n316047 );
xor ( n25623 , n316023 , n316048 );
buf ( n316050 , n25623 );
buf ( n316051 , n316050 );
xor ( n25626 , n315965 , n316051 );
buf ( n316053 , n315777 );
not ( n316054 , n316053 );
buf ( n316055 , n305292 );
not ( n316056 , n316055 );
or ( n25631 , n316054 , n316056 );
buf ( n316058 , n850 );
buf ( n316059 , n874 );
xor ( n25634 , n316058 , n316059 );
buf ( n316061 , n25634 );
buf ( n316062 , n316061 );
buf ( n316063 , n305289 );
nand ( n316064 , n316062 , n316063 );
buf ( n316065 , n316064 );
buf ( n316066 , n316065 );
nand ( n25641 , n25631 , n316066 );
buf ( n25642 , n25641 );
buf ( n316069 , n25642 );
buf ( n316070 , n839 );
buf ( n316071 , n886 );
xor ( n316072 , n316070 , n316071 );
buf ( n316073 , n316072 );
buf ( n316074 , n316073 );
not ( n316075 , n316074 );
buf ( n316076 , n311697 );
not ( n316077 , n316076 );
or ( n316078 , n316075 , n316077 );
buf ( n316079 , n304901 );
xor ( n25654 , n886 , n838 );
buf ( n316081 , n25654 );
nand ( n25656 , n316079 , n316081 );
buf ( n316083 , n25656 );
buf ( n316084 , n316083 );
nand ( n316085 , n316078 , n316084 );
buf ( n316086 , n316085 );
buf ( n316087 , n316086 );
xor ( n25662 , n316069 , n316087 );
buf ( n316089 , n305650 );
buf ( n316090 , n849 );
buf ( n316091 , n876 );
xor ( n25666 , n316090 , n316091 );
buf ( n316093 , n25666 );
buf ( n316094 , n316093 );
not ( n316095 , n316094 );
buf ( n316096 , n316095 );
buf ( n316097 , n316096 );
or ( n25672 , n316089 , n316097 );
buf ( n25673 , n305664 );
buf ( n316100 , n876 );
buf ( n316101 , n848 );
xor ( n25676 , n316100 , n316101 );
buf ( n316103 , n25676 );
buf ( n25678 , n316103 );
not ( n316105 , n25678 );
buf ( n316106 , n316105 );
buf ( n316107 , n316106 );
or ( n316108 , n25673 , n316107 );
nand ( n316109 , n25672 , n316108 );
buf ( n316110 , n316109 );
buf ( n316111 , n316110 );
xor ( n25686 , n25662 , n316111 );
buf ( n316113 , n25686 );
buf ( n316114 , n316113 );
xor ( n316115 , n25626 , n316114 );
buf ( n316116 , n316115 );
buf ( n316117 , n316116 );
xor ( n316118 , n315909 , n316117 );
xor ( n25693 , n25289 , n315716 );
buf ( n316120 , n25693 );
buf ( n316121 , n316120 );
not ( n25696 , n316121 );
buf ( n316123 , n311888 );
not ( n25698 , n316123 );
or ( n316125 , n25696 , n25698 );
buf ( n316126 , n310582 );
buf ( n316127 , n315723 );
nand ( n316128 , n316126 , n316127 );
buf ( n316129 , n316128 );
buf ( n316130 , n316129 );
nand ( n316131 , n316125 , n316130 );
buf ( n316132 , n316131 );
buf ( n316133 , n316132 );
not ( n316134 , n316133 );
buf ( n316135 , n888 );
buf ( n316136 , n838 );
and ( n25711 , n316135 , n316136 );
not ( n25712 , n316135 );
buf ( n316139 , n310377 );
and ( n316140 , n25712 , n316139 );
nor ( n25715 , n25711 , n316140 );
buf ( n316142 , n25715 );
buf ( n316143 , n316142 );
not ( n316144 , n316143 );
buf ( n316145 , n311998 );
not ( n25720 , n316145 );
or ( n25721 , n316144 , n25720 );
buf ( n25722 , n305144 );
buf ( n316149 , n25601 );
nand ( n316150 , n25722 , n316149 );
buf ( n316151 , n316150 );
buf ( n316152 , n316151 );
nand ( n25727 , n25721 , n316152 );
buf ( n316154 , n25727 );
buf ( n316155 , n316154 );
buf ( n316156 , n880 );
buf ( n316157 , n846 );
and ( n25732 , n316156 , n316157 );
not ( n25733 , n316156 );
buf ( n25734 , n311024 );
and ( n316161 , n25733 , n25734 );
nor ( n316162 , n25732 , n316161 );
buf ( n316163 , n316162 );
buf ( n316164 , n316163 );
not ( n316165 , n316164 );
buf ( n316166 , n304984 );
not ( n316167 , n316166 );
or ( n316168 , n316165 , n316167 );
buf ( n316169 , n25316 );
buf ( n316170 , n304973 );
nand ( n316171 , n316169 , n316170 );
buf ( n316172 , n316171 );
buf ( n316173 , n316172 );
nand ( n25748 , n316168 , n316173 );
buf ( n316175 , n25748 );
buf ( n316176 , n316175 );
xnor ( n25751 , n316155 , n316176 );
buf ( n316178 , n25751 );
buf ( n316179 , n316178 );
not ( n316180 , n316179 );
or ( n25755 , n316134 , n316180 );
buf ( n316182 , n316178 );
buf ( n316183 , n316132 );
or ( n25758 , n316182 , n316183 );
nand ( n316185 , n25755 , n25758 );
buf ( n316186 , n316185 );
buf ( n316187 , n316186 );
buf ( n316188 , n313215 );
buf ( n316189 , n860 );
buf ( n316190 , n866 );
xor ( n316191 , n316189 , n316190 );
buf ( n316192 , n316191 );
buf ( n316193 , n316192 );
not ( n25768 , n316193 );
buf ( n316195 , n25768 );
buf ( n316196 , n316195 );
or ( n316197 , n316188 , n316196 );
buf ( n316198 , n310472 );
buf ( n316199 , n859 );
buf ( n316200 , n866 );
xor ( n316201 , n316199 , n316200 );
buf ( n316202 , n316201 );
buf ( n316203 , n316202 );
not ( n316204 , n316203 );
buf ( n316205 , n316204 );
buf ( n316206 , n316205 );
or ( n316207 , n316198 , n316206 );
nand ( n316208 , n316197 , n316207 );
buf ( n316209 , n316208 );
buf ( n316210 , n316209 );
buf ( n316211 , n305210 );
buf ( n316212 , n858 );
buf ( n316213 , n868 );
xnor ( n316214 , n316212 , n316213 );
buf ( n316215 , n316214 );
buf ( n316216 , n316215 );
or ( n316217 , n316211 , n316216 );
buf ( n316218 , n305449 );
buf ( n316219 , n25437 );
not ( n316220 , n316219 );
buf ( n316221 , n316220 );
buf ( n316222 , n316221 );
or ( n316223 , n316218 , n316222 );
nand ( n25798 , n316217 , n316223 );
buf ( n316225 , n25798 );
buf ( n316226 , n316225 );
xor ( n316227 , n316210 , n316226 );
buf ( n316228 , n863 );
buf ( n316229 , n865 );
or ( n316230 , n316228 , n316229 );
buf ( n316231 , n866 );
nand ( n316232 , n316230 , n316231 );
buf ( n316233 , n316232 );
buf ( n316234 , n316233 );
buf ( n316235 , n863 );
buf ( n316236 , n865 );
nand ( n316237 , n316235 , n316236 );
buf ( n316238 , n316237 );
buf ( n316239 , n316238 );
buf ( n316240 , n864 );
and ( n316241 , n316234 , n316239 , n316240 );
buf ( n316242 , n316241 );
buf ( n316243 , n316242 );
buf ( n316244 , n895 );
not ( n25819 , n316244 );
buf ( n316246 , n894 );
buf ( n316247 , n832 );
xor ( n25822 , n316246 , n316247 );
buf ( n316249 , n25822 );
buf ( n316250 , n316249 );
not ( n25825 , n316250 );
or ( n25826 , n25819 , n25825 );
buf ( n316253 , n305032 );
buf ( n316254 , n312298 );
nand ( n25829 , n316253 , n316254 );
buf ( n316256 , n25829 );
buf ( n316257 , n316256 );
nand ( n25832 , n25826 , n316257 );
buf ( n316259 , n25832 );
buf ( n316260 , n316259 );
and ( n25835 , n316243 , n316260 );
buf ( n316262 , n25835 );
buf ( n316263 , n316262 );
xor ( n25838 , n316227 , n316263 );
buf ( n316265 , n25838 );
buf ( n316266 , n316265 );
xor ( n316267 , n316187 , n316266 );
xor ( n25842 , n312352 , n312367 );
and ( n25843 , n25842 , n312390 );
and ( n25844 , n312352 , n312367 );
or ( n25845 , n25843 , n25844 );
buf ( n25846 , n25845 );
buf ( n25847 , n25846 );
xor ( n25848 , n312416 , n312445 );
and ( n25849 , n25848 , n312480 );
and ( n316276 , n312416 , n312445 );
or ( n316277 , n25849 , n316276 );
buf ( n316278 , n316277 );
buf ( n316279 , n316278 );
xor ( n25854 , n25847 , n316279 );
xor ( n25855 , n313378 , n313399 );
and ( n25856 , n25855 , n313419 );
and ( n25857 , n313378 , n313399 );
or ( n25858 , n25856 , n25857 );
buf ( n316285 , n25858 );
buf ( n316286 , n316285 );
and ( n316287 , n25854 , n316286 );
and ( n25862 , n25847 , n316279 );
or ( n25863 , n316287 , n25862 );
buf ( n316290 , n25863 );
buf ( n316291 , n316290 );
and ( n316292 , n316267 , n316291 );
and ( n25867 , n316187 , n316266 );
or ( n25868 , n316292 , n25867 );
buf ( n316295 , n25868 );
buf ( n316296 , n316295 );
and ( n316297 , n316118 , n316296 );
and ( n25872 , n315909 , n316117 );
or ( n25873 , n316297 , n25872 );
buf ( n316300 , n25873 );
buf ( n316301 , n316300 );
xor ( n316302 , n315862 , n315877 );
and ( n25877 , n316302 , n315903 );
and ( n25878 , n315862 , n315877 );
or ( n316305 , n25877 , n25878 );
buf ( n316306 , n316305 );
buf ( n316307 , n316306 );
buf ( n316308 , n315986 );
not ( n316309 , n316308 );
buf ( n316310 , n313029 );
not ( n316311 , n316310 );
or ( n316312 , n316309 , n316311 );
buf ( n316313 , n845 );
buf ( n316314 , n878 );
xor ( n316315 , n316313 , n316314 );
buf ( n316316 , n316315 );
buf ( n316317 , n316316 );
buf ( n316318 , n306272 );
nand ( n316319 , n316317 , n316318 );
buf ( n316320 , n316319 );
buf ( n316321 , n316320 );
nand ( n316322 , n316312 , n316321 );
buf ( n316323 , n316322 );
buf ( n316324 , n316323 );
buf ( n316325 , n316103 );
not ( n316326 , n316325 );
buf ( n316327 , n305338 );
not ( n25902 , n316327 );
or ( n316329 , n316326 , n25902 );
xor ( n316330 , n876 , n847 );
buf ( n316331 , n316330 );
buf ( n316332 , n305344 );
nand ( n316333 , n316331 , n316332 );
buf ( n316334 , n316333 );
buf ( n316335 , n316334 );
nand ( n316336 , n316329 , n316335 );
buf ( n316337 , n316336 );
buf ( n316338 , n316337 );
xor ( n316339 , n316324 , n316338 );
buf ( n316340 , n15804 );
buf ( n316341 , n315919 );
not ( n316342 , n316341 );
buf ( n316343 , n316342 );
buf ( n316344 , n316343 );
or ( n316345 , n316340 , n316344 );
buf ( n316346 , n306238 );
buf ( n316347 , n884 );
buf ( n316348 , n839 );
xnor ( n316349 , n316347 , n316348 );
buf ( n316350 , n316349 );
buf ( n316351 , n316350 );
or ( n316352 , n316346 , n316351 );
nand ( n316353 , n316345 , n316352 );
buf ( n316354 , n316353 );
buf ( n316355 , n316354 );
xor ( n316356 , n316339 , n316355 );
buf ( n316357 , n316356 );
buf ( n316358 , n316357 );
xor ( n316359 , n316307 , n316358 );
buf ( n316360 , n315733 );
not ( n25935 , n316360 );
buf ( n316362 , n311226 );
not ( n316363 , n316362 );
or ( n316364 , n25935 , n316363 );
buf ( n316365 , n310582 );
buf ( n316366 , n864 );
buf ( n316367 , n859 );
xor ( n25942 , n316366 , n316367 );
buf ( n316369 , n25942 );
buf ( n316370 , n316369 );
nand ( n25945 , n316365 , n316370 );
buf ( n316372 , n25945 );
buf ( n316373 , n316372 );
nand ( n25948 , n316364 , n316373 );
buf ( n316375 , n25948 );
buf ( n316376 , n316375 );
buf ( n316377 , n866 );
buf ( n316378 , n858 );
and ( n316379 , n316377 , n316378 );
not ( n25954 , n316377 );
buf ( n316381 , n305060 );
and ( n25956 , n25954 , n316381 );
nor ( n25957 , n316379 , n25956 );
buf ( n316384 , n25957 );
buf ( n316385 , n316384 );
not ( n25960 , n316385 );
buf ( n316387 , n310694 );
not ( n25962 , n316387 );
or ( n25963 , n25960 , n25962 );
buf ( n25964 , n311107 );
buf ( n316391 , n866 );
buf ( n316392 , n857 );
xor ( n316393 , n316391 , n316392 );
buf ( n316394 , n316393 );
buf ( n316395 , n316394 );
nand ( n316396 , n25964 , n316395 );
buf ( n316397 , n316396 );
buf ( n316398 , n316397 );
nand ( n25973 , n25963 , n316398 );
buf ( n316400 , n25973 );
buf ( n316401 , n316400 );
xor ( n25976 , n316376 , n316401 );
buf ( n316403 , n304987 );
buf ( n316404 , n315756 );
not ( n25979 , n316404 );
buf ( n316406 , n25979 );
buf ( n316407 , n316406 );
or ( n316408 , n316403 , n316407 );
buf ( n316409 , n311075 );
buf ( n316410 , n843 );
buf ( n316411 , n880 );
xnor ( n25986 , n316410 , n316411 );
buf ( n316413 , n25986 );
buf ( n316414 , n316413 );
or ( n25989 , n316409 , n316414 );
nand ( n25990 , n316408 , n25989 );
buf ( n316417 , n25990 );
buf ( n316418 , n316417 );
xor ( n25993 , n25976 , n316418 );
buf ( n316420 , n25993 );
buf ( n316421 , n316420 );
xor ( n25996 , n316359 , n316421 );
buf ( n316423 , n25996 );
buf ( n316424 , n316423 );
buf ( n316425 , n315955 );
not ( n316426 , n316425 );
buf ( n316427 , n14420 );
not ( n26002 , n316427 );
or ( n26003 , n316426 , n26002 );
buf ( n316430 , n304864 );
xor ( n316431 , n872 , n851 );
buf ( n316432 , n316431 );
nand ( n26007 , n316430 , n316432 );
buf ( n316434 , n26007 );
buf ( n316435 , n316434 );
nand ( n26010 , n26003 , n316435 );
buf ( n316437 , n26010 );
buf ( n316438 , n316437 );
buf ( n316439 , n316061 );
not ( n316440 , n316439 );
buf ( n316441 , n305627 );
not ( n26016 , n316441 );
or ( n26017 , n316440 , n26016 );
buf ( n316444 , n874 );
buf ( n26019 , n849 );
and ( n26020 , n316444 , n26019 );
not ( n26021 , n316444 );
buf ( n316448 , n305596 );
and ( n26023 , n26021 , n316448 );
nor ( n26024 , n26020 , n26023 );
buf ( n316451 , n26024 );
buf ( n26026 , n316451 );
buf ( n316453 , n305289 );
nand ( n26028 , n26026 , n316453 );
buf ( n316455 , n26028 );
buf ( n316456 , n316455 );
nand ( n316457 , n26017 , n316456 );
buf ( n316458 , n316457 );
buf ( n316459 , n316458 );
xor ( n26034 , n316438 , n316459 );
buf ( n316461 , n316041 );
not ( n26036 , n316461 );
buf ( n316463 , n305138 );
not ( n316464 , n316463 );
or ( n316465 , n26036 , n316464 );
buf ( n316466 , n305144 );
buf ( n316467 , n888 );
buf ( n316468 , n835 );
xor ( n26043 , n316467 , n316468 );
buf ( n26044 , n26043 );
buf ( n316471 , n26044 );
nand ( n26046 , n316466 , n316471 );
buf ( n316473 , n26046 );
buf ( n316474 , n316473 );
nand ( n26049 , n316465 , n316474 );
buf ( n316476 , n26049 );
buf ( n316477 , n316476 );
xor ( n26052 , n26034 , n316477 );
buf ( n316479 , n26052 );
buf ( n316480 , n316479 );
and ( n26055 , n315720 , n315721 );
buf ( n316482 , n26055 );
buf ( n316483 , n316482 );
buf ( n26058 , n315932 );
not ( n26059 , n26058 );
buf ( n26060 , n304633 );
not ( n26061 , n26060 );
or ( n26062 , n26059 , n26061 );
buf ( n26063 , n304655 );
buf ( n316490 , n833 );
buf ( n316491 , n890 );
xnor ( n316492 , n316490 , n316491 );
buf ( n316493 , n316492 );
buf ( n316494 , n316493 );
or ( n316495 , n26063 , n316494 );
buf ( n316496 , n316495 );
buf ( n316497 , n316496 );
nand ( n26072 , n26062 , n316497 );
buf ( n316499 , n26072 );
buf ( n316500 , n316499 );
xor ( n26075 , n316483 , n316500 );
buf ( n316502 , n314747 );
buf ( n316503 , n25654 );
not ( n316504 , n316503 );
buf ( n316505 , n316504 );
buf ( n316506 , n316505 );
or ( n26081 , n316502 , n316506 );
buf ( n316508 , n305363 );
buf ( n316509 , n886 );
buf ( n316510 , n837 );
xor ( n26085 , n316509 , n316510 );
buf ( n316512 , n26085 );
buf ( n316513 , n316512 );
not ( n26088 , n316513 );
buf ( n316515 , n26088 );
buf ( n316516 , n316515 );
or ( n26091 , n316508 , n316516 );
nand ( n316518 , n26081 , n26091 );
buf ( n316519 , n316518 );
buf ( n316520 , n316519 );
xor ( n26095 , n26075 , n316520 );
buf ( n316522 , n26095 );
buf ( n316523 , n316522 );
xor ( n316524 , n316480 , n316523 );
buf ( n316525 , n315896 );
not ( n316526 , n316525 );
buf ( n316527 , n304584 );
not ( n26102 , n316527 );
or ( n316529 , n316526 , n26102 );
buf ( n316530 , n304596 );
xor ( n26105 , n882 , n841 );
buf ( n316532 , n26105 );
nand ( n26107 , n316530 , n316532 );
buf ( n316534 , n26107 );
buf ( n316535 , n316534 );
nand ( n316536 , n316529 , n316535 );
buf ( n316537 , n316536 );
buf ( n316538 , n316537 );
buf ( n316539 , n315870 );
not ( n26114 , n316539 );
buf ( n316541 , n305213 );
not ( n26116 , n316541 );
or ( n316543 , n26114 , n26116 );
buf ( n316544 , n305202 );
buf ( n316545 , n868 );
buf ( n316546 , n855 );
and ( n26121 , n316545 , n316546 );
not ( n316548 , n316545 );
buf ( n316549 , n305319 );
and ( n26124 , n316548 , n316549 );
nor ( n316551 , n26121 , n26124 );
buf ( n316552 , n316551 );
buf ( n316553 , n316552 );
nand ( n316554 , n316544 , n316553 );
buf ( n316555 , n316554 );
buf ( n316556 , n316555 );
nand ( n26131 , n316543 , n316556 );
buf ( n316558 , n26131 );
buf ( n316559 , n316558 );
xor ( n316560 , n316538 , n316559 );
buf ( n316561 , n315120 );
buf ( n316562 , n315855 );
not ( n26137 , n316562 );
buf ( n316564 , n26137 );
buf ( n316565 , n316564 );
or ( n26140 , n316561 , n316565 );
buf ( n316567 , n870 );
buf ( n316568 , n853 );
and ( n26143 , n316567 , n316568 );
not ( n26144 , n316567 );
buf ( n316571 , n304956 );
and ( n26146 , n26144 , n316571 );
nor ( n26147 , n26143 , n26146 );
buf ( n316574 , n26147 );
buf ( n316575 , n316574 );
not ( n26150 , n316575 );
buf ( n316577 , n26150 );
buf ( n316578 , n316577 );
buf ( n316579 , n14318 );
or ( n26154 , n316578 , n316579 );
nand ( n26155 , n26140 , n26154 );
buf ( n316582 , n26155 );
buf ( n26157 , n316582 );
xor ( n26158 , n316560 , n26157 );
buf ( n26159 , n26158 );
buf ( n316586 , n26159 );
xor ( n26161 , n316524 , n316586 );
buf ( n316588 , n26161 );
buf ( n316589 , n316588 );
xor ( n316590 , n316424 , n316589 );
buf ( n316591 , n316202 );
not ( n26166 , n316591 );
buf ( n316593 , n310694 );
not ( n26168 , n316593 );
or ( n26169 , n26166 , n26168 );
buf ( n316596 , n311107 );
buf ( n316597 , n316384 );
nand ( n26172 , n316596 , n316597 );
buf ( n316599 , n26172 );
buf ( n316600 , n316599 );
nand ( n26175 , n26169 , n316600 );
buf ( n316602 , n26175 );
buf ( n316603 , n316602 );
buf ( n316604 , n894 );
xor ( n316605 , n316603 , n316604 );
buf ( n316606 , n863 );
buf ( n316607 , n864 );
and ( n316608 , n316606 , n316607 );
buf ( n316609 , n316608 );
buf ( n316610 , n316609 );
buf ( n316611 , n316249 );
not ( n26186 , n316611 );
buf ( n316613 , n305032 );
not ( n316614 , n316613 );
or ( n316615 , n26186 , n316614 );
buf ( n316616 , n894 );
buf ( n316617 , n895 );
nand ( n26192 , n316616 , n316617 );
buf ( n316619 , n26192 );
buf ( n316620 , n316619 );
nand ( n316621 , n316615 , n316620 );
buf ( n316622 , n316621 );
buf ( n316623 , n316622 );
xor ( n26198 , n316610 , n316623 );
buf ( n316625 , n834 );
buf ( n316626 , n892 );
and ( n26201 , n316625 , n316626 );
not ( n316628 , n316625 );
buf ( n316629 , n305566 );
and ( n26204 , n316628 , n316629 );
nor ( n26205 , n26201 , n26204 );
buf ( n316632 , n26205 );
buf ( n316633 , n316632 );
not ( n26208 , n316633 );
buf ( n316635 , n14272 );
not ( n316636 , n316635 );
or ( n26211 , n26208 , n316636 );
buf ( n316638 , n304694 );
buf ( n316639 , n316001 );
nand ( n26214 , n316638 , n316639 );
buf ( n316641 , n26214 );
buf ( n316642 , n316641 );
nand ( n26217 , n26211 , n316642 );
buf ( n316644 , n26217 );
buf ( n316645 , n316644 );
and ( n26220 , n26198 , n316645 );
and ( n316647 , n316610 , n316623 );
or ( n316648 , n26220 , n316647 );
buf ( n316649 , n316648 );
buf ( n316650 , n316649 );
xor ( n26225 , n316605 , n316650 );
buf ( n316652 , n26225 );
buf ( n26227 , n316652 );
buf ( n26228 , n316154 );
not ( n26229 , n26228 );
buf ( n26230 , n316175 );
not ( n26231 , n26230 );
or ( n26232 , n26229 , n26231 );
buf ( n316659 , n316175 );
buf ( n316660 , n316154 );
or ( n316661 , n316659 , n316660 );
buf ( n316662 , n316132 );
nand ( n316663 , n316661 , n316662 );
buf ( n316664 , n316663 );
buf ( n316665 , n316664 );
nand ( n316666 , n26232 , n316665 );
buf ( n316667 , n316666 );
buf ( n316668 , n316667 );
buf ( n316669 , n886 );
buf ( n26244 , n840 );
xor ( n26245 , n316669 , n26244 );
buf ( n316672 , n26245 );
buf ( n316673 , n316672 );
not ( n316674 , n316673 );
buf ( n316675 , n311697 );
not ( n26250 , n316675 );
or ( n316677 , n316674 , n26250 );
buf ( n26252 , n304901 );
buf ( n26253 , n316073 );
nand ( n26254 , n26252 , n26253 );
buf ( n26255 , n26254 );
buf ( n316682 , n26255 );
nand ( n26257 , n316677 , n316682 );
buf ( n26258 , n26257 );
buf ( n316685 , n26258 );
buf ( n316686 , n876 );
buf ( n316687 , n850 );
and ( n316688 , n316686 , n316687 );
not ( n26263 , n316686 );
buf ( n316690 , n304565 );
and ( n316691 , n26263 , n316690 );
nor ( n316692 , n316688 , n316691 );
buf ( n316693 , n316692 );
buf ( n316694 , n316693 );
not ( n26269 , n316694 );
buf ( n316696 , n305338 );
not ( n316697 , n316696 );
or ( n316698 , n26269 , n316697 );
buf ( n316699 , n305344 );
buf ( n316700 , n316093 );
nand ( n316701 , n316699 , n316700 );
buf ( n316702 , n316701 );
buf ( n316703 , n316702 );
nand ( n316704 , n316698 , n316703 );
buf ( n316705 , n316704 );
buf ( n316706 , n316705 );
xor ( n316707 , n316685 , n316706 );
buf ( n316708 , n878 );
buf ( n316709 , n848 );
and ( n26284 , n316708 , n316709 );
not ( n316711 , n316708 );
buf ( n316712 , n304786 );
and ( n26287 , n316711 , n316712 );
nor ( n316714 , n26284 , n26287 );
buf ( n316715 , n316714 );
buf ( n316716 , n316715 );
not ( n26291 , n316716 );
buf ( n316718 , n15836 );
not ( n316719 , n316718 );
or ( n26294 , n26291 , n316719 );
buf ( n316721 , n306272 );
buf ( n316722 , n315976 );
nand ( n26297 , n316721 , n316722 );
buf ( n26298 , n26297 );
buf ( n316725 , n26298 );
nand ( n26300 , n26294 , n316725 );
buf ( n316727 , n26300 );
buf ( n316728 , n316727 );
and ( n316729 , n316707 , n316728 );
and ( n26304 , n316685 , n316706 );
or ( n26305 , n316729 , n26304 );
buf ( n316732 , n26305 );
buf ( n316733 , n316732 );
xor ( n316734 , n316668 , n316733 );
xor ( n26309 , n882 , n844 );
buf ( n316736 , n26309 );
not ( n316737 , n316736 );
buf ( n316738 , n304584 );
not ( n316739 , n316738 );
or ( n316740 , n316737 , n316739 );
buf ( n316741 , n304596 );
buf ( n316742 , n315882 );
nand ( n316743 , n316741 , n316742 );
buf ( n316744 , n316743 );
buf ( n316745 , n316744 );
nand ( n316746 , n316740 , n316745 );
buf ( n316747 , n316746 );
buf ( n316748 , n316747 );
buf ( n316749 , n856 );
buf ( n316750 , n870 );
xor ( n26325 , n316749 , n316750 );
buf ( n316752 , n26325 );
buf ( n316753 , n316752 );
not ( n26328 , n316753 );
buf ( n316755 , n14323 );
not ( n26330 , n316755 );
or ( n316757 , n26328 , n26330 );
buf ( n316758 , n304763 );
buf ( n316759 , n315845 );
nand ( n316760 , n316758 , n316759 );
buf ( n316761 , n316760 );
buf ( n316762 , n316761 );
nand ( n316763 , n316757 , n316762 );
buf ( n316764 , n316763 );
buf ( n316765 , n316764 );
xor ( n316766 , n316748 , n316765 );
buf ( n316767 , n872 );
buf ( n26342 , n854 );
and ( n26343 , n316767 , n26342 );
not ( n316770 , n316767 );
buf ( n316771 , n854 );
not ( n26346 , n316771 );
buf ( n26347 , n26346 );
buf ( n316774 , n26347 );
and ( n316775 , n316770 , n316774 );
nor ( n316776 , n26343 , n316775 );
buf ( n316777 , n316776 );
buf ( n316778 , n316777 );
not ( n26353 , n316778 );
buf ( n316780 , n304851 );
not ( n26355 , n316780 );
or ( n316782 , n26353 , n26355 );
buf ( n316783 , n304864 );
buf ( n316784 , n25519 );
nand ( n316785 , n316783 , n316784 );
buf ( n316786 , n316785 );
buf ( n316787 , n316786 );
nand ( n26362 , n316782 , n316787 );
buf ( n316789 , n26362 );
buf ( n316790 , n316789 );
and ( n316791 , n316766 , n316790 );
and ( n316792 , n316748 , n316765 );
or ( n26367 , n316791 , n316792 );
buf ( n316794 , n26367 );
buf ( n316795 , n316794 );
xor ( n26370 , n316734 , n316795 );
buf ( n316797 , n26370 );
buf ( n316798 , n316797 );
xor ( n26373 , n26227 , n316798 );
xor ( n26374 , n316685 , n316706 );
xor ( n316801 , n26374 , n316728 );
buf ( n316802 , n316801 );
buf ( n316803 , n316802 );
xor ( n316804 , n25358 , n315809 );
xor ( n26379 , n316804 , n315835 );
buf ( n316806 , n26379 );
buf ( n316807 , n316806 );
xor ( n26382 , n316803 , n316807 );
xor ( n26383 , n316748 , n316765 );
xor ( n316810 , n26383 , n316790 );
buf ( n316811 , n316810 );
buf ( n316812 , n316811 );
and ( n316813 , n26382 , n316812 );
and ( n26388 , n316803 , n316807 );
or ( n316815 , n316813 , n26388 );
buf ( n316816 , n316815 );
buf ( n316817 , n316816 );
and ( n26392 , n26373 , n316817 );
and ( n316819 , n26227 , n316798 );
or ( n316820 , n26392 , n316819 );
buf ( n316821 , n316820 );
buf ( n316822 , n316821 );
xor ( n26397 , n316590 , n316822 );
buf ( n316824 , n26397 );
buf ( n316825 , n316824 );
xor ( n316826 , n316243 , n316260 );
buf ( n316827 , n316826 );
buf ( n316828 , n316827 );
xor ( n316829 , n312285 , n312306 );
and ( n26404 , n316829 , n312328 );
and ( n316831 , n312285 , n312306 );
or ( n26406 , n26404 , n316831 );
buf ( n316833 , n26406 );
buf ( n316834 , n316833 );
xor ( n316835 , n316828 , n316834 );
xor ( n316836 , n313318 , n313336 );
and ( n26411 , n316836 , n313357 );
and ( n316838 , n313318 , n313336 );
or ( n316839 , n26411 , n316838 );
buf ( n316840 , n316839 );
buf ( n316841 , n316840 );
and ( n316842 , n316835 , n316841 );
and ( n26417 , n316828 , n316834 );
or ( n316844 , n316842 , n26417 );
buf ( n316845 , n316844 );
buf ( n26420 , n316845 );
buf ( n316847 , n312409 );
not ( n26422 , n316847 );
buf ( n316849 , n304851 );
not ( n316850 , n316849 );
or ( n26425 , n26422 , n316850 );
buf ( n316852 , n304845 );
buf ( n316853 , n316777 );
nand ( n26428 , n316852 , n316853 );
buf ( n316855 , n26428 );
buf ( n316856 , n316855 );
nand ( n316857 , n26425 , n316856 );
buf ( n316858 , n316857 );
buf ( n316859 , n316858 );
not ( n316860 , n316859 );
buf ( n316861 , n312345 );
not ( n316862 , n316861 );
buf ( n316863 , n20629 );
not ( n26438 , n316863 );
or ( n316865 , n316862 , n26438 );
buf ( n316866 , n311052 );
buf ( n316867 , n316752 );
nand ( n316868 , n316866 , n316867 );
buf ( n316869 , n316868 );
buf ( n316870 , n316869 );
nand ( n316871 , n316865 , n316870 );
buf ( n316872 , n316871 );
buf ( n26447 , n316872 );
not ( n26448 , n26447 );
or ( n26449 , n316860 , n26448 );
buf ( n316876 , n316872 );
buf ( n316877 , n316858 );
or ( n316878 , n316876 , n316877 );
buf ( n316879 , n22012 );
not ( n316880 , n316879 );
buf ( n316881 , n304813 );
not ( n26456 , n316881 );
or ( n316883 , n316880 , n26456 );
buf ( n316884 , n304807 );
buf ( n316885 , n315818 );
nand ( n316886 , n316884 , n316885 );
buf ( n316887 , n316886 );
buf ( n316888 , n316887 );
nand ( n316889 , n316883 , n316888 );
buf ( n316890 , n316889 );
buf ( n316891 , n316890 );
nand ( n26466 , n316878 , n316891 );
buf ( n316893 , n26466 );
buf ( n316894 , n316893 );
nand ( n316895 , n26449 , n316894 );
buf ( n316896 , n316895 );
buf ( n316897 , n316896 );
buf ( n316898 , n22803 );
not ( n316899 , n316898 );
buf ( n316900 , n310477 );
not ( n316901 , n316900 );
or ( n26476 , n316899 , n316901 );
buf ( n316903 , n310483 );
buf ( n316904 , n316192 );
nand ( n26479 , n316903 , n316904 );
buf ( n316906 , n26479 );
buf ( n316907 , n316906 );
nand ( n26482 , n26476 , n316907 );
buf ( n316909 , n26482 );
buf ( n316910 , n316909 );
buf ( n316911 , n312360 );
not ( n26486 , n316911 );
buf ( n316913 , n305213 );
not ( n316914 , n316913 );
or ( n26489 , n26486 , n316914 );
buf ( n316916 , n316215 );
not ( n316917 , n316916 );
buf ( n316918 , n305202 );
nand ( n316919 , n316917 , n316918 );
buf ( n316920 , n316919 );
buf ( n316921 , n316920 );
nand ( n316922 , n26489 , n316921 );
buf ( n316923 , n316922 );
buf ( n26498 , n316923 );
xor ( n26499 , n316910 , n26498 );
buf ( n316926 , n312383 );
not ( n316927 , n316926 );
buf ( n316928 , n304584 );
not ( n316929 , n316928 );
or ( n316930 , n316927 , n316929 );
buf ( n316931 , n304596 );
buf ( n316932 , n26309 );
nand ( n316933 , n316931 , n316932 );
buf ( n316934 , n316933 );
buf ( n316935 , n316934 );
nand ( n316936 , n316930 , n316935 );
buf ( n316937 , n316936 );
buf ( n316938 , n316937 );
and ( n316939 , n26499 , n316938 );
and ( n26514 , n316910 , n26498 );
or ( n26515 , n316939 , n26514 );
buf ( n316942 , n26515 );
buf ( n316943 , n316942 );
xor ( n316944 , n316897 , n316943 );
xor ( n26519 , n316610 , n316623 );
xor ( n316946 , n26519 , n316645 );
buf ( n316947 , n316946 );
buf ( n316948 , n316947 );
xor ( n316949 , n316944 , n316948 );
buf ( n316950 , n316949 );
buf ( n316951 , n316950 );
xor ( n316952 , n26420 , n316951 );
xor ( n26527 , n316910 , n26498 );
xor ( n316954 , n26527 , n316938 );
buf ( n316955 , n316954 );
buf ( n316956 , n316955 );
buf ( n316957 , n22985 );
not ( n316958 , n316957 );
buf ( n316959 , n304912 );
not ( n26534 , n316959 );
or ( n316961 , n316958 , n26534 );
buf ( n316962 , n304901 );
buf ( n316963 , n316672 );
nand ( n26538 , n316962 , n316963 );
buf ( n316965 , n26538 );
buf ( n316966 , n316965 );
nand ( n316967 , n316961 , n316966 );
buf ( n316968 , n316967 );
buf ( n316969 , n316968 );
buf ( n316970 , n313310 );
not ( n26545 , n316970 );
buf ( n316972 , n304984 );
not ( n316973 , n316972 );
or ( n26548 , n26545 , n316973 );
buf ( n316975 , n304997 );
buf ( n316976 , n316163 );
nand ( n26551 , n316975 , n316976 );
buf ( n316978 , n26551 );
buf ( n316979 , n316978 );
nand ( n26554 , n26548 , n316979 );
buf ( n316981 , n26554 );
buf ( n316982 , n316981 );
xor ( n26557 , n316969 , n316982 );
buf ( n316984 , n304941 );
buf ( n316985 , n313327 );
or ( n26560 , n316984 , n316985 );
buf ( n316987 , n14523 );
buf ( n316988 , n316715 );
not ( n316989 , n316988 );
buf ( n316990 , n316989 );
buf ( n316991 , n316990 );
or ( n26566 , n316987 , n316991 );
nand ( n316993 , n26560 , n26566 );
buf ( n316994 , n316993 );
buf ( n316995 , n316994 );
xor ( n316996 , n26557 , n316995 );
buf ( n316997 , n316996 );
buf ( n316998 , n316997 );
xor ( n316999 , n316956 , n316998 );
buf ( n317000 , n312320 );
not ( n26575 , n317000 );
buf ( n317002 , n14272 );
not ( n317003 , n317002 );
or ( n317004 , n26575 , n317003 );
buf ( n317005 , n316632 );
buf ( n317006 , n304694 );
nand ( n317007 , n317005 , n317006 );
buf ( n317008 , n317007 );
buf ( n317009 , n317008 );
nand ( n317010 , n317004 , n317009 );
buf ( n317011 , n317010 );
buf ( n317012 , n317011 );
buf ( n317013 , n313352 );
not ( n317014 , n317013 );
buf ( n317015 , n317014 );
buf ( n317016 , n317015 );
not ( n317017 , n317016 );
buf ( n317018 , n305138 );
not ( n26593 , n317018 );
or ( n317020 , n317017 , n26593 );
buf ( n317021 , n316142 );
buf ( n26596 , n305144 );
nand ( n26597 , n317021 , n26596 );
buf ( n26598 , n26597 );
buf ( n317025 , n26598 );
nand ( n26600 , n317020 , n317025 );
buf ( n317027 , n26600 );
buf ( n317028 , n317027 );
xor ( n317029 , n317012 , n317028 );
buf ( n317030 , n311891 );
buf ( n317031 , n311234 );
buf ( n317032 , n863 );
and ( n317033 , n317031 , n317032 );
buf ( n317034 , n305192 );
buf ( n317035 , n864 );
and ( n317036 , n317034 , n317035 );
nor ( n317037 , n317033 , n317036 );
buf ( n317038 , n317037 );
buf ( n317039 , n317038 );
or ( n317040 , n317030 , n317039 );
buf ( n317041 , n311246 );
buf ( n317042 , n316120 );
not ( n317043 , n317042 );
buf ( n317044 , n317043 );
buf ( n317045 , n317044 );
or ( n317046 , n317041 , n317045 );
nand ( n26621 , n317040 , n317046 );
buf ( n317048 , n26621 );
buf ( n317049 , n317048 );
xor ( n26624 , n317029 , n317049 );
buf ( n317051 , n26624 );
buf ( n317052 , n317051 );
and ( n317053 , n316999 , n317052 );
and ( n26628 , n316956 , n316998 );
or ( n317055 , n317053 , n26628 );
buf ( n317056 , n317055 );
buf ( n317057 , n317056 );
and ( n317058 , n316952 , n317057 );
and ( n317059 , n26420 , n316951 );
or ( n26634 , n317058 , n317059 );
buf ( n317061 , n26634 );
buf ( n317062 , n317061 );
xor ( n26637 , n316210 , n316226 );
and ( n26638 , n26637 , n316263 );
and ( n26639 , n316210 , n316226 );
or ( n317066 , n26638 , n26639 );
buf ( n317067 , n317066 );
buf ( n317068 , n317067 );
xor ( n26643 , n316897 , n316943 );
and ( n317070 , n26643 , n316948 );
and ( n26645 , n316897 , n316943 );
or ( n26646 , n317070 , n26645 );
buf ( n317073 , n26646 );
buf ( n26648 , n317073 );
xor ( n26649 , n317068 , n26648 );
xor ( n317076 , n316969 , n316982 );
and ( n317077 , n317076 , n316995 );
and ( n26652 , n316969 , n316982 );
or ( n317079 , n317077 , n26652 );
buf ( n317080 , n317079 );
buf ( n317081 , n317080 );
xor ( n317082 , n317012 , n317028 );
and ( n26657 , n317082 , n317049 );
and ( n317084 , n317012 , n317028 );
or ( n26659 , n26657 , n317084 );
buf ( n317086 , n26659 );
buf ( n317087 , n317086 );
xor ( n317088 , n317081 , n317087 );
buf ( n317089 , n22945 );
not ( n26664 , n317089 );
buf ( n317091 , n305338 );
not ( n317092 , n317091 );
or ( n317093 , n26664 , n317092 );
buf ( n317094 , n305344 );
buf ( n317095 , n316693 );
nand ( n317096 , n317094 , n317095 );
buf ( n317097 , n317096 );
buf ( n317098 , n317097 );
nand ( n26673 , n317093 , n317098 );
buf ( n26674 , n26673 );
buf ( n317101 , n26674 );
buf ( n317102 , n313392 );
not ( n317103 , n317102 );
buf ( n317104 , n305627 );
not ( n26679 , n317104 );
or ( n317106 , n317103 , n26679 );
buf ( n317107 , n305301 );
buf ( n317108 , n25341 );
nand ( n317109 , n317107 , n317108 );
buf ( n317110 , n317109 );
buf ( n317111 , n317110 );
nand ( n317112 , n317106 , n317111 );
buf ( n317113 , n317112 );
buf ( n317114 , n317113 );
xor ( n317115 , n317101 , n317114 );
buf ( n317116 , n304630 );
buf ( n317117 , n312474 );
or ( n317118 , n317116 , n317117 );
buf ( n317119 , n304655 );
buf ( n317120 , n315792 );
not ( n317121 , n317120 );
buf ( n317122 , n317121 );
buf ( n317123 , n317122 );
or ( n26698 , n317119 , n317123 );
nand ( n317125 , n317118 , n26698 );
buf ( n317126 , n317125 );
buf ( n317127 , n317126 );
and ( n317128 , n317115 , n317127 );
and ( n317129 , n317101 , n317114 );
or ( n26704 , n317128 , n317129 );
buf ( n317131 , n26704 );
buf ( n317132 , n317131 );
and ( n26707 , n317088 , n317132 );
and ( n317134 , n317081 , n317087 );
or ( n317135 , n26707 , n317134 );
buf ( n317136 , n317135 );
buf ( n317137 , n317136 );
xor ( n317138 , n26649 , n317137 );
buf ( n317139 , n317138 );
buf ( n317140 , n317139 );
xor ( n317141 , n317062 , n317140 );
xor ( n26716 , n26227 , n316798 );
xor ( n317143 , n26716 , n316817 );
buf ( n317144 , n317143 );
buf ( n317145 , n317144 );
and ( n317146 , n317141 , n317145 );
and ( n317147 , n317062 , n317140 );
or ( n317148 , n317146 , n317147 );
buf ( n317149 , n317148 );
buf ( n317150 , n317149 );
xor ( n317151 , n316301 , n316825 );
xor ( n26726 , n317151 , n317150 );
buf ( n317153 , n26726 );
xor ( n317154 , n316301 , n316825 );
and ( n26729 , n317154 , n317150 );
and ( n317156 , n316301 , n316825 );
or ( n317157 , n26729 , n317156 );
buf ( n317158 , n317157 );
xor ( n26733 , n314982 , n314988 );
and ( n26734 , n26733 , n314995 );
and ( n317161 , n314982 , n314988 );
or ( n317162 , n26734 , n317161 );
buf ( n317163 , n317162 );
buf ( n317164 , n317163 );
xor ( n317165 , n315005 , n315050 );
and ( n26740 , n317165 , n315106 );
and ( n26741 , n315005 , n315050 );
or ( n26742 , n26740 , n26741 );
buf ( n317169 , n26742 );
buf ( n317170 , n317169 );
xor ( n317171 , n317164 , n317170 );
xor ( n317172 , n315008 , n315029 );
and ( n26747 , n317172 , n315047 );
and ( n317174 , n315008 , n315029 );
or ( n317175 , n26747 , n317174 );
buf ( n317176 , n317175 );
buf ( n317177 , n317176 );
xor ( n26752 , n315174 , n315191 );
and ( n26753 , n26752 , n24782 );
and ( n317180 , n315174 , n315191 );
or ( n317181 , n26753 , n317180 );
buf ( n26756 , n317181 );
xor ( n26757 , n317177 , n26756 );
and ( n317184 , n314840 , n314841 );
buf ( n317185 , n317184 );
buf ( n317186 , n317185 );
buf ( n317187 , n315170 );
not ( n317188 , n317187 );
buf ( n317189 , n317188 );
buf ( n317190 , n317189 );
not ( n317191 , n317190 );
buf ( n317192 , n14323 );
not ( n317193 , n317192 );
or ( n317194 , n317191 , n317193 );
buf ( n317195 , n840 );
buf ( n317196 , n870 );
xnor ( n317197 , n317195 , n317196 );
buf ( n317198 , n317197 );
buf ( n317199 , n317198 );
not ( n26774 , n317199 );
buf ( n317201 , n311052 );
nand ( n317202 , n26774 , n317201 );
buf ( n317203 , n317202 );
buf ( n317204 , n317203 );
nand ( n26779 , n317194 , n317204 );
buf ( n26780 , n26779 );
buf ( n26781 , n26780 );
xor ( n26782 , n317186 , n26781 );
buf ( n317209 , n305650 );
buf ( n317210 , n315204 );
or ( n26785 , n317209 , n317210 );
buf ( n317212 , n305664 );
buf ( n317213 , n876 );
buf ( n317214 , n310658 );
and ( n26789 , n317213 , n317214 );
not ( n317216 , n317213 );
buf ( n317217 , n834 );
and ( n26792 , n317216 , n317217 );
nor ( n26793 , n26789 , n26792 );
buf ( n317220 , n26793 );
buf ( n317221 , n317220 );
or ( n317222 , n317212 , n317221 );
nand ( n26797 , n26785 , n317222 );
buf ( n317224 , n26797 );
buf ( n317225 , n317224 );
xor ( n317226 , n26782 , n317225 );
buf ( n317227 , n317226 );
buf ( n317228 , n317227 );
xor ( n317229 , n26757 , n317228 );
buf ( n317230 , n317229 );
buf ( n317231 , n317230 );
xor ( n317232 , n317171 , n317231 );
buf ( n317233 , n317232 );
buf ( n317234 , n317233 );
xor ( n317235 , n315174 , n315191 );
xor ( n26810 , n317235 , n24782 );
and ( n317237 , n315214 , n26810 );
xor ( n317238 , n315174 , n315191 );
xor ( n26813 , n317238 , n24782 );
and ( n26814 , n315237 , n26813 );
and ( n317241 , n315214 , n315237 );
or ( n26816 , n317237 , n26814 , n317241 );
buf ( n317243 , n26816 );
buf ( n317244 , n304938 );
buf ( n317245 , n315042 );
or ( n317246 , n317244 , n317245 );
buf ( n317247 , n14523 );
buf ( n317248 , n878 );
buf ( n317249 , n20700 );
and ( n317250 , n317248 , n317249 );
not ( n26825 , n317248 );
buf ( n317252 , n832 );
and ( n317253 , n26825 , n317252 );
nor ( n317254 , n317250 , n317253 );
buf ( n317255 , n317254 );
buf ( n317256 , n317255 );
or ( n317257 , n317247 , n317256 );
nand ( n317258 , n317246 , n317257 );
buf ( n317259 , n317258 );
buf ( n317260 , n304976 );
not ( n26835 , n317260 );
buf ( n317262 , n304987 );
not ( n317263 , n317262 );
or ( n26838 , n26835 , n317263 );
buf ( n317265 , n880 );
nand ( n26840 , n26838 , n317265 );
buf ( n26841 , n26840 );
xor ( n317268 , n317259 , n26841 );
buf ( n317269 , n306340 );
buf ( n317270 , n315098 );
or ( n317271 , n317269 , n317270 );
buf ( n317272 , n306346 );
buf ( n317273 , n315090 );
buf ( n317274 , n836 );
and ( n26849 , n317273 , n317274 );
buf ( n317276 , n311204 );
buf ( n317277 , n874 );
and ( n26852 , n317276 , n317277 );
nor ( n317279 , n26849 , n26852 );
buf ( n317280 , n317279 );
buf ( n317281 , n317280 );
or ( n317282 , n317272 , n317281 );
nand ( n317283 , n317271 , n317282 );
buf ( n317284 , n317283 );
xor ( n317285 , n317268 , n317284 );
buf ( n317286 , n315022 );
not ( n26861 , n317286 );
buf ( n317288 , n304851 );
not ( n26863 , n317288 );
or ( n317290 , n26861 , n26863 );
buf ( n317291 , n304845 );
buf ( n317292 , n872 );
buf ( n317293 , n838 );
and ( n26868 , n317292 , n317293 );
not ( n317295 , n317292 );
buf ( n317296 , n310377 );
and ( n26871 , n317295 , n317296 );
nor ( n26872 , n26868 , n26871 );
buf ( n317299 , n26872 );
buf ( n317300 , n317299 );
nand ( n317301 , n317291 , n317300 );
buf ( n317302 , n317301 );
buf ( n317303 , n317302 );
nand ( n26878 , n317290 , n317303 );
buf ( n317305 , n26878 );
buf ( n317306 , n317305 );
buf ( n317307 , n310691 );
buf ( n317308 , n315077 );
or ( n26883 , n317307 , n317308 );
buf ( n317310 , n313224 );
buf ( n317311 , n844 );
buf ( n317312 , n313871 );
and ( n317313 , n317311 , n317312 );
not ( n26888 , n317311 );
buf ( n317315 , n866 );
and ( n317316 , n26888 , n317315 );
nor ( n26891 , n317313 , n317316 );
buf ( n317318 , n26891 );
buf ( n317319 , n317318 );
or ( n26894 , n317310 , n317319 );
nand ( n317321 , n26883 , n26894 );
buf ( n317322 , n317321 );
buf ( n317323 , n317322 );
xor ( n317324 , n317306 , n317323 );
buf ( n317325 , n311891 );
buf ( n317326 , n315060 );
or ( n317327 , n317325 , n317326 );
buf ( n317328 , n311246 );
buf ( n317329 , n311234 );
buf ( n317330 , n846 );
and ( n317331 , n317329 , n317330 );
buf ( n317332 , n311024 );
buf ( n317333 , n864 );
and ( n317334 , n317332 , n317333 );
nor ( n26909 , n317331 , n317334 );
buf ( n317336 , n26909 );
buf ( n317337 , n317336 );
or ( n317338 , n317328 , n317337 );
nand ( n26913 , n317327 , n317338 );
buf ( n26914 , n26913 );
buf ( n317341 , n26914 );
xor ( n26916 , n317324 , n317341 );
buf ( n317343 , n26916 );
buf ( n317344 , n310726 );
buf ( n317345 , n315183 );
or ( n317346 , n317344 , n317345 );
buf ( n317347 , n305449 );
buf ( n317348 , n310521 );
buf ( n317349 , n842 );
and ( n317350 , n317348 , n317349 );
buf ( n317351 , n304610 );
buf ( n317352 , n868 );
and ( n26927 , n317351 , n317352 );
nor ( n317354 , n317350 , n26927 );
buf ( n317355 , n317354 );
buf ( n317356 , n317355 );
or ( n26931 , n317347 , n317356 );
nand ( n317358 , n317346 , n26931 );
buf ( n317359 , n317358 );
buf ( n317360 , n317359 );
buf ( n317361 , n314978 );
xor ( n317362 , n317360 , n317361 );
xor ( n26937 , n315069 , n315082 );
and ( n317364 , n26937 , n315103 );
and ( n317365 , n315069 , n315082 );
or ( n26940 , n317364 , n317365 );
buf ( n317367 , n26940 );
buf ( n317368 , n317367 );
xor ( n26943 , n317362 , n317368 );
buf ( n317370 , n26943 );
xor ( n317371 , n317343 , n317370 );
xor ( n26946 , n317285 , n317371 );
buf ( n317373 , n26946 );
xor ( n317374 , n317243 , n317373 );
xor ( n26949 , n24544 , n314998 );
and ( n317376 , n26949 , n315109 );
and ( n317377 , n24544 , n314998 );
or ( n26952 , n317376 , n317377 );
buf ( n317379 , n26952 );
buf ( n317380 , n317379 );
xor ( n317381 , n317374 , n317380 );
buf ( n317382 , n317381 );
buf ( n317383 , n317382 );
xor ( n317384 , n315162 , n315240 );
and ( n317385 , n317384 , n315261 );
and ( n26960 , n315162 , n315240 );
or ( n317387 , n317385 , n26960 );
buf ( n317388 , n317387 );
buf ( n317389 , n317388 );
xor ( n317390 , n317234 , n317383 );
xor ( n317391 , n317390 , n317389 );
buf ( n317392 , n317391 );
xor ( n317393 , n317234 , n317383 );
and ( n26968 , n317393 , n317389 );
and ( n317395 , n317234 , n317383 );
or ( n26970 , n26968 , n317395 );
buf ( n317397 , n26970 );
xor ( n317398 , n306177 , n306196 );
xor ( n317399 , n317398 , n306369 );
buf ( n317400 , n317399 );
buf ( n317401 , n317400 );
xor ( n317402 , n315482 , n315486 );
and ( n26977 , n317402 , n315576 );
and ( n317404 , n315482 , n315486 );
or ( n317405 , n26977 , n317404 );
buf ( n317406 , n317405 );
buf ( n317407 , n317406 );
xor ( n317408 , n314699 , n314703 );
xor ( n317409 , n317408 , n314797 );
buf ( n317410 , n317409 );
buf ( n317411 , n317410 );
xor ( n317412 , n317401 , n317407 );
xor ( n317413 , n317412 , n317411 );
buf ( n317414 , n317413 );
xor ( n317415 , n317401 , n317407 );
and ( n317416 , n317415 , n317411 );
and ( n26991 , n317401 , n317407 );
or ( n317418 , n317416 , n26991 );
buf ( n317419 , n317418 );
xor ( n26994 , n317177 , n26756 );
and ( n317421 , n26994 , n317228 );
and ( n26996 , n317177 , n26756 );
or ( n317423 , n317421 , n26996 );
buf ( n317424 , n317423 );
buf ( n317425 , n317424 );
xor ( n317426 , n317360 , n317361 );
and ( n317427 , n317426 , n317368 );
and ( n27002 , n317360 , n317361 );
or ( n317429 , n317427 , n27002 );
buf ( n317430 , n317429 );
buf ( n317431 , n317430 );
xor ( n317432 , n317425 , n317431 );
xor ( n27007 , n317186 , n26781 );
and ( n317434 , n27007 , n317225 );
and ( n27009 , n317186 , n26781 );
or ( n317436 , n317434 , n27009 );
buf ( n317437 , n317436 );
buf ( n317438 , n317437 );
xor ( n317439 , n317306 , n317323 );
and ( n317440 , n317439 , n317341 );
and ( n27015 , n317306 , n317323 );
or ( n317442 , n317440 , n27015 );
buf ( n317443 , n317442 );
buf ( n317444 , n317443 );
xor ( n317445 , n317438 , n317444 );
xor ( n27020 , n317259 , n26841 );
and ( n27021 , n27020 , n317284 );
and ( n27022 , n317259 , n26841 );
or ( n317449 , n27021 , n27022 );
buf ( n317450 , n317449 );
xor ( n27025 , n317445 , n317450 );
buf ( n317452 , n27025 );
buf ( n317453 , n317452 );
xor ( n27028 , n317432 , n317453 );
buf ( n317455 , n27028 );
buf ( n317456 , n317455 );
buf ( n317457 , n313215 );
buf ( n317458 , n317318 );
or ( n27033 , n317457 , n317458 );
buf ( n317460 , n313224 );
buf ( n317461 , n866 );
buf ( n317462 , n305117 );
and ( n27037 , n317461 , n317462 );
not ( n27038 , n317461 );
buf ( n317465 , n843 );
and ( n27040 , n27038 , n317465 );
nor ( n27041 , n27037 , n27040 );
buf ( n317468 , n27041 );
buf ( n317469 , n317468 );
or ( n27044 , n317460 , n317469 );
nand ( n27045 , n27033 , n27044 );
buf ( n317472 , n27045 );
buf ( n317473 , n310726 );
buf ( n317474 , n317355 );
or ( n27049 , n317473 , n317474 );
buf ( n317476 , n305205 );
buf ( n317477 , n310521 );
buf ( n317478 , n841 );
and ( n317479 , n317477 , n317478 );
buf ( n317480 , n310600 );
buf ( n317481 , n868 );
and ( n27056 , n317480 , n317481 );
nor ( n317483 , n317479 , n27056 );
buf ( n317484 , n317483 );
buf ( n317485 , n317484 );
or ( n27060 , n317476 , n317485 );
nand ( n317487 , n27049 , n27060 );
buf ( n317488 , n317487 );
xor ( n27063 , n317472 , n317488 );
buf ( n317490 , n15836 );
buf ( n317491 , n317255 );
not ( n317492 , n317491 );
buf ( n317493 , n317492 );
buf ( n317494 , n317493 );
and ( n317495 , n317490 , n317494 );
buf ( n317496 , n306272 );
buf ( n317497 , n878 );
and ( n317498 , n317496 , n317497 );
nor ( n317499 , n317495 , n317498 );
buf ( n317500 , n317499 );
xor ( n27075 , n27063 , n317500 );
buf ( n317502 , n847 );
buf ( n317503 , n864 );
and ( n27078 , n317502 , n317503 );
buf ( n317505 , n27078 );
buf ( n317506 , n317505 );
buf ( n317507 , n317299 );
not ( n317508 , n317507 );
buf ( n317509 , n304851 );
not ( n27084 , n317509 );
or ( n317511 , n317508 , n27084 );
buf ( n317512 , n304864 );
buf ( n317513 , n872 );
buf ( n317514 , n837 );
and ( n317515 , n317513 , n317514 );
not ( n317516 , n317513 );
buf ( n317517 , n313757 );
and ( n317518 , n317516 , n317517 );
nor ( n317519 , n317515 , n317518 );
buf ( n317520 , n317519 );
buf ( n317521 , n317520 );
nand ( n27096 , n317512 , n317521 );
buf ( n317523 , n27096 );
buf ( n317524 , n317523 );
nand ( n317525 , n317511 , n317524 );
buf ( n317526 , n317525 );
buf ( n317527 , n317526 );
xor ( n317528 , n317506 , n317527 );
buf ( n317529 , n311891 );
buf ( n317530 , n317336 );
or ( n317531 , n317529 , n317530 );
buf ( n317532 , n311246 );
buf ( n317533 , n845 );
buf ( n317534 , n311234 );
and ( n317535 , n317533 , n317534 );
not ( n317536 , n317533 );
buf ( n317537 , n864 );
and ( n317538 , n317536 , n317537 );
nor ( n317539 , n317535 , n317538 );
buf ( n317540 , n317539 );
buf ( n317541 , n317540 );
or ( n317542 , n317532 , n317541 );
nand ( n27117 , n317531 , n317542 );
buf ( n317544 , n27117 );
buf ( n317545 , n317544 );
xor ( n27120 , n317528 , n317545 );
buf ( n317547 , n27120 );
buf ( n317548 , n314219 );
buf ( n317549 , n317198 );
or ( n317550 , n317548 , n317549 );
buf ( n27125 , n304760 );
buf ( n317552 , n870 );
buf ( n317553 , n14992 );
and ( n317554 , n317552 , n317553 );
not ( n317555 , n317552 );
buf ( n317556 , n839 );
and ( n27131 , n317555 , n317556 );
nor ( n317558 , n317554 , n27131 );
buf ( n317559 , n317558 );
buf ( n317560 , n317559 );
or ( n317561 , n27125 , n317560 );
nand ( n27136 , n317550 , n317561 );
buf ( n317563 , n27136 );
buf ( n27138 , n317563 );
buf ( n317565 , n306340 );
buf ( n317566 , n317280 );
or ( n317567 , n317565 , n317566 );
buf ( n27142 , n305298 );
buf ( n317569 , n874 );
buf ( n317570 , n21261 );
and ( n317571 , n317569 , n317570 );
not ( n27146 , n317569 );
buf ( n317573 , n835 );
and ( n317574 , n27146 , n317573 );
nor ( n27149 , n317571 , n317574 );
buf ( n317576 , n27149 );
buf ( n317577 , n317576 );
or ( n27152 , n27142 , n317577 );
nand ( n317579 , n317567 , n27152 );
buf ( n317580 , n317579 );
buf ( n317581 , n317580 );
xor ( n317582 , n27138 , n317581 );
buf ( n317583 , n305650 );
buf ( n317584 , n317220 );
or ( n317585 , n317583 , n317584 );
buf ( n317586 , n305664 );
buf ( n317587 , n876 );
buf ( n317588 , n310964 );
and ( n27163 , n317587 , n317588 );
not ( n317590 , n317587 );
buf ( n317591 , n833 );
and ( n27166 , n317590 , n317591 );
nor ( n27167 , n27163 , n27166 );
buf ( n317594 , n27167 );
buf ( n317595 , n317594 );
or ( n317596 , n317586 , n317595 );
nand ( n27171 , n317585 , n317596 );
buf ( n317598 , n27171 );
buf ( n317599 , n317598 );
xor ( n317600 , n317582 , n317599 );
buf ( n317601 , n317600 );
xor ( n27176 , n317547 , n317601 );
xor ( n27177 , n27075 , n27176 );
buf ( n317604 , n27177 );
xor ( n317605 , n317259 , n26841 );
xor ( n317606 , n317605 , n317284 );
and ( n27181 , n317343 , n317606 );
xor ( n317608 , n317259 , n26841 );
xor ( n27183 , n317608 , n317284 );
and ( n317610 , n317370 , n27183 );
and ( n27185 , n317343 , n317370 );
or ( n317612 , n27181 , n317610 , n27185 );
buf ( n317613 , n317612 );
xor ( n27188 , n317604 , n317613 );
xor ( n317615 , n317164 , n317170 );
and ( n27190 , n317615 , n317231 );
and ( n317617 , n317164 , n317170 );
or ( n27192 , n27190 , n317617 );
buf ( n317619 , n27192 );
buf ( n317620 , n317619 );
xor ( n27195 , n27188 , n317620 );
buf ( n317622 , n27195 );
buf ( n317623 , n317622 );
xor ( n317624 , n317243 , n317373 );
and ( n27199 , n317624 , n317380 );
and ( n317626 , n317243 , n317373 );
or ( n27201 , n27199 , n317626 );
buf ( n317628 , n27201 );
buf ( n317629 , n317628 );
xor ( n317630 , n317456 , n317623 );
xor ( n27205 , n317630 , n317629 );
buf ( n317632 , n27205 );
xor ( n317633 , n317456 , n317623 );
and ( n27208 , n317633 , n317629 );
and ( n317635 , n317456 , n317623 );
or ( n27210 , n27208 , n317635 );
buf ( n317637 , n27210 );
xor ( n317638 , n316424 , n316589 );
and ( n317639 , n317638 , n316822 );
and ( n27214 , n316424 , n316589 );
or ( n317641 , n317639 , n27214 );
buf ( n317642 , n317641 );
buf ( n317643 , n317642 );
xor ( n317644 , n316376 , n316401 );
and ( n317645 , n317644 , n316418 );
and ( n317646 , n316376 , n316401 );
or ( n27221 , n317645 , n317646 );
buf ( n317648 , n27221 );
buf ( n317649 , n317648 );
and ( n317650 , n315730 , n315731 );
buf ( n317651 , n317650 );
buf ( n317652 , n317651 );
buf ( n27227 , n316330 );
not ( n27228 , n27227 );
buf ( n317655 , n305338 );
not ( n27230 , n317655 );
or ( n317657 , n27228 , n27230 );
buf ( n317658 , n305344 );
buf ( n317659 , n312010 );
nand ( n317660 , n317658 , n317659 );
buf ( n317661 , n317660 );
buf ( n317662 , n317661 );
nand ( n317663 , n317657 , n317662 );
buf ( n317664 , n317663 );
buf ( n317665 , n317664 );
xor ( n317666 , n317652 , n317665 );
buf ( n317667 , n316316 );
not ( n27242 , n317667 );
buf ( n317669 , n15836 );
not ( n317670 , n317669 );
or ( n317671 , n27242 , n317670 );
buf ( n317672 , n306272 );
buf ( n317673 , n312162 );
nand ( n317674 , n317672 , n317673 );
buf ( n317675 , n317674 );
buf ( n317676 , n317675 );
nand ( n317677 , n317671 , n317676 );
buf ( n317678 , n317677 );
buf ( n317679 , n317678 );
xor ( n27254 , n317666 , n317679 );
buf ( n317681 , n27254 );
buf ( n317682 , n317681 );
xor ( n317683 , n317649 , n317682 );
buf ( n27258 , n304697 );
not ( n317685 , n27258 );
buf ( n317686 , n317685 );
buf ( n317687 , n317686 );
not ( n317688 , n317687 );
buf ( n317689 , n305489 );
not ( n317690 , n317689 );
or ( n317691 , n317688 , n317690 );
buf ( n317692 , n892 );
nand ( n317693 , n317691 , n317692 );
buf ( n317694 , n317693 );
buf ( n317695 , n317694 );
buf ( n317696 , n316512 );
not ( n27271 , n317696 );
buf ( n317698 , n304912 );
not ( n317699 , n317698 );
or ( n27274 , n27271 , n317699 );
buf ( n317701 , n304901 );
buf ( n317702 , n312207 );
nand ( n317703 , n317701 , n317702 );
buf ( n317704 , n317703 );
buf ( n317705 , n317704 );
nand ( n317706 , n27274 , n317705 );
buf ( n317707 , n317706 );
buf ( n317708 , n317707 );
xor ( n317709 , n317695 , n317708 );
buf ( n317710 , n304630 );
buf ( n317711 , n316493 );
or ( n317712 , n317710 , n317711 );
buf ( n317713 , n304655 );
buf ( n317714 , n311978 );
not ( n27289 , n317714 );
buf ( n317716 , n27289 );
buf ( n317717 , n317716 );
or ( n27292 , n317713 , n317717 );
nand ( n317719 , n317712 , n27292 );
buf ( n317720 , n317719 );
buf ( n317721 , n317720 );
xor ( n317722 , n317709 , n317721 );
buf ( n317723 , n317722 );
buf ( n317724 , n317723 );
xor ( n317725 , n317683 , n317724 );
buf ( n317726 , n317725 );
buf ( n317727 , n317726 );
buf ( n27302 , n26044 );
not ( n27303 , n27302 );
buf ( n27304 , n311998 );
not ( n27305 , n27304 );
or ( n27306 , n27303 , n27305 );
buf ( n27307 , n305144 );
buf ( n27308 , n21566 );
nand ( n27309 , n27307 , n27308 );
buf ( n27310 , n27309 );
buf ( n27311 , n27310 );
nand ( n27312 , n27306 , n27311 );
buf ( n27313 , n27312 );
buf ( n317740 , n27313 );
buf ( n317741 , n26105 );
not ( n317742 , n317741 );
buf ( n317743 , n304584 );
not ( n27318 , n317743 );
or ( n317745 , n317742 , n27318 );
buf ( n317746 , n304596 );
buf ( n317747 , n21651 );
nand ( n27322 , n317746 , n317747 );
buf ( n317749 , n27322 );
buf ( n317750 , n317749 );
nand ( n27325 , n317745 , n317750 );
buf ( n317752 , n27325 );
buf ( n317753 , n317752 );
xor ( n27328 , n317740 , n317753 );
buf ( n317755 , n316574 );
not ( n27330 , n317755 );
buf ( n317757 , n14323 );
not ( n317758 , n317757 );
or ( n27333 , n27330 , n317758 );
buf ( n317760 , n304763 );
buf ( n317761 , n312190 );
nand ( n27336 , n317760 , n317761 );
buf ( n317763 , n27336 );
buf ( n317764 , n317763 );
nand ( n317765 , n27333 , n317764 );
buf ( n317766 , n317765 );
buf ( n317767 , n317766 );
xor ( n317768 , n27328 , n317767 );
buf ( n317769 , n317768 );
buf ( n317770 , n317769 );
buf ( n317771 , n316451 );
not ( n27346 , n317771 );
buf ( n317773 , n305292 );
not ( n317774 , n317773 );
or ( n27349 , n27346 , n317774 );
buf ( n317776 , n305289 );
buf ( n317777 , n312056 );
nand ( n27352 , n317776 , n317777 );
buf ( n317779 , n27352 );
buf ( n317780 , n317779 );
nand ( n317781 , n27349 , n317780 );
buf ( n317782 , n317781 );
buf ( n317783 , n317782 );
buf ( n317784 , n316350 );
not ( n317785 , n317784 );
buf ( n317786 , n317785 );
buf ( n317787 , n317786 );
not ( n27362 , n317787 );
buf ( n317789 , n304813 );
not ( n317790 , n317789 );
or ( n317791 , n27362 , n317790 );
buf ( n317792 , n304807 );
buf ( n317793 , n312032 );
nand ( n27368 , n317792 , n317793 );
buf ( n317795 , n27368 );
buf ( n317796 , n317795 );
nand ( n27371 , n317791 , n317796 );
buf ( n317798 , n27371 );
buf ( n27373 , n317798 );
xor ( n27374 , n317783 , n27373 );
buf ( n317801 , n304854 );
buf ( n317802 , n316431 );
not ( n27377 , n317802 );
buf ( n317804 , n27377 );
buf ( n317805 , n317804 );
or ( n317806 , n317801 , n317805 );
not ( n317807 , n304845 );
buf ( n317808 , n317807 );
buf ( n317809 , n21674 );
or ( n27384 , n317808 , n317809 );
nand ( n27385 , n317806 , n27384 );
buf ( n317812 , n27385 );
buf ( n317813 , n317812 );
xor ( n27388 , n27374 , n317813 );
buf ( n317815 , n27388 );
buf ( n317816 , n317815 );
xor ( n317817 , n317770 , n317816 );
buf ( n317818 , n316394 );
not ( n317819 , n317818 );
buf ( n317820 , n310694 );
not ( n27395 , n317820 );
or ( n317822 , n317819 , n27395 );
buf ( n317823 , n311107 );
buf ( n317824 , n21713 );
nand ( n27399 , n317823 , n317824 );
buf ( n317826 , n27399 );
buf ( n317827 , n317826 );
nand ( n317828 , n317822 , n317827 );
buf ( n317829 , n317828 );
buf ( n317830 , n317829 );
buf ( n317831 , n316552 );
not ( n27406 , n317831 );
buf ( n317833 , n305213 );
not ( n317834 , n317833 );
or ( n27409 , n27406 , n317834 );
buf ( n317836 , n305219 );
buf ( n317837 , n312122 );
nand ( n27412 , n317836 , n317837 );
buf ( n317839 , n27412 );
buf ( n317840 , n317839 );
nand ( n27415 , n27409 , n317840 );
buf ( n27416 , n27415 );
buf ( n317843 , n27416 );
xor ( n27418 , n317830 , n317843 );
buf ( n317845 , n304987 );
buf ( n317846 , n316413 );
or ( n317847 , n317845 , n317846 );
buf ( n317848 , n311075 );
buf ( n317849 , n312233 );
or ( n317850 , n317848 , n317849 );
nand ( n317851 , n317847 , n317850 );
buf ( n317852 , n317851 );
buf ( n317853 , n317852 );
xor ( n27428 , n27418 , n317853 );
buf ( n317855 , n27428 );
buf ( n317856 , n317855 );
xor ( n317857 , n317817 , n317856 );
buf ( n317858 , n317857 );
buf ( n317859 , n317858 );
xor ( n317860 , n317727 , n317859 );
buf ( n317861 , n894 );
not ( n317862 , n317861 );
buf ( n317863 , n317862 );
buf ( n317864 , n317863 );
buf ( n317865 , n316015 );
not ( n27440 , n317865 );
buf ( n317867 , n14272 );
not ( n27442 , n317867 );
or ( n317869 , n27440 , n27442 );
buf ( n27444 , n305430 );
buf ( n317871 , n892 );
nand ( n317872 , n27444 , n317871 );
buf ( n317873 , n317872 );
buf ( n317874 , n317873 );
nand ( n317875 , n317869 , n317874 );
buf ( n317876 , n317875 );
buf ( n317877 , n317876 );
not ( n317878 , n317877 );
buf ( n317879 , n317878 );
buf ( n317880 , n317879 );
xor ( n317881 , n317864 , n317880 );
xor ( n317882 , n315719 , n315740 );
and ( n27457 , n317882 , n315763 );
and ( n317884 , n315719 , n315740 );
or ( n317885 , n27457 , n317884 );
buf ( n317886 , n317885 );
buf ( n317887 , n317886 );
and ( n27462 , n317881 , n317887 );
and ( n27463 , n317864 , n317880 );
or ( n27464 , n27462 , n27463 );
buf ( n317891 , n27464 );
buf ( n317892 , n317891 );
buf ( n317893 , n317876 );
buf ( n317894 , n316369 );
not ( n317895 , n317894 );
buf ( n317896 , n311888 );
not ( n27471 , n317896 );
or ( n317898 , n317895 , n27471 );
buf ( n317899 , n310582 );
xor ( n317900 , n311880 , n311881 );
buf ( n317901 , n317900 );
buf ( n317902 , n317901 );
nand ( n317903 , n317899 , n317902 );
buf ( n317904 , n317903 );
buf ( n317905 , n317904 );
nand ( n317906 , n317898 , n317905 );
buf ( n317907 , n317906 );
buf ( n317908 , n317907 );
xor ( n317909 , n317893 , n317908 );
xor ( n317910 , n316483 , n316500 );
and ( n317911 , n317910 , n316520 );
and ( n317912 , n316483 , n316500 );
or ( n27487 , n317911 , n317912 );
buf ( n317914 , n27487 );
buf ( n317915 , n317914 );
xor ( n27490 , n317909 , n317915 );
buf ( n317917 , n27490 );
buf ( n317918 , n317917 );
xor ( n27493 , n317892 , n317918 );
xor ( n317920 , n316069 , n316087 );
and ( n317921 , n317920 , n316111 );
and ( n27496 , n316069 , n316087 );
or ( n317923 , n317921 , n27496 );
buf ( n317924 , n317923 );
buf ( n317925 , n317924 );
xor ( n27500 , n315993 , n316022 );
and ( n317927 , n27500 , n316048 );
and ( n317928 , n315993 , n316022 );
or ( n27503 , n317927 , n317928 );
buf ( n317930 , n27503 );
buf ( n27505 , n317930 );
xor ( n27506 , n317925 , n27505 );
xor ( n317933 , n315926 , n315940 );
and ( n27508 , n317933 , n315962 );
and ( n27509 , n315926 , n315940 );
or ( n27510 , n27508 , n27509 );
buf ( n317937 , n27510 );
buf ( n317938 , n317937 );
and ( n317939 , n27506 , n317938 );
and ( n27514 , n317925 , n27505 );
or ( n27515 , n317939 , n27514 );
buf ( n317942 , n27515 );
buf ( n317943 , n317942 );
xor ( n317944 , n27493 , n317943 );
buf ( n317945 , n317944 );
buf ( n317946 , n317945 );
xor ( n317947 , n317860 , n317946 );
buf ( n317948 , n317947 );
buf ( n317949 , n317948 );
xor ( n27524 , n317068 , n26648 );
and ( n317951 , n27524 , n317137 );
and ( n317952 , n317068 , n26648 );
or ( n27527 , n317951 , n317952 );
buf ( n317954 , n27527 );
buf ( n317955 , n317954 );
xor ( n27530 , n317864 , n317880 );
xor ( n317957 , n27530 , n317887 );
buf ( n317958 , n317957 );
buf ( n317959 , n317958 );
xor ( n27534 , n315766 , n315840 );
and ( n317961 , n27534 , n315906 );
and ( n317962 , n315766 , n315840 );
or ( n27537 , n317961 , n317962 );
buf ( n317964 , n27537 );
buf ( n317965 , n317964 );
xor ( n317966 , n317959 , n317965 );
xor ( n27541 , n315965 , n316051 );
and ( n27542 , n27541 , n316114 );
and ( n27543 , n315965 , n316051 );
or ( n317970 , n27542 , n27543 );
buf ( n317971 , n317970 );
buf ( n317972 , n317971 );
xor ( n27547 , n317966 , n317972 );
buf ( n317974 , n27547 );
buf ( n317975 , n317974 );
xor ( n27550 , n317955 , n317975 );
xor ( n317977 , n316603 , n316604 );
and ( n27552 , n317977 , n316650 );
and ( n27553 , n316603 , n316604 );
or ( n317980 , n27552 , n27553 );
buf ( n317981 , n317980 );
buf ( n317982 , n317981 );
xor ( n27557 , n316668 , n316733 );
and ( n317984 , n27557 , n316795 );
and ( n317985 , n316668 , n316733 );
or ( n27560 , n317984 , n317985 );
buf ( n317987 , n27560 );
buf ( n317988 , n317987 );
xor ( n317989 , n317982 , n317988 );
xor ( n27564 , n317925 , n27505 );
xor ( n317991 , n27564 , n317938 );
buf ( n317992 , n317991 );
buf ( n317993 , n317992 );
xor ( n27568 , n317989 , n317993 );
buf ( n317995 , n27568 );
buf ( n317996 , n317995 );
and ( n317997 , n27550 , n317996 );
and ( n317998 , n317955 , n317975 );
or ( n27573 , n317997 , n317998 );
buf ( n318000 , n27573 );
buf ( n318001 , n318000 );
xor ( n27576 , n317643 , n317949 );
xor ( n318003 , n27576 , n318001 );
buf ( n318004 , n318003 );
xor ( n318005 , n317643 , n317949 );
and ( n27580 , n318005 , n318001 );
and ( n318007 , n317643 , n317949 );
or ( n27582 , n27580 , n318007 );
buf ( n318009 , n27582 );
xor ( n318010 , n317081 , n317087 );
xor ( n27585 , n318010 , n317132 );
buf ( n318012 , n27585 );
buf ( n318013 , n318012 );
xor ( n27588 , n316803 , n316807 );
xor ( n27589 , n27588 , n316812 );
buf ( n318016 , n27589 );
buf ( n318017 , n318016 );
xor ( n27592 , n318013 , n318017 );
xor ( n27593 , n317101 , n317114 );
xor ( n27594 , n27593 , n317127 );
buf ( n318021 , n27594 );
buf ( n318022 , n318021 );
xor ( n27597 , n316890 , n316872 );
buf ( n318024 , n27597 );
buf ( n318025 , n316858 );
xor ( n27600 , n318024 , n318025 );
buf ( n318027 , n27600 );
buf ( n318028 , n318027 );
xor ( n318029 , n318022 , n318028 );
xor ( n318030 , n313272 , n313278 );
and ( n27605 , n318030 , n313285 );
and ( n318032 , n313272 , n313278 );
or ( n27607 , n27605 , n318032 );
buf ( n318034 , n27607 );
buf ( n318035 , n318034 );
and ( n318036 , n318029 , n318035 );
and ( n318037 , n318022 , n318028 );
or ( n27612 , n318036 , n318037 );
buf ( n318039 , n27612 );
buf ( n318040 , n318039 );
and ( n318041 , n27592 , n318040 );
and ( n27616 , n318013 , n318017 );
or ( n318043 , n318041 , n27616 );
buf ( n318044 , n318043 );
buf ( n318045 , n318044 );
xor ( n27620 , n315909 , n316117 );
xor ( n318047 , n27620 , n316296 );
buf ( n318048 , n318047 );
buf ( n318049 , n318048 );
xor ( n27624 , n316187 , n316266 );
xor ( n27625 , n27624 , n316291 );
buf ( n318052 , n27625 );
buf ( n27627 , n318052 );
xor ( n318054 , n313237 , n313240 );
and ( n27629 , n318054 , n313247 );
and ( n318056 , n313237 , n313240 );
or ( n318057 , n27629 , n318056 );
buf ( n318058 , n318057 );
buf ( n318059 , n318058 );
xor ( n318060 , n316828 , n316834 );
xor ( n27635 , n318060 , n316841 );
buf ( n318062 , n27635 );
buf ( n318063 , n318062 );
xor ( n27638 , n318059 , n318063 );
xor ( n318065 , n25847 , n316279 );
xor ( n318066 , n318065 , n316286 );
buf ( n318067 , n318066 );
buf ( n318068 , n318067 );
and ( n318069 , n27638 , n318068 );
and ( n27644 , n318059 , n318063 );
or ( n318071 , n318069 , n27644 );
buf ( n318072 , n318071 );
buf ( n318073 , n318072 );
xor ( n318074 , n27627 , n318073 );
xor ( n27649 , n312331 , n312393 );
and ( n318076 , n27649 , n312483 );
and ( n27651 , n312331 , n312393 );
or ( n318078 , n318076 , n27651 );
buf ( n318079 , n318078 );
buf ( n318080 , n318079 );
xor ( n318081 , n313301 , n313360 );
and ( n318082 , n318081 , n313422 );
and ( n27657 , n313301 , n313360 );
or ( n318084 , n318082 , n27657 );
buf ( n318085 , n318084 );
buf ( n318086 , n318085 );
xor ( n318087 , n318080 , n318086 );
xor ( n27662 , n316956 , n316998 );
xor ( n318089 , n27662 , n317052 );
buf ( n318090 , n318089 );
buf ( n318091 , n318090 );
and ( n318092 , n318087 , n318091 );
and ( n27667 , n318080 , n318086 );
or ( n318094 , n318092 , n27667 );
buf ( n318095 , n318094 );
buf ( n318096 , n318095 );
and ( n318097 , n318074 , n318096 );
and ( n27672 , n27627 , n318073 );
or ( n318099 , n318097 , n27672 );
buf ( n318100 , n318099 );
buf ( n318101 , n318100 );
xor ( n318102 , n318045 , n318049 );
xor ( n27677 , n318102 , n318101 );
buf ( n318104 , n27677 );
xor ( n318105 , n318045 , n318049 );
and ( n318106 , n318105 , n318101 );
and ( n318107 , n318045 , n318049 );
or ( n27682 , n318106 , n318107 );
buf ( n318109 , n27682 );
xor ( n318110 , n26420 , n316951 );
xor ( n27685 , n318110 , n317057 );
buf ( n318112 , n27685 );
buf ( n318113 , n318112 );
xor ( n27688 , n318013 , n318017 );
xor ( n318115 , n27688 , n318040 );
buf ( n318116 , n318115 );
buf ( n318117 , n318116 );
xor ( n318118 , n27627 , n318073 );
xor ( n27693 , n318118 , n318096 );
buf ( n318120 , n27693 );
buf ( n318121 , n318120 );
xor ( n27696 , n318113 , n318117 );
xor ( n27697 , n27696 , n318121 );
buf ( n318124 , n27697 );
xor ( n318125 , n318113 , n318117 );
and ( n318126 , n318125 , n318121 );
and ( n27701 , n318113 , n318117 );
or ( n318128 , n318126 , n27701 );
buf ( n318129 , n318128 );
xor ( n27704 , n311949 , n311953 );
xor ( n318131 , n27704 , n312267 );
buf ( n318132 , n318131 );
xor ( n27707 , n311935 , n311939 );
xor ( n27708 , n27707 , n311944 );
buf ( n318135 , n27708 );
buf ( n27710 , n318135 );
xor ( n318137 , n311874 , n311878 );
xor ( n318138 , n318137 , n311930 );
buf ( n318139 , n318138 );
not ( n318140 , n318139 );
xor ( n318141 , n311621 , n311642 );
xor ( n27716 , n318141 , n311656 );
buf ( n318143 , n27716 );
buf ( n318144 , n318143 );
xor ( n27719 , n311808 , n311820 );
xor ( n318146 , n27719 , n311837 );
buf ( n318147 , n318146 );
buf ( n318148 , n318147 );
xor ( n318149 , n318144 , n318148 );
xor ( n318150 , n21458 , n311904 );
xor ( n27725 , n318150 , n311925 );
buf ( n318152 , n27725 );
buf ( n318153 , n318152 );
and ( n318154 , n318149 , n318153 );
and ( n318155 , n318144 , n318148 );
or ( n27730 , n318154 , n318155 );
buf ( n318157 , n27730 );
not ( n318158 , n318157 );
nand ( n27733 , n318140 , n318158 );
not ( n318160 , n27733 );
buf ( n318161 , n311729 );
buf ( n318162 , n21253 );
xnor ( n318163 , n318161 , n318162 );
buf ( n318164 , n318163 );
buf ( n318165 , n318164 );
buf ( n318166 , n21281 );
xnor ( n318167 , n318165 , n318166 );
buf ( n318168 , n318167 );
buf ( n318169 , n318168 );
and ( n318170 , n316366 , n316367 );
buf ( n318171 , n318170 );
buf ( n318172 , n318171 );
buf ( n318173 , n317901 );
not ( n318174 , n318173 );
buf ( n318175 , n310576 );
not ( n27750 , n318175 );
or ( n318177 , n318174 , n27750 );
buf ( n318178 , n311896 );
not ( n27753 , n318178 );
buf ( n318180 , n310582 );
nand ( n318181 , n27753 , n318180 );
buf ( n318182 , n318181 );
buf ( n318183 , n318182 );
nand ( n27758 , n318177 , n318183 );
buf ( n318185 , n27758 );
buf ( n318186 , n318185 );
xor ( n318187 , n318172 , n318186 );
buf ( n318188 , n311990 );
not ( n27763 , n318188 );
buf ( n318190 , n27763 );
buf ( n318191 , n318190 );
and ( n318192 , n318187 , n318191 );
and ( n27767 , n318172 , n318186 );
or ( n27768 , n318192 , n27767 );
buf ( n318195 , n27768 );
buf ( n318196 , n318195 );
xor ( n318197 , n318169 , n318196 );
xor ( n27772 , n317652 , n317665 );
and ( n318199 , n27772 , n317679 );
and ( n318200 , n317652 , n317665 );
or ( n27775 , n318199 , n318200 );
buf ( n318202 , n27775 );
buf ( n27777 , n318202 );
xor ( n318204 , n317695 , n317708 );
and ( n318205 , n318204 , n317721 );
and ( n27780 , n317695 , n317708 );
or ( n318207 , n318205 , n27780 );
buf ( n318208 , n318207 );
buf ( n318209 , n318208 );
xor ( n318210 , n27777 , n318209 );
xor ( n27785 , n317783 , n27373 );
and ( n27786 , n27785 , n317813 );
and ( n318213 , n317783 , n27373 );
or ( n318214 , n27786 , n318213 );
buf ( n318215 , n318214 );
buf ( n318216 , n318215 );
and ( n318217 , n318210 , n318216 );
and ( n318218 , n27777 , n318209 );
or ( n27793 , n318217 , n318218 );
buf ( n318220 , n27793 );
buf ( n318221 , n318220 );
and ( n27796 , n318197 , n318221 );
and ( n318223 , n318169 , n318196 );
or ( n318224 , n27796 , n318223 );
buf ( n318225 , n318224 );
not ( n318226 , n318225 );
or ( n318227 , n318160 , n318226 );
nand ( n27802 , n318139 , n318157 );
nand ( n318229 , n318227 , n27802 );
buf ( n318230 , n318229 );
xor ( n27805 , n311969 , n311973 );
xor ( n318232 , n27805 , n312262 );
buf ( n318233 , n318232 );
buf ( n318234 , n318233 );
xor ( n318235 , n27710 , n318230 );
xor ( n318236 , n318235 , n318234 );
buf ( n318237 , n318236 );
xor ( n27812 , n27710 , n318230 );
and ( n318239 , n27812 , n318234 );
and ( n318240 , n27710 , n318230 );
or ( n27815 , n318239 , n318240 );
buf ( n318242 , n27815 );
xor ( n318243 , n318059 , n318063 );
xor ( n27818 , n318243 , n318068 );
buf ( n318245 , n27818 );
buf ( n318246 , n318245 );
xor ( n27821 , n318080 , n318086 );
xor ( n27822 , n27821 , n318091 );
buf ( n318249 , n27822 );
buf ( n318250 , n318249 );
xor ( n318251 , n312486 , n312752 );
and ( n27826 , n318251 , n312995 );
and ( n27827 , n312486 , n312752 );
or ( n27828 , n27826 , n27827 );
buf ( n27829 , n27828 );
buf ( n318256 , n27829 );
xor ( n27831 , n318246 , n318250 );
xor ( n27832 , n27831 , n318256 );
buf ( n318259 , n27832 );
xor ( n27834 , n318246 , n318250 );
and ( n318261 , n27834 , n318256 );
and ( n318262 , n318246 , n318250 );
or ( n27837 , n318261 , n318262 );
buf ( n318264 , n27837 );
xor ( n27839 , n313266 , n313428 );
and ( n27840 , n27839 , n313435 );
and ( n318267 , n313266 , n313428 );
or ( n27842 , n27840 , n318267 );
buf ( n318269 , n27842 );
buf ( n318270 , n317500 );
not ( n27845 , n318270 );
buf ( n318272 , n27845 );
xor ( n318273 , n317506 , n317527 );
and ( n318274 , n318273 , n317545 );
and ( n27849 , n317506 , n317527 );
or ( n318276 , n318274 , n27849 );
buf ( n318277 , n318276 );
xor ( n27852 , n318272 , n318277 );
xor ( n318279 , n27138 , n317581 );
and ( n318280 , n318279 , n317599 );
and ( n27855 , n27138 , n317581 );
or ( n318282 , n318280 , n27855 );
buf ( n318283 , n318282 );
xor ( n318284 , n27852 , n318283 );
xor ( n27859 , n317472 , n317488 );
and ( n318286 , n27859 , n317500 );
and ( n27861 , n317472 , n317488 );
or ( n27862 , n318286 , n27861 );
xor ( n318289 , n317438 , n317444 );
and ( n318290 , n318289 , n317450 );
and ( n318291 , n317438 , n317444 );
or ( n27866 , n318290 , n318291 );
buf ( n318293 , n27866 );
xor ( n318294 , n27862 , n318293 );
xor ( n27869 , n318284 , n318294 );
buf ( n318296 , n27869 );
xor ( n318297 , n317604 , n317613 );
and ( n27872 , n318297 , n317620 );
and ( n318299 , n317604 , n317613 );
or ( n27874 , n27872 , n318299 );
buf ( n318301 , n27874 );
buf ( n318302 , n318301 );
buf ( n318303 , n846 );
buf ( n318304 , n864 );
and ( n318305 , n318303 , n318304 );
buf ( n318306 , n318305 );
buf ( n318307 , n318306 );
buf ( n318308 , n317559 );
not ( n27883 , n318308 );
buf ( n318310 , n27883 );
buf ( n318311 , n318310 );
not ( n318312 , n318311 );
buf ( n318313 , n304754 );
not ( n27888 , n318313 );
or ( n318315 , n318312 , n27888 );
buf ( n318316 , n304763 );
buf ( n318317 , n870 );
buf ( n318318 , n838 );
and ( n318319 , n318317 , n318318 );
not ( n27894 , n318317 );
buf ( n318321 , n310377 );
and ( n27896 , n27894 , n318321 );
nor ( n318323 , n318319 , n27896 );
buf ( n318324 , n318323 );
buf ( n318325 , n318324 );
nand ( n318326 , n318316 , n318325 );
buf ( n318327 , n318326 );
buf ( n318328 , n318327 );
nand ( n318329 , n318315 , n318328 );
buf ( n318330 , n318329 );
buf ( n318331 , n318330 );
xor ( n318332 , n318307 , n318331 );
buf ( n318333 , n311891 );
buf ( n318334 , n317540 );
or ( n27909 , n318333 , n318334 );
buf ( n318336 , n311246 );
buf ( n318337 , n844 );
buf ( n318338 , n864 );
xnor ( n318339 , n318337 , n318338 );
buf ( n318340 , n318339 );
buf ( n318341 , n318340 );
or ( n318342 , n318336 , n318341 );
nand ( n27917 , n27909 , n318342 );
buf ( n318344 , n27917 );
buf ( n318345 , n318344 );
xor ( n318346 , n318332 , n318345 );
buf ( n318347 , n318346 );
buf ( n318348 , n317468 );
not ( n318349 , n318348 );
buf ( n318350 , n318349 );
buf ( n318351 , n318350 );
not ( n318352 , n318351 );
buf ( n318353 , n310694 );
not ( n27928 , n318353 );
or ( n318355 , n318352 , n27928 );
buf ( n27930 , n310483 );
buf ( n318357 , n866 );
buf ( n318358 , n842 );
and ( n318359 , n318357 , n318358 );
not ( n318360 , n318357 );
buf ( n318361 , n304610 );
and ( n318362 , n318360 , n318361 );
nor ( n318363 , n318359 , n318362 );
buf ( n318364 , n318363 );
buf ( n318365 , n318364 );
nand ( n27940 , n27930 , n318365 );
buf ( n318367 , n27940 );
buf ( n318368 , n318367 );
nand ( n27943 , n318355 , n318368 );
buf ( n318370 , n27943 );
buf ( n318371 , n318370 );
buf ( n318372 , n317576 );
not ( n318373 , n318372 );
buf ( n318374 , n318373 );
buf ( n318375 , n318374 );
not ( n27950 , n318375 );
buf ( n318377 , n305627 );
not ( n318378 , n318377 );
or ( n27953 , n27950 , n318378 );
buf ( n318380 , n315090 );
buf ( n318381 , n834 );
and ( n318382 , n318380 , n318381 );
buf ( n318383 , n310658 );
buf ( n318384 , n874 );
and ( n27959 , n318383 , n318384 );
nor ( n318386 , n318382 , n27959 );
buf ( n318387 , n318386 );
buf ( n318388 , n318387 );
not ( n27963 , n318388 );
buf ( n318390 , n305301 );
nand ( n318391 , n27963 , n318390 );
buf ( n318392 , n318391 );
buf ( n318393 , n318392 );
nand ( n27968 , n27953 , n318393 );
buf ( n318395 , n27968 );
buf ( n318396 , n318395 );
xor ( n318397 , n318371 , n318396 );
buf ( n318398 , n310726 );
buf ( n318399 , n317484 );
or ( n27974 , n318398 , n318399 );
buf ( n318401 , n305205 );
buf ( n318402 , n310521 );
buf ( n318403 , n840 );
and ( n318404 , n318402 , n318403 );
buf ( n318405 , n305261 );
buf ( n318406 , n868 );
and ( n318407 , n318405 , n318406 );
nor ( n318408 , n318404 , n318407 );
buf ( n318409 , n318408 );
buf ( n318410 , n318409 );
or ( n318411 , n318401 , n318410 );
nand ( n27986 , n27974 , n318411 );
buf ( n318413 , n27986 );
buf ( n318414 , n318413 );
xor ( n27989 , n318397 , n318414 );
buf ( n318416 , n27989 );
xor ( n318417 , n318347 , n318416 );
buf ( n318418 , n14523 );
not ( n318419 , n318418 );
buf ( n318420 , n304941 );
not ( n318421 , n318420 );
or ( n318422 , n318419 , n318421 );
buf ( n318423 , n878 );
nand ( n318424 , n318422 , n318423 );
buf ( n318425 , n318424 );
buf ( n318426 , n318425 );
buf ( n318427 , n317520 );
not ( n28002 , n318427 );
buf ( n318429 , n304851 );
not ( n318430 , n318429 );
or ( n318431 , n28002 , n318430 );
buf ( n318432 , n836 );
buf ( n318433 , n872 );
xnor ( n318434 , n318432 , n318433 );
buf ( n318435 , n318434 );
buf ( n318436 , n318435 );
not ( n28011 , n318436 );
buf ( n318438 , n304845 );
nand ( n28013 , n28011 , n318438 );
buf ( n318440 , n28013 );
buf ( n318441 , n318440 );
nand ( n318442 , n318431 , n318441 );
buf ( n318443 , n318442 );
buf ( n318444 , n318443 );
xor ( n318445 , n318426 , n318444 );
buf ( n318446 , n305650 );
buf ( n318447 , n317594 );
or ( n318448 , n318446 , n318447 );
buf ( n28023 , n305664 );
buf ( n318450 , n876 );
buf ( n318451 , n20700 );
and ( n318452 , n318450 , n318451 );
not ( n28027 , n318450 );
buf ( n318454 , n832 );
and ( n28029 , n28027 , n318454 );
nor ( n318456 , n318452 , n28029 );
buf ( n318457 , n318456 );
buf ( n318458 , n318457 );
or ( n318459 , n28023 , n318458 );
nand ( n318460 , n318448 , n318459 );
buf ( n318461 , n318460 );
buf ( n318462 , n318461 );
xor ( n318463 , n318445 , n318462 );
buf ( n318464 , n318463 );
xor ( n28039 , n318417 , n318464 );
xor ( n318466 , n317472 , n317488 );
xor ( n318467 , n318466 , n317500 );
and ( n28042 , n317547 , n318467 );
xor ( n318469 , n317472 , n317488 );
xor ( n318470 , n318469 , n317500 );
and ( n28045 , n317601 , n318470 );
and ( n318472 , n317547 , n317601 );
or ( n318473 , n28042 , n28045 , n318472 );
xor ( n318474 , n317425 , n317431 );
and ( n28049 , n318474 , n317453 );
and ( n318476 , n317425 , n317431 );
or ( n28051 , n28049 , n318476 );
buf ( n318478 , n28051 );
xor ( n318479 , n318473 , n318478 );
xor ( n318480 , n28039 , n318479 );
buf ( n318481 , n318480 );
xor ( n28056 , n318296 , n318302 );
xor ( n318483 , n28056 , n318481 );
buf ( n318484 , n318483 );
xor ( n28059 , n318296 , n318302 );
and ( n318486 , n28059 , n318481 );
and ( n318487 , n318296 , n318302 );
or ( n28062 , n318486 , n318487 );
buf ( n318489 , n28062 );
buf ( n318490 , n305289 );
not ( n318491 , n318490 );
buf ( n28066 , n305192 );
nor ( n28067 , n318491 , n28066 );
buf ( n28068 , n28067 );
buf ( n318495 , n28068 );
buf ( n318496 , n894 );
buf ( n318497 , n844 );
xor ( n28072 , n318496 , n318497 );
buf ( n318499 , n28072 );
buf ( n318500 , n318499 );
not ( n318501 , n318500 );
buf ( n318502 , n305881 );
not ( n28077 , n318502 );
buf ( n28078 , n28077 );
buf ( n318505 , n28078 );
not ( n28080 , n318505 );
or ( n318507 , n318501 , n28080 );
buf ( n318508 , n315411 );
buf ( n318509 , n895 );
nand ( n318510 , n318508 , n318509 );
buf ( n318511 , n318510 );
buf ( n318512 , n318511 );
nand ( n28087 , n318507 , n318512 );
buf ( n318514 , n28087 );
buf ( n318515 , n318514 );
xor ( n318516 , n318495 , n318515 );
buf ( n318517 , n888 );
buf ( n318518 , n850 );
and ( n318519 , n318517 , n318518 );
not ( n318520 , n318517 );
buf ( n318521 , n304565 );
and ( n28096 , n318520 , n318521 );
nor ( n318523 , n318519 , n28096 );
buf ( n318524 , n318523 );
buf ( n318525 , n318524 );
not ( n318526 , n318525 );
buf ( n318527 , n305138 );
not ( n28102 , n318527 );
or ( n318529 , n318526 , n28102 );
buf ( n318530 , n305144 );
buf ( n318531 , n315495 );
nand ( n318532 , n318530 , n318531 );
buf ( n318533 , n318532 );
buf ( n318534 , n318533 );
nand ( n318535 , n318529 , n318534 );
buf ( n318536 , n318535 );
buf ( n318537 , n318536 );
and ( n28112 , n318516 , n318537 );
and ( n28113 , n318495 , n318515 );
or ( n318540 , n28112 , n28113 );
buf ( n318541 , n318540 );
buf ( n318542 , n318541 );
buf ( n318543 , n862 );
buf ( n318544 , n876 );
xor ( n318545 , n318543 , n318544 );
buf ( n318546 , n318545 );
buf ( n318547 , n318546 );
not ( n318548 , n318547 );
buf ( n318549 , n305338 );
not ( n318550 , n318549 );
or ( n318551 , n318548 , n318550 );
buf ( n318552 , n305344 );
buf ( n318553 , n315347 );
nand ( n28128 , n318552 , n318553 );
buf ( n318555 , n28128 );
buf ( n318556 , n318555 );
nand ( n28131 , n318551 , n318556 );
buf ( n318558 , n28131 );
buf ( n28133 , n318558 );
buf ( n318560 , n848 );
buf ( n318561 , n890 );
xor ( n318562 , n318560 , n318561 );
buf ( n318563 , n318562 );
buf ( n318564 , n318563 );
not ( n318565 , n318564 );
buf ( n318566 , n304633 );
not ( n28141 , n318566 );
or ( n318568 , n318565 , n28141 );
buf ( n28143 , n304658 );
buf ( n318570 , n25029 );
nand ( n318571 , n28143 , n318570 );
buf ( n318572 , n318571 );
buf ( n318573 , n318572 );
nand ( n28148 , n318568 , n318573 );
buf ( n318575 , n28148 );
buf ( n318576 , n318575 );
xor ( n28151 , n28133 , n318576 );
buf ( n318578 , n314747 );
buf ( n318579 , n852 );
buf ( n318580 , n886 );
xnor ( n318581 , n318579 , n318580 );
buf ( n318582 , n318581 );
buf ( n318583 , n318582 );
or ( n318584 , n318578 , n318583 );
buf ( n318585 , n305363 );
buf ( n318586 , n315392 );
or ( n318587 , n318585 , n318586 );
nand ( n28162 , n318584 , n318587 );
buf ( n318589 , n28162 );
buf ( n318590 , n318589 );
and ( n318591 , n28151 , n318590 );
and ( n318592 , n28133 , n318576 );
or ( n28167 , n318591 , n318592 );
buf ( n318594 , n28167 );
buf ( n318595 , n318594 );
xor ( n28170 , n318542 , n318595 );
xor ( n318597 , n315425 , n315446 );
xor ( n318598 , n318597 , n315469 );
buf ( n318599 , n318598 );
buf ( n318600 , n318599 );
and ( n318601 , n28170 , n318600 );
and ( n28176 , n318542 , n318595 );
or ( n28177 , n318601 , n28176 );
buf ( n318604 , n28177 );
buf ( n318605 , n318604 );
xor ( n318606 , n315343 , n24979 );
xor ( n318607 , n318606 , n315474 );
buf ( n318608 , n318607 );
buf ( n318609 , n318608 );
xor ( n318610 , n318605 , n318609 );
buf ( n318611 , n882 );
buf ( n318612 , n856 );
and ( n318613 , n318611 , n318612 );
not ( n28188 , n318611 );
buf ( n318615 , n15582 );
and ( n28190 , n28188 , n318615 );
nor ( n28191 , n318613 , n28190 );
buf ( n318618 , n28191 );
buf ( n318619 , n318618 );
not ( n28194 , n318619 );
buf ( n318621 , n304584 );
not ( n28196 , n318621 );
or ( n28197 , n28194 , n28196 );
buf ( n318624 , n315593 );
not ( n318625 , n318624 );
buf ( n318626 , n304596 );
nand ( n28201 , n318625 , n318626 );
buf ( n318628 , n28201 );
buf ( n318629 , n318628 );
nand ( n318630 , n28197 , n318629 );
buf ( n318631 , n318630 );
buf ( n318632 , n318631 );
buf ( n318633 , n884 );
buf ( n318634 , n854 );
xor ( n28209 , n318633 , n318634 );
buf ( n318636 , n28209 );
buf ( n318637 , n318636 );
not ( n28212 , n318637 );
buf ( n318639 , n304813 );
not ( n318640 , n318639 );
or ( n28215 , n28212 , n318640 );
buf ( n318642 , n304807 );
buf ( n318643 , n315433 );
nand ( n28218 , n318642 , n318643 );
buf ( n28219 , n28218 );
buf ( n318646 , n28219 );
nand ( n318647 , n28215 , n318646 );
buf ( n318648 , n318647 );
buf ( n318649 , n318648 );
xor ( n28224 , n318632 , n318649 );
buf ( n318651 , n863 );
buf ( n318652 , n877 );
or ( n318653 , n318651 , n318652 );
buf ( n318654 , n878 );
nand ( n318655 , n318653 , n318654 );
buf ( n318656 , n318655 );
buf ( n318657 , n318656 );
buf ( n318658 , n863 );
buf ( n318659 , n877 );
nand ( n28234 , n318658 , n318659 );
buf ( n318661 , n28234 );
buf ( n318662 , n318661 );
buf ( n318663 , n876 );
and ( n318664 , n318657 , n318662 , n318663 );
buf ( n318665 , n318664 );
buf ( n318666 , n318665 );
xor ( n318667 , n894 , n845 );
buf ( n28242 , n318667 );
not ( n28243 , n28242 );
buf ( n28244 , n28078 );
not ( n28245 , n28244 );
or ( n28246 , n28243 , n28245 );
buf ( n28247 , n318499 );
buf ( n28248 , n895 );
nand ( n28249 , n28247 , n28248 );
buf ( n28250 , n28249 );
buf ( n28251 , n28250 );
nand ( n28252 , n28246 , n28251 );
buf ( n28253 , n28252 );
buf ( n318680 , n28253 );
and ( n28255 , n318666 , n318680 );
buf ( n318682 , n28255 );
buf ( n318683 , n318682 );
and ( n318684 , n28224 , n318683 );
and ( n28259 , n318632 , n318649 );
or ( n318686 , n318684 , n28259 );
buf ( n318687 , n318686 );
buf ( n318688 , n318687 );
xor ( n28263 , n315361 , n315382 );
xor ( n318690 , n28263 , n315400 );
buf ( n318691 , n318690 );
buf ( n318692 , n318691 );
xor ( n318693 , n318688 , n318692 );
xor ( n28268 , n315508 , n315525 );
xor ( n28269 , n28268 , n315546 );
buf ( n318696 , n28269 );
buf ( n318697 , n318696 );
and ( n318698 , n318693 , n318697 );
and ( n28273 , n318688 , n318692 );
or ( n28274 , n318698 , n28273 );
buf ( n318701 , n28274 );
buf ( n318702 , n318701 );
and ( n318703 , n318610 , n318702 );
and ( n28278 , n318605 , n318609 );
or ( n318705 , n318703 , n28278 );
buf ( n318706 , n318705 );
buf ( n318707 , n318706 );
xor ( n28282 , n315583 , n315587 );
xor ( n28283 , n28282 , n315666 );
buf ( n318710 , n28283 );
buf ( n318711 , n318710 );
xor ( n28286 , n315551 , n315555 );
xor ( n318713 , n28286 , n315560 );
buf ( n318714 , n318713 );
buf ( n318715 , n318714 );
xor ( n28290 , n318711 , n318715 );
xor ( n318717 , n25178 , n315607 );
xor ( n28292 , n318717 , n315661 );
buf ( n318719 , n28292 );
buf ( n318720 , n318719 );
xor ( n318721 , n318542 , n318595 );
xor ( n318722 , n318721 , n318600 );
buf ( n318723 , n318722 );
buf ( n318724 , n318723 );
xor ( n318725 , n318720 , n318724 );
buf ( n318726 , n892 );
buf ( n318727 , n847 );
and ( n318728 , n318726 , n318727 );
not ( n318729 , n318726 );
buf ( n318730 , n315972 );
and ( n28305 , n318729 , n318730 );
nor ( n318732 , n318728 , n28305 );
buf ( n318733 , n318732 );
buf ( n318734 , n318733 );
not ( n318735 , n318734 );
buf ( n318736 , n14272 );
not ( n28311 , n318736 );
or ( n318738 , n318735 , n28311 );
buf ( n28313 , n315609 );
buf ( n318740 , n304694 );
nand ( n318741 , n28313 , n318740 );
buf ( n318742 , n318741 );
buf ( n318743 , n318742 );
nand ( n28318 , n318738 , n318743 );
buf ( n318745 , n28318 );
buf ( n318746 , n318745 );
not ( n28321 , n318746 );
buf ( n318748 , n314747 );
buf ( n318749 , n853 );
buf ( n318750 , n886 );
xnor ( n28325 , n318749 , n318750 );
buf ( n318752 , n28325 );
buf ( n318753 , n318752 );
or ( n28328 , n318748 , n318753 );
buf ( n318755 , n305363 );
buf ( n318756 , n318582 );
or ( n28331 , n318755 , n318756 );
nand ( n318758 , n28328 , n28331 );
buf ( n318759 , n318758 );
buf ( n318760 , n318759 );
not ( n318761 , n318760 );
or ( n28336 , n28321 , n318761 );
buf ( n318763 , n318759 );
buf ( n318764 , n318745 );
or ( n318765 , n318763 , n318764 );
buf ( n318766 , n876 );
buf ( n318767 , n863 );
and ( n318768 , n318766 , n318767 );
not ( n28343 , n318766 );
buf ( n318770 , n305192 );
and ( n318771 , n28343 , n318770 );
nor ( n28346 , n318768 , n318771 );
buf ( n318773 , n28346 );
buf ( n318774 , n318773 );
not ( n318775 , n318774 );
buf ( n318776 , n305338 );
not ( n28351 , n318776 );
or ( n318778 , n318775 , n28351 );
buf ( n318779 , n305344 );
buf ( n318780 , n318546 );
nand ( n318781 , n318779 , n318780 );
buf ( n318782 , n318781 );
buf ( n318783 , n318782 );
nand ( n28358 , n318778 , n318783 );
buf ( n28359 , n28358 );
buf ( n28360 , n28359 );
nand ( n28361 , n318765 , n28360 );
buf ( n28362 , n28361 );
buf ( n318789 , n28362 );
nand ( n28364 , n28336 , n318789 );
buf ( n28365 , n28364 );
xor ( n318792 , n880 , n859 );
buf ( n318793 , n318792 );
not ( n318794 , n318793 );
buf ( n318795 , n304984 );
not ( n28370 , n318795 );
or ( n318797 , n318794 , n28370 );
buf ( n318798 , n315648 );
not ( n318799 , n318798 );
buf ( n318800 , n304973 );
nand ( n318801 , n318799 , n318800 );
buf ( n318802 , n318801 );
buf ( n318803 , n318802 );
nand ( n318804 , n318797 , n318803 );
buf ( n318805 , n318804 );
buf ( n318806 , n318805 );
buf ( n318807 , n851 );
buf ( n318808 , n888 );
xnor ( n318809 , n318807 , n318808 );
buf ( n318810 , n318809 );
buf ( n318811 , n318810 );
not ( n28386 , n318811 );
buf ( n318813 , n28386 );
buf ( n318814 , n318813 );
not ( n318815 , n318814 );
buf ( n318816 , n305138 );
not ( n28391 , n318816 );
or ( n318818 , n318815 , n28391 );
buf ( n318819 , n305144 );
buf ( n318820 , n318524 );
nand ( n318821 , n318819 , n318820 );
buf ( n318822 , n318821 );
buf ( n318823 , n318822 );
nand ( n318824 , n318818 , n318823 );
buf ( n318825 , n318824 );
buf ( n318826 , n318825 );
xor ( n28401 , n318806 , n318826 );
buf ( n318828 , n878 );
buf ( n28403 , n861 );
xor ( n28404 , n318828 , n28403 );
buf ( n318831 , n28404 );
buf ( n318832 , n318831 );
not ( n318833 , n318832 );
buf ( n318834 , n318833 );
buf ( n318835 , n318834 );
buf ( n318836 , n304938 );
or ( n318837 , n318835 , n318836 );
buf ( n318838 , n14523 );
buf ( n318839 , n315626 );
or ( n28414 , n318838 , n318839 );
nand ( n318841 , n318837 , n28414 );
buf ( n318842 , n318841 );
buf ( n318843 , n318842 );
and ( n318844 , n28401 , n318843 );
and ( n318845 , n318806 , n318826 );
or ( n318846 , n318844 , n318845 );
buf ( n318847 , n318846 );
xor ( n318848 , n28365 , n318847 );
buf ( n318849 , n855 );
buf ( n318850 , n884 );
xor ( n318851 , n318849 , n318850 );
buf ( n318852 , n318851 );
buf ( n318853 , n318852 );
not ( n28428 , n318853 );
buf ( n318855 , n310401 );
not ( n318856 , n318855 );
or ( n28431 , n28428 , n318856 );
buf ( n318858 , n304819 );
buf ( n318859 , n318636 );
nand ( n28434 , n318858 , n318859 );
buf ( n28435 , n28434 );
buf ( n318862 , n28435 );
nand ( n318863 , n28431 , n318862 );
buf ( n318864 , n318863 );
buf ( n318865 , n318864 );
buf ( n318866 , n890 );
buf ( n318867 , n849 );
and ( n318868 , n318866 , n318867 );
not ( n318869 , n318866 );
buf ( n28444 , n305596 );
and ( n318871 , n318869 , n28444 );
nor ( n28446 , n318868 , n318871 );
buf ( n28447 , n28446 );
buf ( n318874 , n28447 );
not ( n318875 , n318874 );
buf ( n318876 , n304633 );
not ( n318877 , n318876 );
or ( n318878 , n318875 , n318877 );
buf ( n318879 , n304658 );
buf ( n318880 , n318563 );
nand ( n318881 , n318879 , n318880 );
buf ( n318882 , n318881 );
buf ( n318883 , n318882 );
nand ( n318884 , n318878 , n318883 );
buf ( n318885 , n318884 );
buf ( n28460 , n318885 );
xor ( n28461 , n318865 , n28460 );
buf ( n318888 , n857 );
buf ( n28463 , n882 );
xor ( n28464 , n318888 , n28463 );
buf ( n28465 , n28464 );
buf ( n318892 , n28465 );
not ( n28467 , n318892 );
buf ( n318894 , n304584 );
not ( n318895 , n318894 );
or ( n28470 , n28467 , n318895 );
buf ( n318897 , n304596 );
buf ( n28472 , n318618 );
nand ( n28473 , n318897 , n28472 );
buf ( n318900 , n28473 );
buf ( n318901 , n318900 );
nand ( n28476 , n28470 , n318901 );
buf ( n318903 , n28476 );
buf ( n318904 , n318903 );
and ( n28479 , n28461 , n318904 );
and ( n28480 , n318865 , n28460 );
or ( n28481 , n28479 , n28480 );
buf ( n318908 , n28481 );
and ( n28483 , n318848 , n318908 );
and ( n318910 , n28365 , n318847 );
or ( n318911 , n28483 , n318910 );
buf ( n318912 , n318911 );
and ( n28487 , n318725 , n318912 );
and ( n28488 , n318720 , n318724 );
or ( n28489 , n28487 , n28488 );
buf ( n318916 , n28489 );
buf ( n318917 , n318916 );
and ( n318918 , n28290 , n318917 );
and ( n28493 , n318711 , n318715 );
or ( n28494 , n318918 , n28493 );
buf ( n318921 , n28494 );
buf ( n318922 , n318921 );
xor ( n318923 , n315302 , n315305 );
xor ( n318924 , n318923 , n315478 );
xor ( n28499 , n315670 , n315676 );
xor ( n318926 , n318924 , n28499 );
buf ( n318927 , n318926 );
xor ( n318928 , n318707 , n318922 );
xor ( n28503 , n318928 , n318927 );
buf ( n318930 , n28503 );
xor ( n318931 , n318707 , n318922 );
and ( n318932 , n318931 , n318927 );
and ( n28507 , n318707 , n318922 );
or ( n318934 , n318932 , n28507 );
buf ( n318935 , n318934 );
xor ( n318936 , n318605 , n318609 );
xor ( n28511 , n318936 , n318702 );
buf ( n318938 , n28511 );
buf ( n318939 , n318938 );
xor ( n28514 , n318711 , n318715 );
xor ( n318941 , n28514 , n318917 );
buf ( n318942 , n318941 );
buf ( n318943 , n318942 );
xor ( n28518 , n318688 , n318692 );
xor ( n318945 , n28518 , n318697 );
buf ( n318946 , n318945 );
buf ( n318947 , n318946 );
xor ( n318948 , n28133 , n318576 );
xor ( n318949 , n318948 , n318590 );
buf ( n318950 , n318949 );
buf ( n318951 , n318950 );
xor ( n318952 , n318495 , n318515 );
xor ( n318953 , n318952 , n318537 );
buf ( n318954 , n318953 );
buf ( n318955 , n318954 );
xor ( n318956 , n318951 , n318955 );
xor ( n28531 , n25196 , n315642 );
xor ( n318958 , n28531 , n315656 );
buf ( n318959 , n318958 );
buf ( n318960 , n318959 );
and ( n318961 , n318956 , n318960 );
and ( n28536 , n318951 , n318955 );
or ( n318963 , n318961 , n28536 );
buf ( n318964 , n318963 );
buf ( n318965 , n318964 );
xor ( n318966 , n318947 , n318965 );
xor ( n318967 , n318720 , n318724 );
xor ( n318968 , n318967 , n318912 );
buf ( n318969 , n318968 );
buf ( n318970 , n318969 );
and ( n318971 , n318966 , n318970 );
and ( n28546 , n318947 , n318965 );
or ( n318973 , n318971 , n28546 );
buf ( n318974 , n318973 );
buf ( n318975 , n318974 );
xor ( n318976 , n318939 , n318943 );
xor ( n318977 , n318976 , n318975 );
buf ( n318978 , n318977 );
xor ( n318979 , n318939 , n318943 );
and ( n318980 , n318979 , n318975 );
and ( n28555 , n318939 , n318943 );
or ( n318982 , n318980 , n28555 );
buf ( n318983 , n318982 );
xor ( n28558 , n318666 , n318680 );
buf ( n28559 , n28558 );
buf ( n318986 , n28559 );
buf ( n318987 , n305344 );
buf ( n318988 , n863 );
and ( n318989 , n318987 , n318988 );
buf ( n318990 , n318989 );
buf ( n318991 , n318990 );
buf ( n318992 , n894 );
buf ( n318993 , n846 );
xor ( n28568 , n318992 , n318993 );
buf ( n318995 , n28568 );
buf ( n318996 , n318995 );
not ( n28571 , n318996 );
buf ( n318998 , n28078 );
not ( n28573 , n318998 );
or ( n319000 , n28571 , n28573 );
buf ( n28575 , n318667 );
buf ( n319002 , n895 );
nand ( n319003 , n28575 , n319002 );
buf ( n319004 , n319003 );
buf ( n319005 , n319004 );
nand ( n319006 , n319000 , n319005 );
buf ( n319007 , n319006 );
buf ( n319008 , n319007 );
xor ( n319009 , n318991 , n319008 );
buf ( n319010 , n306283 );
xnor ( n319011 , n888 , n852 );
buf ( n319012 , n319011 );
or ( n319013 , n319010 , n319012 );
buf ( n319014 , n15861 );
buf ( n319015 , n318810 );
or ( n319016 , n319014 , n319015 );
nand ( n319017 , n319013 , n319016 );
buf ( n319018 , n319017 );
buf ( n319019 , n319018 );
and ( n319020 , n319009 , n319019 );
and ( n28595 , n318991 , n319008 );
or ( n319022 , n319020 , n28595 );
buf ( n319023 , n319022 );
buf ( n319024 , n319023 );
xor ( n319025 , n318986 , n319024 );
buf ( n319026 , n880 );
buf ( n319027 , n860 );
xor ( n28602 , n319026 , n319027 );
buf ( n319029 , n28602 );
buf ( n319030 , n319029 );
not ( n319031 , n319030 );
buf ( n319032 , n305098 );
not ( n28607 , n319032 );
or ( n319034 , n319031 , n28607 );
buf ( n319035 , n304997 );
buf ( n319036 , n318792 );
nand ( n319037 , n319035 , n319036 );
buf ( n319038 , n319037 );
buf ( n319039 , n319038 );
nand ( n319040 , n319034 , n319039 );
buf ( n319041 , n319040 );
buf ( n319042 , n319041 );
not ( n28617 , n319042 );
not ( n319044 , n306272 );
not ( n319045 , n318831 );
or ( n28620 , n319044 , n319045 );
and ( n319047 , n862 , n878 );
not ( n28622 , n862 );
and ( n319049 , n28622 , n310371 );
nor ( n28624 , n319047 , n319049 );
not ( n28625 , n28624 );
or ( n319052 , n304941 , n28625 );
nand ( n28627 , n28620 , n319052 );
buf ( n319054 , n28627 );
not ( n28629 , n319054 );
or ( n319056 , n28617 , n28629 );
buf ( n319057 , n28627 );
buf ( n319058 , n319041 );
or ( n319059 , n319057 , n319058 );
buf ( n319060 , n892 );
buf ( n319061 , n848 );
and ( n319062 , n319060 , n319061 );
not ( n28637 , n319060 );
buf ( n319064 , n304786 );
and ( n28639 , n28637 , n319064 );
nor ( n28640 , n319062 , n28639 );
buf ( n319067 , n28640 );
buf ( n319068 , n319067 );
not ( n28643 , n319068 );
buf ( n319070 , n14272 );
not ( n319071 , n319070 );
or ( n28646 , n28643 , n319071 );
buf ( n319073 , n305430 );
buf ( n319074 , n318733 );
nand ( n28649 , n319073 , n319074 );
buf ( n319076 , n28649 );
buf ( n319077 , n319076 );
nand ( n319078 , n28646 , n319077 );
buf ( n319079 , n319078 );
buf ( n319080 , n319079 );
nand ( n319081 , n319059 , n319080 );
buf ( n319082 , n319081 );
buf ( n319083 , n319082 );
nand ( n319084 , n319056 , n319083 );
buf ( n319085 , n319084 );
buf ( n319086 , n319085 );
and ( n28661 , n319025 , n319086 );
and ( n28662 , n318986 , n319024 );
or ( n319089 , n28661 , n28662 );
buf ( n319090 , n319089 );
buf ( n319091 , n319090 );
xor ( n319092 , n318632 , n318649 );
xor ( n319093 , n319092 , n318683 );
buf ( n319094 , n319093 );
buf ( n319095 , n319094 );
xor ( n319096 , n319091 , n319095 );
buf ( n319097 , n856 );
buf ( n319098 , n884 );
xor ( n319099 , n319097 , n319098 );
buf ( n319100 , n319099 );
buf ( n319101 , n319100 );
not ( n319102 , n319101 );
buf ( n319103 , n304813 );
not ( n28678 , n319103 );
or ( n319105 , n319102 , n28678 );
buf ( n319106 , n304819 );
buf ( n319107 , n318852 );
nand ( n319108 , n319106 , n319107 );
buf ( n319109 , n319108 );
buf ( n319110 , n319109 );
nand ( n319111 , n319105 , n319110 );
buf ( n319112 , n319111 );
buf ( n319113 , n319112 );
buf ( n319114 , n854 );
buf ( n319115 , n886 );
xor ( n319116 , n319114 , n319115 );
buf ( n319117 , n319116 );
buf ( n319118 , n319117 );
not ( n319119 , n319118 );
buf ( n319120 , n304912 );
not ( n319121 , n319120 );
or ( n319122 , n319119 , n319121 );
buf ( n319123 , n318752 );
not ( n28698 , n319123 );
buf ( n319125 , n304901 );
nand ( n319126 , n28698 , n319125 );
buf ( n319127 , n319126 );
buf ( n319128 , n319127 );
nand ( n28703 , n319122 , n319128 );
buf ( n319130 , n28703 );
buf ( n319131 , n319130 );
or ( n319132 , n319113 , n319131 );
buf ( n319133 , n890 );
buf ( n319134 , n850 );
and ( n28709 , n319133 , n319134 );
not ( n28710 , n319133 );
buf ( n28711 , n304565 );
and ( n319138 , n28710 , n28711 );
nor ( n28713 , n28709 , n319138 );
buf ( n28714 , n28713 );
buf ( n319141 , n28714 );
not ( n28716 , n319141 );
buf ( n319143 , n304633 );
not ( n319144 , n319143 );
or ( n28719 , n28716 , n319144 );
buf ( n319146 , n304658 );
buf ( n319147 , n28447 );
nand ( n28722 , n319146 , n319147 );
buf ( n319149 , n28722 );
buf ( n319150 , n319149 );
nand ( n319151 , n28719 , n319150 );
buf ( n319152 , n319151 );
buf ( n319153 , n319152 );
nand ( n319154 , n319132 , n319153 );
buf ( n319155 , n319154 );
buf ( n319156 , n319155 );
buf ( n319157 , n319112 );
buf ( n319158 , n319130 );
nand ( n28733 , n319157 , n319158 );
buf ( n28734 , n28733 );
buf ( n319161 , n28734 );
nand ( n28736 , n319156 , n319161 );
buf ( n28737 , n28736 );
buf ( n28738 , n28737 );
xor ( n319165 , n318865 , n28460 );
xor ( n319166 , n319165 , n318904 );
buf ( n319167 , n319166 );
buf ( n319168 , n319167 );
xor ( n319169 , n28738 , n319168 );
xor ( n28744 , n318806 , n318826 );
xor ( n319171 , n28744 , n318843 );
buf ( n319172 , n319171 );
buf ( n319173 , n319172 );
and ( n28748 , n319169 , n319173 );
and ( n319175 , n28738 , n319168 );
or ( n319176 , n28748 , n319175 );
buf ( n319177 , n319176 );
buf ( n319178 , n319177 );
and ( n319179 , n319096 , n319178 );
and ( n28754 , n319091 , n319095 );
or ( n319181 , n319179 , n28754 );
buf ( n319182 , n319181 );
buf ( n319183 , n319182 );
xor ( n319184 , n318951 , n318955 );
xor ( n28759 , n319184 , n318960 );
buf ( n319186 , n28759 );
xor ( n319187 , n28365 , n318847 );
xor ( n319188 , n319187 , n318908 );
and ( n28763 , n319186 , n319188 );
xor ( n28764 , n319091 , n319095 );
xor ( n319191 , n28764 , n319178 );
buf ( n319192 , n319191 );
xor ( n28767 , n28365 , n318847 );
xor ( n28768 , n28767 , n318908 );
and ( n28769 , n319192 , n28768 );
and ( n319196 , n319186 , n319192 );
or ( n319197 , n28763 , n28769 , n319196 );
buf ( n319198 , n319197 );
xor ( n319199 , n318947 , n318965 );
xor ( n319200 , n319199 , n318970 );
buf ( n319201 , n319200 );
buf ( n319202 , n319201 );
xor ( n319203 , n319183 , n319198 );
xor ( n28778 , n319203 , n319202 );
buf ( n319205 , n28778 );
xor ( n28780 , n319183 , n319198 );
and ( n319207 , n28780 , n319202 );
and ( n319208 , n319183 , n319198 );
or ( n319209 , n319207 , n319208 );
buf ( n319210 , n319209 );
buf ( n319211 , n305381 );
buf ( n319212 , n858 );
buf ( n319213 , n882 );
xnor ( n319214 , n319212 , n319213 );
buf ( n319215 , n319214 );
buf ( n319216 , n319215 );
or ( n319217 , n319211 , n319216 );
buf ( n28792 , n14959 );
buf ( n319219 , n28465 );
not ( n319220 , n319219 );
buf ( n319221 , n319220 );
buf ( n319222 , n319221 );
or ( n28797 , n28792 , n319222 );
nand ( n319224 , n319217 , n28797 );
buf ( n319225 , n319224 );
buf ( n319226 , n319225 );
buf ( n319227 , n863 );
buf ( n319228 , n879 );
or ( n319229 , n319227 , n319228 );
buf ( n319230 , n880 );
nand ( n28805 , n319229 , n319230 );
buf ( n28806 , n28805 );
buf ( n319233 , n28806 );
buf ( n319234 , n863 );
buf ( n319235 , n879 );
nand ( n319236 , n319234 , n319235 );
buf ( n319237 , n319236 );
buf ( n319238 , n319237 );
buf ( n319239 , n878 );
and ( n28814 , n319233 , n319238 , n319239 );
buf ( n319241 , n28814 );
buf ( n28816 , n895 );
not ( n28817 , n28816 );
buf ( n28818 , n318995 );
not ( n28819 , n28818 );
or ( n28820 , n28817 , n28819 );
buf ( n319247 , n305881 );
buf ( n319248 , n894 );
buf ( n319249 , n847 );
xnor ( n319250 , n319248 , n319249 );
buf ( n319251 , n319250 );
buf ( n319252 , n319251 );
or ( n319253 , n319247 , n319252 );
nand ( n319254 , n28820 , n319253 );
buf ( n319255 , n319254 );
and ( n319256 , n319241 , n319255 );
buf ( n319257 , n319256 );
xor ( n319258 , n319226 , n319257 );
xor ( n28833 , n880 , n861 );
buf ( n319260 , n28833 );
not ( n28835 , n319260 );
buf ( n319262 , n305098 );
not ( n319263 , n319262 );
or ( n28838 , n28835 , n319263 );
buf ( n319265 , n304973 );
buf ( n28840 , n319029 );
nand ( n28841 , n319265 , n28840 );
buf ( n319268 , n28841 );
buf ( n319269 , n319268 );
nand ( n319270 , n28838 , n319269 );
buf ( n319271 , n319270 );
buf ( n319272 , n319271 );
buf ( n319273 , n878 );
buf ( n319274 , n863 );
and ( n28849 , n319273 , n319274 );
not ( n28850 , n319273 );
buf ( n319277 , n305192 );
and ( n319278 , n28850 , n319277 );
nor ( n28853 , n28849 , n319278 );
buf ( n319280 , n28853 );
buf ( n319281 , n319280 );
not ( n319282 , n319281 );
buf ( n319283 , n313029 );
not ( n28858 , n319283 );
or ( n28859 , n319282 , n28858 );
buf ( n319286 , n306272 );
buf ( n319287 , n28624 );
nand ( n28862 , n319286 , n319287 );
buf ( n319289 , n28862 );
buf ( n319290 , n319289 );
nand ( n319291 , n28859 , n319290 );
buf ( n319292 , n319291 );
buf ( n319293 , n319292 );
xor ( n28868 , n319272 , n319293 );
buf ( n319295 , n305135 );
buf ( n319296 , n888 );
buf ( n319297 , n304956 );
and ( n319298 , n319296 , n319297 );
not ( n28873 , n319296 );
buf ( n319300 , n853 );
and ( n319301 , n28873 , n319300 );
nor ( n28876 , n319298 , n319301 );
buf ( n319303 , n28876 );
buf ( n319304 , n319303 );
or ( n319305 , n319295 , n319304 );
buf ( n319306 , n15861 );
buf ( n319307 , n319011 );
or ( n319308 , n319306 , n319307 );
nand ( n319309 , n319305 , n319308 );
buf ( n319310 , n319309 );
buf ( n319311 , n319310 );
and ( n319312 , n28868 , n319311 );
and ( n319313 , n319272 , n319293 );
or ( n28888 , n319312 , n319313 );
buf ( n319315 , n28888 );
buf ( n319316 , n319315 );
and ( n28891 , n319258 , n319316 );
and ( n319318 , n319226 , n319257 );
or ( n319319 , n28891 , n319318 );
buf ( n319320 , n319319 );
buf ( n319321 , n319320 );
buf ( n319322 , n318759 );
not ( n319323 , n319322 );
buf ( n319324 , n28359 );
buf ( n319325 , n318745 );
xnor ( n28900 , n319324 , n319325 );
buf ( n319327 , n28900 );
buf ( n319328 , n319327 );
not ( n319329 , n319328 );
or ( n319330 , n319323 , n319329 );
buf ( n319331 , n319327 );
buf ( n319332 , n318759 );
or ( n28907 , n319331 , n319332 );
nand ( n28908 , n319330 , n28907 );
buf ( n319335 , n28908 );
buf ( n319336 , n319335 );
xor ( n28911 , n319321 , n319336 );
xor ( n28912 , n318986 , n319024 );
xor ( n28913 , n28912 , n319086 );
buf ( n319340 , n28913 );
buf ( n319341 , n319340 );
and ( n28916 , n28911 , n319341 );
and ( n319343 , n319321 , n319336 );
or ( n28918 , n28916 , n319343 );
buf ( n319345 , n28918 );
buf ( n319346 , n319345 );
xor ( n28921 , n318991 , n319008 );
xor ( n319348 , n28921 , n319019 );
buf ( n319349 , n319348 );
buf ( n319350 , n319349 );
buf ( n319351 , n849 );
buf ( n319352 , n892 );
xnor ( n319353 , n319351 , n319352 );
buf ( n319354 , n319353 );
buf ( n319355 , n319354 );
not ( n319356 , n319355 );
buf ( n319357 , n319356 );
buf ( n319358 , n319357 );
not ( n28933 , n319358 );
buf ( n319360 , n14272 );
not ( n28935 , n319360 );
or ( n28936 , n28933 , n28935 );
buf ( n319363 , n305430 );
buf ( n28938 , n319067 );
nand ( n28939 , n319363 , n28938 );
buf ( n319366 , n28939 );
buf ( n319367 , n319366 );
nand ( n28942 , n28936 , n319367 );
buf ( n319369 , n28942 );
buf ( n319370 , n319369 );
buf ( n319371 , n890 );
buf ( n319372 , n305532 );
and ( n319373 , n319371 , n319372 );
not ( n28948 , n319371 );
buf ( n319375 , n851 );
and ( n28950 , n28948 , n319375 );
nor ( n319377 , n319373 , n28950 );
buf ( n319378 , n319377 );
buf ( n319379 , n319378 );
not ( n28954 , n319379 );
buf ( n319381 , n28954 );
buf ( n319382 , n319381 );
not ( n28957 , n319382 );
buf ( n319384 , n304633 );
not ( n319385 , n319384 );
or ( n319386 , n28957 , n319385 );
buf ( n319387 , n304658 );
buf ( n319388 , n28714 );
nand ( n319389 , n319387 , n319388 );
buf ( n319390 , n319389 );
buf ( n319391 , n319390 );
nand ( n319392 , n319386 , n319391 );
buf ( n319393 , n319392 );
buf ( n319394 , n319393 );
xor ( n319395 , n319370 , n319394 );
buf ( n319396 , n314747 );
buf ( n319397 , n886 );
buf ( n319398 , n855 );
xnor ( n319399 , n319397 , n319398 );
buf ( n319400 , n319399 );
buf ( n319401 , n319400 );
or ( n28976 , n319396 , n319401 );
buf ( n319403 , n305363 );
buf ( n319404 , n319117 );
not ( n319405 , n319404 );
buf ( n319406 , n319405 );
buf ( n319407 , n319406 );
or ( n28982 , n319403 , n319407 );
nand ( n28983 , n28976 , n28982 );
buf ( n319410 , n28983 );
buf ( n319411 , n319410 );
and ( n28986 , n319395 , n319411 );
and ( n28987 , n319370 , n319394 );
or ( n319414 , n28986 , n28987 );
buf ( n319415 , n319414 );
buf ( n319416 , n319415 );
xor ( n28991 , n319350 , n319416 );
buf ( n319418 , n319130 );
not ( n28993 , n319418 );
xnor ( n28994 , n319152 , n319112 );
buf ( n319421 , n28994 );
not ( n319422 , n319421 );
or ( n28997 , n28993 , n319422 );
buf ( n319424 , n28994 );
buf ( n319425 , n319130 );
or ( n319426 , n319424 , n319425 );
nand ( n29001 , n28997 , n319426 );
buf ( n29002 , n29001 );
buf ( n319429 , n29002 );
and ( n29004 , n28991 , n319429 );
and ( n319431 , n319350 , n319416 );
or ( n29006 , n29004 , n319431 );
buf ( n319433 , n29006 );
buf ( n319434 , n319433 );
xor ( n319435 , n319079 , n319041 );
xor ( n29010 , n319435 , n28627 );
buf ( n319437 , n29010 );
buf ( n319438 , n304581 );
buf ( n319439 , n882 );
buf ( n319440 , n859 );
xnor ( n319441 , n319439 , n319440 );
buf ( n319442 , n319441 );
buf ( n319443 , n319442 );
or ( n319444 , n319438 , n319443 );
buf ( n319445 , n14959 );
buf ( n319446 , n319215 );
or ( n319447 , n319445 , n319446 );
nand ( n319448 , n319444 , n319447 );
buf ( n319449 , n319448 );
buf ( n319450 , n319449 );
buf ( n319451 , n15804 );
buf ( n319452 , n884 );
buf ( n29027 , n305939 );
and ( n29028 , n319452 , n29027 );
not ( n319455 , n319452 );
buf ( n319456 , n857 );
and ( n29031 , n319455 , n319456 );
nor ( n319458 , n29028 , n29031 );
buf ( n319459 , n319458 );
buf ( n319460 , n319459 );
or ( n319461 , n319451 , n319460 );
buf ( n319462 , n310909 );
buf ( n319463 , n319100 );
not ( n29038 , n319463 );
buf ( n29039 , n29038 );
buf ( n319466 , n29039 );
or ( n29041 , n319462 , n319466 );
nand ( n319468 , n319461 , n29041 );
buf ( n319469 , n319468 );
buf ( n319470 , n319469 );
xor ( n319471 , n319450 , n319470 );
xor ( n319472 , n319241 , n319255 );
buf ( n319473 , n319472 );
and ( n319474 , n319471 , n319473 );
and ( n319475 , n319450 , n319470 );
or ( n29050 , n319474 , n319475 );
buf ( n319477 , n29050 );
buf ( n319478 , n319477 );
xor ( n29053 , n319437 , n319478 );
xor ( n319480 , n319226 , n319257 );
xor ( n29055 , n319480 , n319316 );
buf ( n319482 , n29055 );
buf ( n319483 , n319482 );
and ( n319484 , n29053 , n319483 );
and ( n319485 , n319437 , n319478 );
or ( n29060 , n319484 , n319485 );
buf ( n319487 , n29060 );
buf ( n29062 , n319487 );
xor ( n29063 , n319434 , n29062 );
xor ( n319490 , n28738 , n319168 );
xor ( n319491 , n319490 , n319173 );
buf ( n319492 , n319491 );
buf ( n319493 , n319492 );
and ( n319494 , n29063 , n319493 );
and ( n29069 , n319434 , n29062 );
or ( n29070 , n319494 , n29069 );
buf ( n319497 , n29070 );
buf ( n319498 , n319497 );
xor ( n319499 , n28365 , n318847 );
xor ( n29074 , n319499 , n318908 );
xor ( n319501 , n319186 , n319192 );
xor ( n29076 , n29074 , n319501 );
buf ( n319503 , n29076 );
xor ( n29078 , n319346 , n319498 );
xor ( n29079 , n29078 , n319503 );
buf ( n319506 , n29079 );
xor ( n319507 , n319346 , n319498 );
and ( n319508 , n319507 , n319503 );
and ( n29083 , n319346 , n319498 );
or ( n319510 , n319508 , n29083 );
buf ( n319511 , n319510 );
xor ( n29086 , n317062 , n317140 );
xor ( n319513 , n29086 , n317145 );
buf ( n319514 , n319513 );
xor ( n29089 , n317959 , n317965 );
and ( n319516 , n29089 , n317972 );
and ( n319517 , n317959 , n317965 );
or ( n319518 , n319516 , n319517 );
buf ( n319519 , n319518 );
buf ( n29094 , n319519 );
xor ( n29095 , n317982 , n317988 );
and ( n319522 , n29095 , n317993 );
and ( n319523 , n317982 , n317988 );
or ( n29098 , n319522 , n319523 );
buf ( n319525 , n29098 );
buf ( n319526 , n319525 );
xor ( n29101 , n316307 , n316358 );
and ( n319528 , n29101 , n316421 );
and ( n319529 , n316307 , n316358 );
or ( n29104 , n319528 , n319529 );
buf ( n319531 , n29104 );
buf ( n319532 , n319531 );
xor ( n29107 , n316324 , n316338 );
and ( n319534 , n29107 , n316355 );
and ( n319535 , n316324 , n316338 );
or ( n29110 , n319534 , n319535 );
buf ( n319537 , n29110 );
buf ( n319538 , n319537 );
xor ( n29113 , n316438 , n316459 );
and ( n319540 , n29113 , n316477 );
and ( n319541 , n316438 , n316459 );
or ( n319542 , n319540 , n319541 );
buf ( n319543 , n319542 );
buf ( n319544 , n319543 );
xor ( n319545 , n319538 , n319544 );
xor ( n29120 , n316538 , n316559 );
and ( n319547 , n29120 , n26157 );
and ( n319548 , n316538 , n316559 );
or ( n29123 , n319547 , n319548 );
buf ( n319550 , n29123 );
buf ( n29125 , n319550 );
xor ( n29126 , n319545 , n29125 );
buf ( n319553 , n29126 );
buf ( n319554 , n319553 );
xor ( n319555 , n319532 , n319554 );
xor ( n319556 , n316480 , n316523 );
and ( n29131 , n319556 , n316586 );
and ( n319558 , n316480 , n316523 );
or ( n29133 , n29131 , n319558 );
buf ( n319560 , n29133 );
buf ( n319561 , n319560 );
xor ( n319562 , n319555 , n319561 );
buf ( n319563 , n319562 );
buf ( n319564 , n319563 );
xor ( n319565 , n29094 , n319526 );
xor ( n319566 , n319565 , n319564 );
buf ( n319567 , n319566 );
xor ( n29142 , n29094 , n319526 );
and ( n319569 , n29142 , n319564 );
and ( n319570 , n29094 , n319526 );
or ( n319571 , n319569 , n319570 );
buf ( n319572 , n319571 );
buf ( n319573 , n310691 );
buf ( n319574 , n866 );
buf ( n319575 , n841 );
xnor ( n319576 , n319574 , n319575 );
buf ( n319577 , n319576 );
buf ( n319578 , n319577 );
or ( n319579 , n319573 , n319578 );
buf ( n319580 , n310472 );
buf ( n319581 , n840 );
buf ( n319582 , n866 );
xnor ( n29157 , n319581 , n319582 );
buf ( n319584 , n29157 );
buf ( n319585 , n319584 );
or ( n319586 , n319580 , n319585 );
nand ( n29161 , n319579 , n319586 );
buf ( n29162 , n29161 );
buf ( n319589 , n311891 );
buf ( n319590 , n843 );
buf ( n319591 , n864 );
xnor ( n29166 , n319590 , n319591 );
buf ( n319593 , n29166 );
buf ( n319594 , n319593 );
or ( n29169 , n319589 , n319594 );
buf ( n319596 , n311246 );
buf ( n319597 , n311234 );
buf ( n319598 , n842 );
and ( n319599 , n319597 , n319598 );
buf ( n319600 , n304610 );
buf ( n319601 , n864 );
and ( n29176 , n319600 , n319601 );
nor ( n319603 , n319599 , n29176 );
buf ( n319604 , n319603 );
buf ( n319605 , n319604 );
or ( n319606 , n319596 , n319605 );
nand ( n319607 , n29169 , n319606 );
buf ( n319608 , n319607 );
xor ( n319609 , n29162 , n319608 );
buf ( n319610 , n305650 );
buf ( n319611 , n318457 );
or ( n319612 , n319610 , n319611 );
buf ( n319613 , n305664 );
buf ( n319614 , n876 );
not ( n319615 , n319614 );
buf ( n319616 , n319615 );
buf ( n319617 , n319616 );
or ( n319618 , n319613 , n319617 );
nand ( n319619 , n319612 , n319618 );
buf ( n319620 , n319619 );
xor ( n29195 , n319609 , n319620 );
buf ( n319622 , n844 );
buf ( n319623 , n864 );
and ( n29198 , n319622 , n319623 );
buf ( n319625 , n29198 );
buf ( n29200 , n319625 );
buf ( n319627 , n835 );
buf ( n319628 , n872 );
xor ( n319629 , n319627 , n319628 );
buf ( n319630 , n319629 );
buf ( n319631 , n319630 );
not ( n319632 , n319631 );
buf ( n319633 , n304851 );
not ( n29208 , n319633 );
or ( n319635 , n319632 , n29208 );
buf ( n319636 , n872 );
buf ( n319637 , n834 );
xnor ( n319638 , n319636 , n319637 );
buf ( n319639 , n319638 );
buf ( n319640 , n319639 );
not ( n29215 , n319640 );
buf ( n319642 , n304864 );
nand ( n319643 , n29215 , n319642 );
buf ( n319644 , n319643 );
buf ( n319645 , n319644 );
nand ( n29220 , n319635 , n319645 );
buf ( n29221 , n29220 );
buf ( n29222 , n29221 );
xor ( n29223 , n29200 , n29222 );
buf ( n319650 , n305210 );
buf ( n319651 , n310521 );
buf ( n319652 , n839 );
and ( n319653 , n319651 , n319652 );
buf ( n319654 , n14992 );
buf ( n319655 , n868 );
and ( n319656 , n319654 , n319655 );
nor ( n319657 , n319653 , n319656 );
buf ( n319658 , n319657 );
buf ( n319659 , n319658 );
or ( n319660 , n319650 , n319659 );
buf ( n319661 , n305205 );
buf ( n319662 , n310521 );
buf ( n319663 , n838 );
and ( n319664 , n319662 , n319663 );
buf ( n319665 , n310377 );
buf ( n319666 , n868 );
and ( n319667 , n319665 , n319666 );
nor ( n29242 , n319664 , n319667 );
buf ( n29243 , n29242 );
buf ( n319670 , n29243 );
or ( n29245 , n319661 , n319670 );
nand ( n319672 , n319660 , n29245 );
buf ( n319673 , n319672 );
buf ( n319674 , n319673 );
xor ( n319675 , n29223 , n319674 );
buf ( n319676 , n319675 );
buf ( n319677 , n319620 );
not ( n319678 , n319677 );
buf ( n319679 , n319678 );
buf ( n319680 , n319679 );
buf ( n319681 , n311891 );
buf ( n319682 , n318340 );
or ( n29257 , n319681 , n319682 );
buf ( n319684 , n311246 );
buf ( n319685 , n319593 );
or ( n29260 , n319684 , n319685 );
nand ( n319687 , n29257 , n29260 );
buf ( n319688 , n319687 );
buf ( n319689 , n319688 );
xor ( n319690 , n319680 , n319689 );
xor ( n319691 , n318426 , n318444 );
and ( n29266 , n319691 , n318462 );
and ( n319693 , n318426 , n318444 );
or ( n319694 , n29266 , n319693 );
buf ( n319695 , n319694 );
buf ( n319696 , n319695 );
and ( n319697 , n319690 , n319696 );
and ( n29272 , n319680 , n319689 );
or ( n319699 , n319697 , n29272 );
buf ( n319700 , n319699 );
xor ( n319701 , n319676 , n319700 );
xor ( n29276 , n29195 , n319701 );
buf ( n319703 , n29276 );
buf ( n319704 , n318364 );
not ( n319705 , n319704 );
buf ( n319706 , n310694 );
not ( n319707 , n319706 );
or ( n319708 , n319705 , n319707 );
buf ( n319709 , n319577 );
not ( n319710 , n319709 );
buf ( n29285 , n310483 );
nand ( n29286 , n319710 , n29285 );
buf ( n29287 , n29286 );
buf ( n319714 , n29287 );
nand ( n319715 , n319708 , n319714 );
buf ( n319716 , n319715 );
buf ( n319717 , n319716 );
buf ( n319718 , n304854 );
buf ( n319719 , n318435 );
or ( n29294 , n319718 , n319719 );
buf ( n319721 , n14439 );
buf ( n319722 , n319630 );
not ( n29297 , n319722 );
buf ( n319724 , n29297 );
buf ( n319725 , n319724 );
or ( n29300 , n319721 , n319725 );
nand ( n319727 , n29294 , n29300 );
buf ( n319728 , n319727 );
buf ( n319729 , n319728 );
xor ( n319730 , n319717 , n319729 );
buf ( n319731 , n310726 );
buf ( n319732 , n318409 );
or ( n319733 , n319731 , n319732 );
buf ( n29308 , n305449 );
buf ( n319735 , n319658 );
or ( n319736 , n29308 , n319735 );
nand ( n319737 , n319733 , n319736 );
buf ( n319738 , n319737 );
buf ( n319739 , n319738 );
and ( n319740 , n319730 , n319739 );
and ( n29315 , n319717 , n319729 );
or ( n29316 , n319740 , n29315 );
buf ( n319743 , n29316 );
buf ( n319744 , n319743 );
buf ( n319745 , n845 );
buf ( n319746 , n864 );
and ( n319747 , n319745 , n319746 );
buf ( n319748 , n319747 );
buf ( n319749 , n319748 );
buf ( n319750 , n318324 );
not ( n319751 , n319750 );
buf ( n319752 , n14323 );
not ( n319753 , n319752 );
or ( n319754 , n319751 , n319753 );
buf ( n319755 , n837 );
buf ( n319756 , n870 );
xnor ( n29331 , n319755 , n319756 );
buf ( n319758 , n29331 );
buf ( n319759 , n319758 );
not ( n319760 , n319759 );
buf ( n319761 , n311052 );
nand ( n319762 , n319760 , n319761 );
buf ( n319763 , n319762 );
buf ( n319764 , n319763 );
nand ( n319765 , n319754 , n319764 );
buf ( n319766 , n319765 );
buf ( n319767 , n319766 );
xor ( n319768 , n319749 , n319767 );
buf ( n319769 , n306340 );
buf ( n319770 , n318387 );
or ( n319771 , n319769 , n319770 );
buf ( n319772 , n306346 );
buf ( n319773 , n315090 );
buf ( n319774 , n833 );
and ( n29349 , n319773 , n319774 );
buf ( n319776 , n310964 );
buf ( n319777 , n874 );
and ( n319778 , n319776 , n319777 );
nor ( n29353 , n29349 , n319778 );
buf ( n29354 , n29353 );
buf ( n319781 , n29354 );
or ( n29356 , n319772 , n319781 );
nand ( n319783 , n319771 , n29356 );
buf ( n319784 , n319783 );
buf ( n319785 , n319784 );
and ( n29360 , n319768 , n319785 );
and ( n29361 , n319749 , n319767 );
or ( n319788 , n29360 , n29361 );
buf ( n319789 , n319788 );
buf ( n319790 , n319789 );
xor ( n29365 , n319744 , n319790 );
buf ( n319792 , n310629 );
buf ( n319793 , n29354 );
or ( n29368 , n319792 , n319793 );
buf ( n319795 , n306346 );
buf ( n319796 , n874 );
buf ( n319797 , n20700 );
and ( n319798 , n319796 , n319797 );
not ( n29373 , n319796 );
buf ( n319800 , n832 );
and ( n29375 , n29373 , n319800 );
nor ( n319802 , n319798 , n29375 );
buf ( n319803 , n319802 );
buf ( n319804 , n319803 );
or ( n319805 , n319795 , n319804 );
nand ( n319806 , n29368 , n319805 );
buf ( n319807 , n319806 );
buf ( n319808 , n319807 );
buf ( n319809 , n315120 );
buf ( n319810 , n319758 );
or ( n319811 , n319809 , n319810 );
buf ( n319812 , n304760 );
buf ( n319813 , n870 );
not ( n319814 , n319813 );
buf ( n319815 , n319814 );
buf ( n319816 , n319815 );
buf ( n319817 , n836 );
and ( n29392 , n319816 , n319817 );
buf ( n319819 , n311204 );
buf ( n319820 , n870 );
and ( n29395 , n319819 , n319820 );
nor ( n319822 , n29392 , n29395 );
buf ( n319823 , n319822 );
buf ( n319824 , n319823 );
or ( n319825 , n319812 , n319824 );
nand ( n319826 , n319811 , n319825 );
buf ( n319827 , n319826 );
buf ( n319828 , n319827 );
xor ( n319829 , n319808 , n319828 );
buf ( n319830 , n305338 );
buf ( n319831 , n305344 );
or ( n319832 , n319830 , n319831 );
buf ( n319833 , n876 );
nand ( n319834 , n319832 , n319833 );
buf ( n319835 , n319834 );
buf ( n319836 , n319835 );
xor ( n319837 , n319829 , n319836 );
buf ( n319838 , n319837 );
buf ( n319839 , n319838 );
xor ( n319840 , n29365 , n319839 );
buf ( n319841 , n319840 );
buf ( n319842 , n319841 );
xor ( n319843 , n318307 , n318331 );
and ( n29418 , n319843 , n318345 );
and ( n29419 , n318307 , n318331 );
or ( n319846 , n29418 , n29419 );
buf ( n319847 , n319846 );
buf ( n319848 , n319847 );
xor ( n319849 , n318371 , n318396 );
and ( n319850 , n319849 , n318414 );
and ( n29425 , n318371 , n318396 );
or ( n319852 , n319850 , n29425 );
buf ( n319853 , n319852 );
buf ( n319854 , n319853 );
xor ( n319855 , n319848 , n319854 );
xor ( n319856 , n319717 , n319729 );
xor ( n319857 , n319856 , n319739 );
buf ( n319858 , n319857 );
buf ( n319859 , n319858 );
and ( n319860 , n319855 , n319859 );
and ( n319861 , n319848 , n319854 );
or ( n29436 , n319860 , n319861 );
buf ( n319863 , n29436 );
buf ( n29438 , n319863 );
xor ( n29439 , n319842 , n29438 );
xor ( n319866 , n319749 , n319767 );
xor ( n319867 , n319866 , n319785 );
buf ( n319868 , n319867 );
buf ( n319869 , n319868 );
xor ( n319870 , n319680 , n319689 );
xor ( n29445 , n319870 , n319696 );
buf ( n319872 , n29445 );
buf ( n319873 , n319872 );
xor ( n29448 , n319869 , n319873 );
xor ( n319875 , n318272 , n318277 );
and ( n319876 , n319875 , n318283 );
and ( n29451 , n318272 , n318277 );
or ( n319878 , n319876 , n29451 );
buf ( n319879 , n319878 );
and ( n29454 , n29448 , n319879 );
and ( n319881 , n319869 , n319873 );
or ( n319882 , n29454 , n319881 );
buf ( n319883 , n319882 );
buf ( n319884 , n319883 );
xor ( n319885 , n29439 , n319884 );
buf ( n319886 , n319885 );
buf ( n319887 , n319886 );
xor ( n319888 , n319848 , n319854 );
xor ( n29463 , n319888 , n319859 );
buf ( n319890 , n29463 );
xor ( n319891 , n318347 , n318416 );
and ( n29466 , n319891 , n318464 );
and ( n319893 , n318347 , n318416 );
or ( n29468 , n29466 , n319893 );
xor ( n29469 , n319890 , n29468 );
xor ( n319896 , n319869 , n319873 );
xor ( n319897 , n319896 , n319879 );
buf ( n319898 , n319897 );
and ( n319899 , n29469 , n319898 );
and ( n319900 , n319890 , n29468 );
or ( n29475 , n319899 , n319900 );
buf ( n319902 , n29475 );
xor ( n319903 , n319703 , n319887 );
xor ( n29478 , n319903 , n319902 );
buf ( n319905 , n29478 );
xor ( n29480 , n319703 , n319887 );
and ( n319907 , n29480 , n319902 );
and ( n319908 , n319703 , n319887 );
or ( n29483 , n319907 , n319908 );
buf ( n319910 , n29483 );
xor ( n29485 , n313250 , n313256 );
and ( n319912 , n29485 , n313263 );
and ( n319913 , n313250 , n313256 );
or ( n29488 , n319912 , n319913 );
buf ( n319915 , n29488 );
buf ( n319916 , n319915 );
xor ( n29491 , n318022 , n318028 );
xor ( n319918 , n29491 , n318035 );
buf ( n319919 , n319918 );
buf ( n319920 , n319919 );
xor ( n319921 , n22862 , n313294 );
and ( n29496 , n319921 , n313425 );
and ( n29497 , n22862 , n313294 );
or ( n319924 , n29496 , n29497 );
buf ( n319925 , n319924 );
buf ( n319926 , n319925 );
xor ( n319927 , n319916 , n319920 );
xor ( n319928 , n319927 , n319926 );
buf ( n319929 , n319928 );
xor ( n319930 , n319916 , n319920 );
and ( n319931 , n319930 , n319926 );
and ( n319932 , n319916 , n319920 );
or ( n319933 , n319931 , n319932 );
buf ( n319934 , n319933 );
xor ( n319935 , n319321 , n319336 );
xor ( n319936 , n319935 , n319341 );
buf ( n319937 , n319936 );
buf ( n319938 , n319937 );
xor ( n29513 , n319272 , n319293 );
xor ( n29514 , n29513 , n319311 );
buf ( n319941 , n29514 );
buf ( n319942 , n319941 );
xor ( n29517 , n319370 , n319394 );
xor ( n319944 , n29517 , n319411 );
buf ( n319945 , n319944 );
buf ( n319946 , n319945 );
xor ( n319947 , n319942 , n319946 );
xor ( n319948 , n319450 , n319470 );
xor ( n29523 , n319948 , n319473 );
buf ( n319950 , n29523 );
buf ( n319951 , n319950 );
and ( n319952 , n319947 , n319951 );
and ( n29527 , n319942 , n319946 );
or ( n29528 , n319952 , n29527 );
buf ( n319955 , n29528 );
buf ( n319956 , n319955 );
buf ( n319957 , n306272 );
buf ( n319958 , n863 );
and ( n319959 , n319957 , n319958 );
buf ( n319960 , n319959 );
buf ( n319961 , n319960 );
buf ( n319962 , n305881 );
buf ( n319963 , n894 );
buf ( n319964 , n848 );
xnor ( n319965 , n319963 , n319964 );
buf ( n319966 , n319965 );
buf ( n319967 , n319966 );
or ( n29542 , n319962 , n319967 );
buf ( n319969 , n15469 );
buf ( n319970 , n319251 );
or ( n29545 , n319969 , n319970 );
nand ( n319972 , n29542 , n29545 );
buf ( n319973 , n319972 );
buf ( n319974 , n319973 );
xor ( n29549 , n319961 , n319974 );
buf ( n319976 , n305561 );
buf ( n319977 , n850 );
buf ( n319978 , n892 );
xnor ( n29553 , n319977 , n319978 );
buf ( n319980 , n29553 );
buf ( n319981 , n319980 );
or ( n29556 , n319976 , n319981 );
buf ( n319983 , n305489 );
buf ( n319984 , n319354 );
or ( n29559 , n319983 , n319984 );
nand ( n29560 , n29556 , n29559 );
buf ( n319987 , n29560 );
buf ( n319988 , n319987 );
and ( n319989 , n29549 , n319988 );
and ( n29564 , n319961 , n319974 );
or ( n29565 , n319989 , n29564 );
buf ( n319992 , n29565 );
buf ( n319993 , n319992 );
buf ( n319994 , n856 );
buf ( n319995 , n886 );
xor ( n319996 , n319994 , n319995 );
buf ( n319997 , n319996 );
buf ( n319998 , n319997 );
not ( n319999 , n319998 );
buf ( n320000 , n304912 );
not ( n320001 , n320000 );
or ( n29576 , n319999 , n320001 );
buf ( n320003 , n319400 );
not ( n29578 , n320003 );
buf ( n320005 , n304901 );
nand ( n320006 , n29578 , n320005 );
buf ( n320007 , n320006 );
buf ( n320008 , n320007 );
nand ( n29583 , n29576 , n320008 );
buf ( n29584 , n29583 );
buf ( n320011 , n29584 );
buf ( n320012 , n862 );
buf ( n320013 , n880 );
xor ( n320014 , n320012 , n320013 );
buf ( n320015 , n320014 );
buf ( n320016 , n320015 );
not ( n320017 , n320016 );
buf ( n320018 , n304984 );
not ( n320019 , n320018 );
or ( n320020 , n320017 , n320019 );
buf ( n320021 , n304973 );
buf ( n320022 , n28833 );
nand ( n29597 , n320021 , n320022 );
buf ( n320024 , n29597 );
buf ( n320025 , n320024 );
nand ( n320026 , n320020 , n320025 );
buf ( n320027 , n320026 );
buf ( n320028 , n320027 );
xor ( n320029 , n320011 , n320028 );
buf ( n320030 , n305135 );
buf ( n320031 , n854 );
buf ( n320032 , n888 );
xnor ( n29607 , n320031 , n320032 );
buf ( n320034 , n29607 );
buf ( n320035 , n320034 );
or ( n320036 , n320030 , n320035 );
buf ( n320037 , n15861 );
buf ( n320038 , n319303 );
or ( n29613 , n320037 , n320038 );
nand ( n29614 , n320036 , n29613 );
buf ( n320041 , n29614 );
buf ( n320042 , n320041 );
and ( n320043 , n320029 , n320042 );
and ( n29618 , n320011 , n320028 );
or ( n320045 , n320043 , n29618 );
buf ( n320046 , n320045 );
buf ( n320047 , n320046 );
xor ( n29622 , n319993 , n320047 );
buf ( n29623 , n860 );
buf ( n320050 , n882 );
xor ( n320051 , n29623 , n320050 );
buf ( n320052 , n320051 );
buf ( n320053 , n320052 );
not ( n29628 , n320053 );
buf ( n320055 , n304584 );
not ( n29630 , n320055 );
or ( n320057 , n29628 , n29630 );
buf ( n320058 , n319442 );
not ( n320059 , n320058 );
buf ( n29634 , n304596 );
nand ( n29635 , n320059 , n29634 );
buf ( n29636 , n29635 );
buf ( n320063 , n29636 );
nand ( n29638 , n320057 , n320063 );
buf ( n29639 , n29638 );
buf ( n29640 , n29639 );
buf ( n320067 , n15804 );
buf ( n320068 , n858 );
buf ( n320069 , n884 );
xnor ( n29644 , n320068 , n320069 );
buf ( n320071 , n29644 );
buf ( n320072 , n320071 );
or ( n320073 , n320067 , n320072 );
buf ( n320074 , n310909 );
buf ( n320075 , n319459 );
or ( n320076 , n320074 , n320075 );
nand ( n320077 , n320073 , n320076 );
buf ( n320078 , n320077 );
buf ( n320079 , n320078 );
xor ( n320080 , n29640 , n320079 );
buf ( n320081 , n304633 );
not ( n320082 , n320081 );
buf ( n320083 , n320082 );
buf ( n320084 , n320083 );
buf ( n320085 , n312467 );
buf ( n320086 , n852 );
and ( n29661 , n320085 , n320086 );
buf ( n320088 , n305168 );
buf ( n320089 , n890 );
and ( n320090 , n320088 , n320089 );
nor ( n320091 , n29661 , n320090 );
buf ( n320092 , n320091 );
buf ( n320093 , n320092 );
or ( n320094 , n320084 , n320093 );
buf ( n320095 , n304655 );
buf ( n320096 , n319378 );
or ( n320097 , n320095 , n320096 );
nand ( n29672 , n320094 , n320097 );
buf ( n29673 , n29672 );
buf ( n320100 , n29673 );
and ( n29675 , n320080 , n320100 );
and ( n320102 , n29640 , n320079 );
or ( n29677 , n29675 , n320102 );
buf ( n320104 , n29677 );
buf ( n320105 , n320104 );
and ( n29680 , n29622 , n320105 );
and ( n320107 , n319993 , n320047 );
or ( n320108 , n29680 , n320107 );
buf ( n320109 , n320108 );
buf ( n320110 , n320109 );
xor ( n320111 , n319956 , n320110 );
xor ( n320112 , n319350 , n319416 );
xor ( n29687 , n320112 , n319429 );
buf ( n320114 , n29687 );
buf ( n320115 , n320114 );
and ( n29690 , n320111 , n320115 );
and ( n320117 , n319956 , n320110 );
or ( n320118 , n29690 , n320117 );
buf ( n320119 , n320118 );
buf ( n320120 , n320119 );
xor ( n320121 , n319434 , n29062 );
xor ( n29696 , n320121 , n319493 );
buf ( n320123 , n29696 );
buf ( n320124 , n320123 );
xor ( n320125 , n319938 , n320120 );
xor ( n29700 , n320125 , n320124 );
buf ( n320127 , n29700 );
xor ( n320128 , n319938 , n320120 );
and ( n320129 , n320128 , n320124 );
and ( n320130 , n319938 , n320120 );
or ( n29705 , n320129 , n320130 );
buf ( n320132 , n29705 );
xor ( n320133 , n319437 , n319478 );
xor ( n29708 , n320133 , n319483 );
buf ( n320135 , n29708 );
buf ( n320136 , n320135 );
buf ( n320137 , n863 );
buf ( n320138 , n881 );
or ( n29713 , n320137 , n320138 );
buf ( n320140 , n882 );
nand ( n29715 , n29713 , n320140 );
buf ( n320142 , n29715 );
buf ( n29717 , n320142 );
buf ( n320144 , n863 );
buf ( n320145 , n881 );
nand ( n320146 , n320144 , n320145 );
buf ( n320147 , n320146 );
buf ( n320148 , n320147 );
buf ( n320149 , n880 );
and ( n29724 , n29717 , n320148 , n320149 );
buf ( n320151 , n29724 );
buf ( n320152 , n320151 );
buf ( n320153 , n305881 );
buf ( n320154 , n894 );
buf ( n320155 , n849 );
xor ( n29730 , n320154 , n320155 );
buf ( n320157 , n29730 );
buf ( n29732 , n320157 );
not ( n320159 , n29732 );
buf ( n320160 , n320159 );
buf ( n320161 , n320160 );
or ( n320162 , n320153 , n320161 );
buf ( n320163 , n319966 );
buf ( n320164 , n15469 );
or ( n320165 , n320163 , n320164 );
nand ( n29740 , n320162 , n320165 );
buf ( n29741 , n29740 );
buf ( n320168 , n29741 );
and ( n320169 , n320152 , n320168 );
buf ( n320170 , n320169 );
buf ( n320171 , n888 );
buf ( n320172 , n855 );
and ( n29747 , n320171 , n320172 );
not ( n320174 , n320171 );
buf ( n320175 , n305319 );
and ( n29750 , n320174 , n320175 );
nor ( n320177 , n29747 , n29750 );
buf ( n320178 , n320177 );
buf ( n320179 , n320178 );
not ( n320180 , n320179 );
buf ( n320181 , n305138 );
not ( n29756 , n320181 );
or ( n320183 , n320180 , n29756 );
buf ( n320184 , n320034 );
not ( n320185 , n320184 );
buf ( n320186 , n305144 );
nand ( n320187 , n320185 , n320186 );
buf ( n320188 , n320187 );
buf ( n320189 , n320188 );
nand ( n320190 , n320183 , n320189 );
buf ( n320191 , n320190 );
buf ( n320192 , n320191 );
buf ( n320193 , n305561 );
buf ( n320194 , n851 );
buf ( n320195 , n892 );
xnor ( n29770 , n320194 , n320195 );
buf ( n320197 , n29770 );
buf ( n320198 , n320197 );
or ( n320199 , n320193 , n320198 );
buf ( n320200 , n305489 );
buf ( n320201 , n319980 );
or ( n320202 , n320200 , n320201 );
nand ( n320203 , n320199 , n320202 );
buf ( n320204 , n320203 );
buf ( n320205 , n320204 );
xor ( n320206 , n320192 , n320205 );
buf ( n320207 , n304987 );
buf ( n320208 , n21800 );
buf ( n320209 , n863 );
and ( n29784 , n320208 , n320209 );
buf ( n320211 , n305192 );
buf ( n320212 , n880 );
and ( n320213 , n320211 , n320212 );
nor ( n29788 , n29784 , n320213 );
buf ( n320215 , n29788 );
buf ( n320216 , n320215 );
or ( n29791 , n320207 , n320216 );
buf ( n320218 , n305000 );
buf ( n320219 , n320015 );
not ( n29794 , n320219 );
buf ( n29795 , n29794 );
buf ( n320222 , n29795 );
or ( n320223 , n320218 , n320222 );
nand ( n29798 , n29791 , n320223 );
buf ( n29799 , n29798 );
buf ( n320226 , n29799 );
and ( n29801 , n320206 , n320226 );
and ( n320228 , n320192 , n320205 );
or ( n320229 , n29801 , n320228 );
buf ( n320230 , n320229 );
xor ( n29805 , n320170 , n320230 );
buf ( n320232 , n15804 );
buf ( n320233 , n884 );
buf ( n320234 , n14447 );
and ( n320235 , n320233 , n320234 );
not ( n320236 , n320233 );
buf ( n320237 , n859 );
and ( n29812 , n320236 , n320237 );
nor ( n320239 , n320235 , n29812 );
buf ( n320240 , n320239 );
buf ( n320241 , n320240 );
or ( n320242 , n320232 , n320241 );
buf ( n29817 , n306238 );
buf ( n320244 , n320071 );
or ( n320245 , n29817 , n320244 );
nand ( n320246 , n320242 , n320245 );
buf ( n320247 , n320246 );
buf ( n320248 , n320247 );
buf ( n320249 , n304630 );
buf ( n320250 , n890 );
buf ( n320251 , n304956 );
and ( n29826 , n320250 , n320251 );
not ( n320253 , n320250 );
buf ( n29828 , n853 );
and ( n320255 , n320253 , n29828 );
nor ( n29830 , n29826 , n320255 );
buf ( n29831 , n29830 );
buf ( n320258 , n29831 );
or ( n29833 , n320249 , n320258 );
buf ( n320260 , n320092 );
buf ( n320261 , n304655 );
or ( n29836 , n320260 , n320261 );
nand ( n320263 , n29833 , n29836 );
buf ( n320264 , n320263 );
buf ( n320265 , n320264 );
xor ( n320266 , n320248 , n320265 );
buf ( n320267 , n313403 );
buf ( n320268 , n857 );
buf ( n320269 , n886 );
xnor ( n29844 , n320268 , n320269 );
buf ( n320271 , n29844 );
buf ( n320272 , n320271 );
or ( n320273 , n320267 , n320272 );
buf ( n320274 , n305363 );
buf ( n320275 , n319997 );
not ( n320276 , n320275 );
buf ( n320277 , n320276 );
buf ( n320278 , n320277 );
or ( n29853 , n320274 , n320278 );
nand ( n29854 , n320273 , n29853 );
buf ( n320281 , n29854 );
buf ( n320282 , n320281 );
and ( n320283 , n320266 , n320282 );
and ( n320284 , n320248 , n320265 );
or ( n29859 , n320283 , n320284 );
buf ( n320286 , n29859 );
and ( n320287 , n29805 , n320286 );
and ( n29862 , n320170 , n320230 );
or ( n29863 , n320287 , n29862 );
buf ( n320290 , n29863 );
xor ( n29865 , n319993 , n320047 );
xor ( n29866 , n29865 , n320105 );
buf ( n320293 , n29866 );
buf ( n320294 , n320293 );
xor ( n29869 , n320290 , n320294 );
xor ( n29870 , n29640 , n320079 );
xor ( n29871 , n29870 , n320100 );
buf ( n320298 , n29871 );
buf ( n320299 , n320298 );
xor ( n29874 , n319961 , n319974 );
xor ( n29875 , n29874 , n319988 );
buf ( n320302 , n29875 );
buf ( n320303 , n320302 );
xor ( n320304 , n320299 , n320303 );
xor ( n29879 , n320011 , n320028 );
xor ( n320306 , n29879 , n320042 );
buf ( n320307 , n320306 );
buf ( n320308 , n320307 );
and ( n320309 , n320304 , n320308 );
and ( n320310 , n320299 , n320303 );
or ( n320311 , n320309 , n320310 );
buf ( n320312 , n320311 );
buf ( n29887 , n320312 );
and ( n29888 , n29869 , n29887 );
and ( n29889 , n320290 , n320294 );
or ( n29890 , n29888 , n29889 );
buf ( n29891 , n29890 );
buf ( n29892 , n29891 );
xor ( n29893 , n319956 , n320110 );
xor ( n320320 , n29893 , n320115 );
buf ( n320321 , n320320 );
buf ( n320322 , n320321 );
xor ( n320323 , n320136 , n29892 );
xor ( n320324 , n320323 , n320322 );
buf ( n320325 , n320324 );
xor ( n320326 , n320136 , n29892 );
and ( n29901 , n320326 , n320322 );
and ( n320328 , n320136 , n29892 );
or ( n29903 , n29901 , n320328 );
buf ( n320330 , n29903 );
xor ( n320331 , n319942 , n319946 );
xor ( n320332 , n320331 , n319951 );
buf ( n320333 , n320332 );
buf ( n320334 , n320333 );
xor ( n320335 , n320152 , n320168 );
buf ( n320336 , n320335 );
buf ( n320337 , n320336 );
buf ( n320338 , n305381 );
buf ( n320339 , n861 );
buf ( n29914 , n882 );
xnor ( n29915 , n320339 , n29914 );
buf ( n29916 , n29915 );
buf ( n320343 , n29916 );
or ( n320344 , n320338 , n320343 );
buf ( n320345 , n14959 );
buf ( n320346 , n320052 );
not ( n320347 , n320346 );
buf ( n320348 , n320347 );
buf ( n320349 , n320348 );
or ( n320350 , n320345 , n320349 );
nand ( n29925 , n320344 , n320350 );
buf ( n320352 , n29925 );
buf ( n320353 , n320352 );
xor ( n320354 , n320337 , n320353 );
buf ( n320355 , n863 );
buf ( n320356 , n304997 );
and ( n320357 , n320355 , n320356 );
buf ( n320358 , n320357 );
buf ( n320359 , n320358 );
buf ( n320360 , n894 );
buf ( n320361 , n850 );
xor ( n320362 , n320360 , n320361 );
buf ( n320363 , n320362 );
buf ( n320364 , n320363 );
not ( n320365 , n320364 );
buf ( n320366 , n28078 );
not ( n29941 , n320366 );
or ( n320368 , n320365 , n29941 );
buf ( n29943 , n320157 );
buf ( n320370 , n895 );
nand ( n29945 , n29943 , n320370 );
buf ( n320372 , n29945 );
buf ( n320373 , n320372 );
nand ( n320374 , n320368 , n320373 );
buf ( n320375 , n320374 );
buf ( n320376 , n320375 );
xor ( n320377 , n320359 , n320376 );
buf ( n320378 , n852 );
buf ( n320379 , n892 );
xnor ( n320380 , n320378 , n320379 );
buf ( n320381 , n320380 );
buf ( n320382 , n320381 );
not ( n29957 , n320382 );
buf ( n320384 , n29957 );
buf ( n320385 , n320384 );
not ( n320386 , n320385 );
buf ( n320387 , n14272 );
not ( n29962 , n320387 );
or ( n320389 , n320386 , n29962 );
buf ( n320390 , n320197 );
not ( n29965 , n320390 );
buf ( n320392 , n305430 );
nand ( n320393 , n29965 , n320392 );
buf ( n320394 , n320393 );
buf ( n320395 , n320394 );
nand ( n320396 , n320389 , n320395 );
buf ( n320397 , n320396 );
buf ( n320398 , n320397 );
and ( n320399 , n320377 , n320398 );
and ( n320400 , n320359 , n320376 );
or ( n29975 , n320399 , n320400 );
buf ( n320402 , n29975 );
buf ( n320403 , n320402 );
and ( n29978 , n320354 , n320403 );
and ( n320405 , n320337 , n320353 );
or ( n320406 , n29978 , n320405 );
buf ( n320407 , n320406 );
xor ( n320408 , n320170 , n320230 );
xor ( n320409 , n320408 , n320286 );
and ( n320410 , n320407 , n320409 );
xor ( n29985 , n320248 , n320265 );
xor ( n320412 , n29985 , n320282 );
buf ( n320413 , n320412 );
buf ( n320414 , n320413 );
buf ( n320415 , n314747 );
buf ( n320416 , n886 );
buf ( n320417 , n305060 );
and ( n320418 , n320416 , n320417 );
not ( n320419 , n320416 );
buf ( n320420 , n858 );
and ( n320421 , n320419 , n320420 );
nor ( n29996 , n320418 , n320421 );
buf ( n320423 , n29996 );
buf ( n320424 , n320423 );
or ( n320425 , n320415 , n320424 );
buf ( n320426 , n305363 );
buf ( n320427 , n320271 );
or ( n320428 , n320426 , n320427 );
nand ( n320429 , n320425 , n320428 );
buf ( n320430 , n320429 );
buf ( n320431 , n320430 );
buf ( n320432 , n304630 );
buf ( n320433 , n890 );
buf ( n320434 , n26347 );
and ( n320435 , n320433 , n320434 );
not ( n30010 , n320433 );
buf ( n320437 , n854 );
and ( n320438 , n30010 , n320437 );
nor ( n30013 , n320435 , n320438 );
buf ( n30014 , n30013 );
buf ( n320441 , n30014 );
or ( n320442 , n320432 , n320441 );
buf ( n320443 , n304655 );
buf ( n320444 , n29831 );
or ( n30019 , n320443 , n320444 );
nand ( n320446 , n320442 , n30019 );
buf ( n320447 , n320446 );
buf ( n320448 , n320447 );
xor ( n30023 , n320431 , n320448 );
buf ( n320450 , n306283 );
buf ( n320451 , n888 );
buf ( n320452 , n15582 );
and ( n320453 , n320451 , n320452 );
not ( n320454 , n320451 );
buf ( n320455 , n856 );
and ( n30030 , n320454 , n320455 );
nor ( n320457 , n320453 , n30030 );
buf ( n320458 , n320457 );
buf ( n320459 , n320458 );
or ( n320460 , n320450 , n320459 );
buf ( n320461 , n15861 );
buf ( n320462 , n320178 );
not ( n320463 , n320462 );
buf ( n320464 , n320463 );
buf ( n320465 , n320464 );
or ( n320466 , n320461 , n320465 );
nand ( n30041 , n320460 , n320466 );
buf ( n30042 , n30041 );
buf ( n320469 , n30042 );
and ( n30044 , n30023 , n320469 );
and ( n320471 , n320431 , n320448 );
or ( n320472 , n30044 , n320471 );
buf ( n320473 , n320472 );
buf ( n320474 , n320473 );
xor ( n320475 , n320414 , n320474 );
xor ( n30050 , n320192 , n320205 );
xor ( n320477 , n30050 , n320226 );
buf ( n320478 , n320477 );
buf ( n320479 , n320478 );
and ( n320480 , n320475 , n320479 );
and ( n320481 , n320414 , n320474 );
or ( n30056 , n320480 , n320481 );
buf ( n320483 , n30056 );
xor ( n320484 , n320170 , n320230 );
xor ( n320485 , n320484 , n320286 );
and ( n320486 , n320483 , n320485 );
and ( n30061 , n320407 , n320483 );
or ( n320488 , n320410 , n320486 , n30061 );
buf ( n320489 , n320488 );
xor ( n30064 , n320290 , n320294 );
xor ( n320491 , n30064 , n29887 );
buf ( n320492 , n320491 );
buf ( n320493 , n320492 );
xor ( n320494 , n320334 , n320489 );
xor ( n320495 , n320494 , n320493 );
buf ( n320496 , n320495 );
xor ( n320497 , n320334 , n320489 );
and ( n320498 , n320497 , n320493 );
and ( n320499 , n320334 , n320489 );
or ( n30074 , n320498 , n320499 );
buf ( n320501 , n30074 );
xor ( n320502 , n29162 , n319608 );
xor ( n320503 , n320502 , n319620 );
and ( n30078 , n319676 , n320503 );
xor ( n320505 , n29162 , n319608 );
xor ( n320506 , n320505 , n319620 );
and ( n30081 , n319700 , n320506 );
and ( n320508 , n319676 , n319700 );
or ( n320509 , n30078 , n30081 , n320508 );
buf ( n320510 , n320509 );
xor ( n30085 , n319744 , n319790 );
and ( n320512 , n30085 , n319839 );
and ( n320513 , n319744 , n319790 );
or ( n30088 , n320512 , n320513 );
buf ( n320515 , n30088 );
buf ( n320516 , n320515 );
xor ( n30091 , n29200 , n29222 );
and ( n320518 , n30091 , n319674 );
and ( n320519 , n29200 , n29222 );
or ( n30094 , n320518 , n320519 );
buf ( n320521 , n30094 );
buf ( n30096 , n320521 );
buf ( n320523 , n305627 );
buf ( n320524 , n319803 );
not ( n320525 , n320524 );
buf ( n320526 , n320525 );
buf ( n320527 , n320526 );
and ( n320528 , n320523 , n320527 );
buf ( n320529 , n305301 );
buf ( n320530 , n874 );
and ( n320531 , n320529 , n320530 );
nor ( n30106 , n320528 , n320531 );
buf ( n320533 , n30106 );
buf ( n320534 , n320533 );
xor ( n320535 , n30096 , n320534 );
xor ( n320536 , n319808 , n319828 );
and ( n320537 , n320536 , n319836 );
and ( n320538 , n319808 , n319828 );
or ( n30113 , n320537 , n320538 );
buf ( n320540 , n30113 );
buf ( n320541 , n320540 );
xor ( n30116 , n320535 , n320541 );
buf ( n320543 , n30116 );
buf ( n320544 , n320543 );
xor ( n320545 , n320516 , n320544 );
buf ( n320546 , n313215 );
buf ( n320547 , n319584 );
or ( n320548 , n320546 , n320547 );
buf ( n320549 , n313224 );
buf ( n320550 , n839 );
buf ( n320551 , n866 );
xnor ( n30126 , n320550 , n320551 );
buf ( n320553 , n30126 );
buf ( n320554 , n320553 );
or ( n320555 , n320549 , n320554 );
nand ( n320556 , n320548 , n320555 );
buf ( n320557 , n320556 );
buf ( n320558 , n320557 );
buf ( n320559 , n304854 );
buf ( n320560 , n319639 );
or ( n30135 , n320559 , n320560 );
buf ( n320562 , n14439 );
buf ( n320563 , n872 );
buf ( n30138 , n310964 );
and ( n30139 , n320563 , n30138 );
not ( n320566 , n320563 );
buf ( n320567 , n833 );
and ( n320568 , n320566 , n320567 );
nor ( n320569 , n30139 , n320568 );
buf ( n320570 , n320569 );
buf ( n320571 , n320570 );
or ( n30146 , n320562 , n320571 );
nand ( n320573 , n30135 , n30146 );
buf ( n320574 , n320573 );
buf ( n320575 , n320574 );
xor ( n30150 , n320558 , n320575 );
buf ( n320577 , n310726 );
buf ( n320578 , n29243 );
or ( n320579 , n320577 , n320578 );
buf ( n320580 , n305449 );
buf ( n320581 , n310521 );
buf ( n320582 , n837 );
and ( n30157 , n320581 , n320582 );
buf ( n320584 , n313757 );
buf ( n320585 , n868 );
and ( n30160 , n320584 , n320585 );
nor ( n30161 , n30157 , n30160 );
buf ( n320588 , n30161 );
buf ( n320589 , n320588 );
or ( n320590 , n320580 , n320589 );
nand ( n320591 , n320579 , n320590 );
buf ( n320592 , n320591 );
buf ( n320593 , n320592 );
xor ( n30168 , n30150 , n320593 );
buf ( n320595 , n30168 );
buf ( n320596 , n320595 );
xor ( n320597 , n29162 , n319608 );
and ( n320598 , n320597 , n319620 );
and ( n30173 , n29162 , n319608 );
or ( n30174 , n320598 , n30173 );
buf ( n320601 , n30174 );
xor ( n320602 , n320596 , n320601 );
buf ( n320603 , n843 );
buf ( n320604 , n864 );
and ( n320605 , n320603 , n320604 );
buf ( n320606 , n320605 );
buf ( n320607 , n320606 );
buf ( n320608 , n314219 );
buf ( n320609 , n319823 );
or ( n30184 , n320608 , n320609 );
buf ( n320611 , n304760 );
buf ( n320612 , n319815 );
buf ( n320613 , n835 );
and ( n320614 , n320612 , n320613 );
buf ( n320615 , n21261 );
buf ( n320616 , n870 );
and ( n320617 , n320615 , n320616 );
nor ( n320618 , n320614 , n320617 );
buf ( n320619 , n320618 );
buf ( n320620 , n320619 );
or ( n320621 , n320611 , n320620 );
nand ( n320622 , n30184 , n320621 );
buf ( n320623 , n320622 );
buf ( n320624 , n320623 );
xor ( n320625 , n320607 , n320624 );
buf ( n320626 , n311891 );
buf ( n320627 , n319604 );
or ( n320628 , n320626 , n320627 );
buf ( n320629 , n311246 );
buf ( n320630 , n311234 );
buf ( n320631 , n841 );
and ( n30206 , n320630 , n320631 );
buf ( n320633 , n310600 );
buf ( n320634 , n864 );
and ( n30209 , n320633 , n320634 );
nor ( n30210 , n30206 , n30209 );
buf ( n320637 , n30210 );
buf ( n320638 , n320637 );
or ( n30213 , n320629 , n320638 );
nand ( n320640 , n320628 , n30213 );
buf ( n320641 , n320640 );
buf ( n320642 , n320641 );
xor ( n320643 , n320625 , n320642 );
buf ( n320644 , n320643 );
buf ( n320645 , n320644 );
xor ( n320646 , n320602 , n320645 );
buf ( n320647 , n320646 );
buf ( n320648 , n320647 );
xor ( n320649 , n320545 , n320648 );
buf ( n320650 , n320649 );
buf ( n320651 , n320650 );
xor ( n320652 , n319842 , n29438 );
and ( n320653 , n320652 , n319884 );
and ( n320654 , n319842 , n29438 );
or ( n30229 , n320653 , n320654 );
buf ( n320656 , n30229 );
buf ( n320657 , n320656 );
xor ( n320658 , n320510 , n320651 );
xor ( n320659 , n320658 , n320657 );
buf ( n320660 , n320659 );
xor ( n30235 , n320510 , n320651 );
and ( n30236 , n30235 , n320657 );
and ( n30237 , n320510 , n320651 );
or ( n320664 , n30236 , n30237 );
buf ( n320665 , n320664 );
xor ( n30240 , n317955 , n317975 );
xor ( n320667 , n30240 , n317996 );
buf ( n320668 , n320667 );
xor ( n30243 , n311588 , n311857 );
xor ( n320670 , n30243 , n311862 );
buf ( n320671 , n320670 );
xor ( n320672 , n317893 , n317908 );
and ( n320673 , n320672 , n317915 );
and ( n30248 , n317893 , n317908 );
or ( n320675 , n320673 , n30248 );
buf ( n320676 , n320675 );
buf ( n320677 , n320676 );
xor ( n320678 , n318172 , n318186 );
xor ( n320679 , n320678 , n318191 );
buf ( n320680 , n320679 );
buf ( n320681 , n320680 );
xor ( n30256 , n320677 , n320681 );
xor ( n30257 , n319538 , n319544 );
and ( n30258 , n30257 , n29125 );
and ( n30259 , n319538 , n319544 );
or ( n30260 , n30258 , n30259 );
buf ( n320687 , n30260 );
buf ( n320688 , n320687 );
xor ( n320689 , n30256 , n320688 );
buf ( n320690 , n320689 );
buf ( n30265 , n320690 );
xor ( n30266 , n27777 , n318209 );
xor ( n320693 , n30266 , n318216 );
buf ( n320694 , n320693 );
buf ( n320695 , n320694 );
xor ( n30270 , n317649 , n317682 );
and ( n320697 , n30270 , n317724 );
and ( n30272 , n317649 , n317682 );
or ( n320699 , n320697 , n30272 );
buf ( n320700 , n320699 );
buf ( n320701 , n320700 );
xor ( n320702 , n320695 , n320701 );
xor ( n30277 , n312009 , n312023 );
xor ( n320704 , n30277 , n312046 );
buf ( n320705 , n320704 );
buf ( n320706 , n320705 );
xor ( n320707 , n317740 , n317753 );
and ( n320708 , n320707 , n317767 );
and ( n30283 , n317740 , n317753 );
or ( n320710 , n320708 , n30283 );
buf ( n320711 , n320710 );
buf ( n320712 , n320711 );
xor ( n30287 , n320706 , n320712 );
xor ( n320714 , n317830 , n317843 );
and ( n30289 , n320714 , n317853 );
and ( n320716 , n317830 , n317843 );
or ( n320717 , n30289 , n320716 );
buf ( n320718 , n320717 );
buf ( n320719 , n320718 );
xor ( n320720 , n30287 , n320719 );
buf ( n320721 , n320720 );
buf ( n320722 , n320721 );
xor ( n320723 , n320702 , n320722 );
buf ( n320724 , n320723 );
buf ( n320725 , n320724 );
xor ( n320726 , n319532 , n319554 );
and ( n30301 , n320726 , n319561 );
and ( n320728 , n319532 , n319554 );
or ( n320729 , n30301 , n320728 );
buf ( n320730 , n320729 );
buf ( n320731 , n320730 );
xor ( n320732 , n30265 , n320725 );
xor ( n30307 , n320732 , n320731 );
buf ( n320734 , n30307 );
xor ( n30309 , n30265 , n320725 );
and ( n320736 , n30309 , n320731 );
and ( n320737 , n30265 , n320725 );
or ( n30312 , n320736 , n320737 );
buf ( n320739 , n30312 );
xor ( n320740 , n320299 , n320303 );
xor ( n30315 , n320740 , n320308 );
buf ( n320742 , n30315 );
buf ( n320743 , n320742 );
xor ( n320744 , n320337 , n320353 );
xor ( n320745 , n320744 , n320403 );
buf ( n320746 , n320745 );
buf ( n320747 , n320746 );
buf ( n320748 , n883 );
buf ( n320749 , n863 );
or ( n320750 , n320748 , n320749 );
buf ( n320751 , n884 );
nand ( n30326 , n320750 , n320751 );
buf ( n320753 , n30326 );
buf ( n320754 , n320753 );
buf ( n320755 , n863 );
buf ( n320756 , n883 );
nand ( n30331 , n320755 , n320756 );
buf ( n30332 , n30331 );
buf ( n320759 , n30332 );
buf ( n320760 , n882 );
and ( n320761 , n320754 , n320759 , n320760 );
buf ( n320762 , n320761 );
buf ( n320763 , n320762 );
buf ( n320764 , n851 );
buf ( n30339 , n894 );
xnor ( n30340 , n320764 , n30339 );
buf ( n320767 , n30340 );
buf ( n30342 , n320767 );
not ( n30343 , n30342 );
buf ( n30344 , n30343 );
buf ( n320771 , n30344 );
not ( n30346 , n320771 );
buf ( n320773 , n28078 );
not ( n320774 , n320773 );
or ( n30349 , n30346 , n320774 );
buf ( n320776 , n320363 );
buf ( n320777 , n895 );
nand ( n30352 , n320776 , n320777 );
buf ( n320779 , n30352 );
buf ( n320780 , n320779 );
nand ( n30355 , n30349 , n320780 );
buf ( n320782 , n30355 );
buf ( n320783 , n320782 );
and ( n30358 , n320763 , n320783 );
buf ( n320785 , n30358 );
buf ( n320786 , n320785 );
buf ( n320787 , n304581 );
buf ( n320788 , n862 );
buf ( n320789 , n882 );
xnor ( n30364 , n320788 , n320789 );
buf ( n320791 , n30364 );
buf ( n320792 , n320791 );
or ( n30367 , n320787 , n320792 );
buf ( n320794 , n14959 );
buf ( n320795 , n29916 );
or ( n320796 , n320794 , n320795 );
nand ( n30371 , n30367 , n320796 );
buf ( n30372 , n30371 );
buf ( n320799 , n30372 );
xor ( n30374 , n320786 , n320799 );
buf ( n320801 , n15804 );
buf ( n320802 , n304827 );
buf ( n320803 , n860 );
and ( n30378 , n320802 , n320803 );
buf ( n320805 , n305241 );
buf ( n320806 , n884 );
and ( n30381 , n320805 , n320806 );
nor ( n320808 , n30378 , n30381 );
buf ( n320809 , n320808 );
buf ( n320810 , n320809 );
or ( n320811 , n320801 , n320810 );
buf ( n320812 , n310909 );
buf ( n320813 , n320240 );
or ( n320814 , n320812 , n320813 );
nand ( n320815 , n320811 , n320814 );
buf ( n320816 , n320815 );
buf ( n320817 , n320816 );
and ( n320818 , n30374 , n320817 );
and ( n30393 , n320786 , n320799 );
or ( n320820 , n320818 , n30393 );
buf ( n320821 , n320820 );
buf ( n320822 , n320821 );
xor ( n320823 , n320747 , n320822 );
xor ( n320824 , n320359 , n320376 );
xor ( n30399 , n320824 , n320398 );
buf ( n320826 , n30399 );
buf ( n320827 , n320826 );
buf ( n320828 , n311275 );
buf ( n320829 , n857 );
buf ( n320830 , n888 );
xnor ( n30405 , n320829 , n320830 );
buf ( n320832 , n30405 );
buf ( n320833 , n320832 );
or ( n320834 , n320828 , n320833 );
buf ( n320835 , n15861 );
buf ( n320836 , n320458 );
or ( n320837 , n320835 , n320836 );
nand ( n30412 , n320834 , n320837 );
buf ( n320839 , n30412 );
buf ( n320840 , n320839 );
buf ( n320841 , n305561 );
and ( n30416 , n892 , n304956 );
not ( n30417 , n892 );
and ( n320844 , n30417 , n853 );
nor ( n30419 , n30416 , n320844 );
buf ( n320846 , n30419 );
or ( n320847 , n320841 , n320846 );
buf ( n320848 , n305489 );
buf ( n320849 , n320381 );
or ( n30424 , n320848 , n320849 );
nand ( n320851 , n320847 , n30424 );
buf ( n320852 , n320851 );
buf ( n320853 , n320852 );
xor ( n320854 , n320840 , n320853 );
buf ( n320855 , n314747 );
buf ( n320856 , n305993 );
buf ( n320857 , n859 );
and ( n320858 , n320856 , n320857 );
buf ( n320859 , n14447 );
buf ( n320860 , n886 );
and ( n320861 , n320859 , n320860 );
nor ( n30436 , n320858 , n320861 );
buf ( n30437 , n30436 );
buf ( n320864 , n30437 );
or ( n30439 , n320855 , n320864 );
buf ( n320866 , n305363 );
buf ( n320867 , n320423 );
or ( n30442 , n320866 , n320867 );
nand ( n320869 , n30439 , n30442 );
buf ( n320870 , n320869 );
buf ( n320871 , n320870 );
and ( n320872 , n320854 , n320871 );
and ( n30447 , n320840 , n320853 );
or ( n320874 , n320872 , n30447 );
buf ( n320875 , n320874 );
buf ( n320876 , n320875 );
xor ( n320877 , n320827 , n320876 );
buf ( n320878 , n882 );
buf ( n320879 , n305192 );
or ( n320880 , n320878 , n320879 );
buf ( n320881 , n305526 );
buf ( n320882 , n863 );
or ( n30457 , n320881 , n320882 );
nand ( n320884 , n320880 , n30457 );
buf ( n320885 , n320884 );
buf ( n320886 , n320885 );
not ( n30461 , n320886 );
buf ( n320888 , n304584 );
not ( n30463 , n320888 );
or ( n30464 , n30461 , n30463 );
buf ( n320891 , n320791 );
not ( n320892 , n320891 );
buf ( n320893 , n304596 );
nand ( n320894 , n320892 , n320893 );
buf ( n320895 , n320894 );
buf ( n320896 , n320895 );
nand ( n320897 , n30464 , n320896 );
buf ( n320898 , n320897 );
buf ( n320899 , n320898 );
buf ( n320900 , n304630 );
buf ( n320901 , n312467 );
buf ( n320902 , n855 );
and ( n320903 , n320901 , n320902 );
buf ( n320904 , n305319 );
buf ( n320905 , n890 );
and ( n30480 , n320904 , n320905 );
nor ( n320907 , n320903 , n30480 );
buf ( n320908 , n320907 );
buf ( n320909 , n320908 );
or ( n320910 , n320900 , n320909 );
buf ( n320911 , n304655 );
buf ( n320912 , n30014 );
or ( n30487 , n320911 , n320912 );
nand ( n320914 , n320910 , n30487 );
buf ( n320915 , n320914 );
buf ( n320916 , n320915 );
xor ( n320917 , n320899 , n320916 );
buf ( n320918 , n15804 );
buf ( n320919 , n861 );
buf ( n320920 , n884 );
xnor ( n30495 , n320919 , n320920 );
buf ( n320922 , n30495 );
buf ( n320923 , n320922 );
or ( n30498 , n320918 , n320923 );
buf ( n320925 , n310909 );
buf ( n320926 , n320809 );
or ( n320927 , n320925 , n320926 );
nand ( n320928 , n30498 , n320927 );
buf ( n320929 , n320928 );
buf ( n320930 , n320929 );
and ( n320931 , n320917 , n320930 );
and ( n320932 , n320899 , n320916 );
or ( n30507 , n320931 , n320932 );
buf ( n320934 , n30507 );
buf ( n320935 , n320934 );
and ( n30510 , n320877 , n320935 );
and ( n320937 , n320827 , n320876 );
or ( n30512 , n30510 , n320937 );
buf ( n320939 , n30512 );
buf ( n320940 , n320939 );
and ( n30515 , n320823 , n320940 );
and ( n320942 , n320747 , n320822 );
or ( n320943 , n30515 , n320942 );
buf ( n320944 , n320943 );
buf ( n320945 , n320944 );
xor ( n320946 , n320170 , n320230 );
xor ( n30521 , n320946 , n320286 );
xor ( n30522 , n320407 , n320483 );
xor ( n320949 , n30521 , n30522 );
buf ( n320950 , n320949 );
xor ( n30525 , n320743 , n320945 );
xor ( n30526 , n30525 , n320950 );
buf ( n320953 , n30526 );
xor ( n30528 , n320743 , n320945 );
and ( n320955 , n30528 , n320950 );
and ( n30530 , n320743 , n320945 );
or ( n30531 , n320955 , n30530 );
buf ( n320958 , n30531 );
xor ( n30533 , n311991 , n312051 );
xor ( n320960 , n30533 , n312116 );
buf ( n320961 , n320960 );
buf ( n320962 , n320961 );
xor ( n30537 , n21752 , n312181 );
xor ( n320964 , n30537 , n312248 );
buf ( n320965 , n320964 );
xor ( n320966 , n320706 , n320712 );
and ( n320967 , n320966 , n320719 );
and ( n30542 , n320706 , n320712 );
or ( n320969 , n320967 , n30542 );
buf ( n320970 , n320969 );
buf ( n320971 , n320970 );
xor ( n30546 , n320962 , n320965 );
xor ( n320973 , n30546 , n320971 );
buf ( n320974 , n320973 );
xor ( n30549 , n320962 , n320965 );
and ( n320976 , n30549 , n320971 );
and ( n30551 , n320962 , n320965 );
or ( n30552 , n320976 , n30551 );
buf ( n320979 , n30552 );
not ( n30554 , n312177 );
nand ( n320981 , n30554 , n312174 );
not ( n30556 , n312152 );
not ( n30557 , n312174 );
nand ( n320984 , n30556 , n30557 , n312138 );
not ( n30559 , n312153 );
nand ( n320986 , n30559 , n312174 );
not ( n320987 , n312152 );
nor ( n320988 , n320987 , n312138 );
nand ( n320989 , n30557 , n320988 );
nand ( n30564 , n320981 , n320984 , n320986 , n320989 );
xor ( n320991 , n312203 , n312220 );
xor ( n320992 , n320991 , n312244 );
buf ( n320993 , n320992 );
xor ( n320994 , n30564 , n320993 );
xor ( n320995 , n312069 , n312090 );
xor ( n30570 , n320995 , n312111 );
buf ( n320997 , n30570 );
and ( n320998 , n320994 , n320997 );
and ( n30573 , n30564 , n320993 );
or ( n30574 , n320998 , n30573 );
buf ( n321001 , n30574 );
xor ( n30576 , n318144 , n318148 );
xor ( n30577 , n30576 , n318153 );
buf ( n321004 , n30577 );
buf ( n321005 , n321004 );
xor ( n321006 , n318169 , n318196 );
xor ( n30581 , n321006 , n318221 );
buf ( n321008 , n30581 );
buf ( n321009 , n321008 );
xor ( n321010 , n321001 , n321005 );
xor ( n30585 , n321010 , n321009 );
buf ( n321012 , n30585 );
xor ( n321013 , n321001 , n321005 );
and ( n30588 , n321013 , n321009 );
and ( n30589 , n321001 , n321005 );
or ( n321016 , n30588 , n30589 );
buf ( n321017 , n321016 );
xor ( n30592 , n317770 , n317816 );
and ( n321019 , n30592 , n317856 );
and ( n30594 , n317770 , n317816 );
or ( n30595 , n321019 , n30594 );
buf ( n321022 , n30595 );
buf ( n321023 , n321022 );
xor ( n30598 , n30564 , n320993 );
xor ( n321025 , n30598 , n320997 );
buf ( n321026 , n321025 );
xor ( n321027 , n317892 , n317918 );
and ( n30602 , n321027 , n317943 );
and ( n321029 , n317892 , n317918 );
or ( n30604 , n30602 , n321029 );
buf ( n321031 , n30604 );
buf ( n321032 , n321031 );
xor ( n30607 , n321023 , n321026 );
xor ( n321034 , n30607 , n321032 );
buf ( n321035 , n321034 );
xor ( n30610 , n321023 , n321026 );
and ( n30611 , n30610 , n321032 );
and ( n321038 , n321023 , n321026 );
or ( n30613 , n30611 , n321038 );
buf ( n321040 , n30613 );
xor ( n30615 , n317727 , n317859 );
and ( n321042 , n30615 , n317946 );
and ( n30617 , n317727 , n317859 );
or ( n30618 , n321042 , n30617 );
buf ( n321045 , n30618 );
xor ( n321046 , n320763 , n320783 );
buf ( n321047 , n321046 );
buf ( n321048 , n321047 );
buf ( n321049 , n305881 );
buf ( n321050 , n894 );
buf ( n321051 , n852 );
xnor ( n321052 , n321050 , n321051 );
buf ( n321053 , n321052 );
buf ( n321054 , n321053 );
or ( n321055 , n321049 , n321054 );
buf ( n321056 , n320767 );
buf ( n321057 , n15469 );
or ( n30632 , n321056 , n321057 );
nand ( n30633 , n321055 , n30632 );
buf ( n321060 , n30633 );
buf ( n321061 , n321060 );
or ( n30636 , n310909 , n320922 );
buf ( n321063 , n862 );
buf ( n321064 , n884 );
xnor ( n321065 , n321063 , n321064 );
buf ( n321066 , n321065 );
buf ( n321067 , n321066 );
not ( n321068 , n321067 );
buf ( n321069 , n304813 );
nand ( n30644 , n321068 , n321069 );
buf ( n321071 , n30644 );
nand ( n321072 , n30636 , n321071 );
buf ( n321073 , n321072 );
xor ( n321074 , n321061 , n321073 );
buf ( n321075 , n314747 );
buf ( n321076 , n305993 );
buf ( n321077 , n860 );
and ( n30652 , n321076 , n321077 );
buf ( n321079 , n305241 );
buf ( n321080 , n886 );
and ( n321081 , n321079 , n321080 );
nor ( n30656 , n30652 , n321081 );
buf ( n321083 , n30656 );
buf ( n321084 , n321083 );
or ( n321085 , n321075 , n321084 );
buf ( n321086 , n305363 );
buf ( n321087 , n30437 );
or ( n30662 , n321086 , n321087 );
nand ( n321089 , n321085 , n30662 );
buf ( n321090 , n321089 );
buf ( n321091 , n321090 );
and ( n321092 , n321074 , n321091 );
and ( n30667 , n321061 , n321073 );
or ( n30668 , n321092 , n30667 );
buf ( n321095 , n30668 );
buf ( n321096 , n321095 );
xor ( n30671 , n321048 , n321096 );
buf ( n30672 , n14959 );
buf ( n30673 , n305192 );
nor ( n30674 , n30672 , n30673 );
buf ( n321101 , n30674 );
buf ( n321102 , n321101 );
buf ( n321103 , n888 );
buf ( n321104 , n858 );
and ( n321105 , n321103 , n321104 );
not ( n321106 , n321103 );
buf ( n321107 , n305060 );
and ( n321108 , n321106 , n321107 );
nor ( n30683 , n321105 , n321108 );
buf ( n321110 , n30683 );
buf ( n321111 , n321110 );
not ( n321112 , n321111 );
buf ( n321113 , n305138 );
not ( n30688 , n321113 );
or ( n321115 , n321112 , n30688 );
buf ( n321116 , n320832 );
not ( n30691 , n321116 );
buf ( n321118 , n305144 );
nand ( n30693 , n30691 , n321118 );
buf ( n321120 , n30693 );
buf ( n321121 , n321120 );
nand ( n321122 , n321115 , n321121 );
buf ( n321123 , n321122 );
buf ( n321124 , n321123 );
xor ( n321125 , n321102 , n321124 );
buf ( n321126 , n15057 );
buf ( n321127 , n892 );
buf ( n321128 , n26347 );
and ( n321129 , n321127 , n321128 );
not ( n30704 , n321127 );
buf ( n321131 , n854 );
and ( n30706 , n30704 , n321131 );
nor ( n321133 , n321129 , n30706 );
buf ( n321134 , n321133 );
buf ( n321135 , n321134 );
or ( n30710 , n321126 , n321135 );
buf ( n321137 , n305489 );
buf ( n321138 , n30419 );
or ( n321139 , n321137 , n321138 );
nand ( n321140 , n30710 , n321139 );
buf ( n321141 , n321140 );
buf ( n321142 , n321141 );
and ( n321143 , n321125 , n321142 );
and ( n30718 , n321102 , n321124 );
or ( n321145 , n321143 , n30718 );
buf ( n321146 , n321145 );
buf ( n321147 , n321146 );
xor ( n30722 , n30671 , n321147 );
buf ( n321149 , n30722 );
buf ( n321150 , n321149 );
xor ( n30725 , n321061 , n321073 );
xor ( n321152 , n30725 , n321091 );
buf ( n321153 , n321152 );
buf ( n321154 , n321153 );
xor ( n30729 , n321102 , n321124 );
xor ( n321156 , n30729 , n321142 );
buf ( n321157 , n321156 );
buf ( n321158 , n321157 );
xor ( n30733 , n321154 , n321158 );
buf ( n321160 , n320083 );
buf ( n321161 , n312467 );
buf ( n321162 , n857 );
and ( n30737 , n321161 , n321162 );
buf ( n321164 , n305939 );
buf ( n321165 , n890 );
and ( n30740 , n321164 , n321165 );
nor ( n321167 , n30737 , n30740 );
buf ( n321168 , n321167 );
buf ( n321169 , n321168 );
or ( n30744 , n321160 , n321169 );
buf ( n321171 , n304655 );
buf ( n321172 , n312467 );
buf ( n321173 , n856 );
and ( n321174 , n321172 , n321173 );
buf ( n321175 , n15582 );
buf ( n321176 , n890 );
and ( n321177 , n321175 , n321176 );
nor ( n30752 , n321174 , n321177 );
buf ( n321179 , n30752 );
buf ( n321180 , n321179 );
or ( n321181 , n321171 , n321180 );
nand ( n321182 , n30744 , n321181 );
buf ( n321183 , n321182 );
buf ( n321184 , n321183 );
buf ( n321185 , n15804 );
buf ( n321186 , n304827 );
buf ( n321187 , n863 );
and ( n321188 , n321186 , n321187 );
buf ( n321189 , n305192 );
buf ( n321190 , n884 );
and ( n321191 , n321189 , n321190 );
nor ( n321192 , n321188 , n321191 );
buf ( n321193 , n321192 );
buf ( n321194 , n321193 );
or ( n30769 , n321185 , n321194 );
buf ( n321196 , n310909 );
buf ( n321197 , n321066 );
or ( n321198 , n321196 , n321197 );
nand ( n30773 , n30769 , n321198 );
buf ( n30774 , n30773 );
buf ( n321201 , n30774 );
xor ( n30776 , n321184 , n321201 );
buf ( n321203 , n863 );
buf ( n321204 , n885 );
or ( n30779 , n321203 , n321204 );
buf ( n321206 , n886 );
nand ( n321207 , n30779 , n321206 );
buf ( n321208 , n321207 );
buf ( n321209 , n321208 );
buf ( n321210 , n863 );
buf ( n321211 , n885 );
nand ( n321212 , n321210 , n321211 );
buf ( n321213 , n321212 );
buf ( n321214 , n321213 );
buf ( n321215 , n884 );
and ( n321216 , n321209 , n321214 , n321215 );
buf ( n321217 , n321216 );
buf ( n321218 , n321217 );
buf ( n321219 , n15057 );
buf ( n321220 , n892 );
buf ( n321221 , n305319 );
and ( n321222 , n321220 , n321221 );
not ( n321223 , n321220 );
buf ( n321224 , n855 );
and ( n321225 , n321223 , n321224 );
nor ( n321226 , n321222 , n321225 );
buf ( n321227 , n321226 );
buf ( n321228 , n321227 );
or ( n321229 , n321219 , n321228 );
buf ( n321230 , n305489 );
buf ( n321231 , n321134 );
or ( n321232 , n321230 , n321231 );
nand ( n321233 , n321229 , n321232 );
buf ( n321234 , n321233 );
buf ( n321235 , n321234 );
xor ( n321236 , n321218 , n321235 );
buf ( n321237 , n321236 );
buf ( n321238 , n321237 );
and ( n321239 , n30776 , n321238 );
and ( n321240 , n321184 , n321201 );
or ( n321241 , n321239 , n321240 );
buf ( n321242 , n321241 );
buf ( n321243 , n321242 );
and ( n321244 , n30733 , n321243 );
and ( n30819 , n321154 , n321158 );
or ( n321246 , n321244 , n30819 );
buf ( n321247 , n321246 );
buf ( n30822 , n321247 );
xor ( n30823 , n320840 , n320853 );
xor ( n321250 , n30823 , n320871 );
buf ( n321251 , n321250 );
buf ( n321252 , n321251 );
xor ( n321253 , n320899 , n320916 );
xor ( n321254 , n321253 , n320930 );
buf ( n321255 , n321254 );
buf ( n321256 , n321255 );
xor ( n321257 , n321252 , n321256 );
buf ( n321258 , n304630 );
buf ( n321259 , n321179 );
or ( n321260 , n321258 , n321259 );
buf ( n321261 , n304655 );
buf ( n321262 , n320908 );
or ( n321263 , n321261 , n321262 );
nand ( n30838 , n321260 , n321263 );
buf ( n321265 , n30838 );
buf ( n30840 , n321265 );
and ( n321267 , n321218 , n321235 );
buf ( n321268 , n321267 );
buf ( n321269 , n321268 );
xor ( n321270 , n30840 , n321269 );
buf ( n321271 , n305881 );
buf ( n321272 , n853 );
buf ( n321273 , n894 );
xnor ( n30848 , n321272 , n321273 );
buf ( n321275 , n30848 );
buf ( n321276 , n321275 );
or ( n321277 , n321271 , n321276 );
buf ( n321278 , n15469 );
buf ( n321279 , n321053 );
or ( n30854 , n321278 , n321279 );
nand ( n321281 , n321277 , n30854 );
buf ( n321282 , n321281 );
buf ( n321283 , n321282 );
buf ( n321284 , n311275 );
buf ( n321285 , n888 );
buf ( n321286 , n859 );
xnor ( n30861 , n321285 , n321286 );
buf ( n321288 , n30861 );
buf ( n321289 , n321288 );
or ( n30864 , n321284 , n321289 );
buf ( n321291 , n15861 );
buf ( n30866 , n321110 );
not ( n321293 , n30866 );
buf ( n321294 , n321293 );
buf ( n321295 , n321294 );
or ( n321296 , n321291 , n321295 );
nand ( n30871 , n30864 , n321296 );
buf ( n30872 , n30871 );
buf ( n321299 , n30872 );
xor ( n30874 , n321283 , n321299 );
buf ( n321301 , n314747 );
buf ( n321302 , n305993 );
buf ( n321303 , n861 );
and ( n30878 , n321302 , n321303 );
buf ( n321305 , n304771 );
buf ( n321306 , n886 );
and ( n30881 , n321305 , n321306 );
nor ( n30882 , n30878 , n30881 );
buf ( n321309 , n30882 );
buf ( n321310 , n321309 );
or ( n321311 , n321301 , n321310 );
buf ( n321312 , n305363 );
buf ( n321313 , n321083 );
or ( n321314 , n321312 , n321313 );
nand ( n321315 , n321311 , n321314 );
buf ( n321316 , n321315 );
buf ( n30891 , n321316 );
and ( n30892 , n30874 , n30891 );
and ( n321319 , n321283 , n321299 );
or ( n321320 , n30892 , n321319 );
buf ( n321321 , n321320 );
buf ( n321322 , n321321 );
and ( n321323 , n321270 , n321322 );
and ( n30898 , n30840 , n321269 );
or ( n321325 , n321323 , n30898 );
buf ( n321326 , n321325 );
buf ( n321327 , n321326 );
xor ( n321328 , n321257 , n321327 );
buf ( n321329 , n321328 );
buf ( n321330 , n321329 );
xor ( n321331 , n321150 , n30822 );
xor ( n321332 , n321331 , n321330 );
buf ( n321333 , n321332 );
xor ( n321334 , n321150 , n30822 );
and ( n30909 , n321334 , n321330 );
and ( n321336 , n321150 , n30822 );
or ( n321337 , n30909 , n321336 );
buf ( n321338 , n321337 );
xor ( n321339 , n321184 , n321201 );
xor ( n321340 , n321339 , n321238 );
buf ( n321341 , n321340 );
buf ( n321342 , n321341 );
buf ( n321343 , n310909 );
buf ( n321344 , n305192 );
nor ( n30919 , n321343 , n321344 );
buf ( n321346 , n30919 );
buf ( n321347 , n321346 );
buf ( n321348 , n888 );
buf ( n321349 , n305241 );
and ( n30924 , n321348 , n321349 );
not ( n30925 , n321348 );
buf ( n321352 , n860 );
and ( n30927 , n30925 , n321352 );
nor ( n30928 , n30924 , n30927 );
buf ( n321355 , n30928 );
buf ( n321356 , n321355 );
not ( n321357 , n321356 );
buf ( n321358 , n321357 );
buf ( n321359 , n321358 );
not ( n321360 , n321359 );
buf ( n321361 , n305138 );
not ( n30936 , n321361 );
or ( n321363 , n321360 , n30936 );
buf ( n321364 , n321288 );
not ( n30939 , n321364 );
buf ( n321366 , n305144 );
nand ( n30941 , n30939 , n321366 );
buf ( n30942 , n30941 );
buf ( n321369 , n30942 );
nand ( n30944 , n321363 , n321369 );
buf ( n30945 , n30944 );
buf ( n321372 , n30945 );
xor ( n30947 , n321347 , n321372 );
buf ( n321374 , n305561 );
buf ( n321375 , n892 );
buf ( n321376 , n15582 );
and ( n321377 , n321375 , n321376 );
not ( n321378 , n321375 );
buf ( n321379 , n856 );
and ( n30954 , n321378 , n321379 );
nor ( n30955 , n321377 , n30954 );
buf ( n30956 , n30955 );
buf ( n321383 , n30956 );
or ( n30958 , n321374 , n321383 );
buf ( n321385 , n305489 );
buf ( n321386 , n321227 );
or ( n30961 , n321385 , n321386 );
nand ( n30962 , n30958 , n30961 );
buf ( n321389 , n30962 );
buf ( n321390 , n321389 );
xor ( n30965 , n30947 , n321390 );
buf ( n321392 , n30965 );
buf ( n30967 , n321392 );
buf ( n321394 , n863 );
buf ( n321395 , n887 );
or ( n321396 , n321394 , n321395 );
buf ( n321397 , n888 );
nand ( n30972 , n321396 , n321397 );
buf ( n30973 , n30972 );
buf ( n321400 , n30973 );
buf ( n321401 , n863 );
buf ( n321402 , n887 );
nand ( n321403 , n321401 , n321402 );
buf ( n321404 , n321403 );
buf ( n321405 , n321404 );
buf ( n321406 , n886 );
and ( n30981 , n321400 , n321405 , n321406 );
buf ( n30982 , n30981 );
buf ( n30983 , n30982 );
buf ( n321410 , n305561 );
buf ( n321411 , n892 );
buf ( n321412 , n305939 );
and ( n321413 , n321411 , n321412 );
not ( n321414 , n321411 );
buf ( n321415 , n857 );
and ( n321416 , n321414 , n321415 );
nor ( n30991 , n321413 , n321416 );
buf ( n321418 , n30991 );
buf ( n321419 , n321418 );
or ( n30994 , n321410 , n321419 );
buf ( n321421 , n305489 );
buf ( n321422 , n30956 );
or ( n30997 , n321421 , n321422 );
nand ( n321424 , n30994 , n30997 );
buf ( n321425 , n321424 );
buf ( n321426 , n321425 );
and ( n321427 , n30983 , n321426 );
buf ( n321428 , n321427 );
buf ( n321429 , n321428 );
xor ( n321430 , n30967 , n321429 );
buf ( n321431 , n311275 );
buf ( n321432 , n888 );
buf ( n31007 , n304771 );
and ( n31008 , n321432 , n31007 );
not ( n321435 , n321432 );
buf ( n321436 , n861 );
and ( n31011 , n321435 , n321436 );
nor ( n321438 , n31008 , n31011 );
buf ( n321439 , n321438 );
buf ( n321440 , n321439 );
or ( n321441 , n321431 , n321440 );
buf ( n321442 , n305130 );
buf ( n321443 , n321355 );
or ( n321444 , n321442 , n321443 );
nand ( n31019 , n321441 , n321444 );
buf ( n31020 , n31019 );
buf ( n31021 , n31020 );
buf ( n321448 , n305881 );
buf ( n321449 , n894 );
not ( n321450 , n321449 );
buf ( n321451 , n855 );
nor ( n31026 , n321450 , n321451 );
buf ( n321453 , n31026 );
buf ( n321454 , n321453 );
buf ( n321455 , n855 );
not ( n31030 , n321455 );
buf ( n321457 , n894 );
nor ( n31032 , n31030 , n321457 );
buf ( n321459 , n31032 );
buf ( n321460 , n321459 );
nor ( n31035 , n321454 , n321460 );
buf ( n31036 , n31035 );
buf ( n321463 , n31036 );
or ( n31038 , n321448 , n321463 );
buf ( n321465 , n854 );
buf ( n321466 , n894 );
xnor ( n321467 , n321465 , n321466 );
buf ( n321468 , n321467 );
buf ( n321469 , n321468 );
buf ( n321470 , n15469 );
or ( n31045 , n321469 , n321470 );
nand ( n31046 , n31038 , n31045 );
buf ( n321473 , n31046 );
buf ( n321474 , n321473 );
xor ( n321475 , n31021 , n321474 );
buf ( n321476 , n313403 );
buf ( n321477 , n305993 );
buf ( n321478 , n863 );
and ( n31053 , n321477 , n321478 );
buf ( n321480 , n305192 );
buf ( n321481 , n886 );
and ( n31056 , n321480 , n321481 );
nor ( n321483 , n31053 , n31056 );
buf ( n321484 , n321483 );
buf ( n321485 , n321484 );
or ( n321486 , n321476 , n321485 );
buf ( n321487 , n305363 );
buf ( n321488 , n305993 );
buf ( n321489 , n862 );
and ( n31064 , n321488 , n321489 );
buf ( n321491 , n304739 );
buf ( n321492 , n886 );
and ( n321493 , n321491 , n321492 );
nor ( n321494 , n31064 , n321493 );
buf ( n321495 , n321494 );
buf ( n321496 , n321495 );
or ( n31071 , n321487 , n321496 );
nand ( n321498 , n321486 , n31071 );
buf ( n321499 , n321498 );
buf ( n321500 , n321499 );
and ( n31075 , n321475 , n321500 );
and ( n321502 , n31021 , n321474 );
or ( n321503 , n31075 , n321502 );
buf ( n321504 , n321503 );
buf ( n321505 , n321504 );
and ( n31080 , n321430 , n321505 );
and ( n321507 , n30967 , n321429 );
or ( n31082 , n31080 , n321507 );
buf ( n321509 , n31082 );
buf ( n321510 , n321509 );
buf ( n321511 , n305881 );
buf ( n321512 , n321468 );
or ( n321513 , n321511 , n321512 );
buf ( n321514 , n321275 );
buf ( n321515 , n15469 );
or ( n321516 , n321514 , n321515 );
nand ( n31091 , n321513 , n321516 );
buf ( n31092 , n31091 );
buf ( n321519 , n31092 );
buf ( n321520 , n304630 );
buf ( n321521 , n312467 );
buf ( n321522 , n858 );
and ( n31097 , n321521 , n321522 );
buf ( n321524 , n305060 );
buf ( n321525 , n890 );
and ( n321526 , n321524 , n321525 );
nor ( n31101 , n31097 , n321526 );
buf ( n321528 , n31101 );
buf ( n321529 , n321528 );
or ( n31104 , n321520 , n321529 );
buf ( n31105 , n304655 );
buf ( n321532 , n321168 );
or ( n321533 , n31105 , n321532 );
nand ( n321534 , n31104 , n321533 );
buf ( n321535 , n321534 );
buf ( n31110 , n321535 );
xor ( n31111 , n321519 , n31110 );
buf ( n321538 , n314747 );
buf ( n321539 , n321495 );
or ( n31114 , n321538 , n321539 );
buf ( n321541 , n305363 );
buf ( n321542 , n321309 );
or ( n321543 , n321541 , n321542 );
nand ( n31118 , n31114 , n321543 );
buf ( n321545 , n31118 );
buf ( n321546 , n321545 );
and ( n321547 , n31111 , n321546 );
and ( n31122 , n321519 , n31110 );
or ( n31123 , n321547 , n31122 );
buf ( n321550 , n31123 );
buf ( n321551 , n321550 );
xor ( n31126 , n321347 , n321372 );
and ( n321553 , n31126 , n321390 );
and ( n321554 , n321347 , n321372 );
or ( n31129 , n321553 , n321554 );
buf ( n321556 , n31129 );
buf ( n321557 , n321556 );
xor ( n31132 , n321551 , n321557 );
xor ( n321559 , n321283 , n321299 );
xor ( n321560 , n321559 , n30891 );
buf ( n321561 , n321560 );
buf ( n321562 , n321561 );
xor ( n321563 , n31132 , n321562 );
buf ( n321564 , n321563 );
buf ( n321565 , n321564 );
xor ( n321566 , n321342 , n321510 );
xor ( n31141 , n321566 , n321565 );
buf ( n321568 , n31141 );
xor ( n321569 , n321342 , n321510 );
and ( n31144 , n321569 , n321565 );
and ( n321571 , n321342 , n321510 );
or ( n31146 , n31144 , n321571 );
buf ( n321573 , n31146 );
xor ( n31148 , n30096 , n320534 );
and ( n321575 , n31148 , n320541 );
and ( n321576 , n30096 , n320534 );
or ( n31151 , n321575 , n321576 );
buf ( n321578 , n31151 );
buf ( n321579 , n321578 );
buf ( n31154 , n320533 );
not ( n321581 , n31154 );
buf ( n321582 , n321581 );
buf ( n321583 , n321582 );
buf ( n321584 , n842 );
buf ( n321585 , n864 );
and ( n321586 , n321584 , n321585 );
buf ( n321587 , n321586 );
buf ( n321588 , n321587 );
xor ( n321589 , n321583 , n321588 );
xor ( n321590 , n320558 , n320575 );
and ( n31165 , n321590 , n320593 );
and ( n321592 , n320558 , n320575 );
or ( n31167 , n31165 , n321592 );
buf ( n321594 , n31167 );
buf ( n321595 , n321594 );
xor ( n31170 , n321589 , n321595 );
buf ( n321597 , n31170 );
buf ( n321598 , n321597 );
xor ( n31173 , n320596 , n320601 );
and ( n31174 , n31173 , n320645 );
and ( n321601 , n320596 , n320601 );
or ( n31176 , n31174 , n321601 );
buf ( n321603 , n31176 );
buf ( n321604 , n321603 );
xor ( n31179 , n321579 , n321598 );
xor ( n321606 , n31179 , n321604 );
buf ( n321607 , n321606 );
xor ( n31182 , n321579 , n321598 );
and ( n31183 , n31182 , n321604 );
and ( n321610 , n321579 , n321598 );
or ( n31185 , n31183 , n321610 );
buf ( n321612 , n31185 );
xor ( n321613 , n320695 , n320701 );
and ( n31188 , n321613 , n320722 );
and ( n321615 , n320695 , n320701 );
or ( n31190 , n31188 , n321615 );
buf ( n321617 , n31190 );
xor ( n321618 , n30840 , n321269 );
xor ( n321619 , n321618 , n321322 );
buf ( n321620 , n321619 );
buf ( n321621 , n321620 );
xor ( n321622 , n321551 , n321557 );
and ( n31197 , n321622 , n321562 );
and ( n31198 , n321551 , n321557 );
or ( n31199 , n31197 , n31198 );
buf ( n31200 , n31199 );
buf ( n31201 , n31200 );
xor ( n31202 , n321154 , n321158 );
xor ( n321629 , n31202 , n321243 );
buf ( n321630 , n321629 );
buf ( n321631 , n321630 );
xor ( n31206 , n321621 , n31201 );
xor ( n321633 , n31206 , n321631 );
buf ( n321634 , n321633 );
xor ( n321635 , n321621 , n31201 );
and ( n321636 , n321635 , n321631 );
and ( n31211 , n321621 , n31201 );
or ( n321638 , n321636 , n31211 );
buf ( n321639 , n321638 );
buf ( n321640 , n313215 );
buf ( n321641 , n313871 );
buf ( n321642 , n835 );
and ( n321643 , n321641 , n321642 );
buf ( n321644 , n21261 );
buf ( n321645 , n866 );
and ( n321646 , n321644 , n321645 );
nor ( n31221 , n321643 , n321646 );
buf ( n31222 , n31221 );
buf ( n321649 , n31222 );
or ( n31224 , n321640 , n321649 );
buf ( n321651 , n313224 );
buf ( n321652 , n313871 );
buf ( n321653 , n834 );
and ( n321654 , n321652 , n321653 );
buf ( n321655 , n310658 );
buf ( n321656 , n866 );
and ( n31231 , n321655 , n321656 );
nor ( n321658 , n321654 , n31231 );
buf ( n321659 , n321658 );
buf ( n321660 , n321659 );
or ( n31235 , n321651 , n321660 );
nand ( n321662 , n31224 , n31235 );
buf ( n321663 , n321662 );
buf ( n321664 , n321663 );
buf ( n31239 , n838 );
buf ( n31240 , n864 );
and ( n31241 , n31239 , n31240 );
buf ( n321668 , n31241 );
buf ( n321669 , n321668 );
xor ( n321670 , n321664 , n321669 );
buf ( n321671 , n310726 );
buf ( n321672 , n310521 );
buf ( n321673 , n834 );
and ( n321674 , n321672 , n321673 );
buf ( n321675 , n310658 );
buf ( n321676 , n868 );
and ( n321677 , n321675 , n321676 );
nor ( n321678 , n321674 , n321677 );
buf ( n321679 , n321678 );
buf ( n321680 , n321679 );
or ( n321681 , n321671 , n321680 );
buf ( n321682 , n305449 );
buf ( n321683 , n310521 );
buf ( n321684 , n833 );
and ( n321685 , n321683 , n321684 );
buf ( n321686 , n310964 );
buf ( n321687 , n868 );
and ( n31262 , n321686 , n321687 );
nor ( n31263 , n321685 , n31262 );
buf ( n321690 , n31263 );
buf ( n321691 , n321690 );
or ( n31266 , n321682 , n321691 );
nand ( n321693 , n321681 , n31266 );
buf ( n321694 , n321693 );
buf ( n321695 , n321694 );
and ( n321696 , n321670 , n321695 );
and ( n321697 , n321664 , n321669 );
or ( n31272 , n321696 , n321697 );
buf ( n321699 , n31272 );
buf ( n321700 , n321699 );
buf ( n321701 , n311891 );
buf ( n321702 , n311234 );
buf ( n321703 , n837 );
and ( n31278 , n321702 , n321703 );
buf ( n321705 , n313757 );
buf ( n321706 , n864 );
and ( n31281 , n321705 , n321706 );
nor ( n321708 , n31278 , n31281 );
buf ( n321709 , n321708 );
buf ( n321710 , n321709 );
or ( n31285 , n321701 , n321710 );
buf ( n321712 , n311246 );
buf ( n321713 , n311234 );
buf ( n321714 , n836 );
and ( n321715 , n321713 , n321714 );
buf ( n321716 , n311204 );
buf ( n321717 , n864 );
and ( n31292 , n321716 , n321717 );
nor ( n31293 , n321715 , n31292 );
buf ( n321720 , n31293 );
buf ( n321721 , n321720 );
or ( n321722 , n321712 , n321721 );
nand ( n31297 , n31285 , n321722 );
buf ( n31298 , n31297 );
buf ( n31299 , n31298 );
buf ( n321726 , n304763 );
buf ( n321727 , n14323 );
or ( n321728 , n321726 , n321727 );
buf ( n321729 , n870 );
nand ( n31304 , n321728 , n321729 );
buf ( n321731 , n31304 );
buf ( n321732 , n321731 );
xor ( n31307 , n31299 , n321732 );
buf ( n321734 , n310726 );
buf ( n321735 , n321690 );
or ( n31310 , n321734 , n321735 );
buf ( n321737 , n305449 );
buf ( n321738 , n310521 );
buf ( n321739 , n832 );
and ( n321740 , n321738 , n321739 );
buf ( n321741 , n20700 );
buf ( n321742 , n868 );
and ( n321743 , n321741 , n321742 );
nor ( n321744 , n321740 , n321743 );
buf ( n321745 , n321744 );
buf ( n321746 , n321745 );
or ( n321747 , n321737 , n321746 );
nand ( n321748 , n31310 , n321747 );
buf ( n321749 , n321748 );
buf ( n31324 , n321749 );
and ( n31325 , n31307 , n31324 );
and ( n31326 , n31299 , n321732 );
or ( n31327 , n31325 , n31326 );
buf ( n31328 , n31327 );
buf ( n31329 , n31328 );
buf ( n321756 , n310726 );
buf ( n321757 , n321745 );
or ( n321758 , n321756 , n321757 );
buf ( n321759 , n305449 );
buf ( n321760 , n310521 );
or ( n321761 , n321759 , n321760 );
nand ( n321762 , n321758 , n321761 );
buf ( n321763 , n321762 );
buf ( n321764 , n321763 );
not ( n31339 , n321764 );
buf ( n321766 , n31339 );
buf ( n321767 , n321766 );
xor ( n31342 , n31329 , n321767 );
buf ( n321769 , n313215 );
buf ( n321770 , n321659 );
or ( n321771 , n321769 , n321770 );
buf ( n321772 , n313224 );
buf ( n321773 , n313871 );
buf ( n321774 , n833 );
and ( n321775 , n321773 , n321774 );
buf ( n321776 , n310964 );
buf ( n321777 , n866 );
and ( n321778 , n321776 , n321777 );
nor ( n31353 , n321775 , n321778 );
buf ( n31354 , n31353 );
buf ( n321781 , n31354 );
or ( n321782 , n321772 , n321781 );
nand ( n321783 , n321771 , n321782 );
buf ( n321784 , n321783 );
buf ( n321785 , n321784 );
buf ( n321786 , n837 );
buf ( n321787 , n864 );
and ( n31362 , n321786 , n321787 );
buf ( n321789 , n31362 );
buf ( n321790 , n321789 );
xor ( n31365 , n321785 , n321790 );
buf ( n321792 , n311891 );
buf ( n321793 , n321720 );
or ( n321794 , n321792 , n321793 );
buf ( n321795 , n311246 );
buf ( n321796 , n311234 );
buf ( n321797 , n835 );
and ( n31372 , n321796 , n321797 );
buf ( n321799 , n21261 );
buf ( n321800 , n864 );
and ( n31375 , n321799 , n321800 );
nor ( n321802 , n31372 , n31375 );
buf ( n321803 , n321802 );
buf ( n321804 , n321803 );
or ( n321805 , n321795 , n321804 );
nand ( n31380 , n321794 , n321805 );
buf ( n321807 , n31380 );
buf ( n321808 , n321807 );
xor ( n31383 , n31365 , n321808 );
buf ( n321810 , n31383 );
buf ( n321811 , n321810 );
xor ( n31386 , n31342 , n321811 );
buf ( n321813 , n31386 );
buf ( n321814 , n321813 );
xor ( n31389 , n321664 , n321669 );
xor ( n31390 , n31389 , n321695 );
buf ( n321817 , n31390 );
buf ( n321818 , n321817 );
buf ( n321819 , n315120 );
buf ( n321820 , n319815 );
buf ( n321821 , n832 );
and ( n321822 , n321820 , n321821 );
buf ( n321823 , n20700 );
buf ( n321824 , n870 );
and ( n321825 , n321823 , n321824 );
nor ( n31400 , n321822 , n321825 );
buf ( n321827 , n31400 );
buf ( n321828 , n321827 );
or ( n31403 , n321819 , n321828 );
buf ( n321830 , n304760 );
buf ( n321831 , n319815 );
or ( n321832 , n321830 , n321831 );
nand ( n31407 , n31403 , n321832 );
buf ( n321834 , n31407 );
buf ( n321835 , n321834 );
buf ( n321836 , n839 );
buf ( n321837 , n864 );
and ( n321838 , n321836 , n321837 );
buf ( n321839 , n321838 );
buf ( n321840 , n321839 );
xor ( n321841 , n321835 , n321840 );
buf ( n321842 , n311891 );
buf ( n321843 , n311234 );
buf ( n321844 , n838 );
and ( n31419 , n321843 , n321844 );
buf ( n321846 , n310377 );
buf ( n321847 , n864 );
and ( n31422 , n321846 , n321847 );
nor ( n321849 , n31419 , n31422 );
buf ( n321850 , n321849 );
buf ( n321851 , n321850 );
or ( n31426 , n321842 , n321851 );
buf ( n321853 , n311246 );
buf ( n321854 , n321709 );
or ( n321855 , n321853 , n321854 );
nand ( n321856 , n31426 , n321855 );
buf ( n321857 , n321856 );
buf ( n321858 , n321857 );
and ( n321859 , n321841 , n321858 );
and ( n31434 , n321835 , n321840 );
or ( n321861 , n321859 , n31434 );
buf ( n321862 , n321861 );
buf ( n321863 , n321862 );
xor ( n321864 , n321818 , n321863 );
xor ( n31439 , n31299 , n321732 );
xor ( n321866 , n31439 , n31324 );
buf ( n321867 , n321866 );
buf ( n321868 , n321867 );
and ( n321869 , n321864 , n321868 );
and ( n321870 , n321818 , n321863 );
or ( n31445 , n321869 , n321870 );
buf ( n321872 , n31445 );
buf ( n321873 , n321872 );
xor ( n321874 , n321700 , n321814 );
xor ( n31449 , n321874 , n321873 );
buf ( n321876 , n31449 );
xor ( n321877 , n321700 , n321814 );
and ( n31452 , n321877 , n321873 );
and ( n321879 , n321700 , n321814 );
or ( n321880 , n31452 , n321879 );
buf ( n321881 , n321880 );
buf ( n321882 , n321694 );
not ( n321883 , n321882 );
buf ( n321884 , n321883 );
buf ( n321885 , n321884 );
buf ( n321886 , n310691 );
buf ( n321887 , n313871 );
buf ( n321888 , n836 );
and ( n31463 , n321887 , n321888 );
buf ( n321890 , n311204 );
buf ( n321891 , n866 );
and ( n31466 , n321890 , n321891 );
nor ( n321893 , n31463 , n31466 );
buf ( n321894 , n321893 );
buf ( n321895 , n321894 );
or ( n31470 , n321886 , n321895 );
buf ( n321897 , n310472 );
buf ( n321898 , n31222 );
or ( n31473 , n321897 , n321898 );
nand ( n321900 , n31470 , n31473 );
buf ( n321901 , n321900 );
buf ( n31476 , n321901 );
xor ( n31477 , n321885 , n31476 );
buf ( n321904 , n311891 );
buf ( n321905 , n864 );
buf ( n321906 , n839 );
xnor ( n321907 , n321905 , n321906 );
buf ( n321908 , n321907 );
buf ( n321909 , n321908 );
or ( n31484 , n321904 , n321909 );
buf ( n321911 , n311246 );
buf ( n321912 , n321850 );
or ( n321913 , n321911 , n321912 );
nand ( n321914 , n31484 , n321913 );
buf ( n321915 , n321914 );
buf ( n321916 , n321915 );
buf ( n321917 , n864 );
buf ( n321918 , n840 );
and ( n321919 , n321917 , n321918 );
buf ( n321920 , n321919 );
buf ( n321921 , n321920 );
xor ( n321922 , n321916 , n321921 );
buf ( n321923 , n310726 );
buf ( n321924 , n310521 );
buf ( n321925 , n835 );
and ( n31500 , n321924 , n321925 );
buf ( n321927 , n21261 );
buf ( n321928 , n868 );
and ( n31503 , n321927 , n321928 );
nor ( n321930 , n31500 , n31503 );
buf ( n321931 , n321930 );
buf ( n321932 , n321931 );
or ( n321933 , n321923 , n321932 );
buf ( n321934 , n305449 );
buf ( n321935 , n321679 );
or ( n321936 , n321934 , n321935 );
nand ( n31511 , n321933 , n321936 );
buf ( n31512 , n31511 );
buf ( n321939 , n31512 );
and ( n31514 , n321922 , n321939 );
and ( n321941 , n321916 , n321921 );
or ( n321942 , n31514 , n321941 );
buf ( n321943 , n321942 );
buf ( n321944 , n321943 );
and ( n31519 , n31477 , n321944 );
and ( n321946 , n321885 , n31476 );
or ( n321947 , n31519 , n321946 );
buf ( n321948 , n321947 );
buf ( n321949 , n321948 );
xor ( n321950 , n321818 , n321863 );
xor ( n31525 , n321950 , n321868 );
buf ( n321952 , n31525 );
buf ( n321953 , n321952 );
buf ( n321954 , n310691 );
buf ( n321955 , n313871 );
buf ( n321956 , n837 );
and ( n321957 , n321955 , n321956 );
buf ( n321958 , n313757 );
buf ( n321959 , n866 );
and ( n321960 , n321958 , n321959 );
nor ( n31535 , n321957 , n321960 );
buf ( n31536 , n31535 );
buf ( n321963 , n31536 );
or ( n321964 , n321954 , n321963 );
buf ( n321965 , n313224 );
buf ( n321966 , n321894 );
or ( n31541 , n321965 , n321966 );
nand ( n31542 , n321964 , n31541 );
buf ( n321969 , n31542 );
buf ( n321970 , n315120 );
buf ( n321971 , n319815 );
buf ( n321972 , n833 );
and ( n31547 , n321971 , n321972 );
buf ( n321974 , n310964 );
buf ( n321975 , n870 );
and ( n31550 , n321974 , n321975 );
nor ( n321977 , n31547 , n31550 );
buf ( n321978 , n321977 );
buf ( n321979 , n321978 );
or ( n321980 , n321970 , n321979 );
buf ( n321981 , n304760 );
buf ( n321982 , n321827 );
or ( n321983 , n321981 , n321982 );
nand ( n321984 , n321980 , n321983 );
buf ( n321985 , n321984 );
xor ( n321986 , n321969 , n321985 );
buf ( n321987 , n304851 );
buf ( n321988 , n304845 );
or ( n321989 , n321987 , n321988 );
buf ( n321990 , n872 );
nand ( n31565 , n321989 , n321990 );
buf ( n31566 , n31565 );
and ( n321993 , n321986 , n31566 );
and ( n321994 , n321969 , n321985 );
or ( n31569 , n321993 , n321994 );
buf ( n321996 , n31569 );
xor ( n321997 , n321835 , n321840 );
xor ( n321998 , n321997 , n321858 );
buf ( n321999 , n321998 );
buf ( n322000 , n321999 );
xor ( n322001 , n321996 , n322000 );
xor ( n322002 , n321885 , n31476 );
xor ( n31577 , n322002 , n321944 );
buf ( n322004 , n31577 );
buf ( n322005 , n322004 );
and ( n31580 , n322001 , n322005 );
and ( n322007 , n321996 , n322000 );
or ( n322008 , n31580 , n322007 );
buf ( n322009 , n322008 );
buf ( n322010 , n322009 );
xor ( n31585 , n321949 , n321953 );
xor ( n31586 , n31585 , n322010 );
buf ( n322013 , n31586 );
xor ( n31588 , n321949 , n321953 );
and ( n322015 , n31588 , n322010 );
and ( n31590 , n321949 , n321953 );
or ( n322017 , n322015 , n31590 );
buf ( n322018 , n322017 );
xor ( n31593 , n320516 , n320544 );
and ( n322020 , n31593 , n320648 );
and ( n322021 , n320516 , n320544 );
or ( n31596 , n322020 , n322021 );
buf ( n322023 , n31596 );
xor ( n322024 , n312121 , n312252 );
xor ( n31599 , n322024 , n312257 );
buf ( n322026 , n31599 );
xor ( n322027 , n320677 , n320681 );
and ( n31602 , n322027 , n320688 );
and ( n31603 , n320677 , n320681 );
or ( n322030 , n31602 , n31603 );
buf ( n322031 , n322030 );
xor ( n31606 , n321519 , n31110 );
xor ( n322033 , n31606 , n321546 );
buf ( n322034 , n322033 );
buf ( n322035 , n322034 );
buf ( n322036 , n305881 );
buf ( n322037 , n856 );
buf ( n322038 , n894 );
xnor ( n322039 , n322037 , n322038 );
buf ( n322040 , n322039 );
buf ( n322041 , n322040 );
or ( n322042 , n322036 , n322041 );
buf ( n322043 , n31036 );
buf ( n322044 , n15469 );
or ( n322045 , n322043 , n322044 );
nand ( n31620 , n322042 , n322045 );
buf ( n322047 , n31620 );
buf ( n322048 , n322047 );
buf ( n31623 , n305363 );
buf ( n322050 , n305192 );
nor ( n322051 , n31623 , n322050 );
buf ( n322052 , n322051 );
buf ( n322053 , n322052 );
xor ( n31628 , n322048 , n322053 );
buf ( n322055 , n305135 );
buf ( n322056 , n888 );
not ( n31631 , n322056 );
buf ( n322058 , n31631 );
buf ( n322059 , n322058 );
buf ( n322060 , n862 );
and ( n31635 , n322059 , n322060 );
buf ( n322062 , n304739 );
buf ( n322063 , n888 );
and ( n322064 , n322062 , n322063 );
nor ( n322065 , n31635 , n322064 );
buf ( n322066 , n322065 );
buf ( n322067 , n322066 );
or ( n322068 , n322055 , n322067 );
buf ( n322069 , n15861 );
buf ( n322070 , n321439 );
or ( n31645 , n322069 , n322070 );
nand ( n322072 , n322068 , n31645 );
buf ( n322073 , n322072 );
buf ( n322074 , n322073 );
and ( n322075 , n31628 , n322074 );
and ( n322076 , n322048 , n322053 );
or ( n31651 , n322075 , n322076 );
buf ( n322078 , n31651 );
buf ( n322079 , n322078 );
buf ( n322080 , n304630 );
buf ( n322081 , n312467 );
buf ( n322082 , n859 );
and ( n322083 , n322081 , n322082 );
buf ( n322084 , n14447 );
buf ( n322085 , n890 );
and ( n322086 , n322084 , n322085 );
nor ( n322087 , n322083 , n322086 );
buf ( n322088 , n322087 );
buf ( n322089 , n322088 );
or ( n322090 , n322080 , n322089 );
buf ( n322091 , n304655 );
buf ( n322092 , n321528 );
or ( n322093 , n322091 , n322092 );
nand ( n322094 , n322090 , n322093 );
buf ( n322095 , n322094 );
buf ( n322096 , n322095 );
xor ( n322097 , n322079 , n322096 );
xor ( n31672 , n30983 , n321426 );
buf ( n322099 , n31672 );
buf ( n322100 , n322099 );
and ( n322101 , n322097 , n322100 );
and ( n322102 , n322079 , n322096 );
or ( n31677 , n322101 , n322102 );
buf ( n322104 , n31677 );
buf ( n322105 , n322104 );
xor ( n31680 , n30967 , n321429 );
xor ( n322107 , n31680 , n321505 );
buf ( n322108 , n322107 );
buf ( n322109 , n322108 );
xor ( n322110 , n322035 , n322105 );
xor ( n322111 , n322110 , n322109 );
buf ( n322112 , n322111 );
xor ( n322113 , n322035 , n322105 );
and ( n322114 , n322113 , n322109 );
and ( n31689 , n322035 , n322105 );
or ( n322116 , n322114 , n31689 );
buf ( n322117 , n322116 );
xor ( n31692 , n320747 , n320822 );
xor ( n322119 , n31692 , n320940 );
buf ( n322120 , n322119 );
xor ( n322121 , n321583 , n321588 );
and ( n322122 , n322121 , n321595 );
and ( n31697 , n321583 , n321588 );
or ( n322124 , n322122 , n31697 );
buf ( n322125 , n322124 );
buf ( n322126 , n322125 );
buf ( n322127 , n315120 );
buf ( n322128 , n319815 );
buf ( n322129 , n834 );
and ( n322130 , n322128 , n322129 );
buf ( n322131 , n310658 );
buf ( n322132 , n870 );
and ( n31707 , n322131 , n322132 );
nor ( n322134 , n322130 , n31707 );
buf ( n322135 , n322134 );
buf ( n322136 , n322135 );
or ( n322137 , n322127 , n322136 );
buf ( n322138 , n304760 );
buf ( n322139 , n321978 );
or ( n31714 , n322138 , n322139 );
nand ( n31715 , n322137 , n31714 );
buf ( n322142 , n31715 );
buf ( n322143 , n322142 );
not ( n322144 , n322143 );
buf ( n322145 , n322144 );
buf ( n322146 , n322145 );
buf ( n322147 , n841 );
buf ( n322148 , n864 );
and ( n31723 , n322147 , n322148 );
buf ( n322150 , n31723 );
buf ( n322151 , n322150 );
xor ( n31726 , n322146 , n322151 );
buf ( n322153 , n310726 );
buf ( n322154 , n310521 );
buf ( n322155 , n836 );
and ( n31730 , n322154 , n322155 );
buf ( n322157 , n311204 );
buf ( n322158 , n868 );
and ( n31733 , n322157 , n322158 );
nor ( n322160 , n31730 , n31733 );
buf ( n322161 , n322160 );
buf ( n322162 , n322161 );
or ( n31737 , n322153 , n322162 );
buf ( n322164 , n305449 );
buf ( n322165 , n321931 );
or ( n31740 , n322164 , n322165 );
nand ( n322167 , n31737 , n31740 );
buf ( n322168 , n322167 );
buf ( n322169 , n322168 );
xor ( n322170 , n31726 , n322169 );
buf ( n322171 , n322170 );
buf ( n31746 , n322171 );
xor ( n31747 , n320607 , n320624 );
and ( n322174 , n31747 , n320642 );
and ( n322175 , n320607 , n320624 );
or ( n31750 , n322174 , n322175 );
buf ( n322177 , n31750 );
buf ( n322178 , n305627 );
buf ( n322179 , n305289 );
or ( n322180 , n322178 , n322179 );
buf ( n322181 , n874 );
nand ( n31756 , n322180 , n322181 );
buf ( n322183 , n31756 );
buf ( n322184 , n304854 );
buf ( n322185 , n320570 );
or ( n322186 , n322184 , n322185 );
buf ( n322187 , n14439 );
buf ( n322188 , n872 );
buf ( n322189 , n832 );
and ( n31764 , n322188 , n322189 );
not ( n31765 , n322188 );
buf ( n322192 , n20700 );
and ( n322193 , n31765 , n322192 );
nor ( n31768 , n31764 , n322193 );
buf ( n31769 , n31768 );
buf ( n322196 , n31769 );
not ( n31771 , n322196 );
buf ( n31772 , n31771 );
buf ( n322199 , n31772 );
or ( n31774 , n322187 , n322199 );
nand ( n322201 , n322186 , n31774 );
buf ( n322202 , n322201 );
xor ( n31777 , n322183 , n322202 );
buf ( n322204 , n310726 );
buf ( n322205 , n320588 );
or ( n31780 , n322204 , n322205 );
buf ( n322207 , n305449 );
buf ( n322208 , n322161 );
or ( n31783 , n322207 , n322208 );
nand ( n322210 , n31780 , n31783 );
buf ( n322211 , n322210 );
xor ( n31786 , n31777 , n322211 );
and ( n31787 , n322177 , n31786 );
buf ( n322214 , n310691 );
buf ( n322215 , n320553 );
or ( n322216 , n322214 , n322215 );
buf ( n322217 , n313224 );
buf ( n322218 , n313871 );
buf ( n322219 , n838 );
and ( n31794 , n322218 , n322219 );
buf ( n322221 , n310377 );
buf ( n322222 , n866 );
and ( n322223 , n322221 , n322222 );
nor ( n31798 , n31794 , n322223 );
buf ( n322225 , n31798 );
buf ( n322226 , n322225 );
or ( n322227 , n322217 , n322226 );
nand ( n322228 , n322216 , n322227 );
buf ( n322229 , n322228 );
buf ( n322230 , n322229 );
buf ( n322231 , n315120 );
buf ( n322232 , n320619 );
or ( n31807 , n322231 , n322232 );
buf ( n322234 , n304760 );
buf ( n322235 , n322135 );
or ( n31810 , n322234 , n322235 );
nand ( n322237 , n31807 , n31810 );
buf ( n322238 , n322237 );
buf ( n322239 , n322238 );
xor ( n31814 , n322230 , n322239 );
xor ( n31815 , n321917 , n321918 );
buf ( n322242 , n31815 );
buf ( n322243 , n322242 );
not ( n31818 , n322243 );
buf ( n322245 , n310582 );
not ( n322246 , n322245 );
or ( n31821 , n31818 , n322246 );
buf ( n322248 , n311891 );
buf ( n322249 , n320637 );
or ( n31824 , n322248 , n322249 );
nand ( n322251 , n31821 , n31824 );
buf ( n322252 , n322251 );
buf ( n322253 , n322252 );
xor ( n322254 , n31814 , n322253 );
buf ( n322255 , n322254 );
xor ( n322256 , n322183 , n322202 );
xor ( n31831 , n322256 , n322211 );
and ( n322258 , n322255 , n31831 );
and ( n322259 , n322177 , n322255 );
or ( n322260 , n31787 , n322258 , n322259 );
buf ( n322261 , n322260 );
xor ( n322262 , n322126 , n31746 );
xor ( n31837 , n322262 , n322261 );
buf ( n322264 , n31837 );
xor ( n322265 , n322126 , n31746 );
and ( n31840 , n322265 , n322261 );
and ( n31841 , n322126 , n31746 );
or ( n31842 , n31840 , n31841 );
buf ( n322269 , n31842 );
xor ( n31844 , n320431 , n320448 );
xor ( n31845 , n31844 , n320469 );
buf ( n322272 , n31845 );
buf ( n322273 , n322272 );
xor ( n322274 , n320786 , n320799 );
xor ( n31849 , n322274 , n320817 );
buf ( n322276 , n31849 );
buf ( n322277 , n322276 );
xor ( n31852 , n321048 , n321096 );
and ( n31853 , n31852 , n321147 );
and ( n31854 , n321048 , n321096 );
or ( n31855 , n31853 , n31854 );
buf ( n322282 , n31855 );
buf ( n322283 , n322282 );
xor ( n31858 , n322273 , n322277 );
xor ( n322285 , n31858 , n322283 );
buf ( n322286 , n322285 );
xor ( n31861 , n322273 , n322277 );
and ( n322288 , n31861 , n322283 );
and ( n31863 , n322273 , n322277 );
or ( n31864 , n322288 , n31863 );
buf ( n322291 , n31864 );
xor ( n31866 , n322183 , n322202 );
and ( n31867 , n31866 , n322211 );
and ( n31868 , n322183 , n322202 );
or ( n31869 , n31867 , n31868 );
buf ( n322296 , n31869 );
xor ( n31871 , n322230 , n322239 );
and ( n322298 , n31871 , n322253 );
and ( n31873 , n322230 , n322239 );
or ( n322300 , n322298 , n31873 );
buf ( n322301 , n322300 );
buf ( n322302 , n322301 );
buf ( n322303 , n322242 );
not ( n31878 , n322303 );
buf ( n322305 , n311888 );
not ( n322306 , n322305 );
or ( n31881 , n31878 , n322306 );
buf ( n322308 , n321908 );
not ( n322309 , n322308 );
buf ( n322310 , n310582 );
nand ( n322311 , n322309 , n322310 );
buf ( n322312 , n322311 );
buf ( n322313 , n322312 );
nand ( n322314 , n31881 , n322313 );
buf ( n322315 , n322314 );
buf ( n31890 , n322315 );
buf ( n322317 , n31769 );
not ( n322318 , n322317 );
buf ( n322319 , n304851 );
not ( n322320 , n322319 );
or ( n31895 , n322318 , n322320 );
buf ( n322322 , n304845 );
buf ( n31897 , n872 );
nand ( n31898 , n322322 , n31897 );
buf ( n31899 , n31898 );
buf ( n322326 , n31899 );
nand ( n31901 , n31895 , n322326 );
buf ( n31902 , n31901 );
buf ( n31903 , n31902 );
xor ( n31904 , n31890 , n31903 );
buf ( n322331 , n310691 );
buf ( n322332 , n322225 );
or ( n31907 , n322331 , n322332 );
buf ( n322334 , n310472 );
buf ( n322335 , n31536 );
or ( n31910 , n322334 , n322335 );
nand ( n31911 , n31907 , n31910 );
buf ( n322338 , n31911 );
buf ( n322339 , n322338 );
xor ( n31914 , n31904 , n322339 );
buf ( n322341 , n31914 );
buf ( n322342 , n322341 );
xor ( n322343 , n322296 , n322302 );
xor ( n322344 , n322343 , n322342 );
buf ( n322345 , n322344 );
xor ( n31920 , n322296 , n322302 );
and ( n322347 , n31920 , n322342 );
and ( n322348 , n322296 , n322302 );
or ( n31923 , n322347 , n322348 );
buf ( n322350 , n31923 );
xor ( n322351 , n321996 , n322000 );
xor ( n31926 , n322351 , n322005 );
buf ( n322353 , n31926 );
xor ( n322354 , n321252 , n321256 );
and ( n31929 , n322354 , n321327 );
and ( n31930 , n321252 , n321256 );
or ( n322357 , n31929 , n31930 );
buf ( n322358 , n322357 );
buf ( n322359 , n304630 );
buf ( n322360 , n312467 );
buf ( n322361 , n860 );
and ( n322362 , n322360 , n322361 );
buf ( n322363 , n305241 );
buf ( n322364 , n890 );
and ( n322365 , n322363 , n322364 );
nor ( n31940 , n322362 , n322365 );
buf ( n31941 , n31940 );
buf ( n322368 , n31941 );
or ( n322369 , n322359 , n322368 );
buf ( n322370 , n304655 );
buf ( n322371 , n322088 );
or ( n322372 , n322370 , n322371 );
nand ( n322373 , n322369 , n322372 );
buf ( n322374 , n322373 );
buf ( n322375 , n322374 );
buf ( n322376 , n305561 );
buf ( n322377 , n892 );
buf ( n322378 , n305060 );
and ( n322379 , n322377 , n322378 );
not ( n31954 , n322377 );
buf ( n322381 , n858 );
and ( n322382 , n31954 , n322381 );
nor ( n31957 , n322379 , n322382 );
buf ( n322384 , n31957 );
buf ( n322385 , n322384 );
or ( n31960 , n322376 , n322385 );
buf ( n322387 , n305489 );
buf ( n322388 , n321418 );
or ( n322389 , n322387 , n322388 );
nand ( n31964 , n31960 , n322389 );
buf ( n31965 , n31964 );
buf ( n322392 , n31965 );
xor ( n31967 , n322375 , n322392 );
buf ( n322394 , n863 );
buf ( n322395 , n889 );
or ( n31970 , n322394 , n322395 );
buf ( n322397 , n890 );
nand ( n31972 , n31970 , n322397 );
buf ( n322399 , n31972 );
buf ( n322400 , n322399 );
buf ( n322401 , n863 );
buf ( n322402 , n889 );
nand ( n31977 , n322401 , n322402 );
buf ( n322404 , n31977 );
buf ( n322405 , n322404 );
buf ( n322406 , n888 );
and ( n31981 , n322400 , n322405 , n322406 );
buf ( n322408 , n31981 );
buf ( n31983 , n322408 );
buf ( n322410 , n305881 );
buf ( n322411 , n894 );
not ( n322412 , n322411 );
buf ( n322413 , n857 );
nor ( n322414 , n322412 , n322413 );
buf ( n322415 , n322414 );
buf ( n322416 , n322415 );
buf ( n322417 , n857 );
not ( n31992 , n322417 );
buf ( n322419 , n894 );
nor ( n31994 , n31992 , n322419 );
buf ( n31995 , n31994 );
buf ( n322422 , n31995 );
nor ( n322423 , n322416 , n322422 );
buf ( n322424 , n322423 );
buf ( n322425 , n322424 );
or ( n322426 , n322410 , n322425 );
buf ( n322427 , n322040 );
buf ( n322428 , n15469 );
or ( n322429 , n322427 , n322428 );
nand ( n32004 , n322426 , n322429 );
buf ( n322431 , n32004 );
buf ( n322432 , n322431 );
and ( n32007 , n31983 , n322432 );
buf ( n322434 , n32007 );
buf ( n322435 , n322434 );
and ( n32010 , n31967 , n322435 );
and ( n322437 , n322375 , n322392 );
or ( n32012 , n32010 , n322437 );
buf ( n322439 , n32012 );
buf ( n322440 , n322439 );
xor ( n32015 , n31021 , n321474 );
xor ( n322442 , n32015 , n321500 );
buf ( n322443 , n322442 );
buf ( n322444 , n322443 );
xor ( n322445 , n322079 , n322096 );
xor ( n32020 , n322445 , n322100 );
buf ( n322447 , n32020 );
buf ( n322448 , n322447 );
xor ( n32023 , n322440 , n322444 );
xor ( n322450 , n32023 , n322448 );
buf ( n322451 , n322450 );
xor ( n32026 , n322440 , n322444 );
and ( n322453 , n32026 , n322448 );
and ( n322454 , n322440 , n322444 );
or ( n32029 , n322453 , n322454 );
buf ( n322456 , n32029 );
xor ( n322457 , n320414 , n320474 );
xor ( n32032 , n322457 , n320479 );
buf ( n322459 , n32032 );
buf ( n322460 , n310694 );
buf ( n322461 , n313871 );
buf ( n322462 , n832 );
and ( n322463 , n322461 , n322462 );
buf ( n322464 , n20700 );
buf ( n322465 , n866 );
and ( n322466 , n322464 , n322465 );
nor ( n322467 , n322463 , n322466 );
buf ( n322468 , n322467 );
buf ( n322469 , n322468 );
not ( n322470 , n322469 );
buf ( n322471 , n322470 );
buf ( n322472 , n322471 );
and ( n32047 , n322460 , n322472 );
buf ( n322474 , n311107 );
buf ( n322475 , n866 );
and ( n322476 , n322474 , n322475 );
nor ( n322477 , n32047 , n322476 );
buf ( n322478 , n322477 );
buf ( n322479 , n322478 );
buf ( n322480 , n311234 );
buf ( n322481 , n21261 );
nor ( n32056 , n322480 , n322481 );
buf ( n322483 , n32056 );
buf ( n322484 , n322483 );
xor ( n32059 , n322479 , n322484 );
buf ( n322486 , n311234 );
buf ( n322487 , n833 );
and ( n32062 , n322486 , n322487 );
buf ( n322489 , n310964 );
buf ( n322490 , n864 );
and ( n32065 , n322489 , n322490 );
nor ( n322492 , n32062 , n32065 );
buf ( n322493 , n322492 );
buf ( n322494 , n322493 );
not ( n322495 , n322494 );
buf ( n322496 , n322495 );
buf ( n322497 , n322496 );
not ( n322498 , n322497 );
buf ( n322499 , n310582 );
not ( n32074 , n322499 );
or ( n322501 , n322498 , n32074 );
buf ( n322502 , n311891 );
buf ( n322503 , n311234 );
buf ( n322504 , n834 );
and ( n32079 , n322503 , n322504 );
buf ( n322506 , n310658 );
buf ( n322507 , n864 );
and ( n32082 , n322506 , n322507 );
nor ( n322509 , n32079 , n32082 );
buf ( n322510 , n322509 );
buf ( n322511 , n322510 );
or ( n322512 , n322502 , n322511 );
nand ( n32087 , n322501 , n322512 );
buf ( n32088 , n32087 );
buf ( n322515 , n32088 );
xor ( n32090 , n32059 , n322515 );
buf ( n322517 , n32090 );
buf ( n322518 , n322517 );
buf ( n322519 , n310691 );
buf ( n322520 , n31354 );
or ( n322521 , n322519 , n322520 );
buf ( n322522 , n313224 );
buf ( n322523 , n322468 );
or ( n322524 , n322522 , n322523 );
nand ( n322525 , n322521 , n322524 );
buf ( n322526 , n322525 );
buf ( n322527 , n311234 );
buf ( n322528 , n311204 );
nor ( n322529 , n322527 , n322528 );
buf ( n322530 , n322529 );
xor ( n322531 , n322526 , n322530 );
buf ( n322532 , n305213 );
buf ( n322533 , n305219 );
or ( n32108 , n322532 , n322533 );
buf ( n322535 , n868 );
nand ( n322536 , n32108 , n322535 );
buf ( n322537 , n322536 );
and ( n32112 , n322531 , n322537 );
and ( n322539 , n322526 , n322530 );
or ( n32114 , n32112 , n322539 );
buf ( n322541 , n32114 );
buf ( n322542 , n321763 );
buf ( n322543 , n311891 );
buf ( n322544 , n321803 );
or ( n32119 , n322543 , n322544 );
buf ( n322546 , n311246 );
buf ( n322547 , n322510 );
or ( n32122 , n322546 , n322547 );
nand ( n32123 , n32119 , n32122 );
buf ( n322550 , n32123 );
buf ( n322551 , n322550 );
xor ( n322552 , n322542 , n322551 );
xor ( n32127 , n321785 , n321790 );
and ( n322554 , n32127 , n321808 );
and ( n322555 , n321785 , n321790 );
or ( n322556 , n322554 , n322555 );
buf ( n322557 , n322556 );
buf ( n322558 , n322557 );
and ( n322559 , n322552 , n322558 );
and ( n32134 , n322542 , n322551 );
or ( n322561 , n322559 , n32134 );
buf ( n322562 , n322561 );
buf ( n322563 , n322562 );
xor ( n322564 , n322518 , n322541 );
xor ( n32139 , n322564 , n322563 );
buf ( n322566 , n32139 );
xor ( n32141 , n322518 , n322541 );
and ( n32142 , n32141 , n322563 );
and ( n322569 , n322518 , n322541 );
or ( n322570 , n32142 , n322569 );
buf ( n322571 , n322570 );
xor ( n322572 , n31329 , n321767 );
and ( n322573 , n322572 , n321811 );
and ( n32148 , n31329 , n321767 );
or ( n322575 , n322573 , n32148 );
buf ( n322576 , n322575 );
xor ( n322577 , n320827 , n320876 );
xor ( n32152 , n322577 , n320935 );
buf ( n322579 , n32152 );
xor ( n322580 , n322479 , n322484 );
and ( n32155 , n322580 , n322515 );
and ( n322582 , n322479 , n322484 );
or ( n32157 , n32155 , n322582 );
buf ( n322584 , n32157 );
buf ( n322585 , n322584 );
buf ( n322586 , n322478 );
not ( n32161 , n322586 );
buf ( n322588 , n32161 );
buf ( n322589 , n322588 );
buf ( n322590 , n310694 );
buf ( n322591 , n310483 );
or ( n32166 , n322590 , n322591 );
buf ( n322593 , n866 );
nand ( n32168 , n32166 , n322593 );
buf ( n32169 , n32168 );
buf ( n322596 , n32169 );
buf ( n322597 , n311234 );
buf ( n322598 , n310658 );
nor ( n322599 , n322597 , n322598 );
buf ( n322600 , n322599 );
buf ( n322601 , n322600 );
xor ( n322602 , n322596 , n322601 );
buf ( n322603 , n311891 );
buf ( n322604 , n322493 );
or ( n322605 , n322603 , n322604 );
buf ( n322606 , n311246 );
buf ( n322607 , n311234 );
buf ( n322608 , n832 );
and ( n32183 , n322607 , n322608 );
buf ( n322610 , n20700 );
buf ( n322611 , n864 );
and ( n32186 , n322610 , n322611 );
nor ( n322613 , n32183 , n32186 );
buf ( n322614 , n322613 );
buf ( n322615 , n322614 );
or ( n32190 , n322606 , n322615 );
nand ( n322617 , n322605 , n32190 );
buf ( n322618 , n322617 );
buf ( n322619 , n322618 );
xor ( n322620 , n322602 , n322619 );
buf ( n322621 , n322620 );
buf ( n322622 , n322621 );
xor ( n322623 , n322585 , n322589 );
xor ( n32198 , n322623 , n322622 );
buf ( n322625 , n32198 );
xor ( n322626 , n322585 , n322589 );
and ( n32201 , n322626 , n322622 );
and ( n32202 , n322585 , n322589 );
or ( n322629 , n32201 , n32202 );
buf ( n322630 , n322629 );
xor ( n32205 , n31890 , n31903 );
and ( n32206 , n32205 , n322339 );
and ( n322633 , n31890 , n31903 );
or ( n322634 , n32206 , n322633 );
buf ( n322635 , n322634 );
buf ( n322636 , n322635 );
buf ( n322637 , n322142 );
xor ( n322638 , n321916 , n321921 );
xor ( n322639 , n322638 , n321939 );
buf ( n322640 , n322639 );
buf ( n322641 , n322640 );
xor ( n32216 , n322636 , n322637 );
xor ( n32217 , n32216 , n322641 );
buf ( n322644 , n32217 );
xor ( n322645 , n322636 , n322637 );
and ( n32220 , n322645 , n322641 );
and ( n322647 , n322636 , n322637 );
or ( n322648 , n32220 , n322647 );
buf ( n322649 , n322648 );
buf ( n322650 , n304630 );
buf ( n322651 , n312467 );
buf ( n322652 , n862 );
and ( n322653 , n322651 , n322652 );
buf ( n322654 , n304739 );
buf ( n322655 , n890 );
and ( n322656 , n322654 , n322655 );
nor ( n322657 , n322653 , n322656 );
buf ( n322658 , n322657 );
buf ( n322659 , n322658 );
or ( n32234 , n322650 , n322659 );
buf ( n322661 , n304655 );
buf ( n322662 , n312467 );
buf ( n322663 , n861 );
and ( n32238 , n322662 , n322663 );
buf ( n322665 , n304771 );
buf ( n322666 , n890 );
and ( n32241 , n322665 , n322666 );
nor ( n322668 , n32238 , n32241 );
buf ( n322669 , n322668 );
buf ( n322670 , n322669 );
or ( n322671 , n322661 , n322670 );
nand ( n322672 , n32234 , n322671 );
buf ( n322673 , n322672 );
buf ( n322674 , n322673 );
buf ( n322675 , n863 );
buf ( n322676 , n891 );
or ( n322677 , n322675 , n322676 );
buf ( n322678 , n892 );
nand ( n32253 , n322677 , n322678 );
buf ( n322680 , n32253 );
buf ( n322681 , n322680 );
buf ( n322682 , n863 );
buf ( n322683 , n891 );
nand ( n322684 , n322682 , n322683 );
buf ( n322685 , n322684 );
buf ( n322686 , n322685 );
buf ( n322687 , n890 );
and ( n32262 , n322681 , n322686 , n322687 );
buf ( n322689 , n32262 );
buf ( n322690 , n322689 );
buf ( n322691 , n305881 );
buf ( n322692 , n894 );
buf ( n322693 , n14447 );
and ( n322694 , n322692 , n322693 );
not ( n32269 , n322692 );
buf ( n322696 , n859 );
and ( n322697 , n32269 , n322696 );
nor ( n32272 , n322694 , n322697 );
buf ( n322699 , n32272 );
buf ( n322700 , n322699 );
or ( n32275 , n322691 , n322700 );
buf ( n322702 , n894 );
not ( n322703 , n322702 );
buf ( n322704 , n858 );
nor ( n322705 , n322703 , n322704 );
buf ( n322706 , n322705 );
buf ( n322707 , n322706 );
buf ( n322708 , n858 );
not ( n322709 , n322708 );
buf ( n322710 , n894 );
nor ( n322711 , n322709 , n322710 );
buf ( n322712 , n322711 );
buf ( n322713 , n322712 );
nor ( n322714 , n322707 , n322713 );
buf ( n322715 , n322714 );
buf ( n322716 , n322715 );
buf ( n322717 , n15469 );
or ( n32292 , n322716 , n322717 );
nand ( n322719 , n32275 , n32292 );
buf ( n322720 , n322719 );
buf ( n322721 , n322720 );
and ( n32296 , n322690 , n322721 );
buf ( n322723 , n32296 );
buf ( n32298 , n322723 );
buf ( n322725 , n305881 );
buf ( n322726 , n322715 );
or ( n322727 , n322725 , n322726 );
buf ( n322728 , n322424 );
buf ( n322729 , n15469 );
or ( n322730 , n322728 , n322729 );
nand ( n322731 , n322727 , n322730 );
buf ( n322732 , n322731 );
buf ( n322733 , n322732 );
buf ( n322734 , n305144 );
buf ( n322735 , n863 );
and ( n32310 , n322734 , n322735 );
buf ( n322737 , n32310 );
buf ( n322738 , n322737 );
xor ( n32313 , n322733 , n322738 );
buf ( n322740 , n15057 );
buf ( n322741 , n305566 );
buf ( n322742 , n860 );
and ( n322743 , n322741 , n322742 );
buf ( n32318 , n305241 );
buf ( n322745 , n892 );
and ( n322746 , n32318 , n322745 );
nor ( n322747 , n322743 , n322746 );
buf ( n322748 , n322747 );
buf ( n322749 , n322748 );
or ( n322750 , n322740 , n322749 );
buf ( n322751 , n305489 );
buf ( n322752 , n892 );
buf ( n322753 , n14447 );
and ( n32328 , n322752 , n322753 );
not ( n322755 , n322752 );
buf ( n322756 , n859 );
and ( n32331 , n322755 , n322756 );
nor ( n322758 , n32328 , n32331 );
buf ( n322759 , n322758 );
buf ( n322760 , n322759 );
or ( n322761 , n322751 , n322760 );
nand ( n322762 , n322750 , n322761 );
buf ( n322763 , n322762 );
buf ( n322764 , n322763 );
xor ( n322765 , n32313 , n322764 );
buf ( n322766 , n322765 );
buf ( n322767 , n322766 );
xor ( n32342 , n322674 , n32298 );
xor ( n322769 , n32342 , n322767 );
buf ( n322770 , n322769 );
xor ( n322771 , n322674 , n32298 );
and ( n322772 , n322771 , n322767 );
and ( n32347 , n322674 , n32298 );
or ( n322774 , n322772 , n32347 );
buf ( n322775 , n322774 );
xor ( n32350 , n322542 , n322551 );
xor ( n322777 , n32350 , n322558 );
buf ( n322778 , n322777 );
buf ( n322779 , n311891 );
buf ( n322780 , n322614 );
or ( n322781 , n322779 , n322780 );
buf ( n322782 , n311246 );
buf ( n322783 , n311234 );
or ( n322784 , n322782 , n322783 );
nand ( n32359 , n322781 , n322784 );
buf ( n32360 , n32359 );
buf ( n32361 , n32360 );
buf ( n32362 , n833 );
buf ( n32363 , n864 );
nand ( n32364 , n32362 , n32363 );
buf ( n32365 , n32364 );
buf ( n322792 , n32365 );
xor ( n32367 , n322596 , n322601 );
and ( n322794 , n32367 , n322619 );
and ( n32369 , n322596 , n322601 );
or ( n32370 , n322794 , n32369 );
buf ( n322797 , n32370 );
buf ( n322798 , n322797 );
xor ( n32373 , n32361 , n322792 );
xor ( n322800 , n32373 , n322798 );
buf ( n322801 , n322800 );
xor ( n32376 , n32361 , n322792 );
and ( n322803 , n32376 , n322798 );
and ( n322804 , n32361 , n322792 );
or ( n32379 , n322803 , n322804 );
buf ( n322806 , n32379 );
buf ( n322807 , n305561 );
buf ( n322808 , n322759 );
or ( n322809 , n322807 , n322808 );
buf ( n322810 , n305489 );
buf ( n322811 , n322384 );
or ( n322812 , n322810 , n322811 );
nand ( n32387 , n322809 , n322812 );
buf ( n322814 , n32387 );
buf ( n32389 , n322814 );
buf ( n322816 , n322058 );
buf ( n322817 , n863 );
and ( n322818 , n322816 , n322817 );
buf ( n32393 , n305192 );
buf ( n322820 , n888 );
and ( n322821 , n32393 , n322820 );
nor ( n322822 , n322818 , n322821 );
buf ( n322823 , n322822 );
buf ( n322824 , n322823 );
buf ( n322825 , n305135 );
or ( n322826 , n322824 , n322825 );
buf ( n322827 , n15861 );
buf ( n322828 , n322066 );
or ( n322829 , n322827 , n322828 );
nand ( n322830 , n322826 , n322829 );
buf ( n322831 , n322830 );
buf ( n322832 , n322831 );
buf ( n322833 , n320083 );
buf ( n322834 , n322669 );
or ( n322835 , n322833 , n322834 );
buf ( n322836 , n304655 );
buf ( n322837 , n31941 );
or ( n32412 , n322836 , n322837 );
nand ( n322839 , n322835 , n32412 );
buf ( n322840 , n322839 );
buf ( n322841 , n322840 );
xor ( n322842 , n32389 , n322832 );
xor ( n322843 , n322842 , n322841 );
buf ( n322844 , n322843 );
xor ( n322845 , n32389 , n322832 );
and ( n322846 , n322845 , n322841 );
and ( n32421 , n32389 , n322832 );
or ( n322848 , n322846 , n32421 );
buf ( n322849 , n322848 );
xor ( n32424 , n322375 , n322392 );
xor ( n322851 , n32424 , n322435 );
buf ( n322852 , n322851 );
xor ( n32427 , n322146 , n322151 );
and ( n322854 , n32427 , n322169 );
and ( n322855 , n322146 , n322151 );
or ( n32430 , n322854 , n322855 );
buf ( n322857 , n32430 );
buf ( n322858 , n311234 );
buf ( n322859 , n20700 );
nor ( n322860 , n322858 , n322859 );
buf ( n322861 , n322860 );
buf ( n322862 , n322861 );
buf ( n322863 , n32365 );
not ( n322864 , n322863 );
buf ( n322865 , n322864 );
buf ( n322866 , n322865 );
buf ( n322867 , n311246 );
not ( n32442 , n322867 );
buf ( n322869 , n311891 );
not ( n32444 , n322869 );
or ( n322871 , n32442 , n32444 );
buf ( n322872 , n864 );
nand ( n32447 , n322871 , n322872 );
buf ( n322874 , n32447 );
buf ( n322875 , n322874 );
xor ( n322876 , n322862 , n322866 );
xor ( n322877 , n322876 , n322875 );
buf ( n322878 , n322877 );
xor ( n32453 , n322862 , n322866 );
and ( n32454 , n32453 , n322875 );
and ( n322881 , n322862 , n322866 );
or ( n32456 , n32454 , n322881 );
buf ( n322883 , n32456 );
xor ( n322884 , n322048 , n322053 );
xor ( n32459 , n322884 , n322074 );
buf ( n322886 , n32459 );
xor ( n32461 , n322733 , n322738 );
and ( n322888 , n32461 , n322764 );
and ( n322889 , n322733 , n322738 );
or ( n32464 , n322888 , n322889 );
buf ( n322891 , n32464 );
xor ( n322892 , n322690 , n322721 );
buf ( n322893 , n322892 );
xor ( n32468 , n31983 , n322432 );
buf ( n322895 , n32468 );
buf ( n322896 , n863 );
buf ( n322897 , n893 );
or ( n322898 , n322896 , n322897 );
buf ( n322899 , n894 );
nand ( n322900 , n322898 , n322899 );
buf ( n322901 , n322900 );
buf ( n32476 , n322901 );
buf ( n322903 , n863 );
buf ( n322904 , n893 );
nand ( n322905 , n322903 , n322904 );
buf ( n322906 , n322905 );
buf ( n322907 , n322906 );
buf ( n322908 , n892 );
and ( n322909 , n32476 , n322907 , n322908 );
buf ( n322910 , n322909 );
buf ( n322911 , n322910 );
buf ( n322912 , n305029 );
buf ( n322913 , n894 );
not ( n32488 , n322913 );
buf ( n322915 , n861 );
nor ( n32490 , n32488 , n322915 );
buf ( n322917 , n32490 );
buf ( n322918 , n322917 );
buf ( n322919 , n861 );
not ( n32494 , n322919 );
buf ( n322921 , n894 );
nor ( n32496 , n32494 , n322921 );
buf ( n322923 , n32496 );
buf ( n322924 , n322923 );
nor ( n32499 , n322918 , n322924 );
buf ( n322926 , n32499 );
buf ( n322927 , n322926 );
or ( n322928 , n322912 , n322927 );
buf ( n322929 , n894 );
not ( n32504 , n322929 );
buf ( n322931 , n860 );
nor ( n32506 , n32504 , n322931 );
buf ( n322933 , n32506 );
buf ( n322934 , n322933 );
buf ( n322935 , n860 );
not ( n32510 , n322935 );
buf ( n322937 , n894 );
nor ( n32512 , n32510 , n322937 );
buf ( n322939 , n32512 );
buf ( n322940 , n322939 );
nor ( n32515 , n322934 , n322940 );
buf ( n322942 , n32515 );
buf ( n322943 , n322942 );
buf ( n322944 , n15469 );
or ( n32519 , n322943 , n322944 );
nand ( n32520 , n322928 , n32519 );
buf ( n322947 , n32520 );
buf ( n322948 , n322947 );
xor ( n32523 , n322911 , n322948 );
buf ( n322950 , n32523 );
and ( n32525 , n322911 , n322948 );
buf ( n322952 , n32525 );
buf ( n322953 , n312467 );
buf ( n322954 , n863 );
and ( n322955 , n322953 , n322954 );
buf ( n322956 , n305192 );
buf ( n322957 , n890 );
and ( n32532 , n322956 , n322957 );
nor ( n32533 , n322955 , n32532 );
buf ( n322960 , n32533 );
buf ( n322961 , n322960 );
buf ( n322962 , n304630 );
buf ( n322963 , n304655 );
buf ( n322964 , n322658 );
or ( n32539 , n322961 , n322962 );
or ( n322966 , n322963 , n322964 );
nand ( n322967 , n32539 , n322966 );
buf ( n322968 , n322967 );
buf ( n32543 , n305192 );
buf ( n322970 , n28078 );
buf ( n322971 , n862 );
buf ( n322972 , n894 );
xor ( n32547 , n322971 , n322972 );
buf ( n322974 , n32547 );
buf ( n322975 , n322974 );
buf ( n322976 , n895 );
nand ( n322977 , n322975 , n322976 );
buf ( n322978 , n322977 );
buf ( n322979 , n322978 );
not ( n322980 , n32543 );
not ( n322981 , n322970 );
or ( n322982 , n322980 , n322981 );
nand ( n32557 , n322982 , n322979 );
buf ( n322984 , n32557 );
buf ( n322985 , n322974 );
buf ( n322986 , n28078 );
buf ( n322987 , n322926 );
not ( n322988 , n322987 );
buf ( n322989 , n895 );
nand ( n322990 , n322988 , n322989 );
buf ( n322991 , n322990 );
buf ( n322992 , n322991 );
not ( n322993 , n322985 );
not ( n322994 , n322986 );
or ( n32569 , n322993 , n322994 );
nand ( n322996 , n32569 , n322992 );
buf ( n322997 , n322996 );
buf ( n322998 , n305430 );
buf ( n322999 , n863 );
and ( n32574 , n322998 , n322999 );
buf ( n323001 , n32574 );
buf ( n323002 , n305566 );
buf ( n323003 , n862 );
and ( n323004 , n323002 , n323003 );
buf ( n32579 , n304739 );
buf ( n323006 , n892 );
and ( n323007 , n32579 , n323006 );
nor ( n323008 , n323004 , n323007 );
buf ( n323009 , n323008 );
buf ( n323010 , n323009 );
buf ( n323011 , n305430 );
not ( n32586 , n323010 );
nand ( n323013 , n32586 , n323011 );
buf ( n323014 , n323013 );
not ( n32589 , n305191 );
nand ( n32590 , n32589 , n895 );
buf ( n323017 , n32590 );
buf ( n323018 , n894 );
and ( n323019 , n323017 , n323018 );
buf ( n323020 , n323019 );
buf ( n323021 , n305192 );
buf ( n323022 , n892 );
buf ( n323023 , n305566 );
buf ( n323024 , n863 );
or ( n323025 , n323021 , n323022 );
or ( n323026 , n323023 , n323024 );
nand ( n323027 , n323025 , n323026 );
buf ( n323028 , n323027 );
buf ( n323029 , n305566 );
buf ( n323030 , n861 );
buf ( n323031 , n304771 );
buf ( n323032 , n892 );
and ( n323033 , n323029 , n323030 );
and ( n32608 , n323031 , n323032 );
nor ( n323035 , n323033 , n32608 );
buf ( n323036 , n323035 );
buf ( n323037 , n32590 );
not ( n323038 , n323037 );
buf ( n323039 , n323038 );
buf ( n323040 , n323001 );
buf ( n323041 , n322997 );
and ( n32616 , n831 , n307445 );
not ( n323043 , n831 );
buf ( n323044 , n889 );
buf ( n323045 , n307435 );
xor ( n323046 , n323044 , n323045 );
buf ( n323047 , n307440 );
and ( n32622 , n323046 , n323047 );
and ( n323049 , n323044 , n323045 );
or ( n323050 , n32622 , n323049 );
buf ( n323051 , n323050 );
and ( n323052 , n323043 , n323051 );
or ( n323053 , n32616 , n323052 );
not ( n32628 , n831 );
not ( n323055 , n307428 );
or ( n323056 , n32628 , n323055 );
not ( n323057 , n831 );
nand ( n32632 , n19722 , n323057 );
nand ( n323059 , n323056 , n32632 );
nand ( n323060 , n323053 , n323059 );
or ( n323061 , n323059 , n323053 );
nand ( n32636 , n323060 , n323061 );
and ( n323063 , n831 , n303406 );
not ( n32638 , n831 );
and ( n32639 , n32638 , n310169 );
or ( n323066 , n323063 , n32639 );
not ( n323067 , n323066 );
not ( n32642 , n831 );
xor ( n323069 , n323044 , n323045 );
xor ( n323070 , n323069 , n323047 );
buf ( n323071 , n323070 );
and ( n323072 , n32642 , n323071 );
not ( n323073 , n32642 );
and ( n32648 , n323073 , n17022 );
nor ( n323075 , n323072 , n32648 );
nand ( n323076 , n323067 , n323075 );
not ( n32651 , n323076 );
and ( n323078 , n831 , n307422 );
not ( n32653 , n831 );
and ( n323080 , n32653 , n310202 );
or ( n323081 , n323078 , n323080 );
not ( n323082 , n323081 );
and ( n323083 , n831 , n307417 );
not ( n32658 , n831 );
buf ( n323085 , n891 );
buf ( n32660 , n307297 );
xor ( n32661 , n323085 , n32660 );
buf ( n323088 , n307302 );
xor ( n323089 , n32661 , n323088 );
buf ( n323090 , n323089 );
and ( n323091 , n32658 , n323090 );
nor ( n323092 , n323083 , n323091 );
not ( n32667 , n323092 );
not ( n32668 , n32667 );
or ( n32669 , n323082 , n32668 );
nand ( n32670 , n307408 , n831 );
not ( n32671 , n32670 );
nand ( n323098 , n310197 , n323057 );
not ( n323099 , n323098 );
or ( n32674 , n32671 , n323099 );
and ( n323101 , n831 , n307384 );
not ( n323102 , n831 );
and ( n32677 , n323102 , n310213 );
or ( n323104 , n323101 , n32677 );
not ( n323105 , n323104 );
buf ( n323106 , n831 );
not ( n32681 , n323106 );
buf ( n323108 , n307366 );
not ( n32683 , n323108 );
or ( n32684 , n32681 , n32683 );
buf ( n323111 , n831 );
not ( n323112 , n323111 );
buf ( n323113 , n310227 );
nand ( n323114 , n323112 , n323113 );
buf ( n323115 , n323114 );
buf ( n323116 , n323115 );
nand ( n323117 , n32684 , n323116 );
buf ( n323118 , n323117 );
not ( n32693 , n323118 );
not ( n323120 , n32693 );
and ( n323121 , n831 , n307335 );
not ( n323122 , n831 );
and ( n32697 , n323122 , n310208 );
nor ( n323124 , n323121 , n32697 );
not ( n323125 , n323124 );
or ( n32700 , n323120 , n323125 );
not ( n323127 , n831 );
not ( n323128 , n307370 );
or ( n32703 , n323127 , n323128 );
nand ( n32704 , n310222 , n323057 );
nand ( n323131 , n32703 , n32704 );
and ( n32706 , n831 , n307377 );
or ( n32707 , n32706 , C0 );
and ( n323134 , n323131 , n32707 );
nand ( n323135 , n32700 , n323134 );
not ( n32710 , n323124 );
nand ( n32711 , n32710 , n323118 );
nand ( n32712 , n323105 , n323135 , n32711 );
nand ( n32713 , n32674 , n32712 );
not ( n32714 , n32713 );
not ( n323141 , n32711 );
not ( n323142 , n323135 );
or ( n32717 , n323141 , n323142 );
nand ( n323144 , n32717 , n323104 );
not ( n323145 , n323144 );
or ( n32720 , n32714 , n323145 );
not ( n32721 , n323081 );
nand ( n32722 , n32721 , n323092 );
nand ( n32723 , n32720 , n32722 );
nand ( n323150 , n32669 , n32723 );
not ( n323151 , n323150 );
not ( n32726 , n831 );
nand ( n32727 , n32726 , n310164 );
nand ( n32728 , n307258 , n831 );
not ( n32729 , n831 );
not ( n323156 , n307307 );
or ( n323157 , n32729 , n323156 );
xor ( n32732 , n323085 , n32660 );
and ( n32733 , n32732 , n323088 );
and ( n32734 , n323085 , n32660 );
or ( n32735 , n32733 , n32734 );
buf ( n32736 , n32735 );
nand ( n323163 , n32736 , n5980 );
nand ( n32738 , n323157 , n323163 );
not ( n32739 , n32738 );
nand ( n32740 , n32727 , n32728 , n32739 );
not ( n323167 , n32740 );
or ( n323168 , n323151 , n323167 );
not ( n32743 , n32738 );
not ( n323170 , n32743 );
not ( n323171 , n310164 );
not ( n32746 , n831 );
and ( n32747 , n323171 , n32746 );
not ( n32748 , n307258 );
and ( n32749 , n32748 , n831 );
nor ( n32750 , n32747 , n32749 );
nand ( n323177 , n323170 , n32750 );
nand ( n323178 , n323168 , n323177 );
not ( n32753 , n323178 );
or ( n323180 , n32651 , n32753 );
not ( n323181 , n323075 );
nand ( n32756 , n323181 , n323066 );
nand ( n32757 , n323180 , n32756 );
not ( n32758 , n32757 );
and ( n32759 , n32636 , n32758 );
not ( n32760 , n32636 );
and ( n323187 , n32760 , n32757 );
nor ( n323188 , n32759 , n323187 );
buf ( n323189 , n323188 );
xor ( n323190 , n323040 , n323041 );
xor ( n32765 , n323190 , n323189 );
buf ( n323192 , n32765 );
xor ( n32767 , n323040 , n323041 );
and ( n32768 , n32767 , n323189 );
and ( n32769 , n323040 , n323041 );
or ( n323196 , n32768 , n32769 );
buf ( n323197 , n323196 );
buf ( n323198 , n323028 );
not ( n32773 , n323198 );
buf ( n323200 , n14272 );
not ( n32775 , n323200 );
or ( n32776 , n32773 , n32775 );
buf ( n323203 , n323014 );
nand ( n32778 , n32776 , n323203 );
buf ( n323205 , n32778 );
buf ( n323206 , n323205 );
buf ( n323207 , n322950 );
not ( n32782 , n323061 );
not ( n32783 , n32757 );
or ( n323210 , n32782 , n32783 );
nand ( n323211 , n323210 , n323060 );
not ( n32786 , n831 );
not ( n32787 , n307237 );
or ( n32788 , n32786 , n32787 );
not ( n32789 , n831 );
nand ( n323216 , n32789 , n310155 );
nand ( n323217 , n32788 , n323216 );
not ( n32792 , n323217 );
nand ( n32793 , n303570 , n831 );
nand ( n32794 , n310125 , n32642 );
nand ( n323221 , n32792 , n32793 , n32794 );
not ( n323222 , n32794 );
not ( n32797 , n32793 );
or ( n323224 , n323222 , n32797 );
nand ( n323225 , n323224 , n323217 );
nand ( n32800 , n323221 , n323225 );
xnor ( n32801 , n323211 , n32800 );
buf ( n323228 , n32801 );
xor ( n32803 , n323206 , n323207 );
xor ( n32804 , n32803 , n323228 );
buf ( n323231 , n32804 );
xor ( n323232 , n323206 , n323207 );
and ( n32807 , n323232 , n323228 );
and ( n32808 , n323206 , n323207 );
or ( n32809 , n32807 , n32808 );
buf ( n32810 , n32809 );
buf ( n323237 , n304658 );
buf ( n323238 , n863 );
and ( n323239 , n323237 , n323238 );
buf ( n323240 , n323239 );
buf ( n323241 , n305881 );
buf ( n323242 , n322942 );
or ( n323243 , n323241 , n323242 );
buf ( n323244 , n322699 );
buf ( n323245 , n15469 );
or ( n32820 , n323244 , n323245 );
nand ( n32821 , n323243 , n32820 );
buf ( n323248 , n32821 );
xor ( n32823 , n323240 , n323248 );
buf ( n323250 , n15057 );
buf ( n323251 , n323009 );
or ( n32826 , n323250 , n323251 );
buf ( n323253 , n305489 );
buf ( n323254 , n323036 );
or ( n32829 , n323253 , n323254 );
nand ( n32830 , n32826 , n32829 );
buf ( n323257 , n32830 );
and ( n32832 , n32823 , n323257 );
and ( n32833 , n323240 , n323248 );
or ( n32834 , n32832 , n32833 );
buf ( n323261 , n32834 );
buf ( n323262 , n305561 );
buf ( n323263 , n323036 );
or ( n32838 , n323262 , n323263 );
buf ( n323265 , n305489 );
buf ( n323266 , n322748 );
or ( n32841 , n323265 , n323266 );
nand ( n32842 , n32838 , n32841 );
buf ( n323269 , n32842 );
buf ( n323270 , n323269 );
xor ( n32845 , n322968 , n323270 );
xor ( n323272 , n32845 , n322893 );
buf ( n323273 , n323272 );
not ( n32848 , n323211 );
buf ( n32849 , n323057 );
not ( n32850 , n32849 );
not ( n323277 , n310119 );
or ( n32852 , n32850 , n323277 );
nand ( n32853 , n303566 , n831 );
nand ( n323280 , n32852 , n32853 );
and ( n32855 , n831 , n303279 );
not ( n323282 , n831 );
and ( n32857 , n323282 , n310130 );
or ( n32858 , n32855 , n32857 );
or ( n323285 , n323280 , n32858 );
nand ( n323286 , n323285 , n323221 );
not ( n32861 , n323286 );
not ( n323288 , n32861 );
or ( n323289 , n32848 , n323288 );
nand ( n32864 , n323280 , n32858 );
nand ( n323291 , n32864 , n323225 );
nand ( n323292 , n323291 , n323285 );
buf ( n323293 , n323292 );
nand ( n32868 , n323289 , n323293 );
not ( n323295 , n32868 );
not ( n32870 , n295148 );
and ( n32871 , n831 , n303562 );
not ( n323298 , n831 );
xor ( n323299 , n295059 , n295060 );
xor ( n32874 , n323299 , n295062 );
buf ( n323301 , n32874 );
and ( n323302 , n323298 , n323301 );
nor ( n32877 , n32871 , n323302 );
nor ( n323304 , n32870 , n32877 );
not ( n323305 , n323304 );
not ( n32880 , n295148 );
nand ( n323307 , n32877 , n32880 );
nand ( n32882 , n323305 , n323307 );
not ( n323309 , n32882 );
or ( n32884 , n323295 , n323309 );
or ( n32885 , n32868 , n32882 );
nand ( n32886 , n32884 , n32885 );
buf ( n323313 , n32886 );
xor ( n323314 , n323261 , n323273 );
xor ( n32889 , n323314 , n323313 );
buf ( n323316 , n32889 );
xor ( n323317 , n323261 , n323273 );
and ( n32892 , n323317 , n323313 );
and ( n323319 , n323261 , n323273 );
or ( n323320 , n32892 , n323319 );
buf ( n323321 , n323320 );
xor ( n32896 , n322968 , n323270 );
and ( n32897 , n32896 , n322893 );
and ( n323324 , n322968 , n323270 );
or ( n323325 , n32897 , n323324 );
buf ( n323326 , n323325 );
buf ( n323327 , n322770 );
not ( n323328 , n323307 );
not ( n32903 , n32868 );
or ( n32904 , n323328 , n32903 );
nand ( n323331 , n32904 , n323305 );
nor ( n32906 , n310108 , n831 );
nor ( n323333 , n307194 , n296412 );
or ( n323334 , n32906 , n323333 );
not ( n323335 , n4640 );
nand ( n32910 , n323334 , n323335 );
not ( n323337 , n323335 );
nor ( n32912 , n32906 , n323333 );
nand ( n32913 , n323337 , n32912 );
nand ( n323340 , n32910 , n32913 );
not ( n323341 , n323340 );
and ( n32916 , n323331 , n323341 );
not ( n323343 , n323331 );
and ( n323344 , n323343 , n323340 );
nor ( n32919 , n32916 , n323344 );
buf ( n323346 , n32919 );
xor ( n323347 , n323326 , n323327 );
xor ( n323348 , n323347 , n323346 );
buf ( n323349 , n323348 );
xor ( n323350 , n323326 , n323327 );
and ( n32925 , n323350 , n323346 );
and ( n32926 , n323326 , n323327 );
or ( n323353 , n32925 , n32926 );
buf ( n323354 , n323353 );
buf ( n323355 , n322775 );
xor ( n323356 , n322895 , n322891 );
xor ( n323357 , n323356 , n322844 );
buf ( n323358 , n323357 );
not ( n323359 , n323307 );
nor ( n323360 , n323292 , n323359 );
buf ( n32935 , n323304 );
or ( n323362 , n323360 , n32935 );
nand ( n32937 , n323362 , n32910 );
not ( n323364 , n323286 );
nand ( n32939 , n323364 , n323211 , n323307 , n32910 );
nand ( n32940 , n32937 , n32939 , n32913 );
buf ( n323367 , n32940 );
not ( n323368 , n310102 );
not ( n32943 , n32849 );
or ( n323370 , n323368 , n32943 );
nand ( n323371 , n307171 , n831 );
nand ( n32946 , n323370 , n323371 );
not ( n323373 , n32946 );
and ( n323374 , n831 , n307187 );
not ( n32949 , n831 );
and ( n323376 , n32949 , n310113 );
or ( n323377 , n323374 , n323376 );
not ( n32952 , n323377 );
nand ( n32953 , n323373 , n32952 );
nand ( n32954 , n323377 , n32946 );
nand ( n323381 , n32953 , n32954 );
xnor ( n323382 , n323367 , n323381 );
buf ( n323383 , n323382 );
xor ( n32958 , n323355 , n323358 );
xor ( n323385 , n32958 , n323383 );
buf ( n323386 , n323385 );
xor ( n32961 , n323355 , n323358 );
and ( n32962 , n32961 , n323383 );
and ( n32963 , n323355 , n323358 );
or ( n323390 , n32962 , n32963 );
buf ( n323391 , n323390 );
xor ( n32966 , n322895 , n322891 );
and ( n32967 , n32966 , n322844 );
and ( n32968 , n322895 , n322891 );
or ( n323395 , n32967 , n32968 );
buf ( n323396 , n323395 );
xor ( n32971 , n322886 , n322849 );
xor ( n32972 , n32971 , n322852 );
buf ( n323399 , n32972 );
not ( n323400 , n323367 );
not ( n32975 , n32953 );
or ( n323402 , n323400 , n32975 );
nand ( n323403 , n323402 , n32954 );
not ( n32978 , n309969 );
not ( n323405 , n831 );
not ( n323406 , n303558 );
or ( n32981 , n323405 , n323406 );
nand ( n32982 , n310094 , n32642 );
nand ( n32983 , n32981 , n32982 );
not ( n32984 , n32983 );
nand ( n323411 , n32978 , n32984 );
nand ( n323412 , n32983 , n309969 );
and ( n32987 , n323411 , n323412 );
xor ( n32988 , n323403 , n32987 );
buf ( n323415 , n32988 );
xor ( n323416 , n323396 , n323399 );
xor ( n323417 , n323416 , n323415 );
buf ( n323418 , n323417 );
xor ( n323419 , n323396 , n323399 );
and ( n323420 , n323419 , n323415 );
and ( n32995 , n323396 , n323399 );
or ( n323422 , n323420 , n32995 );
buf ( n323423 , n323422 );
xor ( n32998 , n322886 , n322849 );
and ( n323425 , n32998 , n322852 );
and ( n323426 , n322886 , n322849 );
or ( n33001 , n323425 , n323426 );
buf ( n323428 , n33001 );
buf ( n323429 , n322451 );
not ( n33004 , n307128 );
not ( n33005 , n831 );
or ( n33006 , n33004 , n33005 );
nand ( n33007 , n310085 , n32642 );
nand ( n33008 , n33006 , n33007 );
and ( n33009 , n831 , n307134 );
not ( n33010 , n831 );
and ( n323437 , n33010 , n310099 );
or ( n33012 , n33009 , n323437 );
nand ( n323439 , n33008 , n33012 );
buf ( n323440 , n323439 );
not ( n33015 , n33008 );
not ( n33016 , n33012 );
nand ( n33017 , n33015 , n33016 );
buf ( n33018 , n33017 );
and ( n33019 , n323440 , n33018 );
and ( n323446 , n32953 , n323411 );
not ( n323447 , n323446 );
not ( n33022 , n323367 );
or ( n323449 , n323447 , n33022 );
not ( n323450 , n323412 );
not ( n33025 , n32954 );
or ( n33026 , n323450 , n33025 );
nand ( n33027 , n33026 , n323411 );
buf ( n33028 , n33027 );
nand ( n33029 , n323449 , n33028 );
xor ( n33030 , n33019 , n33029 );
buf ( n33031 , n33030 );
xor ( n33032 , n323428 , n323429 );
xor ( n33033 , n33032 , n33031 );
buf ( n323460 , n33033 );
xor ( n323461 , n323428 , n323429 );
and ( n323462 , n323461 , n33031 );
and ( n33037 , n323428 , n323429 );
or ( n33038 , n323462 , n33037 );
buf ( n323465 , n33038 );
buf ( n323466 , n322117 );
buf ( n323467 , n321568 );
buf ( n323468 , n831 );
not ( n323469 , n323468 );
buf ( n323470 , n307031 );
not ( n323471 , n323470 );
or ( n33046 , n323469 , n323471 );
buf ( n323473 , n831 );
not ( n323474 , n323473 );
buf ( n323475 , n310082 );
nand ( n33050 , n323474 , n323475 );
buf ( n323477 , n33050 );
buf ( n323478 , n323477 );
nand ( n33053 , n33046 , n323478 );
buf ( n323480 , n33053 );
buf ( n323481 , n323480 );
not ( n33056 , n323481 );
not ( n323483 , n303514 );
not ( n323484 , n831 );
or ( n33059 , n323483 , n323484 );
buf ( n323486 , n32642 );
nand ( n323487 , n310216 , n323486 );
nand ( n33062 , n33059 , n323487 );
buf ( n323489 , n33062 );
not ( n33064 , n323489 );
nand ( n323491 , n33056 , n33064 );
nand ( n33066 , n323480 , n33062 );
nand ( n33067 , n323491 , n33066 );
not ( n323494 , n292343 );
and ( n323495 , n323057 , n310077 );
not ( n33070 , n323057 );
and ( n323497 , n33070 , n307122 );
nor ( n323498 , n323495 , n323497 );
nand ( n33073 , n323494 , n323498 );
nand ( n323500 , n32940 , n323446 , n33017 , n33073 );
nand ( n323501 , n323439 , n33027 );
nand ( n33076 , n323501 , n33017 , n33073 );
not ( n33077 , n323498 );
nand ( n33078 , n292343 , n33077 );
nand ( n323505 , n323500 , n33076 , n33078 );
buf ( n323506 , n323505 );
xnor ( n33081 , n33067 , n323506 );
buf ( n323508 , n33081 );
xor ( n33083 , n323466 , n323467 );
xor ( n323510 , n33083 , n323508 );
buf ( n323511 , n323510 );
xor ( n33086 , n323466 , n323467 );
and ( n323513 , n33086 , n323508 );
and ( n323514 , n323466 , n323467 );
or ( n33089 , n323513 , n323514 );
buf ( n323516 , n33089 );
buf ( n323517 , n321573 );
buf ( n323518 , n321634 );
not ( n323519 , n323491 );
not ( n323520 , n323505 );
or ( n323521 , n323519 , n323520 );
nand ( n33096 , n323521 , n33066 );
not ( n323523 , n301147 );
not ( n33098 , n323523 );
and ( n33099 , n323057 , n310186 );
not ( n323526 , n323057 );
and ( n323527 , n323526 , n307013 );
nor ( n33102 , n33099 , n323527 );
not ( n323529 , n33102 );
nand ( n323530 , n33098 , n323529 );
nand ( n33105 , n33102 , n323523 );
buf ( n323532 , n33105 );
nand ( n323533 , n323530 , n323532 );
xnor ( n33108 , n33096 , n323533 );
buf ( n323535 , n33108 );
xor ( n33110 , n323517 , n323518 );
xor ( n323537 , n33110 , n323535 );
buf ( n323538 , n323537 );
xor ( n33113 , n323517 , n323518 );
and ( n323540 , n33113 , n323535 );
and ( n323541 , n323517 , n323518 );
or ( n33116 , n323540 , n323541 );
buf ( n323543 , n33116 );
buf ( n323544 , n321639 );
buf ( n323545 , n321333 );
and ( n323546 , n5980 , n310191 );
not ( n323547 , n5980 );
and ( n33122 , n323547 , n307042 );
nor ( n33123 , n323546 , n33122 );
and ( n33124 , n831 , n13082 );
not ( n323551 , n831 );
and ( n323552 , n323551 , n310158 );
nor ( n33127 , n33124 , n323552 );
nand ( n323554 , n33123 , n33127 );
buf ( n323555 , n323554 );
not ( n33130 , n323555 );
nor ( n33131 , n33123 , n33127 );
buf ( n33132 , n33131 );
nor ( n323559 , n33130 , n33132 );
and ( n323560 , n831 , n307031 );
not ( n33135 , n831 );
and ( n33136 , n33135 , n310082 );
or ( n33137 , n323560 , n33136 );
or ( n33138 , n33137 , n323489 );
nand ( n323565 , n33138 , n323532 );
not ( n323566 , n323565 );
not ( n33141 , n323566 );
not ( n33142 , n323506 );
or ( n33143 , n33141 , n33142 );
not ( n323570 , n33105 );
and ( n323571 , n33062 , n323480 );
not ( n33146 , n323571 );
or ( n33147 , n323570 , n33146 );
nand ( n33148 , n33147 , n323530 );
not ( n323575 , n33148 );
nand ( n323576 , n33143 , n323575 );
xor ( n33151 , n323559 , n323576 );
buf ( n323578 , n33151 );
xor ( n323579 , n323544 , n323545 );
xor ( n33154 , n323579 , n323578 );
buf ( n323581 , n33154 );
xor ( n33156 , n323544 , n323545 );
and ( n323583 , n33156 , n323578 );
and ( n323584 , n323544 , n323545 );
or ( n33159 , n323583 , n323584 );
buf ( n323586 , n33159 );
buf ( n323587 , n321338 );
xor ( n323588 , n322579 , n322358 );
xor ( n33163 , n323588 , n322286 );
buf ( n323590 , n33163 );
not ( n323591 , n323576 );
and ( n323592 , n831 , n303476 );
not ( n33167 , n831 );
and ( n33168 , n33167 , n310139 );
nor ( n33169 , n323592 , n33168 );
not ( n33170 , n831 );
not ( n33171 , n303971 );
or ( n323598 , n33170 , n33171 );
nand ( n323599 , n323598 , n310055 );
not ( n33174 , n323599 );
nand ( n323601 , n33169 , n33174 );
and ( n323602 , n32849 , n310139 );
not ( n33177 , n32849 );
and ( n33178 , n33177 , n303476 );
or ( n33179 , n323602 , n33178 );
not ( n33180 , n33174 );
nand ( n33181 , n33179 , n33180 );
nand ( n323608 , n323601 , n33181 );
nor ( n323609 , n323608 , n33132 );
nand ( n33184 , n323591 , n323609 );
and ( n33185 , n323555 , n323608 );
nand ( n33186 , n33185 , n323576 );
and ( n323613 , n323608 , n33132 );
nor ( n323614 , n323608 , n323555 , n33132 );
nor ( n33189 , n323613 , n323614 );
nand ( n33190 , n33184 , n33186 , n33189 );
buf ( n323617 , n33190 );
xor ( n323618 , n323587 , n323590 );
xor ( n323619 , n323618 , n323617 );
buf ( n323620 , n323619 );
xor ( n33195 , n323587 , n323590 );
and ( n33196 , n33195 , n323617 );
and ( n33197 , n323587 , n323590 );
or ( n33198 , n33196 , n33197 );
buf ( n33199 , n33198 );
buf ( n33200 , n314814 );
buf ( n323627 , n306543 );
not ( n33202 , n16359 );
and ( n323629 , n831 , n306799 );
not ( n323630 , n831 );
buf ( n323631 , n864 );
buf ( n323632 , n304554 );
xor ( n33207 , n323631 , n323632 );
buf ( n323634 , n306794 );
and ( n323635 , n33207 , n323634 );
and ( n323636 , n323631 , n323632 );
or ( n33211 , n323635 , n323636 );
buf ( n323638 , n33211 );
and ( n33213 , n323630 , n323638 );
nor ( n323640 , n323629 , n33213 );
nor ( n323641 , n33202 , n323640 );
buf ( n33216 , n323641 );
not ( n323643 , n33216 );
not ( n323644 , n16359 );
nand ( n33219 , n323644 , n323640 );
nand ( n33220 , n323643 , n33219 );
not ( n33221 , n33220 );
and ( n323648 , n831 , n307058 );
not ( n323649 , n831 );
xor ( n33224 , n872 , n296375 );
xor ( n323651 , n33224 , n296396 );
and ( n323652 , n323649 , n323651 );
nor ( n33227 , n323648 , n323652 );
buf ( n323654 , n831 );
not ( n33229 , n323654 );
buf ( n33230 , n293580 );
not ( n33231 , n33230 );
or ( n33232 , n33229 , n33231 );
buf ( n323659 , n293596 );
nand ( n33234 , n33232 , n323659 );
buf ( n323661 , n33234 );
not ( n33236 , n323661 );
nand ( n323663 , n33227 , n33236 );
not ( n323664 , n831 );
not ( n33239 , n307075 );
or ( n323666 , n323664 , n33239 );
not ( n323667 , n831 );
not ( n323668 , n874 );
not ( n323669 , n307068 );
nand ( n33244 , n323668 , n323669 );
not ( n323671 , n33244 );
not ( n323672 , n14130 );
or ( n33247 , n323671 , n323672 );
not ( n323674 , n323669 );
nand ( n323675 , n323674 , n874 );
nand ( n33250 , n33247 , n323675 );
nand ( n323677 , n323667 , n33250 );
nand ( n323678 , n323666 , n323677 );
not ( n33253 , n323678 );
and ( n323680 , n323057 , n310088 );
not ( n323681 , n323057 );
and ( n33256 , n323681 , n307062 );
nor ( n323683 , n323680 , n33256 );
nand ( n33258 , n33253 , n323683 );
and ( n323685 , n323663 , n33258 );
not ( n33260 , n7951 );
not ( n323687 , n33260 );
not ( n33262 , n874 );
not ( n33263 , n323669 );
or ( n323690 , n33262 , n33263 );
not ( n323691 , n874 );
nand ( n33266 , n323691 , n307068 );
nand ( n323693 , n323690 , n33266 );
and ( n323694 , n323693 , n14130 );
not ( n33269 , n323693 );
not ( n323696 , n14130 );
and ( n323697 , n33269 , n323696 );
nor ( n323698 , n323694 , n323697 );
not ( n33273 , n323698 );
not ( n33274 , n831 );
and ( n323701 , n33273 , n33274 );
nor ( n33276 , n307089 , n323486 );
nor ( n323703 , n323701 , n33276 );
nor ( n323704 , n323687 , n323703 );
not ( n33279 , n5980 );
not ( n33280 , n310144 );
or ( n323707 , n33279 , n33280 );
nand ( n323708 , n307085 , n831 );
nand ( n33283 , n323707 , n323708 );
not ( n33284 , n33283 );
nand ( n323711 , n307080 , n831 );
nand ( n323712 , n310116 , n323486 );
nand ( n33287 , n33284 , n323711 , n323712 );
not ( n33288 , n33287 );
nor ( n33289 , n323704 , n33288 );
not ( n33290 , n33174 );
and ( n323717 , n32849 , n310139 );
not ( n323718 , n32849 );
and ( n33293 , n323718 , n303476 );
nor ( n33294 , n323717 , n33293 );
not ( n33295 , n33294 );
or ( n33296 , n33290 , n33295 );
nand ( n33297 , n33296 , n323554 );
nor ( n323724 , n323565 , n33297 );
nand ( n33299 , n323685 , n33289 , n323505 , n323724 );
not ( n33300 , n33297 );
nand ( n33301 , n33300 , n33148 );
nand ( n323728 , n323601 , n33131 );
nand ( n323729 , n323728 , n33181 );
not ( n33304 , n323729 );
not ( n33305 , n323057 );
not ( n33306 , n323698 );
or ( n323733 , n33305 , n33306 );
nand ( n323734 , n307089 , n831 );
nand ( n33309 , n323733 , n323734 );
nand ( n33310 , n33309 , n7951 );
nand ( n33311 , n323711 , n323712 );
nand ( n323738 , n33311 , n33283 );
nand ( n33313 , n33301 , n33304 , n33310 , n323738 );
not ( n33314 , n33287 );
nand ( n33315 , n33314 , n33310 );
not ( n33316 , n33260 );
nor ( n33317 , n33316 , n323703 );
not ( n33318 , n33317 );
nand ( n323745 , n33313 , n323685 , n33315 , n33318 );
buf ( n323746 , n323663 );
not ( n33321 , n831 );
not ( n33322 , n307075 );
or ( n33323 , n33321 , n33322 );
nand ( n33324 , n33323 , n323677 );
not ( n323751 , n33324 );
buf ( n323752 , n32642 );
and ( n33327 , n323752 , n310088 );
not ( n33328 , n323752 );
and ( n33329 , n33328 , n307062 );
nor ( n323756 , n33327 , n33329 );
nor ( n323757 , n323751 , n323756 );
and ( n33332 , n323746 , n323757 );
not ( n33333 , n293599 );
buf ( n33334 , n33227 );
nor ( n33335 , n33333 , n33334 );
nor ( n323762 , n33332 , n33335 );
nand ( n323763 , n33299 , n323745 , n323762 );
and ( n33338 , n323486 , n310133 );
not ( n33339 , n323486 );
and ( n33340 , n33339 , n306943 );
nor ( n323767 , n33338 , n33340 );
not ( n323768 , n323767 );
not ( n33343 , n303205 );
not ( n323770 , n33343 );
or ( n323771 , n323768 , n323770 );
not ( n33346 , n296366 );
buf ( n323773 , n866 );
buf ( n323774 , n306907 );
xor ( n33349 , n323773 , n323774 );
buf ( n323776 , n306936 );
xor ( n33351 , n33349 , n323776 );
buf ( n323778 , n33351 );
and ( n323779 , n323486 , n323778 );
not ( n33354 , n323486 );
and ( n33355 , n33354 , n306937 );
nor ( n33356 , n323779 , n33355 );
nand ( n33357 , n33346 , n33356 );
nand ( n33358 , n323771 , n33357 );
not ( n33359 , n33358 );
and ( n33360 , n323486 , n310071 );
not ( n323787 , n323486 );
and ( n33362 , n323787 , n306869 );
nor ( n323789 , n33360 , n33362 );
not ( n33364 , n831 );
not ( n323791 , n306885 );
or ( n33366 , n33364 , n323791 );
nand ( n33367 , n33366 , n310068 );
not ( n323794 , n33367 );
nand ( n323795 , n323789 , n323794 );
xor ( n33370 , n310057 , n310058 );
xor ( n33371 , n33370 , n310060 );
buf ( n323798 , n33371 );
and ( n33373 , n323486 , n323798 );
not ( n33374 , n323486 );
and ( n33375 , n33374 , n306889 );
nor ( n33376 , n33373 , n33375 );
not ( n33377 , n294735 );
nand ( n33378 , n33376 , n33377 );
nand ( n33379 , n323795 , n33378 );
not ( n33380 , n33379 );
not ( n323807 , n5982 );
not ( n33382 , n831 );
not ( n33383 , n303421 );
or ( n33384 , n33382 , n33383 );
nand ( n33385 , n310175 , n323486 );
nand ( n33386 , n33384 , n33385 );
not ( n33387 , n33386 );
nand ( n33388 , n323807 , n33387 );
xor ( n33389 , n294722 , n294723 );
xor ( n33390 , n33389 , n294725 );
buf ( n323817 , n33390 );
and ( n33392 , n323752 , n323817 );
not ( n33393 , n323752 );
and ( n33394 , n33393 , n306861 );
nor ( n33395 , n33392 , n33394 );
buf ( n323822 , n831 );
not ( n33397 , n323822 );
buf ( n323824 , n303965 );
not ( n323825 , n323824 );
or ( n33400 , n33397 , n323825 );
buf ( n323827 , n310180 );
buf ( n323828 , n296412 );
nand ( n323829 , n323827 , n323828 );
buf ( n323830 , n323829 );
buf ( n323831 , n323830 );
nand ( n33406 , n33400 , n323831 );
buf ( n323833 , n33406 );
not ( n33408 , n323833 );
nand ( n323835 , n33395 , n33408 );
nand ( n323836 , n33388 , n323835 );
not ( n33411 , n323836 );
and ( n33412 , n33359 , n33380 , n33411 );
not ( n33413 , n306968 );
not ( n323840 , n323752 );
nand ( n323841 , n33413 , n323840 );
not ( n33416 , n323841 );
buf ( n323843 , n865 );
buf ( n323844 , n306961 );
xor ( n323845 , n323843 , n323844 );
buf ( n323846 , n306957 );
xor ( n33421 , n323845 , n323846 );
buf ( n323848 , n33421 );
not ( n33423 , n323848 );
nand ( n33424 , n33423 , n323752 );
not ( n323851 , n33424 );
or ( n33426 , n33416 , n323851 );
not ( n33427 , n296412 );
xor ( n33428 , n323773 , n323774 );
and ( n33429 , n33428 , n323776 );
and ( n33430 , n323773 , n323774 );
or ( n33431 , n33429 , n33430 );
buf ( n323858 , n33431 );
not ( n323859 , n323858 );
or ( n33434 , n33427 , n323859 );
nand ( n33435 , n16545 , n831 );
nand ( n323862 , n33434 , n33435 );
not ( n323863 , n323862 );
nand ( n33438 , n33426 , n323863 );
xor ( n33439 , n323631 , n323632 );
xor ( n33440 , n33439 , n323634 );
buf ( n323867 , n33440 );
and ( n33442 , n32849 , n323867 );
not ( n323869 , n32849 );
buf ( n33444 , n306951 );
and ( n33445 , n323869 , n33444 );
nor ( n323872 , n33442 , n33445 );
not ( n323873 , n831 );
not ( n33448 , n306964 );
or ( n33449 , n323873 , n33448 );
xor ( n33450 , n323843 , n323844 );
and ( n33451 , n33450 , n323846 );
and ( n33452 , n323843 , n323844 );
or ( n323879 , n33451 , n33452 );
buf ( n323880 , n323879 );
not ( n33455 , n831 );
nand ( n33456 , n323880 , n33455 );
nand ( n33457 , n33449 , n33456 );
not ( n323884 , n33457 );
nand ( n323885 , n323872 , n323884 );
and ( n33460 , n33438 , n323885 );
nand ( n33461 , n323763 , n33412 , n33460 );
not ( n323888 , n323789 );
buf ( n323889 , n33367 );
nand ( n33464 , n323888 , n323889 );
not ( n33465 , n33377 );
and ( n33466 , n5980 , n323798 );
not ( n323893 , n5980 );
and ( n323894 , n323893 , n306889 );
or ( n33469 , n33466 , n323894 );
nand ( n33470 , n33465 , n33469 );
nand ( n33471 , n33464 , n33470 );
not ( n323898 , n33471 );
not ( n323899 , n323795 );
not ( n33474 , n323899 );
not ( n323901 , n33474 );
or ( n33476 , n323898 , n323901 );
not ( n33477 , n33408 );
not ( n33478 , n33395 );
or ( n323905 , n33477 , n33478 );
nand ( n323906 , n33376 , n33377 );
nand ( n33481 , n323905 , n323906 );
not ( n33482 , n33481 );
not ( n33483 , n323833 );
and ( n33484 , n5980 , n323817 );
not ( n323911 , n5980 );
and ( n33486 , n323911 , n306861 );
nor ( n33487 , n33484 , n33486 );
not ( n33488 , n33487 );
not ( n323915 , n33488 );
or ( n323916 , n33483 , n323915 );
nand ( n33491 , n5982 , n33386 );
nand ( n33492 , n323916 , n33491 );
nand ( n33493 , n33482 , n33492 , n33474 );
nand ( n323920 , n33476 , n33493 );
buf ( n323921 , n33359 );
nand ( n33496 , n323920 , n323921 , n33460 );
not ( n33497 , n296366 );
nand ( n33498 , n33497 , n33356 );
not ( n33499 , n303205 );
nor ( n323926 , n33499 , n323767 );
and ( n323927 , n33498 , n323926 );
not ( n33502 , n296366 );
nor ( n33503 , n33502 , n33356 );
nor ( n323930 , n323927 , n33503 );
nand ( n323931 , n323841 , n33424 );
not ( n33506 , n323931 );
buf ( n33507 , n323862 );
nand ( n33508 , n33506 , n33507 );
nand ( n323935 , n323867 , n32849 );
not ( n323936 , n323935 );
not ( n33511 , n32849 );
nand ( n33512 , n33511 , n33444 );
not ( n33513 , n33512 );
or ( n323940 , n323936 , n33513 );
buf ( n323941 , n33457 );
nand ( n33516 , n323940 , n323941 );
nand ( n33517 , n323930 , n33508 , n33516 );
not ( n33518 , n323935 );
not ( n323945 , n33512 );
or ( n323946 , n33518 , n323945 );
nand ( n33521 , n323946 , n323941 );
not ( n33522 , n33438 );
and ( n33523 , n33521 , n33522 );
not ( n323950 , n323885 );
nor ( n33525 , n33523 , n323950 );
nand ( n33526 , n33517 , n33525 );
nand ( n33527 , n33461 , n33496 , n33526 );
buf ( n33528 , n33527 );
not ( n33529 , n33528 );
or ( n33530 , n33221 , n33529 );
or ( n33531 , n33220 , n33528 );
nand ( n33532 , n33530 , n33531 );
buf ( n323959 , n33532 );
xor ( n33534 , n33200 , n323627 );
xor ( n33535 , n33534 , n323959 );
buf ( n323962 , n33535 );
xor ( n33537 , n33200 , n323627 );
and ( n33538 , n33537 , n323959 );
and ( n33539 , n33200 , n323627 );
or ( n33540 , n33538 , n33539 );
buf ( n323967 , n33540 );
buf ( n323968 , n313441 );
buf ( n323969 , n24026 );
or ( n33544 , n16425 , n306852 );
nand ( n33545 , n306852 , n16425 );
and ( n33546 , n33544 , n33545 );
not ( n33547 , n831 );
not ( n33548 , n306832 );
or ( n33549 , n33547 , n33548 );
not ( n33550 , n831 );
nand ( n33551 , n33550 , n306781 , n306738 );
nand ( n33552 , n33549 , n33551 );
not ( n33553 , n33552 );
not ( n33554 , n306807 );
not ( n33555 , n306822 );
or ( n33556 , n33554 , n33555 );
nand ( n33557 , n33556 , n306826 );
not ( n33558 , n33557 );
nand ( n33559 , n33553 , n33558 );
not ( n33560 , n33559 );
not ( n33561 , n33219 );
nor ( n33562 , n33560 , n33561 );
not ( n33563 , n33562 );
not ( n33564 , n33527 );
or ( n33565 , n33563 , n33564 );
not ( n33566 , n323641 );
not ( n33567 , n33552 );
nand ( n33568 , n33567 , n33558 );
not ( n33569 , n33568 );
or ( n33570 , n33566 , n33569 );
nand ( n33571 , n33552 , n33557 );
nand ( n33572 , n33570 , n33571 );
not ( n33573 , n33572 );
nand ( n33574 , n33565 , n33573 );
not ( n324001 , n306847 );
nand ( n324002 , n306848 , n324001 );
and ( n33577 , n33574 , n324002 );
nor ( n33578 , n33577 , n17077 );
xnor ( n33579 , n33546 , n33578 );
buf ( n324006 , n33579 );
xor ( n324007 , n323968 , n323969 );
xor ( n324008 , n324007 , n324006 );
buf ( n324009 , n324008 );
xor ( n33584 , n323968 , n323969 );
and ( n33585 , n33584 , n324006 );
and ( n33586 , n323968 , n323969 );
or ( n33587 , n33585 , n33586 );
buf ( n324014 , n33587 );
buf ( n324015 , n315295 );
buf ( n324016 , n317392 );
not ( n33591 , n831 );
not ( n33592 , n304011 );
or ( n33593 , n33591 , n33592 );
nand ( n324020 , n33593 , n310037 );
not ( n33595 , n324020 );
not ( n33596 , n17486 );
not ( n33597 , n831 );
or ( n324024 , n33596 , n33597 );
nand ( n33599 , n310297 , n323752 );
nand ( n33600 , n324024 , n33599 );
not ( n33601 , n33600 );
nand ( n33602 , n33595 , n33601 );
not ( n33603 , n831 );
not ( n33604 , n18033 );
or ( n33605 , n33603 , n33604 );
nand ( n33606 , n310263 , n323486 );
nand ( n33607 , n33605 , n33606 );
or ( n33608 , n297875 , n33607 );
buf ( n33609 , n33608 );
nand ( n33610 , n33602 , n33609 );
not ( n33611 , n33610 );
not ( n33612 , n831 );
not ( n324039 , n308450 );
or ( n33614 , n33612 , n324039 );
nand ( n33615 , n310293 , n5980 );
nand ( n33616 , n33614 , n33615 );
or ( n33617 , n33616 , n309986 );
not ( n324044 , n831 );
not ( n33619 , n308268 );
or ( n33620 , n324044 , n33619 );
nand ( n33621 , n310261 , n323486 );
nand ( n33622 , n33620 , n33621 );
or ( n33623 , n11959 , n33622 );
nand ( n33624 , n33611 , n33617 , n33623 );
not ( n324051 , n33624 );
not ( n33626 , n324051 );
nand ( n33627 , n33461 , n33496 , n33526 );
nand ( n324054 , n307700 , n831 );
nand ( n324055 , n310277 , n5980 );
nand ( n33630 , n324054 , n324055 );
not ( n33631 , n33630 );
not ( n324058 , n831 );
not ( n324059 , n17277 );
or ( n33634 , n324058 , n324059 );
nand ( n33635 , n307610 , n307547 , n296412 );
nand ( n33636 , n33634 , n33635 );
not ( n33637 , n33636 );
nand ( n324064 , n33631 , n33637 );
not ( n324065 , n307616 );
and ( n33640 , n831 , n10413 );
not ( n33641 , n831 );
and ( n33642 , n33641 , n300850 );
nor ( n324069 , n33640 , n33642 );
nand ( n324070 , n324065 , n324069 );
buf ( n324071 , n831 );
not ( n324072 , n324071 );
buf ( n324073 , n303958 );
not ( n33648 , n324073 );
or ( n33649 , n324072 , n33648 );
buf ( n324076 , n831 );
not ( n33651 , n324076 );
buf ( n324078 , n310305 );
nand ( n324079 , n33651 , n324078 );
buf ( n324080 , n324079 );
buf ( n324081 , n324080 );
nand ( n324082 , n33649 , n324081 );
buf ( n324083 , n324082 );
not ( n33658 , n324083 );
not ( n33659 , n307523 );
nand ( n324086 , n33658 , n33659 );
not ( n324087 , n16254 );
nand ( n33662 , n831 , n306684 );
nand ( n33663 , n310303 , n32849 );
nand ( n33664 , n324087 , n33662 , n33663 );
and ( n324091 , n324064 , n324070 , n324086 , n33664 );
nand ( n33666 , n33219 , n33568 );
not ( n33667 , n324001 );
not ( n33668 , n306848 );
or ( n33669 , n33667 , n33668 );
nand ( n33670 , n33669 , n33544 );
nor ( n33671 , n33666 , n33670 );
and ( n33672 , n324091 , n33671 );
buf ( n33673 , n17503 );
not ( n33674 , n831 );
not ( n33675 , n307919 );
or ( n33676 , n33674 , n33675 );
and ( n324103 , n307685 , n307667 );
nand ( n324104 , n324103 , n296412 );
nand ( n33679 , n33676 , n324104 );
not ( n324106 , n33679 );
nand ( n324107 , n33673 , n324106 );
not ( n33682 , n831 );
not ( n324109 , n307938 );
or ( n33684 , n33682 , n324109 );
nand ( n33685 , n33684 , n19614 );
not ( n324112 , n33685 );
and ( n324113 , n323752 , n310273 );
not ( n33688 , n323752 );
and ( n324115 , n33688 , n307941 );
nor ( n324116 , n324113 , n324115 );
nand ( n33691 , n324112 , n324116 );
not ( n324118 , n296412 );
not ( n33693 , n310279 );
or ( n33694 , n324118 , n33693 );
not ( n33695 , n17266 );
and ( n33696 , n307630 , n831 );
nand ( n33697 , n33695 , n33696 );
nand ( n33698 , n33694 , n33697 );
not ( n33699 , n33698 );
not ( n33700 , n831 );
not ( n33701 , n307688 );
or ( n324128 , n33700 , n33701 );
xor ( n33703 , n307667 , n307685 );
nand ( n324130 , n33703 , n323752 );
nand ( n324131 , n324128 , n324130 );
not ( n33706 , n324131 );
nand ( n324133 , n33699 , n33706 );
nand ( n33708 , n324107 , n33691 , n324133 );
not ( n33709 , n33708 );
not ( n324136 , n831 );
not ( n324137 , n307986 );
or ( n33712 , n324136 , n324137 );
nand ( n324139 , n310269 , n5980 );
nand ( n324140 , n33712 , n324139 );
not ( n33715 , n324140 );
not ( n324142 , n302177 );
nand ( n33717 , n33715 , n324142 );
not ( n324144 , n307968 );
nand ( n33719 , n12541 , n302978 , n324144 );
buf ( n324146 , n831 );
not ( n324147 , n324146 );
buf ( n324148 , n307991 );
not ( n33723 , n324148 );
or ( n324150 , n324147 , n33723 );
buf ( n324151 , n831 );
not ( n33726 , n324151 );
buf ( n324153 , n310271 );
nand ( n324154 , n33726 , n324153 );
buf ( n324155 , n324154 );
buf ( n324156 , n324155 );
nand ( n324157 , n324150 , n324156 );
buf ( n324158 , n324157 );
not ( n324159 , n831 );
not ( n33734 , n307994 );
or ( n33735 , n324159 , n33734 );
nand ( n324162 , n310265 , n5980 );
nand ( n324163 , n33735 , n324162 );
or ( n33738 , n324158 , n324163 );
nand ( n324165 , n307971 , n831 );
nand ( n324166 , n310319 , n323752 );
nand ( n33741 , n324165 , n324166 , n17546 );
and ( n324168 , n33717 , n33719 , n33738 , n33741 );
not ( n324169 , n831 );
not ( n33744 , n307955 );
or ( n33745 , n324169 , n33744 );
nand ( n33746 , n310299 , n5980 );
nand ( n324173 , n33745 , n33746 );
or ( n324174 , n324173 , n12698 );
and ( n33749 , n33709 , n324168 , n324174 );
nand ( n324176 , n33627 , n33672 , n33749 );
nand ( n33751 , n33717 , n33719 , n33738 , n33741 );
not ( n33752 , n33751 );
not ( n324179 , n33630 );
not ( n324180 , n33636 );
and ( n33755 , n324179 , n324180 );
nor ( n324182 , n324173 , n12698 );
nor ( n324183 , n33755 , n324182 );
nand ( n33758 , n33752 , n33709 , n324183 );
not ( n324185 , n33758 );
and ( n33760 , n831 , n303958 );
not ( n33761 , n831 );
and ( n324188 , n33761 , n310305 );
or ( n324189 , n33760 , n324188 );
not ( n33764 , n324189 );
not ( n324191 , n307523 );
nor ( n324192 , n324191 , C0 );
not ( n33767 , n324192 );
or ( n324194 , n33764 , n33767 );
not ( n324195 , n831 );
not ( n324196 , n306684 );
or ( n33771 , n324195 , n324196 );
nand ( n324198 , n33771 , n33663 );
nand ( n324199 , n324198 , n16254 );
nand ( n33774 , n324194 , n324199 );
nand ( n324201 , n33658 , n33659 );
nand ( n33776 , n324201 , n324070 );
not ( n33777 , n33776 );
nand ( n324204 , n33774 , n33777 );
not ( n324205 , n324055 );
not ( n33780 , n324054 );
or ( n324207 , n324205 , n33780 );
nand ( n324208 , n324207 , n33636 );
nand ( n33783 , n300856 , n307616 );
nand ( n324210 , n324208 , n33783 );
not ( n33785 , n17077 );
not ( n324212 , n33544 );
or ( n324213 , n33785 , n324212 );
nand ( n33788 , n324213 , n33545 );
nor ( n324215 , n324210 , n33788 );
not ( n324216 , n33670 );
nand ( n33791 , n33572 , n324216 );
nand ( n324218 , n324204 , n324215 , n33791 );
nand ( n33793 , n33777 , n33774 );
nand ( n33794 , n324086 , n33664 , n324070 );
not ( n324221 , n324210 );
nand ( n324222 , n33793 , n33794 , n324221 );
nand ( n33797 , n324185 , n324218 , n324222 );
nand ( n324224 , n33673 , n324106 );
not ( n324225 , n324224 );
nor ( n33800 , n33706 , n33699 );
not ( n324227 , n33800 );
or ( n33802 , n324225 , n324227 );
and ( n324229 , n32849 , n307930 );
not ( n324230 , n32849 );
and ( n33805 , n324230 , n307930 );
or ( n324232 , n324229 , n33805 );
buf ( n33807 , n33679 );
nand ( n33808 , n324232 , n33807 );
nand ( n33809 , n33802 , n33808 );
buf ( n324236 , n33691 );
nand ( n33811 , n33809 , n324236 );
and ( n324238 , n32849 , n310273 );
not ( n33813 , n32849 );
and ( n33814 , n33813 , n307941 );
or ( n324241 , n324238 , n33814 );
nand ( n324242 , n324241 , n33685 );
not ( n33817 , n324242 );
and ( n324244 , n12698 , n324173 );
nor ( n324245 , n33817 , n324244 );
nand ( n33820 , n33811 , n324245 );
nor ( n324247 , n33751 , n324182 );
and ( n324248 , n33820 , n324247 );
nor ( n324249 , n302177 , n324140 );
buf ( n324250 , n831 );
not ( n33825 , n324250 );
buf ( n324252 , n307991 );
not ( n324253 , n324252 );
or ( n33828 , n33825 , n324253 );
buf ( n324255 , n324155 );
nand ( n33830 , n33828 , n324255 );
buf ( n324257 , n33830 );
nor ( n324258 , n324257 , n324163 );
nor ( n324259 , n324249 , n324258 );
not ( n33834 , n324259 );
not ( n324261 , n33741 );
not ( n324262 , n12551 );
nor ( n33837 , n324144 , n324262 );
not ( n324264 , n33837 );
or ( n324265 , n324261 , n324264 );
not ( n33840 , n17547 );
nand ( n324267 , n324165 , n324166 );
nand ( n324268 , n33840 , n324267 );
nand ( n33843 , n324265 , n324268 );
not ( n324270 , n33843 );
or ( n324271 , n33834 , n324270 );
nor ( n33846 , n324142 , n324258 );
buf ( n324273 , n324140 );
and ( n33848 , n33846 , n324273 );
nand ( n33849 , n324158 , n324163 );
not ( n324276 , n33849 );
nor ( n324277 , n33848 , n324276 );
nand ( n33852 , n324271 , n324277 );
nor ( n324279 , n324248 , n33852 );
nand ( n324280 , n33797 , n324279 );
not ( n33855 , n324280 );
nand ( n324282 , n324176 , n33855 );
not ( n324283 , n324282 );
or ( n33858 , n33626 , n324283 );
not ( n33859 , n33617 );
not ( n33860 , n33623 );
not ( n324287 , n33608 );
nand ( n33862 , n324020 , n33600 );
not ( n33863 , n33862 );
not ( n33864 , n33863 );
or ( n324291 , n324287 , n33864 );
not ( n324292 , n5980 );
not ( n33867 , n297871 );
or ( n324294 , n324292 , n33867 );
nand ( n324295 , n324294 , n7446 );
buf ( n33870 , n33607 );
nand ( n324297 , n324295 , n33870 );
nand ( n33872 , n324291 , n324297 );
not ( n33873 , n33872 );
or ( n324300 , n33860 , n33873 );
nand ( n324301 , n11959 , n33622 );
nand ( n33876 , n324300 , n324301 );
not ( n324303 , n33876 );
or ( n324304 , n33859 , n324303 );
nand ( n33879 , n309986 , n33616 );
nand ( n324306 , n324304 , n33879 );
not ( n324307 , n324306 );
nand ( n33882 , n33858 , n324307 );
not ( n33883 , n296412 );
not ( n33884 , n310295 );
or ( n33885 , n33883 , n33884 );
nand ( n33886 , n831 , n308469 );
nand ( n33887 , n33885 , n33886 );
not ( n324314 , n831 );
not ( n33889 , n308638 );
or ( n324316 , n324314 , n33889 );
buf ( n324317 , n308475 );
buf ( n324318 , n308637 );
xor ( n324319 , n324317 , n324318 );
buf ( n324320 , n324319 );
nand ( n33895 , n324320 , n5980 );
nand ( n33896 , n324316 , n33895 );
and ( n33897 , n33887 , n33896 );
not ( n33898 , n33897 );
or ( n324325 , n33887 , n33896 );
nand ( n33900 , n33898 , n324325 );
not ( n33901 , n33900 );
and ( n33902 , n33882 , n33901 );
not ( n324329 , n33882 );
and ( n324330 , n324329 , n33900 );
nor ( n33905 , n33902 , n324330 );
buf ( n324332 , n33905 );
xor ( n33907 , n324015 , n324016 );
xor ( n33908 , n33907 , n324332 );
buf ( n324335 , n33908 );
xor ( n33910 , n324015 , n324016 );
and ( n33911 , n33910 , n324332 );
and ( n324338 , n324015 , n324016 );
or ( n33913 , n33911 , n324338 );
buf ( n324340 , n33913 );
buf ( n324341 , n322984 );
nand ( n33916 , n323076 , n32756 );
xnor ( n33917 , n323178 , n33916 );
buf ( n324344 , n33917 );
xor ( n324345 , n324341 , n324344 );
buf ( n324346 , n324345 );
and ( n33921 , n324341 , n324344 );
buf ( n324348 , n33921 );
buf ( n324349 , n322566 );
xor ( n33924 , n322526 , n322530 );
xor ( n324351 , n33924 , n322537 );
and ( n33926 , n322778 , n324351 );
xor ( n33927 , n322526 , n322530 );
xor ( n324354 , n33927 , n322537 );
and ( n324355 , n322576 , n324354 );
and ( n33930 , n322778 , n322576 );
or ( n324357 , n33926 , n324355 , n33930 );
buf ( n324358 , n324357 );
xor ( n33933 , n324349 , n324358 );
buf ( n324360 , n33933 );
and ( n33935 , n324349 , n324358 );
buf ( n324362 , n33935 );
buf ( n324363 , n322625 );
buf ( n324364 , n322571 );
xor ( n33939 , n324363 , n324364 );
buf ( n324366 , n33939 );
and ( n33941 , n324363 , n324364 );
buf ( n324368 , n33941 );
buf ( n324369 , n322801 );
buf ( n324370 , n322630 );
xor ( n33945 , n324369 , n324370 );
buf ( n324372 , n33945 );
and ( n33947 , n324369 , n324370 );
buf ( n324374 , n33947 );
buf ( n324375 , n322806 );
buf ( n324376 , n322878 );
xor ( n33951 , n324375 , n324376 );
buf ( n324378 , n33951 );
and ( n33953 , n831 , n308842 );
not ( n33954 , n831 );
and ( n33955 , n324317 , n324318 );
buf ( n324382 , n33955 );
and ( n33957 , n33954 , n324382 );
or ( n33958 , n33953 , n33957 );
not ( n324385 , n33958 );
and ( n33960 , n831 , n18413 );
not ( n33961 , n831 );
and ( n33962 , n33961 , n310257 );
nor ( n324389 , n33960 , n33962 );
nand ( n324390 , n324385 , n324389 );
not ( n33965 , n296412 );
not ( n33966 , n310259 );
or ( n33967 , n33965 , n33966 );
nand ( n324394 , n309709 , n831 );
nand ( n324395 , n33967 , n324394 );
not ( n33970 , n831 );
not ( n33971 , n309721 );
or ( n33972 , n33970 , n33971 );
nand ( n324399 , n310251 , n323486 );
nand ( n324400 , n33972 , n324399 );
or ( n33975 , n324395 , n324400 );
and ( n33976 , n324325 , n324390 , n33975 );
not ( n33977 , n33610 );
not ( n324404 , n309793 );
nor ( n33979 , n324404 , C0 );
not ( n33980 , n831 );
not ( n33981 , n309795 );
or ( n33982 , n33980 , n33981 );
not ( n33983 , n831 );
nand ( n33984 , n33983 , n310253 );
nand ( n324411 , n33982 , n33984 );
or ( n33986 , n33979 , n324411 );
and ( n33987 , n33623 , n33986 );
and ( n33988 , n33977 , n33987 , n33617 );
buf ( n33989 , n309531 );
not ( n324416 , n831 );
not ( n324417 , n309533 );
or ( n33992 , n324416 , n324417 );
nand ( n324419 , n310245 , n323057 );
nand ( n33994 , n33992 , n324419 );
or ( n324421 , n33989 , n33994 );
not ( n33996 , n309562 );
nor ( n33997 , n33996 , C0 );
not ( n33998 , n5980 );
not ( n33999 , n19128 );
or ( n324426 , n33998 , n33999 );
nand ( n34001 , n19128 , n831 );
nand ( n34002 , n324426 , n34001 );
or ( n34003 , n33997 , n34002 );
and ( n34004 , n324421 , n34003 );
nand ( n34005 , n33976 , n33988 , n34004 );
not ( n34006 , n310287 );
not ( n34007 , n323486 );
or ( n324434 , n34006 , n34007 );
nand ( n34009 , n309386 , n831 );
nand ( n34010 , n324434 , n34009 );
not ( n34011 , n296412 );
not ( n34012 , n310247 );
or ( n324439 , n34011 , n34012 );
nand ( n34014 , n309305 , n831 );
nand ( n34015 , n324439 , n34014 );
nor ( n34016 , n34010 , n34015 );
nor ( n324443 , n34005 , n34016 );
nand ( n324444 , n324176 , n33855 );
buf ( n34019 , n324444 );
nand ( n34020 , n324443 , n34019 );
not ( n34021 , n34016 );
not ( n324448 , n34021 );
not ( n34023 , n34004 );
not ( n34024 , n324411 );
not ( n34025 , n33979 );
and ( n34026 , n34024 , n34025 );
nand ( n324453 , n324325 , n324390 , n33975 );
nor ( n34028 , n34026 , n324453 );
not ( n34029 , n34028 );
not ( n34030 , n33617 );
not ( n34031 , n33876 );
or ( n34032 , n34030 , n34031 );
nand ( n324459 , n34032 , n33879 );
not ( n34034 , n324459 );
or ( n34035 , n34029 , n34034 );
nand ( n34036 , n33979 , n324411 );
nand ( n34037 , n324395 , n324400 );
nand ( n34038 , n33897 , n324390 );
not ( n34039 , n324389 );
nand ( n34040 , n34039 , n33958 );
nand ( n34041 , n34036 , n34037 , n34038 , n34040 );
not ( n34042 , n33975 );
and ( n34043 , n34042 , n34037 , n34036 );
nor ( n34044 , n33979 , n324411 );
nor ( n34045 , n34043 , n34044 );
nand ( n34046 , n34041 , n34045 );
nand ( n34047 , n34035 , n34046 );
not ( n34048 , n34047 );
or ( n34049 , n34023 , n34048 );
and ( n34050 , n34002 , n33997 );
and ( n34051 , n34050 , n324421 );
and ( n34052 , n33989 , n33994 );
nor ( n34053 , n34051 , n34052 );
nand ( n34054 , n34049 , n34053 );
not ( n34055 , n34054 );
or ( n34056 , n324448 , n34055 );
nand ( n34057 , n34015 , n34010 );
nand ( n34058 , n34056 , n34057 );
not ( n34059 , n34058 );
nand ( n34060 , n34020 , n34059 );
not ( n34061 , n322345 );
not ( n34062 , n321612 );
not ( n34063 , n34062 );
or ( n34064 , n34061 , n34063 );
not ( n34065 , n322345 );
nand ( n34066 , n321612 , n34065 );
nand ( n34067 , n34064 , n34066 );
not ( n34068 , n322264 );
and ( n34069 , n34067 , n34068 );
not ( n34070 , n34067 );
and ( n34071 , n34070 , n322264 );
nor ( n34072 , n34069 , n34071 );
xor ( n34073 , n322183 , n322202 );
xor ( n34074 , n34073 , n322211 );
xor ( n34075 , n322177 , n322255 );
xor ( n34076 , n34074 , n34075 );
not ( n34077 , n34076 );
not ( n34078 , n321607 );
or ( n34079 , n34077 , n34078 );
not ( n34080 , n34076 );
not ( n34081 , n34080 );
not ( n34082 , n321607 );
not ( n34083 , n34082 );
or ( n34084 , n34081 , n34083 );
nand ( n34085 , n34084 , n322023 );
nand ( n34086 , n34079 , n34085 );
not ( n34087 , n34086 );
nand ( n34088 , n34072 , n34087 );
and ( n34089 , n831 , n309389 );
not ( n34090 , n831 );
and ( n34091 , n34090 , n310289 );
or ( n34092 , n34089 , n34091 );
and ( n34093 , n831 , n309461 );
not ( n34094 , n831 );
and ( n34095 , n34094 , n310309 );
or ( n324522 , n34093 , n34095 );
nor ( n324523 , n34092 , n324522 );
not ( n34098 , n324523 );
nand ( n324525 , n34092 , n324522 );
nand ( n324526 , n34098 , n324525 );
and ( n34101 , n34088 , n324526 );
nand ( n324528 , n34060 , n34101 );
not ( n34103 , n324526 );
nand ( n34104 , n34103 , n34088 );
nor ( n324531 , n34058 , n34104 );
and ( n324532 , n324531 , n34020 );
not ( n34107 , n34072 );
and ( n324534 , n34107 , n34086 );
nor ( n324535 , n324532 , n324534 );
and ( n34110 , n324528 , n324535 );
not ( n324537 , n34110 );
not ( n34112 , n33976 );
nand ( n324539 , n33617 , n33977 , n33987 );
nor ( n324540 , n34112 , n324539 );
not ( n34115 , n324523 );
and ( n324542 , n34021 , n34004 , n34115 );
and ( n324543 , n324540 , n324542 );
not ( n34118 , n324543 );
nand ( n324545 , n324176 , n33855 );
not ( n34120 , n324545 );
or ( n34121 , n34118 , n34120 );
not ( n324548 , n34028 );
not ( n324549 , n324459 );
or ( n34124 , n324548 , n324549 );
nand ( n324551 , n34124 , n34046 );
and ( n324552 , n324551 , n324542 );
not ( n34127 , n34115 );
not ( n324554 , n34015 );
not ( n34129 , n34010 );
or ( n34130 , n324554 , n34129 );
or ( n34131 , n34053 , n34016 );
nand ( n324558 , n34130 , n34131 );
not ( n324559 , n324558 );
or ( n34134 , n34127 , n324559 );
nand ( n324561 , n34134 , n324525 );
nor ( n34136 , n324552 , n324561 );
nand ( n324563 , n34121 , n34136 );
buf ( n324564 , n324563 );
not ( n324565 , n5980 );
not ( n324566 , n310311 );
or ( n34141 , n324565 , n324566 );
nand ( n324568 , n309575 , n831 );
nand ( n324569 , n34141 , n324568 );
not ( n324570 , n831 );
not ( n34145 , n309640 );
or ( n324572 , n324570 , n34145 );
nand ( n34147 , n310315 , n5980 );
nand ( n324574 , n324572 , n34147 );
or ( n324575 , n324569 , n324574 );
nand ( n34150 , n324569 , n324574 );
nand ( n324577 , n324575 , n34150 );
not ( n324578 , n324577 );
not ( n34153 , n324578 );
nand ( n324580 , n34062 , n34065 );
not ( n34155 , n324580 );
not ( n34156 , n322264 );
or ( n324583 , n34155 , n34156 );
nand ( n324584 , n321612 , n322345 );
nand ( n34159 , n324583 , n324584 );
xor ( n324586 , n321969 , n321985 );
xor ( n324587 , n324586 , n31566 );
xor ( n34162 , n322857 , n322644 );
xor ( n324589 , n324587 , n34162 );
xor ( n34164 , n322350 , n324589 );
xor ( n34165 , n34164 , n322269 );
and ( n34166 , n34159 , n34165 );
not ( n34167 , n34159 );
not ( n34168 , n34165 );
and ( n34169 , n34167 , n34168 );
nor ( n34170 , n34166 , n34169 );
not ( n324597 , n34170 );
or ( n324598 , n34153 , n324597 );
or ( n34173 , n34170 , n324578 );
nand ( n324600 , n324598 , n34173 );
and ( n34175 , n324564 , n324600 );
not ( n34176 , n324564 );
not ( n34177 , n324577 );
not ( n34178 , n34170 );
or ( n34179 , n34177 , n34178 );
or ( n34180 , n34170 , n324577 );
nand ( n34181 , n34179 , n34180 );
and ( n34182 , n34176 , n34181 );
or ( n34183 , n34175 , n34182 );
nand ( n34184 , n324537 , n34183 );
not ( n34185 , n34183 );
nand ( n34186 , n34110 , n34185 );
nand ( n34187 , n34184 , n34186 );
buf ( n324614 , n34187 );
buf ( n324615 , n34187 );
not ( n34190 , n324615 );
buf ( n324617 , n34190 );
buf ( n324618 , n324617 );
and ( n324619 , n34072 , n34086 );
not ( n34194 , n34072 );
and ( n34195 , n34194 , n34087 );
nor ( n34196 , n324619 , n34195 );
not ( n324623 , n324526 );
and ( n34198 , n34196 , n324623 );
not ( n324625 , n34196 );
and ( n34200 , n324625 , n324526 );
or ( n34201 , n34198 , n34200 );
not ( n324628 , n34201 );
and ( n34203 , n34060 , n324628 );
not ( n34204 , n34060 );
and ( n34205 , n34204 , n34201 );
nor ( n324632 , n34203 , n34205 );
buf ( n34207 , n34054 );
not ( n34208 , n34207 );
not ( n34209 , n34005 );
nand ( n324636 , n34209 , n34019 );
nand ( n324637 , n34208 , n324636 );
not ( n34212 , n324637 );
not ( n34213 , n320665 );
not ( n34214 , n34076 );
not ( n34215 , n34082 );
or ( n34216 , n34214 , n34215 );
nand ( n34217 , n321607 , n34080 );
nand ( n324644 , n34216 , n34217 );
not ( n324645 , n322023 );
and ( n34220 , n324644 , n324645 );
not ( n34221 , n324644 );
and ( n34222 , n34221 , n322023 );
nor ( n324649 , n34220 , n34222 );
nand ( n34224 , n34213 , n324649 );
not ( n34225 , n34224 );
nand ( n324652 , n34021 , n34057 );
nor ( n324653 , n34225 , n324652 );
nand ( n34228 , n34212 , n324653 );
not ( n34229 , n324652 );
not ( n324656 , n34229 );
nand ( n324657 , n324656 , n324637 , n34224 );
not ( n34232 , n324649 );
nand ( n34233 , n320665 , n34232 );
and ( n324660 , n34228 , n324657 , n34233 );
nand ( n324661 , n324632 , n324660 );
buf ( n324662 , n324661 );
buf ( n34237 , n324662 );
buf ( n324664 , n34237 );
buf ( n324665 , n324664 );
not ( n34240 , n324665 );
xor ( n34241 , n318272 , n318277 );
xor ( n324668 , n34241 , n318283 );
and ( n324669 , n27862 , n324668 );
xor ( n324670 , n318272 , n318277 );
xor ( n324671 , n324670 , n318283 );
and ( n34246 , n318293 , n324671 );
and ( n324673 , n27862 , n318293 );
or ( n324674 , n324669 , n34246 , n324673 );
xor ( n34249 , n319890 , n29468 );
xor ( n324676 , n34249 , n319898 );
and ( n34251 , n324674 , n324676 );
xor ( n34252 , n318347 , n318416 );
xor ( n324679 , n34252 , n318464 );
and ( n324680 , n318473 , n324679 );
xor ( n324681 , n318347 , n318416 );
xor ( n34256 , n324681 , n318464 );
and ( n324683 , n318478 , n34256 );
and ( n324684 , n318473 , n318478 );
or ( n34259 , n324680 , n324683 , n324684 );
xor ( n324686 , n319890 , n29468 );
xor ( n324687 , n324686 , n319898 );
and ( n34262 , n34259 , n324687 );
and ( n324689 , n324674 , n34259 );
or ( n324690 , n34251 , n34262 , n324689 );
or ( n324691 , n324690 , n319905 );
not ( n34266 , n324691 );
not ( n324693 , n324540 );
not ( n34268 , n324545 );
or ( n34269 , n324693 , n34268 );
not ( n324696 , n324551 );
nand ( n324697 , n34269 , n324696 );
not ( n324698 , n324697 );
not ( n34273 , n324698 );
not ( n324700 , n34050 );
nand ( n324701 , n324700 , n34003 );
or ( n34276 , n34273 , n324701 );
nand ( n324703 , n34273 , n324701 );
nand ( n324704 , n34276 , n324703 );
not ( n34279 , n324704 );
or ( n324706 , n34266 , n34279 );
nand ( n324707 , n324690 , n319905 );
nand ( n34282 , n324706 , n324707 );
not ( n324709 , n34282 );
not ( n324710 , n34052 );
nand ( n34285 , n324710 , n324421 );
and ( n324712 , n34285 , n34003 );
not ( n34287 , n324712 );
not ( n324714 , n324697 );
or ( n324715 , n34287 , n324714 );
nand ( n324716 , n34285 , n34050 );
not ( n324717 , n324716 );
nor ( n34292 , n34285 , n34003 , n34050 );
nor ( n324719 , n324717 , n34292 );
nand ( n324720 , n324715 , n324719 );
not ( n324721 , n324720 );
nor ( n34296 , n34285 , n34050 );
nand ( n324723 , n324698 , n34296 );
nand ( n324724 , n324721 , n324723 );
not ( n34299 , n324724 );
xnor ( n324726 , n320660 , n319910 );
not ( n324727 , n324726 );
and ( n34302 , n34299 , n324727 );
buf ( n324729 , n324724 );
and ( n34304 , n324729 , n324726 );
nor ( n324731 , n34302 , n34304 );
nand ( n34306 , n324709 , n324731 );
xor ( n34307 , n34076 , n321607 );
xor ( n324734 , n34307 , n324645 );
not ( n324735 , n324734 );
not ( n324736 , n320665 );
or ( n34311 , n324735 , n324736 );
or ( n324738 , n320665 , n324649 );
nand ( n324739 , n34311 , n324738 );
not ( n34314 , n324739 );
and ( n324741 , n324652 , n34314 );
not ( n324742 , n324652 );
not ( n34317 , n324739 );
not ( n324744 , n34317 );
and ( n324745 , n324742 , n324744 );
or ( n324746 , n324741 , n324745 );
and ( n34321 , n324637 , n324746 );
not ( n324748 , n324637 );
not ( n34323 , n324739 );
and ( n34324 , n34229 , n34323 );
not ( n324751 , n34229 );
not ( n324752 , n34317 );
and ( n324753 , n324751 , n324752 );
or ( n34328 , n34324 , n324753 );
and ( n324755 , n324748 , n34328 );
or ( n324756 , n34321 , n324755 );
not ( n34331 , n324756 );
or ( n324758 , n320660 , n319910 );
not ( n324759 , n324758 );
not ( n34334 , n324724 );
or ( n324761 , n324759 , n34334 );
nand ( n324762 , n320660 , n319910 );
nand ( n34337 , n324761 , n324762 );
not ( n34338 , n34337 );
nand ( n324765 , n34331 , n34338 );
nand ( n324766 , n34306 , n324765 );
buf ( n324767 , n324766 );
nor ( n324768 , n34240 , n324767 );
buf ( n324769 , n324768 );
buf ( n324770 , n324769 );
not ( n324771 , n324770 );
xnor ( n34346 , n319905 , n324690 );
not ( n324773 , n34346 );
not ( n34348 , n324704 );
or ( n34349 , n324773 , n34348 );
not ( n324776 , n34273 );
not ( n34351 , n324701 );
nand ( n34352 , n324776 , n34351 );
xor ( n34353 , n319905 , n324690 );
nand ( n324780 , n34352 , n34353 , n324703 );
nand ( n324781 , n34349 , n324780 );
xor ( n34356 , n319890 , n29468 );
xor ( n34357 , n34356 , n319898 );
xor ( n34358 , n324674 , n34259 );
xor ( n324785 , n34357 , n34358 );
or ( n324786 , n318489 , n324785 );
not ( n324787 , n324786 );
not ( n324788 , n34044 );
nand ( n34363 , n324788 , n34036 );
not ( n324790 , n34363 );
and ( n324791 , n324325 , n324390 );
not ( n34366 , n324791 );
nor ( n324793 , n34366 , n33624 );
nand ( n324794 , n324444 , n324793 );
or ( n34369 , n34042 , n324794 );
nand ( n324796 , n324306 , n324791 );
not ( n324797 , n324796 );
not ( n34372 , n34042 );
and ( n324799 , n324797 , n34372 );
and ( n34374 , n34040 , n34038 );
or ( n34375 , n34374 , n34042 );
nand ( n324802 , n34375 , n34037 );
nor ( n324803 , n324799 , n324802 );
nand ( n324804 , n34369 , n324803 );
not ( n34379 , n324804 );
or ( n324806 , n324790 , n34379 );
or ( n324807 , n34042 , n324794 );
not ( n34382 , n34363 );
nand ( n324809 , n324807 , n324803 , n34382 );
nand ( n324810 , n324806 , n324809 );
not ( n34385 , n324810 );
or ( n324812 , n324787 , n34385 );
nand ( n324813 , n318489 , n324785 );
nand ( n34388 , n324812 , n324813 );
nor ( n34389 , n324781 , n34388 );
or ( n324816 , n318484 , n317637 );
not ( n324817 , n324816 );
nand ( n34392 , n33975 , n34037 );
not ( n324819 , n34392 );
and ( n34394 , n324796 , n34374 );
nand ( n324821 , n324794 , n34394 );
and ( n34396 , n324819 , n324821 );
not ( n34397 , n324819 );
not ( n324824 , n324821 );
and ( n324825 , n34397 , n324824 );
nor ( n34400 , n34396 , n324825 );
not ( n324827 , n34400 );
or ( n324828 , n324817 , n324827 );
nand ( n34403 , n318484 , n317637 );
nand ( n324830 , n324828 , n34403 );
xor ( n324831 , n318489 , n324785 );
not ( n34406 , n324831 );
not ( n324833 , n324810 );
not ( n324834 , n324833 );
or ( n34409 , n34406 , n324834 );
not ( n324836 , n324831 );
nand ( n324837 , n324836 , n324810 );
nand ( n324838 , n34409 , n324837 );
nor ( n324839 , n324830 , n324838 );
nor ( n34414 , n34389 , n324839 );
nand ( n324841 , n34040 , n324390 );
xor ( n324842 , n317397 , n317632 );
xor ( n34417 , n324841 , n324842 );
nand ( n324844 , n324051 , n324325 , n324282 );
and ( n34419 , n324306 , n324325 );
nor ( n34420 , n34419 , n33897 );
nand ( n324847 , n324844 , n34420 );
xnor ( n324848 , n34417 , n324847 );
not ( n324849 , n324848 );
not ( n34424 , n324340 );
and ( n324851 , n324849 , n34424 );
xor ( n324852 , n317637 , n318484 );
not ( n34427 , n324852 );
not ( n324854 , n324821 );
or ( n324855 , n34427 , n324854 );
not ( n34430 , n324852 );
nand ( n324857 , n34430 , n324794 , n34394 );
nand ( n324858 , n324855 , n324857 );
and ( n34433 , n324858 , n324819 );
not ( n324860 , n324858 );
and ( n324861 , n324860 , n34392 );
nor ( n34436 , n34433 , n324861 );
nor ( n324863 , n317397 , n317632 );
nor ( n324864 , n324841 , n324863 );
and ( n34439 , n324844 , n34420 , n324864 );
and ( n324866 , n317397 , n317632 );
nor ( n34441 , n34439 , n324866 );
not ( n34442 , n324841 );
nor ( n324869 , n34442 , n324863 );
nand ( n324870 , n324869 , n324847 );
and ( n324871 , n34441 , n324870 );
and ( n34446 , n34436 , n324871 );
nor ( n324873 , n324851 , n34446 );
nand ( n324874 , n34414 , n324873 );
buf ( n34449 , n324874 );
buf ( n324876 , n34449 );
nor ( n324877 , n324771 , n324876 );
buf ( n324878 , n324877 );
buf ( n324879 , n324878 );
not ( n324880 , n324879 );
nand ( n34455 , n33709 , n324174 );
nand ( n34456 , n302978 , n12541 , n324144 );
not ( n324883 , n34456 );
nor ( n324884 , n34455 , n324883 );
not ( n34459 , n324884 );
not ( n324886 , n324216 );
not ( n324887 , n33572 );
or ( n34462 , n324886 , n324887 );
not ( n324889 , n33788 );
nand ( n324890 , n34462 , n324889 );
not ( n34465 , n324890 );
not ( n324892 , n34465 );
not ( n34467 , n324091 );
not ( n34468 , n34467 );
and ( n324895 , n324892 , n34468 );
nand ( n324896 , n33631 , n33637 );
not ( n324897 , n324896 );
buf ( n34472 , n33783 );
nand ( n324899 , n324204 , n34472 );
not ( n324900 , n324899 );
or ( n34475 , n324897 , n324900 );
buf ( n324902 , n324208 );
nand ( n324903 , n34475 , n324902 );
nor ( n34478 , n324895 , n324903 );
nand ( n324905 , n33627 , n33672 );
nand ( n324906 , n34478 , n324905 );
not ( n34481 , n324906 );
or ( n324908 , n34459 , n34481 );
not ( n324909 , n324174 );
not ( n34484 , n324236 );
not ( n324911 , n33809 );
or ( n324912 , n34484 , n324911 );
and ( n34487 , n5980 , n310273 );
not ( n324914 , n5980 );
and ( n34489 , n324914 , n307941 );
or ( n324916 , n34487 , n34489 );
buf ( n34491 , n33685 );
nand ( n34492 , n324916 , n34491 );
nand ( n324919 , n324912 , n34492 );
not ( n324920 , n324919 );
or ( n34495 , n324909 , n324920 );
nand ( n324922 , n12698 , n324173 );
nand ( n324923 , n34495 , n324922 );
and ( n34498 , n324923 , n34456 );
buf ( n324925 , n33837 );
nor ( n324926 , n34498 , n324925 );
nand ( n324927 , n324908 , n324926 );
nand ( n324928 , n324268 , n33741 );
not ( n34503 , n324928 );
and ( n324930 , n324927 , n34503 );
not ( n324931 , n324927 );
and ( n34506 , n324931 , n324928 );
nor ( n324933 , n324930 , n34506 );
xor ( n34508 , n311065 , n311077 );
xor ( n34509 , n34508 , n311090 );
xor ( n324936 , n311957 , n311963 );
xor ( n324937 , n34509 , n324936 );
xor ( n34512 , n320979 , n324937 );
and ( n324939 , n34512 , n322026 );
and ( n324940 , n320979 , n324937 );
or ( n34515 , n324939 , n324940 );
xor ( n324942 , n34515 , n318237 );
not ( n324943 , n318158 );
not ( n34518 , n318139 );
or ( n324945 , n324943 , n34518 );
nand ( n34520 , n318140 , n318157 );
nand ( n324947 , n324945 , n34520 );
and ( n34522 , n324947 , n318225 );
not ( n34523 , n324947 );
not ( n324950 , n318225 );
and ( n324951 , n34523 , n324950 );
nor ( n34526 , n34522 , n324951 );
not ( n324953 , n34526 );
not ( n324954 , n321017 );
nand ( n34529 , n324953 , n324954 );
not ( n324956 , n34529 );
xor ( n324957 , n320979 , n324937 );
xor ( n34532 , n324957 , n322026 );
not ( n324959 , n34532 );
not ( n324960 , n324959 );
not ( n34535 , n324960 );
or ( n324962 , n324956 , n34535 );
and ( n324963 , n321017 , n34526 );
not ( n34538 , n324963 );
nand ( n324965 , n324962 , n34538 );
and ( n324966 , n324942 , n324965 );
and ( n324967 , n34515 , n318237 );
or ( n34542 , n324966 , n324967 );
xor ( n324969 , n320671 , n318132 );
xor ( n324970 , n324969 , n318242 );
xor ( n34545 , n34542 , n324970 );
and ( n34546 , n324933 , n34545 );
not ( n324973 , n324933 );
not ( n34548 , n34545 );
and ( n324975 , n324973 , n34548 );
nor ( n324976 , n34546 , n324975 );
not ( n34551 , n324976 );
xor ( n34552 , n34515 , n318237 );
xor ( n324979 , n34552 , n324965 );
not ( n324980 , n324979 );
not ( n324981 , n321012 );
not ( n34556 , n321040 );
nand ( n34557 , n324981 , n34556 );
not ( n324984 , n34557 );
not ( n34559 , n320739 );
or ( n324986 , n324984 , n34559 );
nand ( n324987 , n321012 , n321040 );
nand ( n34562 , n324986 , n324987 );
not ( n34563 , n34562 );
not ( n324990 , n324954 );
and ( n324991 , n34532 , n324953 );
not ( n34566 , n34532 );
and ( n34567 , n34566 , n34526 );
nor ( n34568 , n324991 , n34567 );
not ( n34569 , n34568 );
not ( n324996 , n34569 );
or ( n324997 , n324990 , n324996 );
or ( n324998 , n34569 , n324954 );
nand ( n34573 , n324997 , n324998 );
not ( n325000 , n34573 );
or ( n325001 , n34563 , n325000 );
not ( n34576 , n322031 );
not ( n325003 , n321617 );
or ( n34578 , n34576 , n325003 );
or ( n325005 , n322031 , n321617 );
nand ( n325006 , n325005 , n320974 );
nand ( n34581 , n34578 , n325006 );
buf ( n325008 , n34581 );
nand ( n34583 , n34562 , n325008 );
nor ( n34584 , n34526 , n324954 );
nand ( n34585 , n324959 , n34584 , n325008 );
nand ( n325012 , n325008 , n324963 , n324960 );
and ( n325013 , n34585 , n325012 );
not ( n325014 , n34529 );
and ( n34589 , n324960 , n325014 , n325008 );
nand ( n325016 , n34526 , n34581 , n324954 );
nor ( n325017 , n324960 , n325016 );
nor ( n34592 , n34589 , n325017 );
and ( n325019 , n34583 , n325013 , n34592 );
nand ( n34594 , n325001 , n325019 );
not ( n34595 , n34594 );
or ( n325022 , n324980 , n34595 );
not ( n325023 , n34455 );
not ( n34598 , n325023 );
not ( n325025 , n324906 );
or ( n34600 , n34598 , n325025 );
not ( n34601 , n324923 );
nand ( n34602 , n34600 , n34601 );
nor ( n325029 , n324883 , n324925 );
or ( n325030 , n34602 , n325029 );
or ( n325031 , n34594 , n324979 );
not ( n34606 , n34602 );
not ( n325033 , n325029 );
or ( n325034 , n34606 , n325033 );
nand ( n34609 , n325030 , n325031 , n325034 );
nand ( n325036 , n325022 , n34609 );
not ( n34611 , n325036 );
nand ( n34612 , n34551 , n34611 );
not ( n325039 , n324335 );
not ( n34614 , n33623 );
nor ( n34615 , n34614 , n33610 );
not ( n325042 , n34615 );
not ( n325043 , n34019 );
or ( n34618 , n325042 , n325043 );
not ( n325045 , n33876 );
nand ( n325046 , n34618 , n325045 );
or ( n34621 , n315290 , n315714 );
not ( n325048 , n34621 );
nand ( n325049 , n33617 , n33879 );
not ( n34624 , n325049 );
or ( n325051 , n325048 , n34624 );
nand ( n34626 , n315290 , n315714 );
nand ( n34627 , n325051 , n34626 );
and ( n325054 , n325046 , n34627 );
not ( n325055 , n325046 );
not ( n34630 , n34621 );
not ( n325057 , n325049 );
not ( n325058 , n325057 );
or ( n325059 , n34630 , n325058 );
nand ( n34634 , n325059 , n34626 );
and ( n325061 , n325055 , n34634 );
or ( n325062 , n325054 , n325061 );
not ( n34637 , n325062 );
nand ( n325064 , n325039 , n34637 );
or ( n325065 , n34542 , n324970 );
not ( n325066 , n325065 );
not ( n34641 , n324933 );
or ( n325068 , n325066 , n34641 );
nand ( n34643 , n34542 , n324970 );
nand ( n34644 , n325068 , n34643 );
not ( n325071 , n34644 );
xor ( n325072 , n320671 , n318132 );
and ( n325073 , n325072 , n318242 );
and ( n34648 , n320671 , n318132 );
or ( n325075 , n325073 , n34648 );
xor ( n325076 , n312275 , n325075 );
not ( n34651 , n325076 );
and ( n325078 , n34456 , n33741 );
and ( n325079 , n325023 , n325078 );
not ( n34654 , n325079 );
not ( n325081 , n324906 );
or ( n325082 , n34654 , n325081 );
and ( n34657 , n324923 , n325078 );
buf ( n325084 , n33843 );
nor ( n34659 , n34657 , n325084 );
nand ( n325086 , n325082 , n34659 );
buf ( n34661 , n324273 );
not ( n34662 , n324142 );
nand ( n325089 , n34661 , n34662 );
not ( n34664 , n324249 );
and ( n325091 , n325089 , n34664 );
and ( n34666 , n325086 , n325091 );
not ( n325093 , n325086 );
not ( n325094 , n34661 );
not ( n34669 , n34662 );
or ( n325096 , n325094 , n34669 );
nand ( n325097 , n325096 , n34664 );
and ( n34672 , n325093 , n325097 );
nor ( n325099 , n34666 , n34672 );
not ( n325100 , n325099 );
not ( n34675 , n325100 );
or ( n325102 , n34651 , n34675 );
not ( n325103 , n325076 );
nand ( n34678 , n325103 , n325099 );
nand ( n325105 , n325102 , n34678 );
not ( n325106 , n325105 );
nand ( n34681 , n325071 , n325106 );
nand ( n34682 , n33609 , n324297 );
and ( n34683 , n34682 , n33602 );
not ( n325110 , n34683 );
not ( n325111 , n34019 );
or ( n34686 , n325110 , n325111 );
or ( n34687 , n34682 , n33863 );
nor ( n34688 , n34019 , n34687 );
or ( n325115 , n34682 , n33602 , n33863 );
nand ( n325116 , n34682 , n33863 );
nand ( n34691 , n325115 , n325116 );
nor ( n325118 , n34688 , n34691 );
nand ( n34693 , n34686 , n325118 );
xor ( n34694 , n314315 , n314380 );
and ( n34695 , n34693 , n34694 );
not ( n34696 , n34693 );
xnor ( n325123 , n314315 , n314380 );
and ( n325124 , n34696 , n325123 );
nor ( n34699 , n34695 , n325124 );
not ( n325126 , n34699 );
not ( n34701 , n314358 );
not ( n34702 , n314375 );
or ( n34703 , n34701 , n34702 );
not ( n34704 , n314358 );
not ( n34705 , n314375 );
and ( n325132 , n34704 , n34705 );
not ( n325133 , n325132 );
and ( n34708 , n33862 , n33602 );
xor ( n325135 , n34708 , n34019 );
nand ( n34710 , n325133 , n325135 );
nand ( n34711 , n34703 , n34710 );
not ( n34712 , n34711 );
nand ( n34713 , n325126 , n34712 );
nand ( n34714 , n34612 , n325064 , n34681 , n34713 );
or ( n325141 , n314315 , n314380 );
not ( n34716 , n325141 );
not ( n34717 , n34693 );
or ( n325144 , n34716 , n34717 );
nand ( n34719 , n314315 , n314380 );
nand ( n34720 , n325144 , n34719 );
not ( n34721 , n34720 );
xor ( n34722 , n315709 , n314320 );
not ( n325149 , n34722 );
not ( n325150 , n325149 );
not ( n34725 , n33977 );
not ( n325152 , n324282 );
or ( n34727 , n34725 , n325152 );
not ( n34728 , n33608 );
not ( n34729 , n33863 );
or ( n325156 , n34728 , n34729 );
nand ( n34731 , n325156 , n324297 );
not ( n325158 , n34731 );
nand ( n34733 , n34727 , n325158 );
nand ( n34734 , n33623 , n324301 );
not ( n325161 , n34734 );
and ( n325162 , n34733 , n325161 );
not ( n34737 , n34733 );
and ( n325164 , n34737 , n34734 );
nor ( n325165 , n325162 , n325164 );
not ( n34740 , n325165 );
or ( n325167 , n325150 , n34740 );
or ( n34742 , n325149 , n325165 );
nand ( n34743 , n325167 , n34742 );
not ( n34744 , n34743 );
nand ( n325171 , n34721 , n34744 );
xor ( n34746 , n34704 , n34705 );
not ( n325173 , n34746 );
not ( n34748 , n325173 );
not ( n34749 , n325135 );
not ( n325176 , n34749 );
or ( n325177 , n34748 , n325176 );
not ( n34752 , n325173 );
nand ( n325179 , n34752 , n325135 );
nand ( n325180 , n325177 , n325179 );
nand ( n34755 , n325023 , n325078 );
not ( n325182 , n34664 );
nor ( n34757 , n34755 , n325182 );
not ( n34758 , n34757 );
not ( n34759 , n324905 );
not ( n325186 , n34759 );
or ( n34761 , n34758 , n325186 );
nand ( n34762 , n34761 , n325089 );
not ( n34763 , n33849 );
nor ( n325190 , n34763 , n324258 );
not ( n325191 , n325190 );
nand ( n34766 , n34762 , n325191 );
not ( n34767 , n314353 );
not ( n34768 , n312280 );
nor ( n34769 , n34767 , n34768 );
not ( n34770 , n34769 );
or ( n34771 , n34467 , n34465 );
not ( n34772 , n324896 );
not ( n34773 , n324899 );
or ( n34774 , n34772 , n34773 );
nand ( n34775 , n34774 , n324902 );
not ( n34776 , n34775 );
nand ( n34777 , n34771 , n34776 );
not ( n34778 , n34777 );
not ( n34779 , n325079 );
or ( n34780 , n34778 , n34779 );
nand ( n34781 , n34780 , n34659 );
nor ( n325208 , n325190 , n325182 );
nand ( n34783 , n34781 , n325208 );
and ( n325210 , n34759 , n34757 );
nand ( n34785 , n325190 , n325089 );
nor ( n325212 , n325210 , n34785 );
not ( n325213 , n325212 );
nand ( n34788 , n34766 , n34770 , n34783 , n325213 );
nor ( n34789 , n325208 , n34769 , n325182 );
and ( n325216 , n34789 , n34766 , n34781 );
nand ( n34791 , n34767 , n34768 );
nor ( n325218 , n34769 , n34791 );
nor ( n34793 , n325216 , n325218 );
nand ( n325220 , n34788 , n34793 );
nand ( n325221 , n325180 , n325220 );
or ( n34796 , n315709 , n314320 );
not ( n34797 , n34796 );
not ( n325224 , n325165 );
or ( n34799 , n34797 , n325224 );
nand ( n325226 , n315709 , n314320 );
nand ( n34801 , n34799 , n325226 );
not ( n34802 , n34801 );
not ( n325229 , n315714 );
not ( n325230 , n315290 );
or ( n34805 , n325229 , n325230 );
or ( n325232 , n315290 , n315714 );
nand ( n325233 , n34805 , n325232 );
not ( n34808 , n325233 );
and ( n325235 , n325057 , n34808 );
not ( n325236 , n325057 );
and ( n325237 , n325236 , n325233 );
nor ( n34812 , n325235 , n325237 );
and ( n325239 , n325046 , n34812 );
not ( n34814 , n325046 );
and ( n34815 , n325049 , n34808 );
not ( n325242 , n325049 );
and ( n325243 , n325242 , n325233 );
nor ( n34818 , n34815 , n325243 );
and ( n325245 , n34814 , n34818 );
or ( n325246 , n325239 , n325245 );
nand ( n34821 , n34802 , n325246 );
not ( n325248 , n312280 );
not ( n325249 , n34767 );
or ( n34824 , n325248 , n325249 );
nand ( n325251 , n34768 , n314353 );
nand ( n34826 , n34824 , n325251 );
not ( n325253 , n34826 );
not ( n34828 , n34781 );
not ( n34829 , n34664 );
or ( n325256 , n34828 , n34829 );
not ( n325257 , n325213 );
nand ( n34832 , n325256 , n325257 );
nand ( n325259 , n34781 , n325208 );
nand ( n325260 , n34762 , n325191 );
nand ( n34835 , n34832 , n325259 , n325260 );
not ( n325262 , n34835 );
or ( n325263 , n325253 , n325262 );
nand ( n34838 , n34832 , n325259 , n325260 );
or ( n325265 , n34838 , n34826 );
nand ( n325266 , n325263 , n325265 );
not ( n325267 , n325099 );
or ( n34842 , n312275 , n325075 );
not ( n325269 , n34842 );
or ( n34844 , n325267 , n325269 );
nand ( n34845 , n312275 , n325075 );
nand ( n325272 , n34844 , n34845 );
not ( n325273 , n325272 );
nand ( n34848 , n325266 , n325273 );
nand ( n325275 , n325171 , n325221 , n34821 , n34848 );
nor ( n325276 , n34714 , n325275 );
not ( n34851 , n325276 );
nand ( n325278 , n324922 , n324174 );
not ( n325279 , n34562 );
not ( n34854 , n325279 );
and ( n325281 , n34581 , n324954 );
not ( n34856 , n34581 );
and ( n34857 , n34856 , n321017 );
nor ( n325284 , n325281 , n34857 );
xor ( n325285 , n325284 , n34568 );
not ( n34860 , n325285 );
or ( n325287 , n34854 , n34860 );
or ( n325288 , n325279 , n325285 );
nand ( n34863 , n325287 , n325288 );
buf ( n325290 , n34863 );
xor ( n34865 , n322031 , n321617 );
xor ( n325292 , n34865 , n320974 );
buf ( n325293 , n325292 );
buf ( n325294 , n321035 );
buf ( n325295 , n321045 );
xor ( n34870 , n325294 , n325295 );
buf ( n325297 , n319572 );
and ( n325298 , n34870 , n325297 );
and ( n34873 , n325294 , n325295 );
or ( n325300 , n325298 , n34873 );
buf ( n325301 , n325300 );
buf ( n325302 , n325301 );
xor ( n325303 , n325293 , n325302 );
and ( n34878 , n321012 , n34556 );
not ( n325305 , n321012 );
and ( n34880 , n325305 , n321040 );
or ( n325307 , n34878 , n34880 );
xor ( n34882 , n325307 , n320739 );
buf ( n325309 , n34882 );
and ( n34884 , n325303 , n325309 );
and ( n34885 , n325293 , n325302 );
or ( n325312 , n34884 , n34885 );
buf ( n325313 , n325312 );
or ( n34888 , n325290 , n325313 );
nand ( n325315 , n325290 , n325313 );
nand ( n325316 , n34888 , n325315 );
xor ( n34891 , n325278 , n325316 );
buf ( n325318 , n33709 );
not ( n325319 , n325318 );
not ( n34894 , n34759 );
or ( n325321 , n325319 , n34894 );
and ( n34896 , n34777 , n325318 );
nor ( n34897 , n34896 , n324919 );
nand ( n325324 , n325321 , n34897 );
xnor ( n325325 , n34891 , n325324 );
not ( n34900 , n33671 );
not ( n325327 , n33527 );
or ( n325328 , n34900 , n325327 );
nand ( n34903 , n325328 , n34465 );
buf ( n325330 , n324133 );
nand ( n34905 , n324224 , n325330 );
nor ( n325332 , n34905 , n34467 );
and ( n325333 , n34903 , n325332 );
not ( n34908 , n325333 );
not ( n325335 , n34905 );
not ( n325336 , n325335 );
not ( n34911 , n34775 );
or ( n34912 , n325336 , n34911 );
buf ( n325339 , n33809 );
not ( n34914 , n325339 );
nand ( n325341 , n34912 , n34914 );
not ( n34916 , n325341 );
xor ( n325343 , n325293 , n325302 );
xor ( n325344 , n325343 , n325309 );
buf ( n325345 , n325344 );
buf ( n325346 , n320734 );
buf ( n325347 , n318009 );
xor ( n34922 , n325346 , n325347 );
xor ( n325349 , n325294 , n325295 );
xor ( n325350 , n325349 , n325297 );
buf ( n325351 , n325350 );
buf ( n325352 , n325351 );
and ( n34927 , n34922 , n325352 );
and ( n325354 , n325346 , n325347 );
or ( n34929 , n34927 , n325354 );
buf ( n325356 , n34929 );
or ( n325357 , n325345 , n325356 );
nand ( n34932 , n324242 , n33691 );
not ( n34933 , n34932 );
and ( n325360 , n325357 , n34933 );
nand ( n34935 , n34908 , n34916 , n325360 );
and ( n325362 , n325357 , n34932 );
nand ( n325363 , n325362 , n325341 );
nand ( n34938 , n325333 , n325362 );
nand ( n34939 , n325345 , n325356 );
and ( n34940 , n34935 , n325363 , n34938 , n34939 );
nand ( n34941 , n325325 , n34940 );
nand ( n34942 , n34908 , n34916 );
not ( n325369 , n325345 );
not ( n34944 , n325356 );
and ( n325371 , n325369 , n34944 );
and ( n325372 , n325345 , n325356 );
nor ( n34947 , n325371 , n325372 );
and ( n34948 , n34947 , n34932 );
not ( n34949 , n34947 );
and ( n34950 , n34949 , n34933 );
nor ( n325377 , n34948 , n34950 );
not ( n325378 , n325377 );
and ( n34953 , n34942 , n325378 );
not ( n34954 , n34942 );
and ( n34955 , n34954 , n325377 );
nor ( n34956 , n34953 , n34955 );
not ( n34957 , n34956 );
buf ( n325384 , n319567 );
buf ( n325385 , n317158 );
xor ( n34960 , n325384 , n325385 );
buf ( n325387 , n318004 );
and ( n325388 , n34960 , n325387 );
and ( n34963 , n325384 , n325385 );
or ( n34964 , n325388 , n34963 );
buf ( n325391 , n34964 );
xor ( n325392 , n325346 , n325347 );
xor ( n325393 , n325392 , n325352 );
buf ( n325394 , n325393 );
or ( n34969 , n325391 , n325394 );
not ( n34970 , n34969 );
nand ( n34971 , n324232 , n33807 );
nand ( n34972 , n34971 , n324107 );
nor ( n325399 , n34970 , n34972 );
not ( n325400 , n325399 );
not ( n325401 , n325330 );
not ( n34976 , n324906 );
or ( n325403 , n325401 , n34976 );
not ( n34978 , n33800 );
nand ( n34979 , n325403 , n34978 );
not ( n325406 , n34979 );
not ( n325407 , n325406 );
or ( n34982 , n325400 , n325407 );
not ( n325409 , n34969 );
not ( n34984 , n34972 );
nor ( n325411 , n325409 , n34984 );
and ( n325412 , n325411 , n34979 );
and ( n34987 , n325391 , n325394 );
nor ( n325414 , n325412 , n34987 );
nand ( n34989 , n34982 , n325414 );
not ( n34990 , n34989 );
nand ( n34991 , n34957 , n34990 );
not ( n34992 , n325278 );
buf ( n34993 , n34992 );
not ( n325420 , n325324 );
nand ( n325421 , n34993 , n325420 );
not ( n34996 , n325421 );
not ( n325423 , n325420 );
not ( n34998 , n34993 );
nand ( n34999 , n325423 , n34998 );
not ( n35000 , n34999 );
or ( n35001 , n34996 , n35000 );
or ( n35002 , n325290 , n325313 );
nand ( n325429 , n35001 , n35002 );
xnor ( n325430 , n34594 , n324979 );
xor ( n35005 , n325033 , n325430 );
xnor ( n325432 , n35005 , n34602 );
nand ( n35007 , n325429 , n325432 , n325315 );
not ( n35008 , n325391 );
not ( n35009 , n325394 );
and ( n35010 , n35008 , n35009 );
and ( n325437 , n325391 , n325394 );
nor ( n325438 , n35010 , n325437 );
not ( n35013 , n325438 );
and ( n325440 , n34972 , n35013 );
not ( n35015 , n34972 );
and ( n325442 , n35015 , n325438 );
nor ( n35017 , n325440 , n325442 );
not ( n35018 , n35017 );
not ( n325445 , n325406 );
or ( n35020 , n35018 , n325445 );
and ( n35021 , n34984 , n35013 );
not ( n35022 , n34984 );
and ( n35023 , n35022 , n325438 );
nor ( n35024 , n35021 , n35023 );
nand ( n325451 , n35024 , n34979 );
nand ( n35026 , n35020 , n325451 );
not ( n35027 , n35026 );
xor ( n35028 , n325384 , n325385 );
xor ( n35029 , n35028 , n325387 );
buf ( n325456 , n35029 );
xor ( n325457 , n320668 , n318109 );
and ( n35032 , n325457 , n317153 );
and ( n35033 , n320668 , n318109 );
or ( n325460 , n35032 , n35033 );
or ( n35035 , n325456 , n325460 );
not ( n35036 , n35035 );
and ( n35037 , n325330 , n34978 );
xor ( n35038 , n35037 , n324906 );
not ( n35039 , n35038 );
or ( n325466 , n35036 , n35039 );
nand ( n325467 , n325456 , n325460 );
nand ( n35042 , n325466 , n325467 );
buf ( n325469 , n35042 );
not ( n325470 , n325469 );
buf ( n325471 , n325470 );
nand ( n35046 , n35027 , n325471 );
nand ( n325473 , n34941 , n34991 , n35007 , n35046 );
not ( n35048 , n325473 );
not ( n35049 , n318129 );
not ( n325476 , n319514 );
nand ( n325477 , n35049 , n325476 );
not ( n35052 , n325477 );
nand ( n325479 , n35052 , n318104 );
not ( n325480 , n325476 );
and ( n35055 , n318129 , n325480 );
nand ( n35056 , n35055 , n318104 );
nor ( n35057 , n318129 , n325476 );
not ( n325484 , n318104 );
nand ( n325485 , n35057 , n325484 );
not ( n325486 , n318129 );
nor ( n35061 , n325486 , n325480 );
nand ( n325488 , n35061 , n325484 );
nand ( n35063 , n325479 , n35056 , n325485 , n325488 );
not ( n325490 , n35063 );
xor ( n325491 , n319934 , n318264 );
and ( n35066 , n325491 , n318124 );
and ( n35067 , n319934 , n318264 );
or ( n325494 , n35066 , n35067 );
not ( n325495 , n325494 );
and ( n35070 , n325490 , n325495 );
and ( n35071 , n35063 , n325494 );
nor ( n325498 , n35070 , n35071 );
nand ( n325499 , n324070 , n34472 );
xnor ( n325500 , n325498 , n325499 );
buf ( n35075 , n324201 );
and ( n35076 , n35075 , n33664 );
not ( n325503 , n35076 );
not ( n35078 , n34903 );
or ( n35079 , n325503 , n35078 );
nand ( n325506 , n33774 , n35075 );
nand ( n325507 , n35079 , n325506 );
and ( n35082 , n325500 , n325507 );
not ( n325509 , n325500 );
not ( n325510 , n325507 );
and ( n35085 , n325509 , n325510 );
nor ( n35086 , n35082 , n35085 );
not ( n35087 , n33664 );
not ( n325514 , n34903 );
or ( n35089 , n35087 , n325514 );
buf ( n325516 , n324199 );
nand ( n325517 , n35089 , n325516 );
not ( n325518 , n325517 );
not ( n325519 , n324189 );
not ( n35094 , n324192 );
or ( n325521 , n325519 , n35094 );
nand ( n325522 , n325521 , n35075 );
xor ( n35097 , n319934 , n318264 );
xor ( n325524 , n35097 , n318124 );
not ( n325525 , n318269 );
not ( n35100 , n319929 );
nand ( n325527 , n325525 , n35100 );
not ( n325528 , n325527 );
not ( n35103 , n318259 );
or ( n35104 , n325528 , n35103 );
nand ( n35105 , n319929 , n318269 );
nand ( n325532 , n35104 , n35105 );
nor ( n35107 , n325524 , n325532 );
nor ( n35108 , n325522 , n35107 );
and ( n35109 , n325518 , n35108 );
and ( n35110 , n325524 , n325532 );
nor ( n35111 , n35109 , n35110 );
not ( n325538 , n35107 );
nand ( n325539 , n325538 , n325522 , n325517 );
nand ( n35114 , n35111 , n325539 );
nand ( n325541 , n35086 , n35114 );
not ( n35116 , n325541 );
xor ( n35117 , n325524 , n325517 );
xor ( n325544 , n325532 , n325522 );
xnor ( n325545 , n35117 , n325544 );
buf ( n325546 , n325545 );
buf ( n35121 , n34903 );
nand ( n325548 , n324199 , n33664 );
xor ( n325549 , n35121 , n325548 );
not ( n325550 , n319929 );
not ( n35125 , n325525 );
or ( n35126 , n325550 , n35125 );
nand ( n35127 , n35100 , n318269 );
nand ( n325554 , n35126 , n35127 );
and ( n35129 , n325554 , n318259 );
not ( n35130 , n325554 );
not ( n325557 , n318259 );
and ( n325558 , n35130 , n325557 );
nor ( n35133 , n35129 , n325558 );
nor ( n35134 , n35133 , n313446 );
or ( n35135 , n325549 , n35134 );
nand ( n35136 , n313446 , n35133 );
nand ( n35137 , n35135 , n35136 );
buf ( n325564 , n35137 );
nand ( n325565 , n325546 , n325564 );
buf ( n325566 , n325565 );
not ( n325567 , n325566 );
or ( n325568 , n35116 , n325567 );
or ( n35143 , n35063 , n325494 );
not ( n35144 , n35143 );
not ( n35145 , n325499 );
not ( n35146 , n325507 );
or ( n325573 , n35145 , n35146 );
or ( n325574 , n325507 , n325499 );
nand ( n35149 , n325573 , n325574 );
not ( n35150 , n35149 );
or ( n35151 , n35144 , n35150 );
nand ( n325578 , n35063 , n325494 );
nand ( n325579 , n35151 , n325578 );
not ( n35154 , n325579 );
nand ( n325581 , n324902 , n324896 );
not ( n35156 , n33794 );
not ( n325583 , n35156 );
not ( n325584 , n34903 );
or ( n35159 , n325583 , n325584 );
buf ( n35160 , n324899 );
not ( n35161 , n35160 );
nand ( n35162 , n35159 , n35161 );
xor ( n325589 , n325581 , n35162 );
xor ( n35164 , n320668 , n318109 );
xor ( n325591 , n35164 , n317153 );
not ( n325592 , n318104 );
not ( n325593 , n325477 );
or ( n35168 , n325592 , n325593 );
nand ( n325595 , n318129 , n325480 );
nand ( n325596 , n35168 , n325595 );
not ( n35171 , n325596 );
or ( n325598 , n325591 , n35171 );
not ( n325599 , n325591 );
or ( n35174 , n325599 , n325596 );
nand ( n35175 , n325598 , n35174 );
xor ( n35176 , n325589 , n35175 );
nand ( n35177 , n35154 , n35176 );
nand ( n325604 , n325568 , n35177 );
not ( n325605 , n35086 );
not ( n35180 , n325605 );
not ( n325607 , n35114 );
not ( n35182 , n325607 );
or ( n325609 , n35180 , n35182 );
xor ( n325610 , n325456 , n325460 );
and ( n35185 , n35038 , n325610 );
not ( n325612 , n35038 );
not ( n35187 , n325610 );
and ( n325614 , n325612 , n35187 );
or ( n35189 , n35185 , n325614 );
not ( n325616 , n35162 );
not ( n325617 , n325581 );
nor ( n35192 , n325599 , n35171 );
nor ( n325619 , n325617 , n35192 );
nand ( n35194 , n325616 , n325619 );
nor ( n35195 , n325581 , n35192 );
nand ( n35196 , n35195 , n35162 );
nand ( n35197 , n325599 , n35171 );
nand ( n35198 , n35194 , n35196 , n35197 );
nand ( n35199 , n35189 , n35198 );
nand ( n325626 , n325609 , n35199 );
nor ( n325627 , n325604 , n325626 );
nand ( n35202 , n35048 , n325627 );
not ( n35203 , n34990 );
not ( n35204 , n34956 );
not ( n35205 , n35204 );
or ( n325632 , n35203 , n35205 );
nand ( n325633 , n35027 , n325471 );
nand ( n35208 , n325632 , n325633 );
not ( n35209 , n35208 );
not ( n35210 , n35199 );
nor ( n325637 , n35154 , n35176 );
not ( n325638 , n325637 );
or ( n325639 , n35210 , n325638 );
or ( n35214 , n35189 , n35198 );
nand ( n325641 , n325639 , n35214 );
not ( n35216 , n325432 );
not ( n35217 , n325315 );
or ( n325644 , n35217 , n35002 );
not ( n325645 , n35217 );
nand ( n35220 , n325645 , n34993 );
or ( n35221 , n35220 , n325420 );
nor ( n325648 , n34993 , n35217 );
nand ( n325649 , n325420 , n325648 );
nand ( n325650 , n325644 , n35221 , n325649 );
not ( n35225 , n325650 );
or ( n35226 , n35216 , n35225 );
nand ( n325653 , n35226 , n34941 );
not ( n35228 , n325653 );
nand ( n35229 , n35209 , n325641 , n35228 );
not ( n325656 , n325432 );
not ( n325657 , n325650 );
nand ( n35232 , n325656 , n325657 );
nand ( n35233 , n35026 , n35042 );
not ( n35234 , n35233 );
nand ( n325661 , n34990 , n35204 );
nand ( n325662 , n35234 , n34941 , n325661 );
not ( n35237 , n34940 );
xnor ( n325664 , n325290 , n325313 );
and ( n325665 , n325324 , n34992 );
not ( n35240 , n325324 );
and ( n325667 , n35240 , n325278 );
nor ( n35242 , n325665 , n325667 );
xnor ( n35243 , n325664 , n35242 );
nand ( n35244 , n35237 , n35243 );
nand ( n35245 , n35232 , n325662 , n35244 );
buf ( n35246 , n35007 );
nand ( n325673 , n35245 , n35246 );
and ( n35248 , n34989 , n34956 );
nand ( n35249 , n35228 , n35248 );
nand ( n35250 , n35202 , n35229 , n325673 , n35249 );
not ( n35251 , n35250 );
or ( n35252 , n34851 , n35251 );
nand ( n35253 , n34644 , n325105 );
nand ( n35254 , n324976 , n325036 );
nand ( n35255 , n35253 , n35254 );
nand ( n325682 , n35255 , n34681 , n34848 , n325221 );
not ( n35257 , n325272 );
nor ( n35258 , n325266 , n35257 );
and ( n325685 , n325221 , n35258 );
nor ( n325686 , n325180 , n325220 );
nor ( n35261 , n325685 , n325686 );
nand ( n35262 , n325682 , n35261 );
not ( n325689 , n325062 );
not ( n325690 , n324335 );
and ( n35265 , n325689 , n325690 );
not ( n35266 , n34801 );
and ( n35267 , n325246 , n35266 );
nor ( n35268 , n35265 , n35267 );
not ( n35269 , n35268 );
nand ( n325696 , n325126 , n34712 );
nand ( n325697 , n325696 , n325171 );
nor ( n35272 , n35269 , n325697 );
and ( n325699 , n35262 , n35272 );
not ( n35274 , n35268 );
not ( n35275 , n34699 );
nor ( n35276 , n35275 , n34712 );
not ( n325703 , n35276 );
nand ( n35278 , n34744 , n34721 );
not ( n35279 , n35278 );
or ( n35280 , n325703 , n35279 );
nand ( n35281 , n34720 , n34743 );
nand ( n325708 , n35280 , n35281 );
not ( n35283 , n325708 );
or ( n35284 , n35274 , n35283 );
not ( n35285 , n324335 );
not ( n35286 , n35285 );
not ( n35287 , n34637 );
and ( n35288 , n35286 , n35287 );
nand ( n325715 , n34637 , n35285 );
nor ( n35290 , n35266 , n325246 );
and ( n35291 , n325715 , n35290 );
nor ( n325718 , n35288 , n35291 );
nand ( n325719 , n35284 , n325718 );
nor ( n35294 , n325699 , n325719 );
nand ( n325721 , n35252 , n35294 );
buf ( n325722 , n325721 );
not ( n35297 , n325722 );
or ( n325724 , n324880 , n35297 );
xor ( n325725 , n322579 , n322358 );
and ( n35300 , n325725 , n322286 );
and ( n325727 , n322579 , n322358 );
or ( n325728 , n35300 , n325727 );
buf ( n325729 , n325728 );
xor ( n325730 , n322459 , n322291 );
xor ( n325731 , n325730 , n322120 );
buf ( n325732 , n325731 );
xor ( n35307 , n325729 , n325732 );
not ( n325734 , n323724 );
not ( n35309 , n323505 );
or ( n35310 , n325734 , n35309 );
not ( n325737 , n33301 );
nand ( n325738 , n323728 , n33181 );
nor ( n35313 , n325737 , n325738 );
nand ( n325740 , n35310 , n35313 );
not ( n325741 , n323738 );
not ( n35316 , n325741 );
nand ( n325743 , n33287 , n35316 );
xnor ( n325744 , n325740 , n325743 );
buf ( n325745 , n325744 );
and ( n325746 , n35307 , n325745 );
and ( n35321 , n325729 , n325732 );
or ( n325748 , n325746 , n35321 );
buf ( n325749 , n325748 );
not ( n35324 , n33287 );
not ( n325751 , n325740 );
or ( n325752 , n35324 , n325751 );
nand ( n35327 , n325752 , n35316 );
buf ( n35328 , n33310 );
nand ( n325755 , n35328 , n33318 );
not ( n325756 , n325755 );
and ( n35331 , n35327 , n325756 );
not ( n35332 , n35327 );
and ( n35333 , n35332 , n325755 );
nor ( n325760 , n35331 , n35333 );
not ( n325761 , n325760 );
xor ( n35336 , n322459 , n322291 );
and ( n35337 , n35336 , n322120 );
and ( n325764 , n322459 , n322291 );
or ( n325765 , n35337 , n325764 );
xor ( n35340 , n320953 , n325765 );
not ( n35341 , n35340 );
and ( n35342 , n325761 , n35341 );
not ( n35343 , n325761 );
and ( n35344 , n35343 , n35340 );
nor ( n325771 , n35342 , n35344 );
or ( n325772 , n325749 , n325771 );
or ( n35347 , n320501 , n320325 );
not ( n35348 , n35347 );
buf ( n35349 , n33258 );
buf ( n35350 , n35349 );
not ( n325777 , n35350 );
not ( n325778 , n33289 );
not ( n35353 , n325740 );
or ( n35354 , n325778 , n35353 );
not ( n35355 , n33310 );
nor ( n35356 , n35316 , n33317 );
nor ( n35357 , n35355 , n35356 );
nand ( n325784 , n35354 , n35357 );
not ( n325785 , n325784 );
or ( n35360 , n325777 , n325785 );
not ( n35361 , n323757 );
nand ( n35362 , n35360 , n35361 );
not ( n325789 , n33335 );
nand ( n325790 , n325789 , n323746 );
not ( n35365 , n325790 );
and ( n35366 , n35362 , n35365 );
not ( n35367 , n35362 );
and ( n325794 , n35367 , n325790 );
nor ( n325795 , n35366 , n325794 );
not ( n35370 , n325795 );
or ( n35371 , n35348 , n35370 );
nand ( n325798 , n320501 , n320325 );
nand ( n325799 , n35371 , n325798 );
not ( n35374 , n325799 );
xor ( n325801 , n320127 , n320330 );
buf ( n325802 , n323745 );
buf ( n35377 , n33299 );
buf ( n325804 , n323762 );
nand ( n35379 , n325802 , n35377 , n325804 );
buf ( n325806 , n35379 );
nand ( n325807 , n33388 , n33491 );
not ( n325808 , n325807 );
and ( n325809 , n325806 , n325808 );
not ( n35384 , n325806 );
and ( n325811 , n35384 , n325807 );
nor ( n325812 , n325809 , n325811 );
not ( n35387 , n325812 );
and ( n325814 , n325801 , n35387 );
not ( n325815 , n325801 );
and ( n35390 , n325815 , n325812 );
nor ( n35391 , n325814 , n35390 );
nand ( n325818 , n35374 , n35391 );
xnor ( n35393 , n320501 , n320325 );
not ( n35394 , n325795 );
and ( n35395 , n35393 , n35394 );
not ( n325822 , n35393 );
and ( n325823 , n325822 , n325795 );
nor ( n35398 , n35395 , n325823 );
not ( n35399 , n35398 );
buf ( n325826 , n320958 );
buf ( n325827 , n320496 );
xor ( n325828 , n325826 , n325827 );
not ( n35403 , n323757 );
nand ( n325830 , n35403 , n35350 );
not ( n325831 , n325830 );
and ( n35406 , n325784 , n325831 );
not ( n35407 , n325784 );
and ( n35408 , n35407 , n325830 );
nor ( n325835 , n35406 , n35408 );
buf ( n325836 , n325835 );
and ( n35411 , n325828 , n325836 );
and ( n325838 , n325826 , n325827 );
or ( n325839 , n35411 , n325838 );
buf ( n325840 , n325839 );
not ( n35415 , n325840 );
nand ( n35416 , n35399 , n35415 );
xor ( n35417 , n325826 , n325827 );
xor ( n325844 , n35417 , n325836 );
buf ( n325845 , n325844 );
buf ( n325846 , n325845 );
or ( n325847 , n320953 , n325765 );
not ( n325848 , n325847 );
not ( n325849 , n325760 );
or ( n35424 , n325848 , n325849 );
nand ( n325851 , n320953 , n325765 );
nand ( n325852 , n35424 , n325851 );
buf ( n325853 , n325852 );
nor ( n325854 , n325846 , n325853 );
buf ( n325855 , n325854 );
not ( n35430 , n325855 );
nand ( n35431 , n325772 , n325818 , n35416 , n35430 );
not ( n35432 , n35431 );
buf ( n325859 , n323418 );
buf ( n35434 , n323391 );
or ( n35435 , n325859 , n35434 );
buf ( n325862 , n35435 );
buf ( n325863 , n325862 );
buf ( n325864 , n323423 );
buf ( n325865 , n323460 );
or ( n35440 , n325864 , n325865 );
buf ( n325867 , n35440 );
buf ( n325868 , n325867 );
and ( n325869 , n325863 , n325868 );
buf ( n325870 , n325869 );
buf ( n325871 , n323316 );
buf ( n325872 , n322952 );
xor ( n325873 , n323240 , n323248 );
xor ( n35448 , n325873 , n323257 );
buf ( n35449 , n35448 );
buf ( n325876 , n35449 );
xor ( n35451 , n325872 , n325876 );
and ( n35452 , n323211 , n323221 );
not ( n35453 , n323225 );
nor ( n325880 , n35452 , n35453 );
nand ( n35455 , n32864 , n323285 );
xor ( n35456 , n325880 , n35455 );
buf ( n325883 , n35456 );
and ( n325884 , n35451 , n325883 );
and ( n35459 , n325872 , n325876 );
or ( n35460 , n325884 , n35459 );
buf ( n325887 , n35460 );
buf ( n325888 , n325887 );
nor ( n35463 , n325871 , n325888 );
buf ( n325890 , n35463 );
buf ( n325891 , n325890 );
xor ( n35466 , n325872 , n325876 );
xor ( n35467 , n35466 , n325883 );
buf ( n325894 , n35467 );
buf ( n325895 , n325894 );
buf ( n325896 , n32810 );
nand ( n35471 , n325895 , n325896 );
buf ( n325898 , n35471 );
buf ( n325899 , n325898 );
or ( n325900 , n325891 , n325899 );
buf ( n325901 , n323316 );
buf ( n325902 , n325887 );
nand ( n35477 , n325901 , n325902 );
buf ( n325904 , n35477 );
buf ( n325905 , n325904 );
nand ( n35480 , n325900 , n325905 );
buf ( n325907 , n35480 );
buf ( n325908 , n325890 );
not ( n35483 , n325908 );
buf ( n325910 , n35483 );
buf ( n325911 , n325910 );
buf ( n325912 , n324348 );
buf ( n325913 , n323192 );
nand ( n35488 , n325912 , n325913 );
buf ( n325915 , n35488 );
not ( n325916 , n325915 );
buf ( n325917 , n323192 );
buf ( n325918 , n324348 );
or ( n35493 , n325917 , n325918 );
buf ( n325920 , n35493 );
buf ( n325921 , n325920 );
buf ( n325922 , n323020 );
buf ( n325923 , n323039 );
nand ( n35498 , n32740 , n323177 );
not ( n325925 , n323150 );
and ( n35500 , n35498 , n325925 );
not ( n35501 , n35498 );
and ( n35502 , n35501 , n323150 );
nor ( n325929 , n35500 , n35502 );
buf ( n325930 , n325929 );
and ( n35505 , n325923 , n325930 );
buf ( n325932 , n35505 );
buf ( n325933 , n325932 );
xor ( n35508 , n325922 , n325933 );
buf ( n325935 , n324346 );
and ( n35510 , n35508 , n325935 );
or ( n35511 , n35510 , C0 );
buf ( n325938 , n35511 );
buf ( n325939 , n325938 );
nand ( n35514 , n325921 , n325939 );
buf ( n325941 , n35514 );
not ( n35516 , n325941 );
or ( n35517 , n325916 , n35516 );
buf ( n325944 , n323231 );
buf ( n325945 , n323197 );
nor ( n35520 , n325944 , n325945 );
buf ( n325947 , n35520 );
not ( n35522 , n325947 );
nand ( n35523 , n35517 , n35522 );
buf ( n325950 , n323197 );
buf ( n325951 , n323231 );
nand ( n35526 , n325950 , n325951 );
buf ( n325953 , n35526 );
nand ( n35528 , n35523 , n325953 );
buf ( n35529 , n35528 );
buf ( n325956 , n325894 );
buf ( n325957 , n32810 );
or ( n35532 , n325956 , n325957 );
buf ( n325959 , n35532 );
buf ( n325960 , n325959 );
and ( n35535 , n325911 , n35529 , n325960 );
buf ( n325962 , n35535 );
or ( n35537 , n325907 , n325962 );
buf ( n325964 , n323386 );
buf ( n325965 , n323354 );
nor ( n35540 , n325964 , n325965 );
buf ( n325967 , n35540 );
buf ( n325968 , n325967 );
buf ( n325969 , n323349 );
buf ( n325970 , n323321 );
nor ( n35545 , n325969 , n325970 );
buf ( n325972 , n35545 );
buf ( n325973 , n325972 );
nor ( n35548 , n325968 , n325973 );
buf ( n325975 , n35548 );
nand ( n35550 , n35537 , n325975 );
buf ( n325977 , n323349 );
buf ( n325978 , n323321 );
nand ( n35553 , n325977 , n325978 );
buf ( n325980 , n35553 );
buf ( n325981 , n325980 );
not ( n35556 , n325981 );
buf ( n325983 , n325967 );
not ( n35558 , n325983 );
and ( n35559 , n35556 , n35558 );
buf ( n325986 , n323386 );
buf ( n325987 , n323354 );
and ( n35562 , n325986 , n325987 );
buf ( n325989 , n35562 );
buf ( n325990 , n325989 );
nor ( n35565 , n35559 , n325990 );
buf ( n325992 , n35565 );
nand ( n35567 , n35550 , n325992 );
nand ( n35568 , n325870 , n35567 );
buf ( n325995 , n323418 );
buf ( n325996 , n323391 );
and ( n35571 , n325995 , n325996 );
buf ( n325998 , n35571 );
not ( n35573 , n325998 );
not ( n35574 , n325867 );
or ( n35575 , n35573 , n35574 );
buf ( n326002 , n323423 );
buf ( n326003 , n323460 );
nand ( n35578 , n326002 , n326003 );
buf ( n326005 , n35578 );
nand ( n35580 , n35575 , n326005 );
not ( n35581 , n35580 );
and ( n35582 , n35568 , n35581 );
or ( n35583 , n322112 , n322456 );
not ( n35584 , n35583 );
and ( n35585 , n33073 , n33078 );
not ( n35586 , n35585 );
and ( n35587 , n33029 , n33018 );
not ( n35588 , n323440 );
nor ( n326015 , n35587 , n35588 );
not ( n35590 , n326015 );
or ( n35591 , n35586 , n35590 );
or ( n35592 , n326015 , n35585 );
nand ( n35593 , n35591 , n35592 );
not ( n35594 , n35593 );
or ( n35595 , n35584 , n35594 );
nand ( n35596 , n322112 , n322456 );
nand ( n35597 , n35595 , n35596 );
buf ( n35598 , n35597 );
not ( n35599 , n35598 );
buf ( n326026 , n35599 );
buf ( n326027 , n326026 );
buf ( n326028 , n323511 );
not ( n326029 , n326028 );
buf ( n326030 , n326029 );
buf ( n326031 , n326030 );
nand ( n35606 , n326027 , n326031 );
buf ( n326033 , n35606 );
xor ( n35608 , n322112 , n322456 );
not ( n35609 , n35608 );
not ( n326036 , n35593 );
or ( n326037 , n35609 , n326036 );
or ( n35612 , n35593 , n35608 );
nand ( n35613 , n326037 , n35612 );
buf ( n326040 , n35613 );
buf ( n326041 , n323465 );
not ( n35616 , n326041 );
buf ( n326043 , n35616 );
buf ( n326044 , n326043 );
nand ( n35619 , n326040 , n326044 );
buf ( n326046 , n35619 );
nand ( n326047 , n326033 , n326046 );
nor ( n35622 , n35582 , n326047 );
buf ( n326049 , n35613 );
buf ( n326050 , n326043 );
nor ( n35625 , n326049 , n326050 );
buf ( n326052 , n35625 );
buf ( n326053 , n326052 );
not ( n326054 , n326053 );
buf ( n326055 , n326033 );
not ( n35630 , n326055 );
or ( n326057 , n326054 , n35630 );
buf ( n35632 , n323511 );
buf ( n326059 , n35597 );
nand ( n35634 , n35632 , n326059 );
buf ( n326061 , n35634 );
buf ( n326062 , n326061 );
nand ( n326063 , n326057 , n326062 );
buf ( n326064 , n326063 );
or ( n35639 , n35622 , n326064 );
xor ( n35640 , n325729 , n325732 );
xor ( n35641 , n35640 , n325745 );
buf ( n35642 , n35641 );
buf ( n326069 , n35642 );
not ( n35644 , n326069 );
buf ( n326071 , n35644 );
buf ( n326072 , n326071 );
buf ( n326073 , n33199 );
not ( n35648 , n326073 );
buf ( n326075 , n35648 );
buf ( n326076 , n326075 );
nand ( n35651 , n326072 , n326076 );
buf ( n326078 , n35651 );
buf ( n326079 , n326078 );
buf ( n326080 , n323620 );
not ( n35655 , n326080 );
buf ( n326082 , n35655 );
buf ( n326083 , n326082 );
buf ( n326084 , n323586 );
not ( n35659 , n326084 );
buf ( n326086 , n35659 );
buf ( n326087 , n326086 );
nand ( n326088 , n326083 , n326087 );
buf ( n326089 , n326088 );
buf ( n326090 , n326089 );
nand ( n35665 , n326079 , n326090 );
buf ( n326092 , n35665 );
not ( n326093 , n323543 );
buf ( n326094 , n326093 );
not ( n35669 , n323581 );
buf ( n326096 , n35669 );
nand ( n35671 , n326094 , n326096 );
buf ( n326098 , n35671 );
buf ( n326099 , n326098 );
buf ( n326100 , n323538 );
not ( n35675 , n326100 );
buf ( n326102 , n35675 );
buf ( n326103 , n326102 );
buf ( n326104 , n323516 );
not ( n35679 , n326104 );
buf ( n326106 , n35679 );
buf ( n326107 , n326106 );
nand ( n35682 , n326103 , n326107 );
buf ( n326109 , n35682 );
buf ( n326110 , n326109 );
nand ( n35685 , n326099 , n326110 );
buf ( n326112 , n35685 );
nor ( n35687 , n326092 , n326112 );
nand ( n35688 , n35639 , n35687 );
buf ( n326115 , n326092 );
not ( n35690 , n326115 );
buf ( n326117 , n35690 );
buf ( n326118 , n326102 );
buf ( n326119 , n326106 );
nor ( n35694 , n326118 , n326119 );
buf ( n326121 , n35694 );
not ( n35696 , n326121 );
not ( n35697 , n326098 );
or ( n35698 , n35696 , n35697 );
nand ( n35699 , n323581 , n323543 );
nand ( n35700 , n35698 , n35699 );
and ( n35701 , n326117 , n35700 );
buf ( n326128 , n326082 );
buf ( n326129 , n326086 );
nor ( n35704 , n326128 , n326129 );
buf ( n326131 , n35704 );
buf ( n326132 , n326131 );
not ( n35707 , n326132 );
buf ( n326134 , n326078 );
not ( n35709 , n326134 );
or ( n35710 , n35707 , n35709 );
buf ( n326137 , n326075 );
buf ( n326138 , n326071 );
or ( n35713 , n326137 , n326138 );
buf ( n326140 , n35713 );
buf ( n326141 , n326140 );
nand ( n35716 , n35710 , n326141 );
buf ( n326143 , n35716 );
nor ( n35718 , n35701 , n326143 );
nand ( n35719 , n35688 , n35718 );
xor ( n35720 , n319205 , n319511 );
buf ( n35721 , n33470 );
buf ( n35722 , n323906 );
nand ( n35723 , n35721 , n35722 );
xor ( n35724 , n35720 , n35723 );
not ( n35725 , n33411 );
not ( n35726 , n35379 );
or ( n35727 , n35725 , n35726 );
buf ( n35728 , n323835 );
not ( n326155 , n33491 );
and ( n326156 , n35728 , n326155 );
nand ( n35731 , n323833 , n33488 );
not ( n35732 , n35731 );
nor ( n35733 , n326156 , n35732 );
nand ( n35734 , n35727 , n35733 );
xnor ( n326161 , n35724 , n35734 );
buf ( n326162 , n326161 );
not ( n35737 , n326162 );
not ( n35738 , n319506 );
not ( n35739 , n320132 );
nand ( n326166 , n35738 , n35739 );
not ( n326167 , n5982 );
nand ( n35742 , n326167 , n33387 );
not ( n326169 , n35742 );
nand ( n35744 , n35377 , n325802 , n325804 );
not ( n35745 , n35744 );
or ( n35746 , n326169 , n35745 );
nand ( n35747 , n35746 , n33491 );
nand ( n35748 , n35728 , n35731 );
not ( n326175 , n35748 );
and ( n35750 , n35747 , n326175 );
not ( n35751 , n35747 );
and ( n35752 , n35751 , n35748 );
nor ( n35753 , n35750 , n35752 );
and ( n326180 , n326166 , n35753 );
and ( n326181 , n319506 , n320132 );
nor ( n35756 , n326180 , n326181 );
buf ( n326183 , n35756 );
nand ( n35758 , n35737 , n326183 );
buf ( n326185 , n35758 );
buf ( n326186 , n326185 );
or ( n326187 , n320127 , n320330 );
not ( n35762 , n326187 );
not ( n35763 , n325812 );
or ( n35764 , n35762 , n35763 );
nand ( n326191 , n320127 , n320330 );
nand ( n326192 , n35764 , n326191 );
or ( n35767 , n319506 , n35739 );
or ( n35768 , n35738 , n320132 );
nand ( n35769 , n35767 , n35768 );
xor ( n326196 , n35769 , n35748 );
xnor ( n35771 , n326196 , n35747 );
or ( n35772 , n326192 , n35771 );
buf ( n326199 , n35772 );
and ( n35774 , n326186 , n326199 );
buf ( n326201 , n35774 );
xnor ( n35776 , n318930 , n318983 );
not ( n35777 , n35776 );
not ( n326204 , n323926 );
nand ( n35779 , n33343 , n323767 );
nand ( n35780 , n326204 , n35779 );
not ( n35781 , n35780 );
or ( n35782 , n35777 , n35781 );
or ( n326209 , n35780 , n35776 );
nand ( n35784 , n35782 , n326209 );
not ( n35785 , n35784 );
not ( n35786 , n33380 );
nor ( n35787 , n35786 , n323836 );
not ( n35788 , n35787 );
not ( n35789 , n35744 );
or ( n35790 , n35788 , n35789 );
not ( n35791 , n323920 );
nand ( n326218 , n35790 , n35791 );
buf ( n35793 , n326218 );
not ( n35794 , n35793 );
or ( n35795 , n35785 , n35794 );
or ( n326222 , n35793 , n35784 );
nand ( n326223 , n35795 , n326222 );
not ( n35798 , n35722 );
not ( n326225 , n35734 );
or ( n326226 , n35798 , n326225 );
nand ( n326227 , n326226 , n35721 );
not ( n35802 , n323899 );
nand ( n326229 , n35802 , n33464 );
nor ( n35804 , n318978 , n319210 );
or ( n35805 , n326227 , n326229 , n35804 );
not ( n326232 , n326229 );
nor ( n326233 , n326232 , n35804 );
and ( n35808 , n326227 , n326233 );
and ( n326235 , n319210 , n318978 );
nor ( n326236 , n35808 , n326235 );
nand ( n326237 , n35805 , n326236 );
nor ( n35812 , n326223 , n326237 );
buf ( n326239 , n35812 );
not ( n326240 , n319205 );
not ( n35815 , n319511 );
or ( n326242 , n326240 , n35815 );
xor ( n326243 , n35734 , n35723 );
nor ( n35818 , n319205 , n319511 );
or ( n326245 , n326243 , n35818 );
nand ( n326246 , n326242 , n326245 );
xor ( n35821 , n319210 , n318978 );
xor ( n326248 , n326229 , n35821 );
xnor ( n326249 , n326248 , n326227 );
nor ( n35824 , n326246 , n326249 );
buf ( n326251 , n35824 );
nor ( n35826 , n326239 , n326251 );
buf ( n326253 , n35826 );
nand ( n326254 , n326201 , n326253 );
not ( n326255 , n326254 );
nand ( n326256 , n35432 , n35719 , n326255 );
nand ( n35831 , n35416 , n325818 );
buf ( n326258 , n35831 );
not ( n326259 , n326258 );
buf ( n326260 , n325855 );
not ( n326261 , n326260 );
buf ( n326262 , n325771 );
buf ( n326263 , n325749 );
nand ( n326264 , n326262 , n326263 );
buf ( n326265 , n326264 );
buf ( n326266 , n326265 );
not ( n326267 , n326266 );
and ( n35842 , n326261 , n326267 );
buf ( n326269 , n325852 );
buf ( n326270 , n325845 );
and ( n35845 , n326269 , n326270 );
buf ( n326272 , n35845 );
buf ( n326273 , n326272 );
nor ( n35848 , n35842 , n326273 );
buf ( n326275 , n35848 );
buf ( n326276 , n326275 );
not ( n35851 , n326276 );
and ( n326278 , n326259 , n35851 );
and ( n326279 , n35398 , n325840 );
not ( n326280 , n326279 );
not ( n35855 , n325818 );
or ( n326282 , n326280 , n35855 );
not ( n326283 , n35391 );
nand ( n35858 , n326283 , n325799 );
nand ( n326285 , n326282 , n35858 );
buf ( n35860 , n326285 );
nor ( n35861 , n326278 , n35860 );
buf ( n35862 , n35861 );
not ( n326289 , n35862 );
and ( n326290 , n326255 , n326289 );
not ( n326291 , n326253 );
buf ( n326292 , n35771 );
buf ( n326293 , n326192 );
and ( n326294 , n326292 , n326293 );
buf ( n326295 , n326294 );
not ( n326296 , n326295 );
not ( n35871 , n326185 );
or ( n35872 , n326296 , n35871 );
buf ( n326299 , n35756 );
not ( n326300 , n326299 );
buf ( n35875 , n326161 );
nand ( n35876 , n326300 , n35875 );
buf ( n35877 , n35876 );
nand ( n326304 , n35872 , n35877 );
not ( n35879 , n326304 );
or ( n326306 , n326291 , n35879 );
buf ( n326307 , n35812 );
not ( n35882 , n326307 );
buf ( n35883 , n35882 );
buf ( n326310 , n35883 );
buf ( n326311 , n326249 );
buf ( n326312 , n326246 );
and ( n35887 , n326311 , n326312 );
buf ( n326314 , n35887 );
buf ( n326315 , n326314 );
and ( n326316 , n326310 , n326315 );
buf ( n326317 , n326237 );
buf ( n326318 , n326223 );
and ( n326319 , n326317 , n326318 );
buf ( n326320 , n326319 );
buf ( n326321 , n326320 );
nor ( n326322 , n326316 , n326321 );
buf ( n326323 , n326322 );
nand ( n326324 , n326306 , n326323 );
nor ( n326325 , n326290 , n326324 );
nand ( n35900 , n326256 , n326325 );
xor ( n326327 , n15083 , n306402 );
and ( n35902 , n326327 , n306540 );
and ( n326329 , n15083 , n306402 );
or ( n326330 , n35902 , n326329 );
buf ( n326331 , n326330 );
or ( n35906 , n314469 , n326331 );
not ( n326333 , n35906 );
not ( n35908 , n33561 );
not ( n35909 , n35908 );
not ( n35910 , n33528 );
or ( n35911 , n35909 , n35910 );
not ( n35912 , n33216 );
nand ( n35913 , n35911 , n35912 );
nand ( n326340 , n33559 , n33571 );
xnor ( n35915 , n35913 , n326340 );
not ( n326342 , n35915 );
or ( n35917 , n326333 , n326342 );
nand ( n35918 , n314469 , n326331 );
nand ( n35919 , n35917 , n35918 );
xor ( n35920 , n314474 , n24021 );
not ( n35921 , n324002 );
nor ( n326348 , n35921 , n17077 );
xor ( n35923 , n33574 , n326348 );
xor ( n35924 , n35920 , n35923 );
or ( n35925 , n35919 , n35924 );
not ( n35926 , n323967 );
xnor ( n35927 , n314469 , n326331 );
xor ( n35928 , n35927 , n326340 );
xnor ( n35929 , n35928 , n35913 );
nand ( n35930 , n35926 , n35929 );
nand ( n326357 , n35925 , n35930 );
not ( n326358 , n326357 );
or ( n35933 , n314809 , n317419 );
not ( n326360 , n35933 );
not ( n326361 , n323950 );
nand ( n35936 , n326361 , n33516 );
not ( n326363 , n35936 );
buf ( n35938 , n33438 );
not ( n35939 , n35938 );
not ( n326366 , n323921 );
not ( n326367 , n326218 );
or ( n35942 , n326366 , n326367 );
buf ( n326369 , n323930 );
nand ( n326370 , n35942 , n326369 );
not ( n35945 , n326370 );
or ( n326372 , n35939 , n35945 );
nand ( n35947 , n326372 , n33508 );
not ( n326374 , n35947 );
or ( n35949 , n326363 , n326374 );
or ( n326376 , n35947 , n35936 );
nand ( n35951 , n35949 , n326376 );
not ( n35952 , n35951 );
or ( n326379 , n326360 , n35952 );
nand ( n326380 , n314809 , n317419 );
nand ( n35955 , n326379 , n326380 );
not ( n326382 , n35955 );
not ( n326383 , n323962 );
and ( n35958 , n326382 , n326383 );
not ( n326385 , n317419 );
not ( n326386 , n314809 );
or ( n326387 , n326385 , n326386 );
or ( n35962 , n314809 , n317419 );
nand ( n326389 , n326387 , n35962 );
xor ( n35964 , n326389 , n35936 );
xor ( n326391 , n35964 , n35947 );
not ( n326392 , n326391 );
or ( n35967 , n315690 , n317414 );
not ( n326394 , n35967 );
nand ( n326395 , n35938 , n33508 );
not ( n326396 , n326395 );
and ( n35971 , n326370 , n326396 );
not ( n326398 , n326370 );
and ( n35973 , n326398 , n326395 );
nor ( n35974 , n35971 , n35973 );
not ( n35975 , n35974 );
or ( n35976 , n326394 , n35975 );
nand ( n35977 , n317414 , n315690 );
nand ( n35978 , n35976 , n35977 );
not ( n35979 , n35978 );
and ( n35980 , n326392 , n35979 );
nor ( n35981 , n35958 , n35980 );
or ( n35982 , n318930 , n318983 );
not ( n35983 , n35982 );
and ( n326410 , n35780 , n35793 );
not ( n326411 , n35780 );
not ( n35986 , n35793 );
and ( n326413 , n326411 , n35986 );
or ( n326414 , n326410 , n326413 );
not ( n35989 , n326414 );
or ( n326416 , n35983 , n35989 );
nand ( n326417 , n318930 , n318983 );
nand ( n35992 , n326416 , n326417 );
not ( n326419 , n35992 );
not ( n35994 , n33503 );
nand ( n326421 , n35994 , n33498 );
nor ( n35996 , n323926 , n326421 );
not ( n35997 , n35996 );
not ( n326424 , n35986 );
or ( n326425 , n35997 , n326424 );
and ( n36000 , n326421 , n35779 );
and ( n326427 , n35793 , n36000 );
not ( n326428 , n323926 );
not ( n36003 , n326421 );
or ( n326430 , n326428 , n36003 );
or ( n326431 , n326421 , n323926 , n35779 );
nand ( n36006 , n326430 , n326431 );
nor ( n36007 , n326427 , n36006 );
nand ( n326434 , n326425 , n36007 );
xnor ( n36009 , n315685 , n318935 );
not ( n326436 , n36009 );
and ( n326437 , n326434 , n326436 );
not ( n36012 , n326434 );
and ( n326439 , n36012 , n36009 );
nor ( n36014 , n326437 , n326439 );
not ( n36015 , n36014 );
and ( n326442 , n326419 , n36015 );
or ( n36017 , n315685 , n318935 );
not ( n326444 , n36017 );
not ( n36019 , n326434 );
or ( n36020 , n326444 , n36019 );
nand ( n326447 , n315685 , n318935 );
nand ( n326448 , n36020 , n326447 );
not ( n36023 , n326448 );
xnor ( n326450 , n317414 , n315690 );
xnor ( n326451 , n326450 , n35974 );
not ( n36026 , n326451 );
and ( n326453 , n36023 , n36026 );
nor ( n326454 , n326442 , n326453 );
nand ( n36029 , n35981 , n326454 );
not ( n326456 , n36029 );
not ( n326457 , n24021 );
not ( n36032 , n314474 );
or ( n326459 , n326457 , n36032 );
or ( n326460 , n314474 , n24021 );
nand ( n36035 , n326460 , n35923 );
nand ( n326462 , n326459 , n36035 );
not ( n326463 , n326462 );
not ( n36038 , n326463 );
buf ( n326465 , n324009 );
not ( n326466 , n326465 );
buf ( n326467 , n326466 );
not ( n36042 , n326467 );
or ( n326469 , n36038 , n36042 );
not ( n326470 , n325548 );
xor ( n36045 , n35133 , n313446 );
not ( n36046 , n36045 );
and ( n326473 , n326470 , n36046 );
and ( n326474 , n325548 , n36045 );
nor ( n36049 , n326473 , n326474 );
not ( n36050 , n36049 );
not ( n326477 , n35121 );
or ( n36052 , n36050 , n326477 );
or ( n36053 , n35121 , n36049 );
nand ( n36054 , n36052 , n36053 );
not ( n36055 , n36054 );
buf ( n326482 , n324014 );
not ( n36057 , n326482 );
buf ( n326484 , n36057 );
nand ( n36059 , n36055 , n326484 );
nand ( n36060 , n326469 , n36059 );
not ( n326487 , n36060 );
nand ( n326488 , n35900 , n326358 , n326456 , n326487 );
not ( n36063 , n35981 );
nor ( n326490 , n326451 , n326448 );
not ( n326491 , n326490 );
not ( n36066 , n326491 );
buf ( n326493 , n35992 );
buf ( n326494 , n36014 );
nand ( n36069 , n326493 , n326494 );
buf ( n36070 , n36069 );
not ( n36071 , n36070 );
not ( n36072 , n36071 );
or ( n326499 , n36066 , n36072 );
buf ( n326500 , n326448 );
buf ( n326501 , n326451 );
nand ( n36076 , n326500 , n326501 );
buf ( n326503 , n36076 );
nand ( n36078 , n326499 , n326503 );
not ( n326505 , n36078 );
or ( n326506 , n36063 , n326505 );
buf ( n326507 , n35955 );
buf ( n326508 , n323962 );
nor ( n36083 , n326507 , n326508 );
buf ( n326510 , n36083 );
not ( n326511 , n326510 );
buf ( n326512 , n326391 );
buf ( n326513 , n35978 );
nand ( n36088 , n326512 , n326513 );
buf ( n326515 , n36088 );
not ( n36090 , n326515 );
and ( n36091 , n326511 , n36090 );
buf ( n326518 , n35955 );
buf ( n326519 , n323962 );
and ( n326520 , n326518 , n326519 );
buf ( n326521 , n326520 );
nor ( n326522 , n36091 , n326521 );
nand ( n326523 , n326506 , n326522 );
nor ( n36098 , n36060 , n326357 );
nand ( n326525 , n326523 , n36098 );
or ( n36100 , n35919 , n35924 );
not ( n36101 , n36100 );
nor ( n326528 , n35926 , n35929 );
not ( n326529 , n326528 );
or ( n36104 , n36101 , n326529 );
nand ( n326531 , n35919 , n35924 );
nand ( n326532 , n36104 , n326531 );
and ( n36107 , n326487 , n326532 );
not ( n326534 , n36059 );
and ( n36109 , n324009 , n326462 );
not ( n36110 , n36109 );
or ( n36111 , n326534 , n36110 );
buf ( n326538 , n326484 );
not ( n36113 , n326538 );
buf ( n326540 , n36054 );
nand ( n36115 , n36113 , n326540 );
buf ( n326542 , n36115 );
nand ( n36117 , n36111 , n326542 );
nor ( n36118 , n36107 , n36117 );
nand ( n36119 , n326488 , n326525 , n36118 );
buf ( n36120 , n36119 );
buf ( n326547 , n36120 );
buf ( n326548 , n35177 );
nand ( n36123 , n35198 , n35189 );
buf ( n326550 , n36123 );
nand ( n36125 , n326548 , n326550 );
buf ( n326552 , n36125 );
buf ( n326553 , n326552 );
buf ( n326554 , n325545 );
buf ( n326555 , n35137 );
or ( n36130 , n326554 , n326555 );
buf ( n36131 , n36130 );
buf ( n36132 , n36131 );
nand ( n326559 , n325607 , n325605 );
buf ( n36134 , n326559 );
nand ( n36135 , n36132 , n36134 );
buf ( n36136 , n36135 );
buf ( n36137 , n36136 );
nor ( n36138 , n326553 , n36137 );
buf ( n36139 , n36138 );
buf ( n36140 , n36139 );
buf ( n326567 , n35048 );
and ( n36142 , n36140 , n326567 );
buf ( n326569 , n36142 );
nand ( n326570 , n326569 , n325276 );
not ( n36145 , n326570 );
buf ( n326572 , n36145 );
buf ( n326573 , n324878 );
and ( n326574 , n326547 , n326572 , n326573 );
not ( n326575 , n324769 );
not ( n36150 , n34414 );
nand ( n36151 , n34436 , n324871 );
not ( n36152 , n36151 );
and ( n326579 , n324848 , n324340 );
not ( n36154 , n326579 );
or ( n36155 , n36152 , n36154 );
not ( n36156 , n34436 );
not ( n36157 , n324871 );
nand ( n36158 , n36156 , n36157 );
nand ( n326585 , n36155 , n36158 );
not ( n36160 , n326585 );
or ( n36161 , n36150 , n36160 );
not ( n36162 , n34389 );
nand ( n36163 , n324838 , n324830 );
not ( n36164 , n36163 );
and ( n36165 , n36162 , n36164 );
nand ( n36166 , n324781 , n34388 );
not ( n326593 , n36166 );
nor ( n36168 , n36165 , n326593 );
nand ( n326595 , n36161 , n36168 );
buf ( n36170 , n326595 );
not ( n326597 , n36170 );
or ( n326598 , n326575 , n326597 );
not ( n36173 , n34282 );
nor ( n326600 , n36173 , n324731 );
buf ( n326601 , n326600 );
not ( n36176 , n326601 );
buf ( n326603 , n324765 );
not ( n36178 , n326603 );
or ( n326605 , n36176 , n36178 );
not ( n36180 , n34317 );
and ( n326607 , n34229 , n36180 );
not ( n326608 , n34229 );
not ( n36183 , n324739 );
and ( n326610 , n326608 , n36183 );
or ( n36185 , n326607 , n326610 );
and ( n36186 , n324637 , n36185 );
not ( n36187 , n324637 );
not ( n36188 , n34317 );
and ( n36189 , n324652 , n36188 );
not ( n36190 , n324652 );
not ( n36191 , n324739 );
and ( n326618 , n36190 , n36191 );
or ( n36193 , n36189 , n326618 );
and ( n36194 , n36187 , n36193 );
or ( n36195 , n36186 , n36194 );
buf ( n326622 , n36195 );
buf ( n36197 , n34337 );
buf ( n326624 , n36197 );
nand ( n36199 , n326622 , n326624 );
buf ( n326626 , n36199 );
buf ( n326627 , n326626 );
nand ( n36202 , n326605 , n326627 );
buf ( n326629 , n36202 );
and ( n36204 , n324664 , n326629 );
nor ( n36205 , n324632 , n324660 );
nor ( n36206 , n36204 , n36205 );
nand ( n36207 , n326598 , n36206 );
buf ( n326634 , n36207 );
nor ( n36209 , n326574 , n326634 );
buf ( n326636 , n36209 );
buf ( n326637 , n326636 );
nand ( n36212 , n325724 , n326637 );
buf ( n326639 , n36212 );
buf ( n326640 , n326639 );
and ( n36215 , n326640 , n324618 );
not ( n36216 , n326640 );
and ( n36217 , n36216 , n324614 );
nor ( n36218 , n36215 , n36217 );
buf ( n326645 , n36218 );
not ( n36220 , n36205 );
nand ( n36221 , n36220 , n324664 );
buf ( n326648 , n36221 );
buf ( n326649 , n36221 );
not ( n36224 , n326649 );
buf ( n326651 , n36224 );
buf ( n326652 , n326651 );
nor ( n36227 , n34449 , n324766 );
buf ( n326654 , n36227 );
not ( n36229 , n326654 );
buf ( n326656 , n325721 );
not ( n36231 , n326656 );
or ( n36232 , n36229 , n36231 );
and ( n36233 , n36120 , n36145 , n36227 );
not ( n36234 , n326600 );
not ( n36235 , n324765 );
or ( n36236 , n36234 , n36235 );
nand ( n36237 , n36236 , n326626 );
not ( n36238 , n36237 );
not ( n36239 , n324766 );
nand ( n36240 , n36239 , n326595 );
nand ( n36241 , n36238 , n36240 );
nor ( n36242 , n36233 , n36241 );
buf ( n326669 , n36242 );
nand ( n36244 , n36232 , n326669 );
buf ( n326671 , n36244 );
buf ( n326672 , n326671 );
and ( n36247 , n326672 , n326652 );
not ( n36248 , n326672 );
and ( n36249 , n36248 , n326648 );
nor ( n36250 , n36247 , n36249 );
buf ( n326677 , n36250 );
buf ( n36252 , n36162 );
nand ( n36253 , n36166 , n36252 );
buf ( n326680 , n36253 );
buf ( n326681 , n36253 );
not ( n36256 , n326681 );
buf ( n326683 , n36256 );
buf ( n326684 , n326683 );
not ( n36259 , n326570 );
buf ( n36260 , n324873 );
not ( n36261 , n324839 );
nand ( n36262 , n36260 , n36261 );
not ( n36263 , n36262 );
nand ( n36264 , n36120 , n36259 , n36263 );
buf ( n326691 , n36264 );
not ( n36266 , n34644 );
not ( n36267 , n325105 );
and ( n36268 , n36266 , n36267 );
and ( n36269 , n325180 , n325220 );
nor ( n36270 , n36268 , n36269 );
nand ( n36271 , n34551 , n34611 );
and ( n36272 , n34848 , n36270 , n36271 );
not ( n36273 , n36272 );
nand ( n36274 , n35202 , n35229 , n325673 , n35249 );
not ( n36275 , n36274 );
or ( n36276 , n36273 , n36275 );
not ( n36277 , n35268 );
not ( n36278 , n325708 );
or ( n36279 , n36277 , n36278 );
nand ( n36280 , n36279 , n325718 );
buf ( n326707 , n325682 );
buf ( n326708 , n35261 );
nand ( n36283 , n326707 , n326708 );
buf ( n326710 , n36283 );
nor ( n36285 , n36280 , n326710 );
nand ( n36286 , n36276 , n36285 );
buf ( n326713 , n36286 );
nor ( n36288 , n36280 , n35272 );
buf ( n326715 , n36288 );
buf ( n326716 , n36262 );
nor ( n36291 , n326715 , n326716 );
buf ( n326718 , n36291 );
buf ( n326719 , n326718 );
nand ( n36294 , n326713 , n326719 );
buf ( n326721 , n36294 );
buf ( n326722 , n326721 );
buf ( n36297 , n326585 );
not ( n36298 , n36297 );
not ( n36299 , n36261 );
or ( n36300 , n36298 , n36299 );
not ( n36301 , n36164 );
nand ( n36302 , n36300 , n36301 );
buf ( n326729 , n36302 );
not ( n36304 , n326729 );
buf ( n326731 , n36304 );
buf ( n326732 , n326731 );
nand ( n36307 , n326691 , n326722 , n326732 );
buf ( n326734 , n36307 );
buf ( n326735 , n326734 );
and ( n36310 , n326735 , n326684 );
not ( n36311 , n326735 );
and ( n36312 , n36311 , n326680 );
nor ( n36313 , n36310 , n36312 );
buf ( n326740 , n36313 );
buf ( n326741 , n324368 );
buf ( n326742 , n324372 );
and ( n36317 , n326741 , n326742 );
buf ( n326744 , n36317 );
buf ( n326745 , n326744 );
buf ( n326746 , n324368 );
buf ( n326747 , n324372 );
nor ( n36322 , n326746 , n326747 );
buf ( n326749 , n36322 );
buf ( n326750 , n326749 );
nor ( n36325 , n326745 , n326750 );
buf ( n326752 , n36325 );
buf ( n326753 , n326752 );
not ( n36328 , n326753 );
buf ( n326755 , n36328 );
buf ( n326756 , n326755 );
buf ( n326757 , n326752 );
and ( n36332 , n831 , n309695 );
not ( n36333 , n831 );
and ( n36334 , n36333 , n310231 );
or ( n36335 , n36332 , n36334 );
and ( n36336 , n831 , n309643 );
not ( n36337 , n831 );
and ( n36338 , n36337 , n310317 );
or ( n36339 , n36336 , n36338 );
and ( n36340 , n36335 , n36339 );
not ( n36341 , n36340 );
nor ( n36342 , n36339 , n36335 );
not ( n36343 , n36342 );
nand ( n36344 , n36341 , n36343 );
not ( n36345 , n322350 );
not ( n36346 , n324589 );
or ( n36347 , n36345 , n36346 );
or ( n36348 , n322350 , n324589 );
nand ( n36349 , n36348 , n322269 );
nand ( n36350 , n36347 , n36349 );
xor ( n36351 , n322649 , n322353 );
xor ( n36352 , n321969 , n321985 );
xor ( n36353 , n36352 , n31566 );
and ( n36354 , n322857 , n36353 );
xor ( n36355 , n321969 , n321985 );
xor ( n36356 , n36355 , n31566 );
and ( n36357 , n322644 , n36356 );
and ( n36358 , n322857 , n322644 );
or ( n36359 , n36354 , n36357 , n36358 );
xor ( n36360 , n36351 , n36359 );
xor ( n36361 , n36350 , n36360 );
xor ( n36362 , n36344 , n36361 );
not ( n36363 , n324575 );
not ( n36364 , n324563 );
or ( n36365 , n36363 , n36364 );
nand ( n36366 , n36365 , n34150 );
xnor ( n36367 , n36362 , n36366 );
not ( n36368 , n34159 );
nand ( n36369 , n36368 , n34168 );
not ( n36370 , n36369 );
nor ( n36371 , n36370 , n324578 );
not ( n36372 , n36371 );
not ( n36373 , n324564 );
or ( n36374 , n36372 , n36373 );
not ( n36375 , n324564 );
not ( n36376 , n36369 );
nor ( n36377 , n36376 , n324577 );
and ( n36378 , n36375 , n36377 );
and ( n36379 , n34165 , n34159 );
nor ( n36380 , n36378 , n36379 );
nand ( n36381 , n36374 , n36380 );
nor ( n36382 , n36367 , n36381 );
not ( n36383 , n36382 );
not ( n36384 , n36366 );
or ( n36385 , n36350 , n36360 );
not ( n36386 , n36385 );
nor ( n36387 , n36386 , n36344 );
nand ( n36388 , n36384 , n36387 );
and ( n36389 , n36385 , n36344 );
nand ( n36390 , n36389 , n36366 );
nand ( n36391 , n36360 , n36350 );
nand ( n36392 , n36388 , n36390 , n36391 );
not ( n36393 , n36392 );
and ( n326820 , n831 , n309733 );
not ( n36395 , n831 );
and ( n36396 , n36395 , n310233 );
or ( n36397 , n326820 , n36396 );
and ( n36398 , n831 , n309765 );
not ( n326825 , n831 );
and ( n326826 , n326825 , n310237 );
or ( n36401 , n36398 , n326826 );
or ( n36402 , n36397 , n36401 );
not ( n36403 , n36402 );
and ( n36404 , n36397 , n36401 );
nor ( n326831 , n36403 , n36404 );
xor ( n326832 , n322649 , n322353 );
and ( n326833 , n326832 , n36359 );
and ( n36408 , n322649 , n322353 );
or ( n326835 , n326833 , n36408 );
xor ( n36410 , n326835 , n322013 );
xor ( n36411 , n326831 , n36410 );
and ( n326838 , n36343 , n324575 );
not ( n36413 , n326838 );
not ( n326840 , n324563 );
or ( n36415 , n36413 , n326840 );
not ( n326842 , n36342 );
not ( n326843 , n34150 );
and ( n36418 , n326842 , n326843 );
nor ( n326845 , n36418 , n36340 );
nand ( n326846 , n36415 , n326845 );
xor ( n36421 , n36411 , n326846 );
not ( n326848 , n36421 );
nand ( n36423 , n36393 , n326848 );
nand ( n326850 , n36383 , n36423 );
or ( n36425 , n326835 , n322013 );
not ( n36426 , n36425 );
not ( n36427 , n36404 );
nand ( n326854 , n36427 , n36402 );
not ( n36429 , n326854 );
and ( n326856 , n326846 , n36429 );
not ( n36431 , n326846 );
and ( n326858 , n36431 , n326854 );
nor ( n36433 , n326856 , n326858 );
not ( n36434 , n36433 );
or ( n326861 , n36426 , n36434 );
nand ( n326862 , n326835 , n322013 );
nand ( n326863 , n326861 , n326862 );
not ( n36438 , n326863 );
not ( n326865 , n36438 );
and ( n326866 , n831 , n310321 );
not ( n36441 , n831 );
and ( n326868 , n36441 , n310239 );
or ( n326869 , n326866 , n326868 );
and ( n36444 , n310241 , n5980 );
xor ( n326871 , n19591 , n19592 );
buf ( n326872 , n326871 );
and ( n36447 , n326872 , n831 );
nor ( n326874 , n36444 , n36447 );
and ( n326875 , n326869 , n326874 );
not ( n36450 , n326869 );
not ( n326877 , n326874 );
and ( n326878 , n36450 , n326877 );
nor ( n326879 , n326875 , n326878 );
not ( n36454 , n321876 );
not ( n326881 , n322018 );
xor ( n36456 , n36454 , n326881 );
xor ( n326883 , n326879 , n36456 );
and ( n326884 , n326838 , n36402 );
and ( n326885 , n324551 , n324542 , n326884 );
not ( n326886 , n326885 );
nand ( n36461 , n324282 , n324543 , n326884 );
not ( n326888 , n326838 );
not ( n326889 , n324561 );
or ( n36464 , n326888 , n326889 );
nand ( n326891 , n36464 , n326845 );
and ( n326892 , n36402 , n326891 );
nor ( n36467 , n326892 , n36404 );
nand ( n36468 , n326886 , n36461 , n36467 );
xnor ( n326895 , n326883 , n36468 );
buf ( n36470 , n326895 );
not ( n326897 , n36470 );
buf ( n326898 , n326897 );
not ( n326899 , n326898 );
or ( n36474 , n326865 , n326899 );
not ( n36475 , n36468 );
and ( n326902 , n36454 , n326881 );
nor ( n326903 , n326879 , n326902 );
nand ( n326904 , n36475 , n326903 );
not ( n36479 , n326902 );
nand ( n326906 , n36479 , n36468 , n326879 );
nand ( n326907 , n322018 , n321876 );
nand ( n36482 , n326904 , n326906 , n326907 );
buf ( n326909 , n36482 );
xor ( n326910 , n322526 , n322530 );
xor ( n36485 , n326910 , n322537 );
xor ( n326912 , n322778 , n322576 );
xor ( n326913 , n36485 , n326912 );
buf ( n326914 , n326913 );
buf ( n326915 , n321881 );
xor ( n36490 , n326914 , n326915 );
buf ( n326917 , n36490 );
buf ( n326918 , n326917 );
or ( n36493 , n326909 , n326918 );
buf ( n326920 , n36493 );
nand ( n326921 , n36474 , n326920 );
nor ( n326922 , n326850 , n326921 );
buf ( n326923 , n326922 );
and ( n326924 , n326914 , n326915 );
buf ( n326925 , n326924 );
buf ( n326926 , n326925 );
buf ( n326927 , n324360 );
or ( n326928 , n326926 , n326927 );
buf ( n326929 , n326928 );
buf ( n326930 , n326929 );
not ( n326931 , n326930 );
buf ( n326932 , n324362 );
buf ( n326933 , n324366 );
nor ( n326934 , n326932 , n326933 );
buf ( n326935 , n326934 );
buf ( n326936 , n326935 );
nor ( n326937 , n326931 , n326936 );
buf ( n326938 , n326937 );
buf ( n326939 , n326938 );
and ( n326940 , n326923 , n326939 );
buf ( n326941 , n326940 );
buf ( n326942 , n326941 );
not ( n36517 , n326942 );
nand ( n36518 , n34306 , n324661 , n34186 , n324765 );
not ( n36519 , n36518 );
not ( n326946 , n36519 );
not ( n326947 , n326595 );
or ( n36522 , n326946 , n326947 );
and ( n326949 , n324661 , n34186 );
and ( n36524 , n326949 , n36237 );
not ( n36525 , n34186 );
not ( n36526 , n36205 );
or ( n36527 , n36525 , n36526 );
nand ( n36528 , n36527 , n34184 );
nor ( n36529 , n36524 , n36528 );
nand ( n36530 , n36522 , n36529 );
buf ( n326957 , n36530 );
not ( n36532 , n326957 );
or ( n36533 , n36517 , n36532 );
buf ( n326960 , n326938 );
not ( n36535 , n326960 );
not ( n36536 , n326921 );
not ( n36537 , n36536 );
and ( n36538 , n36367 , n36381 );
buf ( n326965 , n36538 );
not ( n36540 , n326965 );
not ( n36541 , n36392 );
nand ( n36542 , n36541 , n326848 );
buf ( n326969 , n36542 );
not ( n36544 , n326969 );
or ( n36545 , n36540 , n36544 );
buf ( n326972 , n36421 );
buf ( n326973 , n36392 );
nand ( n36548 , n326972 , n326973 );
buf ( n326975 , n36548 );
buf ( n326976 , n326975 );
nand ( n36551 , n36545 , n326976 );
buf ( n326978 , n36551 );
not ( n36553 , n326978 );
or ( n36554 , n36537 , n36553 );
not ( n36555 , n36425 );
not ( n36556 , n36433 );
or ( n36557 , n36555 , n36556 );
nand ( n36558 , n36557 , n326862 );
buf ( n326985 , n36558 );
buf ( n326986 , n326895 );
and ( n36561 , n326985 , n326986 );
buf ( n326988 , n36561 );
buf ( n326989 , n326988 );
buf ( n326990 , n326920 );
and ( n36565 , n326989 , n326990 );
buf ( n326992 , n36482 );
buf ( n326993 , n326917 );
and ( n36568 , n326992 , n326993 );
buf ( n326995 , n36568 );
buf ( n326996 , n326995 );
nor ( n36571 , n36565 , n326996 );
buf ( n326998 , n36571 );
nand ( n36573 , n36554 , n326998 );
buf ( n327000 , n36573 );
not ( n36575 , n327000 );
or ( n36576 , n36535 , n36575 );
buf ( n327003 , n326925 );
buf ( n327004 , n324360 );
nand ( n36579 , n327003 , n327004 );
buf ( n327006 , n36579 );
buf ( n327007 , n327006 );
not ( n36582 , n327007 );
buf ( n327009 , n326935 );
not ( n36584 , n327009 );
and ( n36585 , n36582 , n36584 );
buf ( n327012 , n324362 );
buf ( n327013 , n324366 );
and ( n36588 , n327012 , n327013 );
buf ( n327015 , n36588 );
buf ( n327016 , n327015 );
nor ( n36591 , n36585 , n327016 );
buf ( n327018 , n36591 );
buf ( n327019 , n327018 );
nand ( n36594 , n36576 , n327019 );
buf ( n327021 , n36594 );
buf ( n327022 , n327021 );
not ( n36597 , n327022 );
buf ( n327024 , n36597 );
buf ( n327025 , n327024 );
nand ( n36600 , n36533 , n327025 );
buf ( n327027 , n36600 );
not ( n36602 , n327027 );
buf ( n327029 , n36286 );
buf ( n327030 , n326941 );
not ( n36605 , n324874 );
nand ( n36606 , n36519 , n36605 );
not ( n36607 , n36606 );
buf ( n327034 , n36607 );
and ( n36609 , n327030 , n327034 );
buf ( n327036 , n36609 );
buf ( n327037 , n327036 );
buf ( n327038 , n36288 );
not ( n36613 , n327038 );
buf ( n327040 , n36613 );
buf ( n327041 , n327040 );
nand ( n36616 , n327029 , n327037 , n327041 );
buf ( n327043 , n36616 );
buf ( n327044 , n327036 );
buf ( n327045 , n36120 );
buf ( n327046 , n36145 );
nand ( n36621 , n327044 , n327045 , n327046 );
buf ( n327048 , n36621 );
nand ( n36623 , n36602 , n327043 , n327048 );
buf ( n327050 , n36623 );
and ( n36625 , n327050 , n326757 );
not ( n36626 , n327050 );
and ( n36627 , n36626 , n326756 );
nor ( n36628 , n36625 , n36627 );
buf ( n327055 , n36628 );
buf ( n327056 , n327015 );
buf ( n327057 , n326935 );
nor ( n36632 , n327056 , n327057 );
buf ( n327059 , n36632 );
buf ( n327060 , n327059 );
not ( n36635 , n327060 );
buf ( n327062 , n36635 );
buf ( n327063 , n327062 );
buf ( n327064 , n327059 );
buf ( n327065 , n326922 );
buf ( n327066 , n326929 );
and ( n36641 , n327065 , n327066 );
buf ( n327068 , n36641 );
buf ( n327069 , n327068 );
not ( n36644 , n327069 );
buf ( n327071 , n36530 );
not ( n36646 , n327071 );
or ( n36647 , n36644 , n36646 );
buf ( n327074 , n326929 );
not ( n36649 , n327074 );
buf ( n327076 , n36573 );
not ( n36651 , n327076 );
or ( n36652 , n36649 , n36651 );
buf ( n327079 , n327006 );
nand ( n36654 , n36652 , n327079 );
buf ( n327081 , n36654 );
buf ( n327082 , n327081 );
not ( n36657 , n327082 );
buf ( n327084 , n36657 );
buf ( n327085 , n327084 );
nand ( n36660 , n36647 , n327085 );
buf ( n327087 , n36660 );
not ( n36662 , n327087 );
buf ( n327089 , n36286 );
and ( n36664 , n36519 , n36605 );
and ( n36665 , n36664 , n327068 );
buf ( n327092 , n36665 );
buf ( n327093 , n327040 );
nand ( n36668 , n327089 , n327092 , n327093 );
buf ( n327095 , n36668 );
buf ( n327096 , n36665 );
buf ( n327097 , n36120 );
buf ( n327098 , n36259 );
nand ( n36673 , n327096 , n327097 , n327098 );
buf ( n327100 , n36673 );
nand ( n36675 , n36662 , n327095 , n327100 );
buf ( n327102 , n36675 );
and ( n36677 , n327102 , n327064 );
not ( n36678 , n327102 );
and ( n36679 , n36678 , n327063 );
nor ( n36680 , n36677 , n36679 );
buf ( n327107 , n36680 );
nand ( n36682 , n35246 , n35232 );
buf ( n327109 , n36682 );
buf ( n327110 , n36682 );
not ( n36685 , n327110 );
buf ( n327112 , n36685 );
buf ( n327113 , n327112 );
buf ( n327114 , n34941 );
buf ( n36689 , n327114 );
buf ( n327116 , n36689 );
not ( n36691 , n327116 );
nor ( n36692 , n36691 , n35208 );
buf ( n327119 , n36692 );
not ( n36694 , n327119 );
buf ( n327121 , n36139 );
not ( n36696 , n327121 );
buf ( n327123 , n36696 );
buf ( n327124 , n327123 );
nor ( n327125 , n36694 , n327124 );
buf ( n327126 , n327125 );
buf ( n327127 , n327126 );
not ( n36702 , n327127 );
buf ( n327129 , n36120 );
not ( n327130 , n327129 );
or ( n327131 , n36702 , n327130 );
not ( n327132 , n325641 );
or ( n36707 , n325604 , n325626 );
nand ( n327134 , n327132 , n36707 );
and ( n327135 , n36692 , n327134 );
not ( n36710 , n327116 );
not ( n327137 , n34991 );
not ( n327138 , n35233 );
not ( n36713 , n327138 );
or ( n327140 , n327137 , n36713 );
buf ( n36715 , n35248 );
not ( n327142 , n36715 );
buf ( n327143 , n327142 );
nand ( n327144 , n327140 , n327143 );
not ( n36719 , n327144 );
or ( n36720 , n36710 , n36719 );
nand ( n327147 , n36720 , n35244 );
nor ( n327148 , n327135 , n327147 );
buf ( n327149 , n327148 );
nand ( n327150 , n327131 , n327149 );
buf ( n327151 , n327150 );
buf ( n327152 , n327151 );
and ( n327153 , n327152 , n327113 );
not ( n36728 , n327152 );
and ( n327155 , n36728 , n327109 );
nor ( n327156 , n327153 , n327155 );
buf ( n327157 , n327156 );
buf ( n327158 , n34848 );
buf ( n327159 , n327158 );
buf ( n327160 , n327159 );
buf ( n327161 , n327160 );
buf ( n327162 , n35258 );
not ( n36737 , n327162 );
buf ( n327164 , n36737 );
buf ( n327165 , n327164 );
nand ( n36740 , n327161 , n327165 );
buf ( n327167 , n36740 );
buf ( n327168 , n327167 );
buf ( n327169 , n327167 );
not ( n36744 , n327169 );
buf ( n327171 , n36744 );
buf ( n327172 , n327171 );
buf ( n327173 , n326569 );
not ( n327174 , n327173 );
buf ( n327175 , n327174 );
buf ( n327176 , n327175 );
nand ( n327177 , n36271 , n34681 );
buf ( n327178 , n327177 );
nor ( n36753 , n327176 , n327178 );
buf ( n327180 , n36753 );
buf ( n327181 , n327180 );
not ( n36756 , n327181 );
buf ( n327183 , n36120 );
not ( n327184 , n327183 );
or ( n327185 , n36756 , n327184 );
buf ( n327186 , n35250 );
buf ( n327187 , n327186 );
buf ( n327188 , n327187 );
buf ( n327189 , n327188 );
buf ( n327190 , n327177 );
not ( n327191 , n327190 );
buf ( n327192 , n327191 );
buf ( n327193 , n327192 );
and ( n327194 , n327189 , n327193 );
buf ( n327195 , n34681 );
not ( n327196 , n327195 );
buf ( n327197 , n327196 );
buf ( n327198 , n327197 );
buf ( n327199 , n35254 );
or ( n36774 , n327198 , n327199 );
buf ( n327201 , n35253 );
nand ( n327202 , n36774 , n327201 );
buf ( n327203 , n327202 );
buf ( n327204 , n327203 );
nor ( n327205 , n327194 , n327204 );
buf ( n327206 , n327205 );
buf ( n327207 , n327206 );
nand ( n327208 , n327185 , n327207 );
buf ( n327209 , n327208 );
buf ( n327210 , n327209 );
and ( n327211 , n327210 , n327172 );
not ( n36786 , n327210 );
and ( n36787 , n36786 , n327168 );
nor ( n36788 , n327211 , n36787 );
buf ( n327215 , n36788 );
or ( n327216 , n324340 , n324848 );
buf ( n327217 , n327216 );
buf ( n327218 , n326579 );
not ( n36793 , n327218 );
buf ( n327220 , n36793 );
buf ( n327221 , n327220 );
nand ( n327222 , n327217 , n327221 );
buf ( n327223 , n327222 );
buf ( n327224 , n327223 );
buf ( n327225 , n327223 );
not ( n327226 , n327225 );
buf ( n327227 , n327226 );
buf ( n327228 , n327227 );
buf ( n327229 , n36145 );
not ( n36804 , n327229 );
buf ( n327231 , n36120 );
not ( n36806 , n327231 );
or ( n327233 , n36804 , n36806 );
not ( n327234 , n325721 );
buf ( n327235 , n327234 );
nand ( n327236 , n327233 , n327235 );
buf ( n327237 , n327236 );
buf ( n327238 , n327237 );
and ( n36813 , n327238 , n327228 );
not ( n327240 , n327238 );
and ( n36815 , n327240 , n327224 );
nor ( n36816 , n36813 , n36815 );
buf ( n327243 , n36816 );
or ( n327244 , n35285 , n34637 );
nand ( n36819 , n327244 , n325715 );
buf ( n327246 , n36819 );
buf ( n327247 , n36819 );
not ( n36822 , n327247 );
buf ( n327249 , n36822 );
buf ( n327250 , n327249 );
not ( n327251 , n34821 );
nor ( n327252 , n327251 , n325697 );
buf ( n327253 , n327252 );
buf ( n327254 , n36272 );
nand ( n327255 , n327253 , n327254 );
buf ( n327256 , n327255 );
buf ( n327257 , n327256 );
buf ( n327258 , n327175 );
nor ( n327259 , n327257 , n327258 );
buf ( n327260 , n327259 );
buf ( n327261 , n327260 );
not ( n327262 , n327261 );
buf ( n327263 , n36120 );
not ( n327264 , n327263 );
or ( n36839 , n327262 , n327264 );
buf ( n327266 , n327256 );
not ( n327267 , n327266 );
buf ( n327268 , n327267 );
buf ( n327269 , n327268 );
buf ( n327270 , n327188 );
and ( n327271 , n327269 , n327270 );
buf ( n327272 , n327252 );
not ( n36847 , n327272 );
buf ( n327274 , n326710 );
not ( n327275 , n327274 );
or ( n36850 , n36847 , n327275 );
nand ( n327277 , n325708 , n34821 );
not ( n327278 , n327277 );
nor ( n327279 , n35266 , n325246 );
nor ( n327280 , n327278 , n327279 );
buf ( n327281 , n327280 );
nand ( n327282 , n36850 , n327281 );
buf ( n327283 , n327282 );
buf ( n327284 , n327283 );
nor ( n327285 , n327271 , n327284 );
buf ( n327286 , n327285 );
buf ( n327287 , n327286 );
nand ( n36862 , n36839 , n327287 );
buf ( n36863 , n36862 );
buf ( n327290 , n36863 );
and ( n327291 , n327290 , n327250 );
not ( n36866 , n327290 );
and ( n327293 , n36866 , n327246 );
nor ( n327294 , n327291 , n327293 );
buf ( n327295 , n327294 );
not ( n36870 , n327279 );
nand ( n327297 , n36870 , n34821 );
buf ( n327298 , n327297 );
buf ( n327299 , n327297 );
not ( n36874 , n327299 );
buf ( n327301 , n36874 );
buf ( n327302 , n327301 );
buf ( n327303 , n36272 );
not ( n327304 , n325697 );
buf ( n327305 , n327304 );
nand ( n36880 , n327303 , n327305 );
buf ( n327307 , n36880 );
buf ( n327308 , n327307 );
buf ( n327309 , n327175 );
nor ( n36884 , n327308 , n327309 );
buf ( n327311 , n36884 );
buf ( n327312 , n327311 );
not ( n36887 , n327312 );
buf ( n327314 , n36120 );
not ( n327315 , n327314 );
or ( n36890 , n36887 , n327315 );
buf ( n327317 , n36274 );
not ( n36892 , n327317 );
buf ( n327319 , n36892 );
buf ( n327320 , n327319 );
not ( n36895 , n327320 );
buf ( n327322 , n36895 );
buf ( n327323 , n327322 );
buf ( n327324 , n327307 );
not ( n36899 , n327324 );
buf ( n327326 , n36899 );
buf ( n327327 , n327326 );
and ( n36902 , n327323 , n327327 );
not ( n36903 , n327304 );
not ( n36904 , n35262 );
or ( n36905 , n36903 , n36904 );
not ( n36906 , n325708 );
nand ( n327333 , n36905 , n36906 );
buf ( n327334 , n327333 );
nor ( n36909 , n36902 , n327334 );
buf ( n327336 , n36909 );
buf ( n327337 , n327336 );
nand ( n327338 , n36890 , n327337 );
buf ( n327339 , n327338 );
buf ( n327340 , n327339 );
and ( n36915 , n327340 , n327302 );
not ( n36916 , n327340 );
and ( n36917 , n36916 , n327298 );
nor ( n327344 , n36915 , n36917 );
buf ( n327345 , n327344 );
buf ( n327346 , n325171 );
buf ( n327347 , n35281 );
nand ( n36922 , n327346 , n327347 );
buf ( n327349 , n36922 );
buf ( n327350 , n327349 );
buf ( n327351 , n327349 );
not ( n36926 , n327351 );
buf ( n327353 , n36926 );
buf ( n327354 , n327353 );
buf ( n327355 , n325696 );
buf ( n36930 , n327355 );
buf ( n327357 , n36930 );
buf ( n327358 , n327357 );
buf ( n327359 , n36272 );
nand ( n36934 , n327358 , n327359 );
buf ( n327361 , n36934 );
buf ( n327362 , n327361 );
buf ( n327363 , n327175 );
nor ( n36938 , n327362 , n327363 );
buf ( n327365 , n36938 );
buf ( n327366 , n327365 );
not ( n36941 , n327366 );
buf ( n327368 , n36120 );
not ( n36943 , n327368 );
or ( n36944 , n36941 , n36943 );
buf ( n327371 , n327322 );
buf ( n327372 , n327361 );
not ( n36947 , n327372 );
buf ( n327374 , n36947 );
buf ( n327375 , n327374 );
and ( n36950 , n327371 , n327375 );
not ( n36951 , n327357 );
not ( n36952 , n326710 );
or ( n36953 , n36951 , n36952 );
buf ( n36954 , n35276 );
not ( n36955 , n36954 );
nand ( n36956 , n36953 , n36955 );
buf ( n327383 , n36956 );
nor ( n36958 , n36950 , n327383 );
buf ( n327385 , n36958 );
buf ( n327386 , n327385 );
nand ( n36961 , n36944 , n327386 );
buf ( n327388 , n36961 );
buf ( n327389 , n327388 );
and ( n36964 , n327389 , n327354 );
not ( n36965 , n327389 );
and ( n36966 , n36965 , n327350 );
nor ( n36967 , n36964 , n36966 );
buf ( n327394 , n36967 );
buf ( n327395 , n325686 );
not ( n36970 , n327395 );
buf ( n327397 , n325221 );
nand ( n36972 , n36970 , n327397 );
buf ( n327399 , n36972 );
buf ( n327400 , n327399 );
buf ( n327401 , n327399 );
not ( n36976 , n327401 );
buf ( n327403 , n36976 );
buf ( n327404 , n327403 );
buf ( n327405 , n327192 );
buf ( n327406 , n327160 );
and ( n36981 , n327405 , n327406 );
buf ( n327408 , n36981 );
buf ( n327409 , n327408 );
not ( n36984 , n327409 );
buf ( n327411 , n327175 );
nor ( n36986 , n36984 , n327411 );
buf ( n327413 , n36986 );
buf ( n327414 , n327413 );
not ( n36989 , n327414 );
buf ( n327416 , n36120 );
not ( n36991 , n327416 );
or ( n36992 , n36989 , n36991 );
not ( n36993 , n327177 );
nand ( n36994 , n36993 , n327160 , n36274 );
not ( n36995 , n36994 );
buf ( n327422 , n327160 );
not ( n36997 , n327422 );
buf ( n327424 , n327203 );
not ( n36999 , n327424 );
or ( n37000 , n36997 , n36999 );
buf ( n327427 , n327164 );
nand ( n37002 , n37000 , n327427 );
buf ( n327429 , n37002 );
nor ( n37004 , n36995 , n327429 );
buf ( n327431 , n37004 );
nand ( n37006 , n36992 , n327431 );
buf ( n327433 , n37006 );
buf ( n327434 , n327433 );
and ( n37009 , n327434 , n327404 );
not ( n37010 , n327434 );
and ( n37011 , n37010 , n327400 );
nor ( n37012 , n37009 , n37011 );
buf ( n327439 , n37012 );
buf ( n327440 , n35177 );
not ( n37015 , n325637 );
buf ( n327442 , n37015 );
nand ( n37017 , n327440 , n327442 );
buf ( n327444 , n37017 );
buf ( n327445 , n327444 );
buf ( n327446 , n327444 );
not ( n37021 , n327446 );
buf ( n327448 , n37021 );
buf ( n327449 , n327448 );
buf ( n327450 , n36136 );
not ( n37025 , n327450 );
buf ( n327452 , n37025 );
buf ( n327453 , n327452 );
not ( n37028 , n327453 );
buf ( n327455 , n36120 );
not ( n37030 , n327455 );
or ( n37031 , n37028 , n37030 );
buf ( n327458 , n325566 );
not ( n37033 , n327458 );
buf ( n327460 , n37033 );
buf ( n327461 , n327460 );
not ( n37036 , n327461 );
buf ( n327463 , n326559 );
not ( n37038 , n327463 );
or ( n37039 , n37036 , n37038 );
buf ( n327466 , n325541 );
nand ( n37041 , n37039 , n327466 );
buf ( n327468 , n37041 );
buf ( n327469 , n327468 );
not ( n37044 , n327469 );
buf ( n327471 , n37044 );
buf ( n327472 , n327471 );
nand ( n37047 , n37031 , n327472 );
buf ( n327474 , n37047 );
buf ( n327475 , n327474 );
and ( n37050 , n327475 , n327449 );
not ( n37051 , n327475 );
and ( n37052 , n37051 , n327445 );
nor ( n37053 , n37050 , n37052 );
buf ( n327480 , n37053 );
buf ( n327481 , n327138 );
not ( n37056 , n327481 );
buf ( n327483 , n37056 );
nand ( n37058 , n327483 , n35046 );
buf ( n327485 , n37058 );
buf ( n327486 , n37058 );
not ( n37061 , n327486 );
buf ( n327488 , n37061 );
buf ( n327489 , n327488 );
buf ( n327490 , n36139 );
not ( n37065 , n327490 );
buf ( n327492 , n36120 );
not ( n37067 , n327492 );
or ( n37068 , n37065 , n37067 );
buf ( n327495 , n327134 );
not ( n37070 , n327495 );
buf ( n327497 , n37070 );
buf ( n327498 , n327497 );
nand ( n327499 , n37068 , n327498 );
buf ( n327500 , n327499 );
buf ( n327501 , n327500 );
and ( n37076 , n327501 , n327489 );
not ( n37077 , n327501 );
and ( n327504 , n37077 , n327485 );
nor ( n327505 , n37076 , n327504 );
buf ( n327506 , n327505 );
buf ( n37081 , n36123 );
buf ( n327508 , n35214 );
nand ( n327509 , n37081 , n327508 );
buf ( n327510 , n327509 );
buf ( n327511 , n327510 );
buf ( n327512 , n327510 );
not ( n37087 , n327512 );
buf ( n327514 , n37087 );
buf ( n327515 , n327514 );
buf ( n327516 , n35177 );
not ( n37091 , n327516 );
buf ( n327518 , n36136 );
nor ( n327519 , n37091 , n327518 );
buf ( n327520 , n327519 );
buf ( n327521 , n327520 );
not ( n327522 , n327521 );
buf ( n327523 , n36120 );
not ( n327524 , n327523 );
or ( n327525 , n327522 , n327524 );
buf ( n327526 , n35177 );
not ( n37101 , n327526 );
buf ( n327528 , n327468 );
not ( n37103 , n327528 );
or ( n327530 , n37101 , n37103 );
buf ( n327531 , n37015 );
nand ( n37106 , n327530 , n327531 );
buf ( n327533 , n37106 );
buf ( n327534 , n327533 );
not ( n327535 , n327534 );
buf ( n327536 , n327535 );
buf ( n327537 , n327536 );
nand ( n327538 , n327525 , n327537 );
buf ( n327539 , n327538 );
buf ( n327540 , n327539 );
and ( n327541 , n327540 , n327515 );
not ( n327542 , n327540 );
and ( n37117 , n327542 , n327511 );
nor ( n327544 , n327541 , n37117 );
buf ( n327545 , n327544 );
buf ( n327546 , n326559 );
buf ( n37121 , n325541 );
nand ( n37122 , n327546 , n37121 );
buf ( n37123 , n37122 );
buf ( n327550 , n37123 );
buf ( n327551 , n37123 );
not ( n327552 , n327551 );
buf ( n327553 , n327552 );
buf ( n327554 , n327553 );
buf ( n327555 , n36131 );
not ( n327556 , n327555 );
buf ( n327557 , n36120 );
not ( n327558 , n327557 );
or ( n327559 , n327556 , n327558 );
buf ( n37134 , n327460 );
not ( n37135 , n37134 );
buf ( n37136 , n37135 );
buf ( n327563 , n37136 );
nand ( n37138 , n327559 , n327563 );
buf ( n327565 , n37138 );
buf ( n327566 , n327565 );
and ( n37141 , n327566 , n327554 );
not ( n37142 , n327566 );
and ( n327569 , n37142 , n327550 );
nor ( n327570 , n37141 , n327569 );
buf ( n327571 , n327570 );
not ( n37146 , n36954 );
nand ( n327573 , n37146 , n327357 );
buf ( n327574 , n327573 );
buf ( n327575 , n327573 );
not ( n327576 , n327575 );
buf ( n327577 , n327576 );
buf ( n327578 , n327577 );
buf ( n327579 , n36272 );
not ( n327580 , n327579 );
buf ( n327581 , n327175 );
nor ( n37156 , n327580 , n327581 );
buf ( n327583 , n37156 );
buf ( n327584 , n327583 );
not ( n37159 , n327584 );
buf ( n327586 , n36120 );
not ( n327587 , n327586 );
or ( n327588 , n37159 , n327587 );
and ( n37163 , n36274 , n36272 );
buf ( n327590 , n37163 );
buf ( n37165 , n35262 );
buf ( n327592 , n37165 );
nor ( n327593 , n327590 , n327592 );
buf ( n327594 , n327593 );
buf ( n327595 , n327594 );
nand ( n327596 , n327588 , n327595 );
buf ( n327597 , n327596 );
buf ( n327598 , n327597 );
and ( n327599 , n327598 , n327578 );
not ( n37174 , n327598 );
and ( n327601 , n37174 , n327574 );
nor ( n327602 , n327599 , n327601 );
buf ( n327603 , n327602 );
buf ( n327604 , n327197 );
not ( n327605 , n327604 );
buf ( n327606 , n35253 );
nand ( n37181 , n327605 , n327606 );
buf ( n327608 , n37181 );
buf ( n327609 , n327608 );
buf ( n327610 , n327608 );
not ( n37185 , n327610 );
buf ( n327612 , n37185 );
buf ( n327613 , n327612 );
buf ( n327614 , n36271 );
not ( n327615 , n327614 );
buf ( n327616 , n327175 );
nor ( n37191 , n327615 , n327616 );
buf ( n327618 , n37191 );
buf ( n327619 , n327618 );
not ( n327620 , n327619 );
buf ( n327621 , n36120 );
not ( n327622 , n327621 );
or ( n327623 , n327620 , n327622 );
buf ( n327624 , n36271 );
not ( n37199 , n327624 );
buf ( n327626 , n35250 );
not ( n327627 , n327626 );
or ( n37202 , n37199 , n327627 );
buf ( n327629 , n35254 );
nand ( n37204 , n37202 , n327629 );
buf ( n327631 , n37204 );
buf ( n327632 , n327631 );
not ( n327633 , n327632 );
buf ( n327634 , n327633 );
buf ( n327635 , n327634 );
nand ( n327636 , n327623 , n327635 );
buf ( n327637 , n327636 );
buf ( n327638 , n327637 );
and ( n37213 , n327638 , n327613 );
not ( n37214 , n327638 );
and ( n37215 , n37214 , n327609 );
nor ( n37216 , n37213 , n37215 );
buf ( n327643 , n37216 );
nand ( n327644 , n327116 , n35244 );
buf ( n327645 , n327644 );
buf ( n327646 , n327644 );
not ( n37221 , n327646 );
buf ( n327648 , n37221 );
buf ( n327649 , n327648 );
not ( n37224 , n35208 );
nand ( n37225 , n37224 , n36139 );
not ( n37226 , n37225 );
buf ( n327653 , n37226 );
not ( n37228 , n327653 );
buf ( n327655 , n36120 );
not ( n327656 , n327655 );
or ( n37231 , n37228 , n327656 );
not ( n37232 , n37224 );
not ( n37233 , n327134 );
or ( n37234 , n37232 , n37233 );
buf ( n327661 , n327144 );
not ( n37236 , n327661 );
buf ( n327663 , n37236 );
nand ( n327664 , n37234 , n327663 );
buf ( n327665 , n327664 );
not ( n37240 , n327665 );
buf ( n327667 , n37240 );
buf ( n327668 , n327667 );
nand ( n327669 , n37231 , n327668 );
buf ( n327670 , n327669 );
buf ( n327671 , n327670 );
and ( n327672 , n327671 , n327649 );
not ( n37247 , n327671 );
and ( n327674 , n37247 , n327645 );
nor ( n327675 , n327672 , n327674 );
buf ( n327676 , n327675 );
nand ( n37251 , n326503 , n326491 );
buf ( n327678 , n37251 );
buf ( n327679 , n37251 );
not ( n327680 , n327679 );
buf ( n327681 , n327680 );
buf ( n327682 , n327681 );
buf ( n327683 , n326325 );
not ( n37258 , n327683 );
nor ( n327685 , n36014 , n35992 );
not ( n327686 , n327685 );
nand ( n37261 , n37258 , n327686 );
buf ( n327688 , n37261 );
nor ( n327689 , n326254 , n35431 );
buf ( n37264 , n327689 );
buf ( n327691 , n37264 );
not ( n327692 , n35719 );
nor ( n37267 , n327692 , n327685 );
buf ( n327694 , n37267 );
nand ( n327695 , n327691 , n327694 );
buf ( n327696 , n327695 );
buf ( n327697 , n327696 );
buf ( n37272 , n36070 );
buf ( n327699 , n37272 );
nand ( n37274 , n327688 , n327697 , n327699 );
buf ( n327701 , n37274 );
buf ( n327702 , n327701 );
and ( n327703 , n327702 , n327682 );
not ( n37278 , n327702 );
and ( n37279 , n37278 , n327678 );
nor ( n327706 , n327703 , n37279 );
buf ( n327707 , n327706 );
nor ( n37282 , n326391 , n35978 );
not ( n327709 , n37282 );
buf ( n327710 , n327709 );
buf ( n327711 , n326515 );
nand ( n37286 , n327710 , n327711 );
buf ( n327713 , n37286 );
buf ( n327714 , n327713 );
buf ( n327715 , n327713 );
not ( n327716 , n327715 );
buf ( n327717 , n327716 );
buf ( n327718 , n327717 );
buf ( n327719 , n326454 );
not ( n37294 , n327719 );
not ( n37295 , n37258 );
or ( n37296 , n37294 , n37295 );
buf ( n37297 , n35719 );
and ( n37298 , n37297 , n327719 );
and ( n327725 , n37298 , n37264 );
nor ( n327726 , n327725 , n36078 );
nand ( n37301 , n37296 , n327726 );
buf ( n327728 , n37301 );
and ( n327729 , n327728 , n327718 );
not ( n37304 , n327728 );
and ( n37305 , n37304 , n327714 );
nor ( n37306 , n327729 , n37305 );
buf ( n327733 , n37306 );
buf ( n327734 , n36059 );
buf ( n37309 , n326542 );
nand ( n37310 , n327734 , n37309 );
buf ( n327737 , n37310 );
buf ( n327738 , n327737 );
buf ( n327739 , n327737 );
not ( n327740 , n327739 );
buf ( n327741 , n327740 );
buf ( n327742 , n327741 );
nand ( n327743 , n326463 , n326467 );
not ( n327744 , n326357 );
and ( n327745 , n327743 , n327744 );
buf ( n327746 , n327745 );
not ( n327747 , n327746 );
not ( n327748 , n326523 );
not ( n37323 , n327748 );
buf ( n327750 , n37323 );
not ( n327751 , n327750 );
or ( n37326 , n327747 , n327751 );
buf ( n327753 , n327743 );
not ( n327754 , n327753 );
buf ( n327755 , n326532 );
not ( n37330 , n327755 );
or ( n37331 , n327754 , n37330 );
buf ( n37332 , n36109 );
not ( n37333 , n37332 );
buf ( n327760 , n37333 );
buf ( n327761 , n327760 );
nand ( n327762 , n37331 , n327761 );
buf ( n327763 , n327762 );
buf ( n327764 , n327763 );
not ( n327765 , n327764 );
buf ( n327766 , n327765 );
buf ( n327767 , n327766 );
nand ( n327768 , n37326 , n327767 );
buf ( n327769 , n327768 );
buf ( n327770 , n327769 );
not ( n327771 , n327770 );
buf ( n327772 , n327771 );
buf ( n327773 , n327772 );
buf ( n327774 , n327745 );
buf ( n327775 , n326456 );
and ( n37350 , n327774 , n327775 );
buf ( n327777 , n37350 );
buf ( n327778 , n327777 );
buf ( n37353 , n326256 );
not ( n327780 , n37353 );
buf ( n327781 , n327780 );
buf ( n327782 , n327781 );
nand ( n327783 , n327778 , n327782 );
buf ( n327784 , n327783 );
buf ( n327785 , n327784 );
buf ( n327786 , n327777 );
buf ( n327787 , n37258 );
nand ( n327788 , n327786 , n327787 );
buf ( n327789 , n327788 );
buf ( n327790 , n327789 );
nand ( n327791 , n327773 , n327785 , n327790 );
buf ( n327792 , n327791 );
buf ( n327793 , n327792 );
and ( n327794 , n327793 , n327742 );
not ( n327795 , n327793 );
and ( n37370 , n327795 , n327738 );
nor ( n37371 , n327794 , n37370 );
buf ( n327798 , n37371 );
buf ( n327799 , n327743 );
buf ( n327800 , n327760 );
nand ( n327801 , n327799 , n327800 );
buf ( n327802 , n327801 );
buf ( n327803 , n327802 );
buf ( n327804 , n327802 );
not ( n37379 , n327804 );
buf ( n327806 , n37379 );
buf ( n327807 , n327806 );
and ( n37382 , n326456 , n326358 );
nand ( n37383 , n37258 , n37382 );
buf ( n327810 , n37383 );
buf ( n327811 , n37382 );
buf ( n327812 , n327781 );
nand ( n37387 , n327811 , n327812 );
buf ( n327814 , n37387 );
buf ( n327815 , n327814 );
buf ( n327816 , n37323 );
buf ( n327817 , n326358 );
and ( n37392 , n327816 , n327817 );
buf ( n327819 , n326532 );
nor ( n37394 , n37392 , n327819 );
buf ( n327821 , n37394 );
buf ( n327822 , n327821 );
nand ( n37397 , n327810 , n327815 , n327822 );
buf ( n327824 , n37397 );
buf ( n327825 , n327824 );
and ( n37400 , n327825 , n327807 );
not ( n37401 , n327825 );
and ( n37402 , n37401 , n327803 );
nor ( n37403 , n37400 , n37402 );
buf ( n327830 , n37403 );
nand ( n37405 , n36100 , n326531 );
buf ( n327832 , n37405 );
buf ( n327833 , n37405 );
not ( n37408 , n327833 );
buf ( n327835 , n37408 );
buf ( n327836 , n327835 );
or ( n37411 , n37258 , n327781 );
buf ( n327838 , n326456 );
buf ( n327839 , n35930 );
and ( n37414 , n327838 , n327839 );
buf ( n327841 , n37414 );
nand ( n37416 , n37411 , n327841 );
and ( n37417 , n37323 , n35930 );
nor ( n37418 , n37417 , n326528 );
nand ( n37419 , n37416 , n37418 );
buf ( n327846 , n37419 );
and ( n37421 , n327846 , n327836 );
not ( n37422 , n327846 );
and ( n37423 , n37422 , n327832 );
nor ( n37424 , n37421 , n37423 );
buf ( n327851 , n37424 );
buf ( n327852 , n326320 );
not ( n37427 , n327852 );
buf ( n327854 , n35883 );
nand ( n37429 , n37427 , n327854 );
buf ( n327856 , n37429 );
buf ( n327857 , n327856 );
buf ( n327858 , n327856 );
not ( n37433 , n327858 );
buf ( n327860 , n37433 );
buf ( n327861 , n327860 );
not ( n37436 , n326304 );
buf ( n327863 , n35824 );
not ( n37438 , n327863 );
buf ( n327865 , n37438 );
not ( n37440 , n327865 );
or ( n37441 , n37436 , n37440 );
buf ( n327868 , n326314 );
not ( n37443 , n327868 );
buf ( n327870 , n37443 );
nand ( n37445 , n37441 , n327870 );
buf ( n327872 , n37445 );
not ( n37447 , n327872 );
buf ( n37448 , n326201 );
and ( n37449 , n37448 , n327865 );
nand ( n37450 , n37297 , n37449 , n35432 );
buf ( n327877 , n37450 );
buf ( n327878 , n37449 );
not ( n37453 , n35862 );
buf ( n327880 , n37453 );
nand ( n37455 , n327878 , n327880 );
buf ( n327882 , n37455 );
buf ( n327883 , n327882 );
nand ( n37458 , n37447 , n327877 , n327883 );
buf ( n327885 , n37458 );
buf ( n327886 , n327885 );
and ( n37461 , n327886 , n327861 );
not ( n37462 , n327886 );
and ( n37463 , n37462 , n327857 );
nor ( n37464 , n37461 , n37463 );
buf ( n327891 , n37464 );
nand ( n37466 , n327686 , n36070 );
buf ( n327893 , n37466 );
buf ( n327894 , n37466 );
not ( n37469 , n327894 );
buf ( n327896 , n37469 );
buf ( n327897 , n327896 );
not ( n37472 , n327689 );
not ( n37473 , n35719 );
or ( n37474 , n37472 , n37473 );
nand ( n37475 , n37474 , n326325 );
buf ( n327902 , n37475 );
and ( n37477 , n327902 , n327897 );
not ( n37478 , n327902 );
and ( n37479 , n37478 , n327893 );
nor ( n37480 , n37477 , n37479 );
buf ( n327907 , n37480 );
buf ( n327908 , n326185 );
buf ( n327909 , n35877 );
nand ( n37484 , n327908 , n327909 );
buf ( n327911 , n37484 );
buf ( n327912 , n327911 );
not ( n37487 , n327912 );
buf ( n327914 , n37487 );
buf ( n327915 , n327914 );
buf ( n327916 , n327911 );
not ( n37491 , n327692 );
nand ( n37492 , n35432 , n35772 );
not ( n37493 , n37492 );
and ( n37494 , n37491 , n37493 );
not ( n37495 , n35772 );
or ( n37496 , n35862 , n37495 );
not ( n37497 , n326295 );
nand ( n37498 , n37496 , n37497 );
nor ( n37499 , n37494 , n37498 );
buf ( n327926 , n37499 );
and ( n37501 , n327926 , n327916 );
not ( n37502 , n327926 );
and ( n37503 , n37502 , n327915 );
nor ( n37504 , n37501 , n37503 );
buf ( n327931 , n37504 );
nand ( n37506 , n325818 , n35858 );
buf ( n327933 , n37506 );
buf ( n327934 , n37506 );
not ( n37509 , n327934 );
buf ( n327936 , n37509 );
buf ( n327937 , n327936 );
buf ( n327938 , n35416 );
not ( n37513 , n325772 );
nor ( n37514 , n37513 , n325855 );
buf ( n327941 , n37514 );
and ( n37516 , n327938 , n327941 );
buf ( n327943 , n37516 );
buf ( n327944 , n327943 );
not ( n37519 , n327944 );
buf ( n327946 , n37297 );
not ( n37521 , n327946 );
or ( n37522 , n37519 , n37521 );
buf ( n327949 , n35416 );
buf ( n327950 , n326275 );
not ( n37525 , n327950 );
buf ( n327952 , n37525 );
buf ( n327953 , n327952 );
and ( n37528 , n327949 , n327953 );
not ( n37529 , n326279 );
buf ( n327956 , n37529 );
not ( n37531 , n327956 );
buf ( n327958 , n37531 );
buf ( n327959 , n327958 );
nor ( n37534 , n37528 , n327959 );
buf ( n327961 , n37534 );
buf ( n327962 , n327961 );
nand ( n37537 , n37522 , n327962 );
buf ( n327964 , n37537 );
buf ( n327965 , n327964 );
and ( n37540 , n327965 , n327937 );
not ( n37541 , n327965 );
and ( n37542 , n37541 , n327933 );
nor ( n37543 , n37540 , n37542 );
buf ( n327970 , n37543 );
buf ( n327971 , n35416 );
buf ( n327972 , n37529 );
nand ( n37547 , n327971 , n327972 );
buf ( n327974 , n37547 );
buf ( n327975 , n327974 );
buf ( n327976 , n327974 );
not ( n37551 , n327976 );
buf ( n327978 , n37551 );
buf ( n327979 , n327978 );
buf ( n327980 , n37514 );
not ( n37555 , n327980 );
buf ( n327982 , n37297 );
not ( n37557 , n327982 );
or ( n37558 , n37555 , n37557 );
buf ( n327985 , n326275 );
nand ( n37560 , n37558 , n327985 );
buf ( n327987 , n37560 );
buf ( n327988 , n327987 );
and ( n37563 , n327988 , n327979 );
not ( n37564 , n327988 );
and ( n37565 , n37564 , n327975 );
nor ( n37566 , n37563 , n37565 );
buf ( n327993 , n37566 );
buf ( n327994 , n325855 );
buf ( n327995 , n326272 );
nor ( n37570 , n327994 , n327995 );
buf ( n327997 , n37570 );
buf ( n327998 , n327997 );
not ( n37573 , n327998 );
buf ( n328000 , n37573 );
buf ( n328001 , n328000 );
buf ( n328002 , n327997 );
buf ( n328003 , n325772 );
not ( n37578 , n328003 );
buf ( n328005 , n37297 );
not ( n37580 , n328005 );
or ( n37581 , n37578 , n37580 );
buf ( n328008 , n326265 );
nand ( n37583 , n37581 , n328008 );
buf ( n328010 , n37583 );
buf ( n328011 , n328010 );
and ( n37586 , n328011 , n328002 );
not ( n37587 , n328011 );
and ( n37588 , n37587 , n328001 );
nor ( n37589 , n37586 , n37588 );
buf ( n328016 , n37589 );
buf ( n328017 , n327865 );
buf ( n328018 , n327870 );
nand ( n37593 , n328017 , n328018 );
buf ( n328020 , n37593 );
buf ( n328021 , n328020 );
not ( n37596 , n328021 );
buf ( n328023 , n37596 );
buf ( n328024 , n328023 );
buf ( n328025 , n328020 );
buf ( n328026 , n37448 );
not ( n328027 , n328026 );
buf ( n328028 , n37453 );
not ( n328029 , n328028 );
or ( n328030 , n328027 , n328029 );
not ( n37605 , n326304 );
buf ( n328032 , n37605 );
nand ( n328033 , n328030 , n328032 );
buf ( n328034 , n328033 );
buf ( n328035 , n328034 );
buf ( n328036 , n327692 );
nand ( n328037 , n35432 , n37448 );
buf ( n328038 , n328037 );
nor ( n37613 , n328036 , n328038 );
buf ( n328040 , n37613 );
buf ( n328041 , n328040 );
nor ( n328042 , n328035 , n328041 );
buf ( n328043 , n328042 );
buf ( n328044 , n328043 );
and ( n328045 , n328044 , n328025 );
not ( n328046 , n328044 );
and ( n37621 , n328046 , n328024 );
nor ( n37622 , n328045 , n37621 );
buf ( n328049 , n37622 );
buf ( n328050 , n326078 );
buf ( n328051 , n326140 );
nand ( n37626 , n328050 , n328051 );
buf ( n37627 , n37626 );
buf ( n328054 , n37627 );
buf ( n328055 , n37627 );
not ( n37630 , n328055 );
buf ( n328057 , n37630 );
buf ( n328058 , n328057 );
not ( n328059 , n35700 );
not ( n37634 , n326089 );
or ( n37635 , n328059 , n37634 );
buf ( n328062 , n326131 );
not ( n37637 , n328062 );
buf ( n328064 , n37637 );
nand ( n37639 , n37635 , n328064 );
buf ( n328066 , n37639 );
not ( n37641 , n328066 );
buf ( n328068 , n326089 );
not ( n37643 , n328068 );
buf ( n328070 , n326112 );
nor ( n37645 , n37643 , n328070 );
buf ( n328072 , n37645 );
buf ( n328073 , n328072 );
not ( n37648 , n35580 );
not ( n37649 , n326047 );
not ( n37650 , n37649 );
or ( n37651 , n37648 , n37650 );
buf ( n328078 , n326064 );
not ( n37653 , n328078 );
buf ( n328080 , n37653 );
nand ( n37655 , n37651 , n328080 );
buf ( n328082 , n37655 );
nand ( n37657 , n328073 , n328082 );
buf ( n328084 , n37657 );
buf ( n328085 , n328084 );
nor ( n37660 , n35568 , n326047 );
buf ( n328087 , n37660 );
buf ( n328088 , n328072 );
nand ( n37663 , n328087 , n328088 );
buf ( n328090 , n37663 );
buf ( n328091 , n328090 );
nand ( n37666 , n37641 , n328085 , n328091 );
buf ( n328093 , n37666 );
buf ( n328094 , n328093 );
and ( n37669 , n328094 , n328058 );
not ( n37670 , n328094 );
and ( n37671 , n37670 , n328054 );
nor ( n37672 , n37669 , n37671 );
buf ( n328099 , n37672 );
buf ( n328100 , n325867 );
buf ( n328101 , n326005 );
nand ( n37676 , n328100 , n328101 );
buf ( n328103 , n37676 );
buf ( n328104 , n328103 );
buf ( n328105 , n328103 );
not ( n328106 , n328105 );
buf ( n328107 , n328106 );
buf ( n328108 , n328107 );
buf ( n328109 , n325862 );
not ( n328110 , n328109 );
buf ( n328111 , n35567 );
not ( n328112 , n328111 );
or ( n37687 , n328110 , n328112 );
buf ( n328114 , n325998 );
not ( n37689 , n328114 );
buf ( n328116 , n37689 );
buf ( n328117 , n328116 );
nand ( n37692 , n37687 , n328117 );
buf ( n37693 , n37692 );
buf ( n328120 , n37693 );
and ( n37695 , n328120 , n328108 );
not ( n37696 , n328120 );
and ( n37697 , n37696 , n328104 );
nor ( n37698 , n37695 , n37697 );
buf ( n328125 , n37698 );
buf ( n328126 , n326098 );
buf ( n328127 , n35699 );
nand ( n37702 , n328126 , n328127 );
buf ( n328129 , n37702 );
buf ( n328130 , n328129 );
buf ( n328131 , n328129 );
not ( n37706 , n328131 );
buf ( n328133 , n37706 );
buf ( n37708 , n328133 );
buf ( n328135 , n37655 );
buf ( n328136 , n326109 );
nand ( n37711 , n328135 , n328136 );
buf ( n328138 , n37711 );
buf ( n328139 , n328138 );
buf ( n328140 , n37649 );
buf ( n328141 , n326109 );
buf ( n328142 , n325870 );
buf ( n328143 , n35567 );
nand ( n328144 , n328140 , n328141 , n328142 , n328143 );
buf ( n328145 , n328144 );
buf ( n37720 , n328145 );
buf ( n328147 , n326121 );
not ( n328148 , n328147 );
buf ( n328149 , n328148 );
buf ( n328150 , n328149 );
nand ( n37725 , n328139 , n37720 , n328150 );
buf ( n328152 , n37725 );
buf ( n328153 , n328152 );
and ( n328154 , n328153 , n37708 );
not ( n328155 , n328153 );
and ( n328156 , n328155 , n328130 );
nor ( n37731 , n328154 , n328156 );
buf ( n328158 , n37731 );
buf ( n328159 , n326046 );
buf ( n328160 , n326052 );
not ( n328161 , n328160 );
buf ( n328162 , n328161 );
buf ( n328163 , n328162 );
nand ( n328164 , n328159 , n328163 );
buf ( n328165 , n328164 );
buf ( n328166 , n328165 );
buf ( n37741 , n328165 );
not ( n328168 , n37741 );
buf ( n328169 , n328168 );
buf ( n37744 , n328169 );
buf ( n328171 , n325870 );
not ( n328172 , n328171 );
buf ( n328173 , n35567 );
not ( n37748 , n328173 );
or ( n328175 , n328172 , n37748 );
buf ( n328176 , n35581 );
nand ( n328177 , n328175 , n328176 );
buf ( n328178 , n328177 );
buf ( n328179 , n328178 );
and ( n328180 , n328179 , n37744 );
not ( n37755 , n328179 );
and ( n328182 , n37755 , n328166 );
nor ( n328183 , n328180 , n328182 );
buf ( n328184 , n328183 );
buf ( n328185 , n325989 );
buf ( n328186 , n325967 );
or ( n37761 , n328185 , n328186 );
buf ( n37762 , n37761 );
buf ( n328189 , n37762 );
buf ( n37764 , n325962 );
buf ( n328191 , n325972 );
not ( n37766 , n328191 );
buf ( n328193 , n37766 );
buf ( n328194 , n328193 );
nand ( n328195 , n37764 , n328194 );
buf ( n328196 , n328195 );
buf ( n328197 , n328196 );
buf ( n328198 , n328193 );
buf ( n37773 , n325907 );
nand ( n37774 , n328198 , n37773 );
buf ( n37775 , n37774 );
buf ( n328202 , n37775 );
buf ( n328203 , n325980 );
nand ( n37778 , n328197 , n328202 , n328203 );
buf ( n328205 , n37778 );
buf ( n328206 , n328205 );
buf ( n328207 , n37762 );
buf ( n328208 , n328205 );
not ( n328209 , n328189 );
not ( n37784 , n328206 );
or ( n328211 , n328209 , n37784 );
or ( n328212 , n328207 , n328208 );
nand ( n328213 , n328211 , n328212 );
buf ( n328214 , n328213 );
buf ( n328215 , n325962 );
buf ( n328216 , n325907 );
nor ( n328217 , n328215 , n328216 );
buf ( n328218 , n328217 );
buf ( n328219 , n328218 );
buf ( n328220 , n328193 );
buf ( n328221 , n325980 );
and ( n328222 , n328220 , n328221 );
buf ( n328223 , n328222 );
buf ( n328224 , n328223 );
buf ( n328225 , n328223 );
buf ( n328226 , n328218 );
not ( n328227 , n328219 );
not ( n328228 , n328224 );
or ( n37803 , n328227 , n328228 );
or ( n328230 , n328225 , n328226 );
nand ( n328231 , n37803 , n328230 );
buf ( n328232 , n328231 );
buf ( n328233 , n325910 );
buf ( n37808 , n325904 );
nand ( n37809 , n328233 , n37808 );
buf ( n37810 , n37809 );
buf ( n328237 , n37810 );
buf ( n328238 , n325959 );
not ( n328239 , n328238 );
buf ( n328240 , n35528 );
not ( n37815 , n328240 );
or ( n328242 , n328239 , n37815 );
buf ( n328243 , n325898 );
nand ( n37818 , n328242 , n328243 );
buf ( n328245 , n37818 );
buf ( n328246 , n328245 );
buf ( n328247 , n37810 );
buf ( n328248 , n328245 );
not ( n328249 , n328237 );
not ( n37824 , n328246 );
or ( n328251 , n328249 , n37824 );
or ( n328252 , n328247 , n328248 );
nand ( n37827 , n328251 , n328252 );
buf ( n328254 , n37827 );
buf ( n328255 , n325721 );
buf ( n328256 , n36607 );
not ( n328257 , n36382 );
nand ( n37832 , n328257 , n36423 );
buf ( n328259 , n37832 );
not ( n328260 , n328259 );
buf ( n328261 , n328260 );
buf ( n328262 , n328261 );
and ( n328263 , n328256 , n328262 );
buf ( n328264 , n328263 );
buf ( n328265 , n328264 );
nand ( n328266 , n328255 , n328265 );
buf ( n328267 , n328266 );
buf ( n328268 , n325721 );
buf ( n328269 , n36607 );
buf ( n328270 , n326863 );
not ( n37845 , n328270 );
buf ( n328272 , n326898 );
nand ( n328273 , n37845 , n328272 );
buf ( n328274 , n328273 );
not ( n328275 , n328274 );
nor ( n328276 , n328275 , n37832 );
buf ( n328277 , n328276 );
and ( n37852 , n328269 , n328277 );
buf ( n328279 , n37852 );
buf ( n328280 , n328279 );
nand ( n328281 , n328268 , n328280 );
buf ( n328282 , n328281 );
buf ( n328283 , n325721 );
buf ( n328284 , n36607 );
not ( n37859 , n36382 );
buf ( n328286 , n37859 );
and ( n328287 , n328284 , n328286 );
buf ( n328288 , n328287 );
buf ( n328289 , n328288 );
nand ( n37864 , n328283 , n328289 );
buf ( n328291 , n37864 );
buf ( n328292 , n325721 );
buf ( n328293 , n326922 );
buf ( n328294 , n328293 );
buf ( n328295 , n328294 );
and ( n37870 , n36607 , n328295 );
buf ( n328297 , n37870 );
nand ( n328298 , n328292 , n328297 );
buf ( n328299 , n328298 );
buf ( n328300 , n325947 );
not ( n37875 , n328300 );
buf ( n328302 , n325953 );
nand ( n37877 , n37875 , n328302 );
buf ( n37878 , n37877 );
buf ( n328305 , n37878 );
buf ( n328306 , n325941 );
buf ( n328307 , n325915 );
nand ( n328308 , n328306 , n328307 );
buf ( n328309 , n328308 );
buf ( n328310 , n328309 );
buf ( n328311 , n328309 );
buf ( n328312 , n37878 );
not ( n37887 , n328305 );
not ( n328314 , n328310 );
or ( n328315 , n37887 , n328314 );
or ( n37890 , n328311 , n328312 );
nand ( n328317 , n328315 , n37890 );
buf ( n328318 , n328317 );
buf ( n328319 , n36286 );
buf ( n328320 , n326922 );
buf ( n328321 , n326938 );
not ( n328322 , n328321 );
buf ( n328323 , n326749 );
nor ( n328324 , n328322 , n328323 );
buf ( n328325 , n328324 );
buf ( n328326 , n328325 );
and ( n328327 , n328320 , n328326 );
buf ( n328328 , n328327 );
and ( n328329 , n36664 , n328328 );
buf ( n328330 , n328329 );
buf ( n328331 , n327040 );
nand ( n328332 , n328319 , n328330 , n328331 );
buf ( n328333 , n328332 );
buf ( n328334 , n36286 );
buf ( n328335 , n36288 );
buf ( n37910 , n34449 );
nor ( n37911 , n328335 , n37910 );
buf ( n328338 , n37911 );
buf ( n328339 , n328338 );
nand ( n37914 , n328334 , n328339 );
buf ( n328341 , n37914 );
buf ( n328342 , n36286 );
buf ( n328343 , n36260 );
not ( n37918 , n328343 );
buf ( n328345 , n36288 );
nor ( n328346 , n37918 , n328345 );
buf ( n328347 , n328346 );
buf ( n328348 , n328347 );
nand ( n37923 , n328342 , n328348 );
buf ( n328350 , n37923 );
not ( n37925 , n324874 );
buf ( n328352 , n34306 );
buf ( n328353 , n328352 );
buf ( n328354 , n328353 );
nand ( n328355 , n37925 , n328354 );
buf ( n328356 , n328355 );
not ( n328357 , n328356 );
buf ( n328358 , n328357 );
buf ( n328359 , n328358 );
not ( n328360 , n328359 );
buf ( n328361 , n35294 );
not ( n37936 , n328361 );
buf ( n37937 , n37936 );
buf ( n328364 , n37937 );
not ( n37939 , n328364 );
or ( n328366 , n328360 , n37939 );
buf ( n328367 , n328354 );
not ( n328368 , n328367 );
buf ( n328369 , n36170 );
not ( n37944 , n328369 );
or ( n328371 , n328368 , n37944 );
buf ( n37946 , n326600 );
not ( n328373 , n37946 );
buf ( n328374 , n328373 );
buf ( n328375 , n328374 );
nand ( n328376 , n328371 , n328375 );
buf ( n328377 , n328376 );
buf ( n328378 , n328377 );
not ( n328379 , n328378 );
buf ( n328380 , n328379 );
buf ( n328381 , n328380 );
nand ( n328382 , n328366 , n328381 );
buf ( n328383 , n328382 );
buf ( n328384 , n328383 );
not ( n328385 , n328384 );
buf ( n328386 , n328385 );
buf ( n328387 , n36240 );
nor ( n328388 , n36528 , n326629 );
buf ( n328389 , n328388 );
nand ( n328390 , n328387 , n328389 );
buf ( n328391 , n328390 );
buf ( n328392 , n328391 );
buf ( n328393 , n328276 );
not ( n37968 , n328393 );
nor ( n37969 , n36528 , n326949 );
buf ( n328396 , n37969 );
nor ( n328397 , n37968 , n328396 );
buf ( n328398 , n328397 );
buf ( n328399 , n328398 );
nand ( n328400 , n326898 , n36438 );
buf ( n328401 , n328400 );
not ( n37976 , n328401 );
buf ( n328403 , n326978 );
not ( n37978 , n328403 );
or ( n37979 , n37976 , n37978 );
buf ( n328406 , n326988 );
not ( n328407 , n328406 );
buf ( n328408 , n328407 );
buf ( n328409 , n328408 );
nand ( n328410 , n37979 , n328409 );
buf ( n328411 , n328410 );
buf ( n328412 , n328411 );
and ( n328413 , n328392 , n328399 );
nor ( n37988 , n328413 , n328412 );
buf ( n37989 , n37988 );
buf ( n328416 , n37937 );
buf ( n328417 , n327216 );
nand ( n328418 , n328416 , n328417 );
buf ( n328419 , n328418 );
buf ( n328420 , n325920 );
buf ( n328421 , n325915 );
nand ( n328422 , n328420 , n328421 );
buf ( n328423 , n328422 );
buf ( n328424 , n328423 );
buf ( n328425 , n325938 );
buf ( n328426 , n325938 );
buf ( n328427 , n328423 );
not ( n38002 , n328424 );
not ( n38003 , n328425 );
or ( n328430 , n38002 , n38003 );
or ( n328431 , n328426 , n328427 );
nand ( n38006 , n328430 , n328431 );
buf ( n328433 , n38006 );
not ( n328434 , n35046 );
not ( n328435 , n327134 );
or ( n38010 , n328434 , n328435 );
nand ( n328437 , n38010 , n327483 );
buf ( n328438 , n328437 );
not ( n38013 , n328438 );
buf ( n328440 , n38013 );
buf ( n328441 , n328325 );
not ( n38016 , n328441 );
buf ( n328443 , n36573 );
not ( n328444 , n328443 );
or ( n38019 , n38016 , n328444 );
buf ( n328446 , n327018 );
not ( n38021 , n328446 );
buf ( n328448 , n326749 );
not ( n328449 , n328448 );
and ( n38024 , n38021 , n328449 );
buf ( n328451 , n326744 );
nor ( n328452 , n38024 , n328451 );
buf ( n328453 , n328452 );
buf ( n328454 , n328453 );
nand ( n38029 , n38019 , n328454 );
buf ( n328456 , n38029 );
buf ( n328457 , n328456 );
not ( n38032 , n328457 );
buf ( n328459 , n38032 );
xor ( n328460 , n325922 , n325933 );
xor ( n38035 , n328460 , n325935 );
buf ( n328462 , n38035 );
buf ( n328463 , n36573 );
not ( n38038 , n328463 );
buf ( n38039 , n38038 );
buf ( n328466 , n35580 );
buf ( n328467 , n326046 );
nand ( n328468 , n328466 , n328467 );
buf ( n328469 , n328468 );
xor ( n38044 , n325923 , n325930 );
buf ( n328471 , n38044 );
buf ( n328472 , n35772 );
buf ( n328473 , n37497 );
nand ( n328474 , n328472 , n328473 );
buf ( n328475 , n328474 );
buf ( n328476 , n328475 );
not ( n328477 , n328476 );
buf ( n328478 , n328477 );
buf ( n328479 , n326109 );
buf ( n328480 , n328149 );
nand ( n38055 , n328479 , n328480 );
buf ( n328482 , n38055 );
buf ( n38057 , n326112 );
not ( n328484 , n38057 );
buf ( n328485 , n328484 );
buf ( n328486 , n328116 );
buf ( n38061 , n325862 );
nand ( n38062 , n328486 , n38061 );
buf ( n38063 , n38062 );
buf ( n328490 , n36131 );
buf ( n328491 , n37136 );
nand ( n328492 , n328490 , n328491 );
buf ( n328493 , n328492 );
buf ( n328494 , n36538 );
not ( n328495 , n328494 );
buf ( n328496 , n328495 );
buf ( n328497 , n326978 );
not ( n38072 , n328497 );
buf ( n328499 , n38072 );
buf ( n328500 , n37660 );
buf ( n328501 , n37655 );
or ( n328502 , n328500 , n328501 );
buf ( n328503 , n328502 );
buf ( n328504 , n328503 );
buf ( n328505 , n328482 );
xnor ( n328506 , n328504 , n328505 );
buf ( n328507 , n328506 );
buf ( n328508 , n324574 );
buf ( n328509 , n324357 );
buf ( n328510 , n322566 );
xor ( n38085 , n328509 , n328510 );
buf ( n328512 , n324569 );
xor ( n328513 , n38085 , n328512 );
buf ( n328514 , n328513 );
buf ( n328515 , n328514 );
buf ( n328516 , n321881 );
buf ( n328517 , n326913 );
xor ( n38092 , n328516 , n328517 );
buf ( n328519 , n34092 );
and ( n328520 , n38092 , n328519 );
and ( n38095 , n328516 , n328517 );
or ( n328522 , n328520 , n38095 );
buf ( n328523 , n328522 );
buf ( n328524 , n328523 );
xor ( n328525 , n328508 , n328515 );
xor ( n328526 , n328525 , n328524 );
buf ( n328527 , n328526 );
xor ( n38102 , n328508 , n328515 );
and ( n38103 , n38102 , n328524 );
and ( n38104 , n328508 , n328515 );
or ( n38105 , n38103 , n38104 );
buf ( n38106 , n38105 );
not ( n328533 , n323767 );
buf ( n328534 , n328533 );
buf ( n328535 , n306542 );
buf ( n328536 , n314814 );
xor ( n38111 , n328535 , n328536 );
buf ( n328538 , n323889 );
and ( n38113 , n38111 , n328538 );
and ( n38114 , n328535 , n328536 );
or ( n328541 , n38113 , n38114 );
buf ( n328542 , n328541 );
buf ( n328543 , n328542 );
buf ( n328544 , n326331 );
buf ( n38119 , n314469 );
xor ( n38120 , n328544 , n38119 );
buf ( n328547 , n12778 );
xor ( n328548 , n38120 , n328547 );
buf ( n328549 , n328548 );
buf ( n328550 , n328549 );
xor ( n328551 , n328534 , n328543 );
xor ( n38126 , n328551 , n328550 );
buf ( n328553 , n38126 );
xor ( n38128 , n328534 , n328543 );
and ( n38129 , n38128 , n328550 );
and ( n38130 , n328534 , n328543 );
or ( n38131 , n38129 , n38130 );
buf ( n328558 , n38131 );
not ( n38133 , n33127 );
buf ( n328560 , n38133 );
buf ( n328561 , n320958 );
buf ( n328562 , n320496 );
xor ( n328563 , n328561 , n328562 );
buf ( n328564 , n10720 );
and ( n38139 , n328563 , n328564 );
and ( n328566 , n328561 , n328562 );
or ( n38141 , n38139 , n328566 );
buf ( n328568 , n38141 );
buf ( n328569 , n328568 );
buf ( n38144 , n320325 );
buf ( n328571 , n320501 );
xor ( n328572 , n38144 , n328571 );
not ( n328573 , n33123 );
buf ( n328574 , n328573 );
xor ( n328575 , n328572 , n328574 );
buf ( n328576 , n328575 );
buf ( n328577 , n328576 );
xor ( n38152 , n328560 , n328569 );
xor ( n38153 , n38152 , n328577 );
buf ( n328580 , n38153 );
xor ( n38155 , n328560 , n328569 );
and ( n38156 , n38155 , n328577 );
and ( n328583 , n328560 , n328569 );
or ( n38158 , n38156 , n328583 );
buf ( n328585 , n38158 );
buf ( n328586 , n33994 );
buf ( n328587 , n328586 );
buf ( n328588 , n322013 );
buf ( n328589 , n326835 );
xor ( n328590 , n328588 , n328589 );
buf ( n328591 , n33989 );
xor ( n38166 , n328590 , n328591 );
buf ( n328593 , n38166 );
buf ( n328594 , n328593 );
buf ( n328595 , n36350 );
buf ( n328596 , n36360 );
xor ( n328597 , n328595 , n328596 );
buf ( n328598 , n34002 );
and ( n328599 , n328597 , n328598 );
and ( n328600 , n328595 , n328596 );
or ( n38175 , n328599 , n328600 );
buf ( n328602 , n38175 );
buf ( n328603 , n328602 );
xor ( n38178 , n328587 , n328594 );
xor ( n328605 , n38178 , n328603 );
buf ( n328606 , n328605 );
xor ( n38181 , n328587 , n328594 );
and ( n38182 , n38181 , n328603 );
and ( n328609 , n328587 , n328594 );
or ( n38184 , n38182 , n328609 );
buf ( n328611 , n38184 );
buf ( n328612 , n322950 );
buf ( n328613 , n323205 );
xor ( n38188 , n328612 , n328613 );
buf ( n328615 , n323104 );
and ( n38190 , n38188 , n328615 );
and ( n328617 , n328612 , n328613 );
or ( n328618 , n38190 , n328617 );
buf ( n328619 , n328618 );
buf ( n328620 , n328619 );
buf ( n328621 , n32667 );
buf ( n328622 , n328621 );
buf ( n328623 , n35448 );
buf ( n328624 , n322952 );
xor ( n328625 , n328623 , n328624 );
buf ( n328626 , n323081 );
xor ( n328627 , n328625 , n328626 );
buf ( n328628 , n328627 );
buf ( n328629 , n328628 );
xor ( n38204 , n328620 , n328622 );
xor ( n328631 , n38204 , n328629 );
buf ( n328632 , n328631 );
xor ( n38207 , n328620 , n328622 );
and ( n328634 , n38207 , n328629 );
and ( n328635 , n328620 , n328622 );
or ( n328636 , n328634 , n328635 );
buf ( n328637 , n328636 );
nand ( n328638 , n33512 , n323935 );
buf ( n328639 , n328638 );
xor ( n38214 , n323862 , n313441 );
and ( n328641 , n38214 , n24026 );
and ( n328642 , n323862 , n313441 );
or ( n38217 , n328641 , n328642 );
buf ( n328644 , n38217 );
buf ( n328645 , n35133 );
buf ( n328646 , n313446 );
xor ( n328647 , n328645 , n328646 );
buf ( n328648 , n323941 );
buf ( n328649 , n328648 );
xor ( n328650 , n328647 , n328649 );
buf ( n328651 , n328650 );
buf ( n328652 , n328651 );
xor ( n328653 , n328639 , n328644 );
xor ( n328654 , n328653 , n328652 );
buf ( n328655 , n328654 );
xor ( n328656 , n328639 , n328644 );
and ( n328657 , n328656 , n328652 );
and ( n38232 , n328639 , n328644 );
or ( n38233 , n328657 , n38232 );
buf ( n328660 , n38233 );
not ( n328661 , n33356 );
buf ( n328662 , n328661 );
buf ( n328663 , n24021 );
buf ( n328664 , n314474 );
xor ( n38239 , n328663 , n328664 );
buf ( n328666 , n5939 );
xor ( n328667 , n38239 , n328666 );
buf ( n328668 , n328667 );
buf ( n328669 , n328668 );
xor ( n38244 , n328544 , n38119 );
and ( n38245 , n38244 , n328547 );
and ( n38246 , n328544 , n38119 );
or ( n38247 , n38245 , n38246 );
buf ( n38248 , n38247 );
buf ( n328675 , n38248 );
xor ( n38250 , n328662 , n328669 );
xor ( n38251 , n38250 , n328675 );
buf ( n328678 , n38251 );
xor ( n38253 , n328662 , n328669 );
and ( n328680 , n38253 , n328675 );
and ( n328681 , n328662 , n328669 );
or ( n38256 , n328680 , n328681 );
buf ( n328683 , n38256 );
buf ( n328684 , n322630 );
buf ( n328685 , n322801 );
xor ( n328686 , n328684 , n328685 );
buf ( n328687 , n36397 );
xor ( n38262 , n328686 , n328687 );
buf ( n328689 , n38262 );
buf ( n328690 , n328689 );
buf ( n328691 , n36401 );
buf ( n328692 , n322571 );
buf ( n38267 , n322625 );
xor ( n38268 , n328692 , n38267 );
buf ( n328695 , n36339 );
and ( n38270 , n38268 , n328695 );
and ( n38271 , n328692 , n38267 );
or ( n38272 , n38270 , n38271 );
buf ( n38273 , n38272 );
buf ( n328700 , n38273 );
xor ( n38275 , n328690 , n328691 );
xor ( n328702 , n38275 , n328700 );
buf ( n328703 , n328702 );
xor ( n328704 , n328690 , n328691 );
and ( n38279 , n328704 , n328700 );
and ( n328706 , n328690 , n328691 );
or ( n328707 , n38279 , n328706 );
buf ( n328708 , n328707 );
buf ( n38283 , n324267 );
buf ( n38284 , n38283 );
buf ( n328711 , n314320 );
buf ( n328712 , n315709 );
xor ( n328713 , n328711 , n328712 );
buf ( n328714 , n17602 );
xor ( n38289 , n328713 , n328714 );
buf ( n328716 , n38289 );
buf ( n328717 , n328716 );
buf ( n328718 , n314315 );
buf ( n328719 , n314380 );
xor ( n38294 , n328718 , n328719 );
buf ( n328721 , n302980 );
and ( n328722 , n38294 , n328721 );
and ( n328723 , n328718 , n328719 );
or ( n38298 , n328722 , n328723 );
buf ( n328725 , n38298 );
buf ( n328726 , n328725 );
xor ( n38301 , n38284 , n328717 );
xor ( n328728 , n38301 , n328726 );
buf ( n328729 , n328728 );
xor ( n38304 , n38284 , n328717 );
and ( n328731 , n38304 , n328726 );
and ( n328732 , n38284 , n328717 );
or ( n38307 , n328731 , n328732 );
buf ( n328734 , n38307 );
not ( n38309 , n33487 );
buf ( n328736 , n38309 );
buf ( n328737 , n315690 );
buf ( n328738 , n317414 );
xor ( n328739 , n328737 , n328738 );
buf ( n328740 , n323833 );
buf ( n328741 , n328740 );
xor ( n328742 , n328739 , n328741 );
buf ( n328743 , n328742 );
buf ( n328744 , n328743 );
buf ( n328745 , n318935 );
buf ( n328746 , n315685 );
xor ( n328747 , n328745 , n328746 );
buf ( n328748 , n296411 );
and ( n38323 , n328747 , n328748 );
and ( n328750 , n328745 , n328746 );
or ( n328751 , n38323 , n328750 );
buf ( n328752 , n328751 );
buf ( n328753 , n328752 );
xor ( n38328 , n328736 , n328744 );
xor ( n328755 , n38328 , n328753 );
buf ( n328756 , n328755 );
xor ( n328757 , n328736 , n328744 );
and ( n328758 , n328757 , n328753 );
and ( n38333 , n328736 , n328744 );
or ( n328760 , n328758 , n38333 );
buf ( n328761 , n328760 );
buf ( n328762 , n307968 );
buf ( n328763 , n328762 );
buf ( n328764 , n314375 );
buf ( n328765 , n314358 );
xor ( n328766 , n328764 , n328765 );
buf ( n328767 , n12699 );
and ( n328768 , n328766 , n328767 );
and ( n328769 , n328764 , n328765 );
or ( n328770 , n328768 , n328769 );
buf ( n328771 , n328770 );
buf ( n328772 , n328771 );
xor ( n328773 , n328718 , n328719 );
xor ( n328774 , n328773 , n328721 );
buf ( n328775 , n328774 );
buf ( n328776 , n328775 );
xor ( n328777 , n328763 , n328772 );
xor ( n38352 , n328777 , n328776 );
buf ( n328779 , n38352 );
xor ( n328780 , n328763 , n328772 );
and ( n328781 , n328780 , n328776 );
and ( n38356 , n328763 , n328772 );
or ( n328783 , n328781 , n38356 );
buf ( n328784 , n328783 );
not ( n38359 , n33387 );
buf ( n328786 , n38359 );
xor ( n328787 , n328745 , n328746 );
xor ( n38362 , n328787 , n328748 );
buf ( n38363 , n38362 );
buf ( n38364 , n38363 );
buf ( n328791 , n318983 );
buf ( n328792 , n318930 );
xor ( n328793 , n328791 , n328792 );
buf ( n328794 , n3172 );
and ( n328795 , n328793 , n328794 );
and ( n328796 , n328791 , n328792 );
or ( n38371 , n328795 , n328796 );
buf ( n328798 , n38371 );
buf ( n328799 , n328798 );
xor ( n328800 , n328786 , n38364 );
xor ( n328801 , n328800 , n328799 );
buf ( n328802 , n328801 );
xor ( n328803 , n328786 , n38364 );
and ( n328804 , n328803 , n328799 );
and ( n38379 , n328786 , n38364 );
or ( n328806 , n328804 , n38379 );
buf ( n328807 , n328806 );
buf ( n38382 , n33334 );
not ( n38383 , n38382 );
buf ( n38384 , n38383 );
buf ( n328811 , n318978 );
buf ( n328812 , n319210 );
xor ( n328813 , n328811 , n328812 );
buf ( n328814 , n323678 );
buf ( n328815 , n328814 );
and ( n328816 , n328813 , n328815 );
and ( n38391 , n328811 , n328812 );
or ( n328818 , n328816 , n38391 );
buf ( n328819 , n328818 );
buf ( n328820 , n328819 );
xor ( n328821 , n328791 , n328792 );
xor ( n328822 , n328821 , n328794 );
buf ( n328823 , n328822 );
buf ( n328824 , n328823 );
xor ( n38399 , n38384 , n328820 );
xor ( n328826 , n38399 , n328824 );
buf ( n328827 , n328826 );
xor ( n38402 , n38384 , n328820 );
and ( n328829 , n38402 , n328824 );
and ( n38404 , n38384 , n328820 );
or ( n328831 , n328829 , n38404 );
buf ( n328832 , n328831 );
buf ( n328833 , n312280 );
buf ( n328834 , n314353 );
xor ( n328835 , n328833 , n328834 );
buf ( n328836 , n34491 );
and ( n328837 , n328835 , n328836 );
and ( n328838 , n328833 , n328834 );
or ( n38413 , n328837 , n328838 );
buf ( n328840 , n38413 );
buf ( n38415 , n328840 );
xor ( n38416 , n328764 , n328765 );
xor ( n328843 , n38416 , n328767 );
buf ( n328844 , n328843 );
buf ( n328845 , n328844 );
buf ( n38420 , n324173 );
not ( n328847 , n38420 );
not ( n38422 , n328847 );
buf ( n328849 , n38422 );
xor ( n38424 , n38415 , n328845 );
xor ( n38425 , n38424 , n328849 );
buf ( n328852 , n38425 );
xor ( n328853 , n38415 , n328845 );
and ( n38428 , n328853 , n328849 );
and ( n328855 , n38415 , n328845 );
or ( n328856 , n38428 , n328855 );
buf ( n328857 , n328856 );
buf ( n328858 , n33309 );
buf ( n328859 , n328858 );
buf ( n328860 , n320132 );
buf ( n38435 , n319506 );
xor ( n38436 , n328860 , n38435 );
buf ( n328863 , n33283 );
buf ( n328864 , n328863 );
and ( n38439 , n38436 , n328864 );
and ( n328866 , n328860 , n38435 );
or ( n328867 , n38439 , n328866 );
buf ( n328868 , n328867 );
buf ( n328869 , n328868 );
buf ( n328870 , n319511 );
buf ( n328871 , n319205 );
xor ( n38446 , n328870 , n328871 );
buf ( n328873 , n298380 );
xor ( n328874 , n38446 , n328873 );
buf ( n328875 , n328874 );
buf ( n328876 , n328875 );
xor ( n38451 , n328859 , n328869 );
xor ( n38452 , n38451 , n328876 );
buf ( n328879 , n38452 );
xor ( n328880 , n328859 , n328869 );
and ( n328881 , n328880 , n328876 );
and ( n38456 , n328859 , n328869 );
or ( n328883 , n328881 , n38456 );
buf ( n328884 , n328883 );
buf ( n328885 , n324522 );
xor ( n38460 , n328516 , n328517 );
xor ( n328887 , n38460 , n328519 );
buf ( n328888 , n328887 );
buf ( n328889 , n328888 );
buf ( n328890 , n322018 );
buf ( n328891 , n321876 );
xor ( n38466 , n328890 , n328891 );
buf ( n328893 , n34015 );
and ( n38468 , n38466 , n328893 );
and ( n328895 , n328890 , n328891 );
or ( n328896 , n38468 , n328895 );
buf ( n328897 , n328896 );
buf ( n328898 , n328897 );
xor ( n38473 , n328885 , n328889 );
xor ( n328900 , n38473 , n328898 );
buf ( n328901 , n328900 );
xor ( n38476 , n328885 , n328889 );
and ( n328903 , n38476 , n328898 );
and ( n328904 , n328885 , n328889 );
or ( n38479 , n328903 , n328904 );
buf ( n328906 , n38479 );
buf ( n38481 , n33311 );
xor ( n328908 , n328860 , n38435 );
xor ( n328909 , n328908 , n328864 );
buf ( n328910 , n328909 );
buf ( n328911 , n328910 );
xor ( n328912 , n320127 , n320330 );
and ( n38487 , n328912 , n33180 );
and ( n328914 , n320127 , n320330 );
or ( n38489 , n38487 , n328914 );
buf ( n328916 , n38489 );
xor ( n328917 , n38481 , n328911 );
xor ( n38492 , n328917 , n328916 );
buf ( n328919 , n38492 );
xor ( n38494 , n38481 , n328911 );
and ( n38495 , n38494 , n328916 );
and ( n38496 , n38481 , n328911 );
or ( n38497 , n38495 , n38496 );
buf ( n328924 , n38497 );
buf ( n328925 , n34010 );
xor ( n38500 , n328890 , n328891 );
xor ( n328927 , n38500 , n328893 );
buf ( n328928 , n328927 );
buf ( n328929 , n328928 );
xor ( n328930 , n328588 , n328589 );
and ( n328931 , n328930 , n328591 );
and ( n328932 , n328588 , n328589 );
or ( n38507 , n328931 , n328932 );
buf ( n328934 , n38507 );
buf ( n328935 , n328934 );
xor ( n38510 , n328925 , n328929 );
xor ( n328937 , n38510 , n328935 );
buf ( n328938 , n328937 );
xor ( n328939 , n328925 , n328929 );
and ( n328940 , n328939 , n328935 );
and ( n328941 , n328925 , n328929 );
or ( n38516 , n328940 , n328941 );
buf ( n328943 , n38516 );
buf ( n328944 , n323489 );
xor ( n38519 , n325728 , n292343 );
and ( n38520 , n38519 , n325731 );
and ( n328947 , n325728 , n292343 );
or ( n328948 , n38520 , n328947 );
buf ( n328949 , n328948 );
buf ( n328950 , n325765 );
buf ( n328951 , n320953 );
xor ( n328952 , n328950 , n328951 );
buf ( n328953 , n323481 );
xor ( n328954 , n328952 , n328953 );
buf ( n328955 , n328954 );
buf ( n328956 , n328955 );
xor ( n328957 , n328944 , n328949 );
xor ( n328958 , n328957 , n328956 );
buf ( n328959 , n328958 );
xor ( n38534 , n328944 , n328949 );
and ( n328961 , n38534 , n328956 );
and ( n328962 , n328944 , n328949 );
or ( n38537 , n328961 , n328962 );
buf ( n328964 , n38537 );
not ( n328965 , n33015 );
buf ( n328966 , n328965 );
buf ( n328967 , n321333 );
buf ( n328968 , n321639 );
xor ( n328969 , n328967 , n328968 );
buf ( n328970 , n309969 );
and ( n38545 , n328969 , n328970 );
and ( n328972 , n328967 , n328968 );
or ( n328973 , n38545 , n328972 );
buf ( n328974 , n328973 );
buf ( n328975 , n328974 );
buf ( n328976 , n321338 );
buf ( n328977 , n33163 );
xor ( n38552 , n328976 , n328977 );
buf ( n328979 , n33012 );
xor ( n328980 , n38552 , n328979 );
buf ( n328981 , n328980 );
buf ( n328982 , n328981 );
xor ( n328983 , n328966 , n328975 );
xor ( n328984 , n328983 , n328982 );
buf ( n328985 , n328984 );
xor ( n328986 , n328966 , n328975 );
and ( n38561 , n328986 , n328982 );
and ( n328988 , n328966 , n328975 );
or ( n328989 , n38561 , n328988 );
buf ( n328990 , n328989 );
not ( n328991 , n32984 );
buf ( n328992 , n328991 );
xor ( n38567 , n328967 , n328968 );
xor ( n328994 , n38567 , n328970 );
buf ( n328995 , n328994 );
buf ( n328996 , n328995 );
buf ( n328997 , n321634 );
buf ( n328998 , n321573 );
xor ( n328999 , n328997 , n328998 );
buf ( n329000 , n323377 );
and ( n329001 , n328999 , n329000 );
and ( n38576 , n328997 , n328998 );
or ( n329003 , n329001 , n38576 );
buf ( n329004 , n329003 );
buf ( n329005 , n329004 );
xor ( n38580 , n328992 , n328996 );
xor ( n329007 , n38580 , n329005 );
buf ( n329008 , n329007 );
xor ( n38583 , n328992 , n328996 );
and ( n329010 , n38583 , n329005 );
and ( n329011 , n328992 , n328996 );
or ( n38586 , n329010 , n329011 );
buf ( n329013 , n38586 );
buf ( n329014 , n33616 );
buf ( n329015 , n319905 );
buf ( n329016 , n324690 );
xor ( n329017 , n329015 , n329016 );
buf ( n329018 , n309986 );
xor ( n329019 , n329017 , n329018 );
buf ( n329020 , n329019 );
buf ( n329021 , n329020 );
buf ( n329022 , n324785 );
buf ( n329023 , n318489 );
xor ( n329024 , n329022 , n329023 );
buf ( n329025 , n11959 );
and ( n38600 , n329024 , n329025 );
and ( n329027 , n329022 , n329023 );
or ( n329028 , n38600 , n329027 );
buf ( n329029 , n329028 );
buf ( n329030 , n329029 );
xor ( n329031 , n329014 , n329021 );
xor ( n329032 , n329031 , n329030 );
buf ( n329033 , n329032 );
xor ( n329034 , n329014 , n329021 );
and ( n329035 , n329034 , n329030 );
and ( n38610 , n329014 , n329021 );
or ( n329037 , n329035 , n38610 );
buf ( n329038 , n329037 );
not ( n329039 , n323373 );
buf ( n329040 , n329039 );
buf ( n329041 , n4640 );
buf ( n329042 , n322117 );
xor ( n329043 , n329041 , n329042 );
buf ( n329044 , n321568 );
and ( n329045 , n329043 , n329044 );
and ( n329046 , n329041 , n329042 );
or ( n38621 , n329045 , n329046 );
buf ( n329048 , n38621 );
buf ( n329049 , n329048 );
xor ( n329050 , n328997 , n328998 );
xor ( n38625 , n329050 , n329000 );
buf ( n329052 , n38625 );
buf ( n329053 , n329052 );
xor ( n38628 , n329040 , n329049 );
xor ( n329055 , n38628 , n329053 );
buf ( n329056 , n329055 );
xor ( n38631 , n329040 , n329049 );
and ( n38632 , n38631 , n329053 );
and ( n329059 , n329040 , n329049 );
or ( n329060 , n38632 , n329059 );
buf ( n329061 , n329060 );
buf ( n329062 , n32912 );
buf ( n329063 , n322456 );
buf ( n329064 , n4721 );
xor ( n329065 , n329063 , n329064 );
buf ( n329066 , n322112 );
and ( n38641 , n329065 , n329066 );
and ( n329068 , n329063 , n329064 );
or ( n329069 , n38641 , n329068 );
buf ( n329070 , n329069 );
buf ( n329071 , n329070 );
xor ( n329072 , n329041 , n329042 );
xor ( n38647 , n329072 , n329044 );
buf ( n329074 , n38647 );
buf ( n329075 , n329074 );
xor ( n38650 , n329062 , n329071 );
xor ( n329077 , n38650 , n329075 );
buf ( n329078 , n329077 );
xor ( n38653 , n329062 , n329071 );
and ( n38654 , n38653 , n329075 );
and ( n329081 , n329062 , n329071 );
or ( n329082 , n38654 , n329081 );
buf ( n329083 , n329082 );
buf ( n329084 , n324192 );
buf ( n329085 , n329084 );
xor ( n38660 , n325356 , n325345 );
buf ( n329087 , n33658 );
not ( n329088 , n329087 );
xor ( n38663 , n38660 , n329088 );
buf ( n329090 , n38663 );
buf ( n329091 , n16254 );
buf ( n329092 , n329091 );
buf ( n329093 , n325391 );
xor ( n329094 , n329092 , n329093 );
buf ( n329095 , n325394 );
and ( n38670 , n329094 , n329095 );
and ( n329097 , n329092 , n329093 );
or ( n329098 , n38670 , n329097 );
buf ( n329099 , n329098 );
buf ( n329100 , n329099 );
xor ( n329101 , n329085 , n329090 );
xor ( n329102 , n329101 , n329100 );
buf ( n329103 , n329102 );
xor ( n329104 , n329085 , n329090 );
and ( n38679 , n329104 , n329100 );
and ( n38680 , n329085 , n329090 );
or ( n329107 , n38679 , n38680 );
buf ( n329108 , n329107 );
not ( n329109 , n32877 );
buf ( n329110 , n329109 );
xor ( n329111 , n329063 , n329064 );
xor ( n329112 , n329111 , n329066 );
buf ( n329113 , n329112 );
buf ( n329114 , n329113 );
buf ( n329115 , n322451 );
buf ( n329116 , n33001 );
xor ( n329117 , n329115 , n329116 );
buf ( n329118 , n32858 );
and ( n329119 , n329117 , n329118 );
and ( n38694 , n329115 , n329116 );
or ( n38695 , n329119 , n38694 );
buf ( n329122 , n38695 );
buf ( n329123 , n329122 );
xor ( n329124 , n329110 , n329114 );
xor ( n38699 , n329124 , n329123 );
buf ( n329126 , n38699 );
xor ( n329127 , n329110 , n329114 );
and ( n38702 , n329127 , n329123 );
and ( n329129 , n329110 , n329114 );
or ( n329130 , n38702 , n329129 );
buf ( n329131 , n329130 );
buf ( n38706 , n323280 );
buf ( n329133 , n38706 );
xor ( n329134 , n323395 , n323217 );
and ( n329135 , n329134 , n32972 );
and ( n38710 , n323395 , n323217 );
or ( n38711 , n329135 , n38710 );
buf ( n329138 , n38711 );
xor ( n329139 , n329115 , n329116 );
xor ( n329140 , n329139 , n329118 );
buf ( n329141 , n329140 );
buf ( n329142 , n329141 );
xor ( n38717 , n329133 , n329138 );
xor ( n329144 , n38717 , n329142 );
buf ( n329145 , n329144 );
xor ( n38720 , n329133 , n329138 );
and ( n329147 , n38720 , n329142 );
and ( n329148 , n329133 , n329138 );
or ( n329149 , n329147 , n329148 );
buf ( n329150 , n329149 );
buf ( n329151 , n33622 );
buf ( n329152 , n7448 );
buf ( n329153 , n317637 );
xor ( n329154 , n329152 , n329153 );
buf ( n329155 , n318484 );
and ( n38730 , n329154 , n329155 );
and ( n329157 , n329152 , n329153 );
or ( n329158 , n38730 , n329157 );
buf ( n329159 , n329158 );
buf ( n329160 , n329159 );
xor ( n329161 , n329022 , n329023 );
xor ( n329162 , n329161 , n329025 );
buf ( n329163 , n329162 );
buf ( n329164 , n329163 );
xor ( n38739 , n329151 , n329160 );
xor ( n38740 , n38739 , n329164 );
buf ( n329167 , n38740 );
xor ( n329168 , n329151 , n329160 );
and ( n329169 , n329168 , n329164 );
and ( n38744 , n329151 , n329160 );
or ( n329171 , n329169 , n38744 );
buf ( n329172 , n329171 );
buf ( n38747 , n323059 );
buf ( n329174 , n38747 );
buf ( n329175 , n323066 );
buf ( n329176 , n323325 );
xor ( n329177 , n329175 , n329176 );
buf ( n329178 , n322770 );
and ( n38753 , n329177 , n329178 );
and ( n329180 , n329175 , n329176 );
or ( n329181 , n38753 , n329180 );
buf ( n329182 , n329181 );
buf ( n329183 , n329182 );
buf ( n329184 , n323053 );
buf ( n329185 , n322775 );
xor ( n329186 , n329184 , n329185 );
buf ( n329187 , n323357 );
xor ( n38762 , n329186 , n329187 );
buf ( n329189 , n38762 );
buf ( n329190 , n329189 );
xor ( n38765 , n329174 , n329183 );
xor ( n329192 , n38765 , n329190 );
buf ( n329193 , n329192 );
xor ( n329194 , n329174 , n329183 );
and ( n38769 , n329194 , n329190 );
and ( n329196 , n329174 , n329183 );
or ( n329197 , n38769 , n329196 );
buf ( n329198 , n329197 );
buf ( n38773 , n16425 );
buf ( n329200 , n325460 );
buf ( n329201 , n325456 );
xor ( n329202 , n329200 , n329201 );
buf ( n38777 , n306852 );
buf ( n329204 , n38777 );
xor ( n329205 , n329202 , n329204 );
buf ( n329206 , n329205 );
buf ( n329207 , n329206 );
buf ( n329208 , n325596 );
buf ( n329209 , n325591 );
xor ( n329210 , n329208 , n329209 );
buf ( n329211 , n16421 );
and ( n329212 , n329210 , n329211 );
and ( n38787 , n329208 , n329209 );
or ( n329214 , n329212 , n38787 );
buf ( n329215 , n329214 );
buf ( n329216 , n329215 );
xor ( n38791 , n38773 , n329207 );
xor ( n329218 , n38791 , n329216 );
buf ( n329219 , n329218 );
xor ( n38794 , n38773 , n329207 );
and ( n38795 , n38794 , n329216 );
and ( n38796 , n38773 , n329207 );
or ( n38797 , n38795 , n38796 );
buf ( n329224 , n38797 );
buf ( n329225 , n323181 );
xor ( n329226 , n32834 , n323272 );
and ( n38801 , n329226 , n32738 );
and ( n38802 , n32834 , n323272 );
or ( n38803 , n38801 , n38802 );
buf ( n329230 , n38803 );
xor ( n329231 , n329175 , n329176 );
xor ( n38806 , n329231 , n329178 );
buf ( n38807 , n38806 );
buf ( n329234 , n38807 );
xor ( n38809 , n329225 , n329230 );
xor ( n38810 , n38809 , n329234 );
buf ( n329237 , n38810 );
xor ( n38812 , n329225 , n329230 );
and ( n329239 , n38812 , n329234 );
and ( n329240 , n329225 , n329230 );
or ( n38815 , n329239 , n329240 );
buf ( n329242 , n38815 );
buf ( n329243 , n32750 );
buf ( n329244 , n329243 );
xor ( n38819 , n328623 , n328624 );
and ( n38820 , n38819 , n328626 );
and ( n38821 , n328623 , n328624 );
or ( n38822 , n38820 , n38821 );
buf ( n329249 , n38822 );
buf ( n329250 , n329249 );
xor ( n329251 , n32834 , n323272 );
xor ( n38826 , n329251 , n32738 );
buf ( n329253 , n38826 );
xor ( n38828 , n329244 , n329250 );
xor ( n329255 , n38828 , n329253 );
buf ( n329256 , n329255 );
xor ( n38831 , n329244 , n329250 );
and ( n329258 , n38831 , n329253 );
and ( n329259 , n329244 , n329250 );
or ( n38834 , n329258 , n329259 );
buf ( n329261 , n38834 );
buf ( n329262 , n36335 );
xor ( n329263 , n328692 , n38267 );
xor ( n38838 , n329263 , n328695 );
buf ( n329265 , n38838 );
buf ( n329266 , n329265 );
xor ( n38841 , n328509 , n328510 );
and ( n329268 , n38841 , n328512 );
and ( n329269 , n328509 , n328510 );
or ( n38844 , n329268 , n329269 );
buf ( n329271 , n38844 );
buf ( n329272 , n329271 );
xor ( n38847 , n329262 , n329266 );
xor ( n329274 , n38847 , n329272 );
buf ( n329275 , n329274 );
xor ( n38850 , n329262 , n329266 );
and ( n329277 , n38850 , n329272 );
and ( n329278 , n329262 , n329266 );
or ( n38853 , n329277 , n329278 );
buf ( n329280 , n38853 );
buf ( n329281 , n33870 );
xor ( n38856 , n324020 , n317632 );
and ( n329283 , n38856 , n317397 );
and ( n329284 , n324020 , n317632 );
or ( n38859 , n329283 , n329284 );
buf ( n329286 , n38859 );
xor ( n329287 , n329152 , n329153 );
xor ( n38862 , n329287 , n329155 );
buf ( n329289 , n38862 );
buf ( n329290 , n329289 );
xor ( n329291 , n329281 , n329286 );
xor ( n329292 , n329291 , n329290 );
buf ( n329293 , n329292 );
xor ( n38868 , n329281 , n329286 );
and ( n38869 , n38868 , n329290 );
and ( n38870 , n329281 , n329286 );
or ( n329297 , n38869 , n38870 );
buf ( n329298 , n329297 );
not ( n38873 , n324001 );
buf ( n329300 , n38873 );
xor ( n329301 , n329208 , n329209 );
xor ( n38876 , n329301 , n329211 );
buf ( n329303 , n38876 );
buf ( n38878 , n329303 );
buf ( n329305 , n325494 );
buf ( n329306 , n35063 );
xor ( n329307 , n329305 , n329306 );
buf ( n329308 , n33552 );
and ( n329309 , n329307 , n329308 );
and ( n329310 , n329305 , n329306 );
or ( n38885 , n329309 , n329310 );
buf ( n329312 , n38885 );
buf ( n329313 , n329312 );
xor ( n38888 , n329300 , n38878 );
xor ( n329315 , n38888 , n329313 );
buf ( n329316 , n329315 );
xor ( n38891 , n329300 , n38878 );
and ( n329318 , n38891 , n329313 );
and ( n329319 , n329300 , n38878 );
or ( n329320 , n329318 , n329319 );
buf ( n329321 , n329320 );
buf ( n329322 , n323118 );
buf ( n329323 , n322997 );
and ( n329324 , n329322 , n329323 );
buf ( n329325 , n329324 );
buf ( n329326 , n329325 );
nand ( n329327 , n323098 , n32670 );
buf ( n329328 , n329327 );
xor ( n329329 , n328612 , n328613 );
xor ( n329330 , n329329 , n328615 );
buf ( n329331 , n329330 );
buf ( n329332 , n329331 );
xor ( n329333 , n329326 , n329328 );
xor ( n38908 , n329333 , n329332 );
buf ( n329335 , n38908 );
xor ( n38910 , n329326 , n329328 );
and ( n38911 , n38910 , n329332 );
and ( n329338 , n329326 , n329328 );
or ( n38913 , n38911 , n329338 );
buf ( n329340 , n38913 );
buf ( n329341 , n310029 );
not ( n38916 , n329341 );
buf ( n329343 , n322883 );
not ( n329344 , n329343 );
and ( n38919 , n38916 , n329344 );
buf ( n329346 , n310029 );
buf ( n329347 , n322883 );
and ( n329348 , n329346 , n329347 );
nor ( n329349 , n38919 , n329348 );
buf ( n329350 , n329349 );
buf ( n329351 , n329350 );
xor ( n329352 , n322806 , n322878 );
and ( n38927 , n329352 , n326869 );
and ( n329354 , n322806 , n322878 );
or ( n38929 , n38927 , n329354 );
xnor ( n38930 , n38929 , n310326 );
buf ( n329357 , n38930 );
buf ( n329358 , n38930 );
buf ( n329359 , n329350 );
not ( n329360 , n329351 );
not ( n329361 , n329357 );
or ( n329362 , n329360 , n329361 );
or ( n38937 , n329358 , n329359 );
nand ( n329364 , n329362 , n38937 );
buf ( n329365 , n329364 );
buf ( n329366 , n32707 );
buf ( n329367 , n323020 );
buf ( n329368 , n322984 );
xor ( n38943 , n329366 , n329367 );
xor ( n329370 , n38943 , n329368 );
buf ( n329371 , n329370 );
xor ( n38946 , n329366 , n329367 );
and ( n329373 , n38946 , n329368 );
and ( n329374 , n329366 , n329367 );
or ( n38949 , n329373 , n329374 );
buf ( n329376 , n38949 );
buf ( n329377 , n315295 );
buf ( n329378 , n317392 );
buf ( n329379 , n324257 );
buf ( n329380 , n329379 );
xor ( n38955 , n329377 , n329378 );
xor ( n329382 , n38955 , n329380 );
buf ( n329383 , n329382 );
xor ( n329384 , n329377 , n329378 );
and ( n38959 , n329384 , n329380 );
and ( n329386 , n329377 , n329378 );
or ( n329387 , n38959 , n329386 );
buf ( n329388 , n329387 );
xor ( n329389 , n328663 , n328664 );
and ( n329390 , n329389 , n328666 );
and ( n38965 , n328663 , n328664 );
or ( n329392 , n329390 , n38965 );
buf ( n329393 , n329392 );
xor ( n329394 , n328811 , n328812 );
xor ( n38969 , n329394 , n328815 );
buf ( n329396 , n38969 );
xor ( n329397 , n328833 , n328834 );
xor ( n38972 , n329397 , n328836 );
buf ( n329399 , n38972 );
xor ( n38974 , n329015 , n329016 );
and ( n38975 , n38974 , n329018 );
and ( n38976 , n329015 , n329016 );
or ( n38977 , n38975 , n38976 );
buf ( n329404 , n38977 );
xor ( n38979 , n328950 , n328951 );
and ( n38980 , n38979 , n328953 );
and ( n38981 , n328950 , n328951 );
or ( n329408 , n38980 , n38981 );
buf ( n329409 , n329408 );
buf ( n329410 , n317419 );
buf ( n329411 , n314809 );
buf ( n329412 , n294736 );
xor ( n329413 , n329410 , n329411 );
xor ( n38988 , n329413 , n329412 );
buf ( n329415 , n38988 );
xor ( n38990 , n329410 , n329411 );
and ( n329417 , n38990 , n329412 );
and ( n329418 , n329410 , n329411 );
or ( n38993 , n329417 , n329418 );
buf ( n329420 , n38993 );
xor ( n38995 , n329200 , n329201 );
and ( n329422 , n38995 , n329204 );
and ( n329423 , n329200 , n329201 );
or ( n38998 , n329422 , n329423 );
buf ( n329425 , n38998 );
xor ( n329426 , n329184 , n329185 );
and ( n39001 , n329426 , n329187 );
and ( n329428 , n329184 , n329185 );
or ( n39003 , n39001 , n329428 );
buf ( n329430 , n39003 );
buf ( n329431 , n315290 );
buf ( n329432 , n315714 );
buf ( n329433 , n11750 );
xor ( n39008 , n329431 , n329432 );
xor ( n329435 , n39008 , n329433 );
buf ( n329436 , n329435 );
xor ( n329437 , n329431 , n329432 );
and ( n329438 , n329437 , n329433 );
and ( n329439 , n329431 , n329432 );
or ( n39014 , n329438 , n329439 );
buf ( n329441 , n39014 );
buf ( n329442 , n325524 );
buf ( n329443 , n325532 );
buf ( n329444 , n16359 );
buf ( n329445 , n329444 );
xor ( n329446 , n329442 , n329443 );
xor ( n329447 , n329446 , n329445 );
buf ( n329448 , n329447 );
xor ( n329449 , n329442 , n329443 );
and ( n39024 , n329449 , n329445 );
and ( n329451 , n329442 , n329443 );
or ( n329452 , n39024 , n329451 );
buf ( n329453 , n329452 );
xor ( n39028 , n328645 , n328646 );
and ( n329455 , n39028 , n328649 );
and ( n329456 , n328645 , n328646 );
or ( n39031 , n329455 , n329456 );
buf ( n329458 , n39031 );
xor ( n39033 , n328684 , n328685 );
and ( n39034 , n39033 , n328687 );
and ( n329461 , n328684 , n328685 );
or ( n39036 , n39034 , n329461 );
buf ( n329463 , n39036 );
xor ( n39038 , n328535 , n328536 );
xor ( n39039 , n39038 , n328538 );
buf ( n329466 , n39039 );
xor ( n39041 , n328870 , n328871 );
and ( n329468 , n39041 , n328873 );
and ( n329469 , n328870 , n328871 );
or ( n39044 , n329468 , n329469 );
buf ( n329471 , n39044 );
xor ( n329472 , n328561 , n328562 );
xor ( n39047 , n329472 , n328564 );
buf ( n329474 , n39047 );
xor ( n39049 , n328737 , n328738 );
and ( n39050 , n39049 , n328741 );
and ( n39051 , n328737 , n328738 );
or ( n39052 , n39050 , n39051 );
buf ( n329479 , n39052 );
xor ( n39054 , n328711 , n328712 );
and ( n39055 , n39054 , n328714 );
and ( n39056 , n328711 , n328712 );
or ( n329483 , n39055 , n39056 );
buf ( n329484 , n329483 );
xor ( n329485 , n329305 , n329306 );
xor ( n329486 , n329485 , n329308 );
buf ( n329487 , n329486 );
xor ( n329488 , n328595 , n328596 );
xor ( n329489 , n329488 , n328598 );
buf ( n329490 , n329489 );
xor ( n329491 , n328976 , n328977 );
and ( n329492 , n329491 , n328979 );
and ( n39067 , n328976 , n328977 );
or ( n329494 , n329492 , n39067 );
buf ( n329495 , n329494 );
xor ( n329496 , n38144 , n328571 );
and ( n39071 , n329496 , n328574 );
and ( n329498 , n38144 , n328571 );
or ( n39073 , n39071 , n329498 );
buf ( n329500 , n39073 );
buf ( n329501 , n329038 );
not ( n329502 , n831 );
not ( n39077 , n308638 );
or ( n329504 , n329502 , n39077 );
nand ( n39079 , n329504 , n33895 );
buf ( n329506 , n39079 );
buf ( n329507 , n329404 );
xor ( n39082 , n329506 , n329507 );
buf ( n329509 , n319910 );
buf ( n329510 , n320660 );
xor ( n39085 , n329509 , n329510 );
buf ( n329512 , n33887 );
buf ( n329513 , n329512 );
xor ( n329514 , n39085 , n329513 );
buf ( n329515 , n329514 );
buf ( n329516 , n329515 );
xor ( n329517 , n39082 , n329516 );
buf ( n329518 , n329517 );
buf ( n329519 , n329518 );
and ( n39094 , n329501 , n329519 );
buf ( n329521 , n39094 );
buf ( n329522 , n329521 );
not ( n39097 , n329522 );
buf ( n329524 , n329518 );
buf ( n329525 , n329038 );
or ( n39100 , n329524 , n329525 );
buf ( n329527 , n39100 );
buf ( n329528 , n329527 );
nand ( n39103 , n39097 , n329528 );
buf ( n329530 , n39103 );
buf ( n39105 , n329530 );
buf ( n329532 , n329530 );
not ( n329533 , n329532 );
buf ( n329534 , n329533 );
buf ( n39109 , n329534 );
buf ( n39110 , n33601 );
not ( n329537 , n39110 );
xor ( n329538 , n329537 , n329388 );
xor ( n39113 , n324020 , n317632 );
xor ( n329540 , n39113 , n317397 );
and ( n39115 , n329538 , n329540 );
and ( n329542 , n329537 , n329388 );
or ( n329543 , n39115 , n329542 );
buf ( n329544 , n329543 );
buf ( n329545 , n329293 );
nor ( n329546 , n329544 , n329545 );
buf ( n329547 , n329546 );
buf ( n329548 , n329547 );
not ( n39123 , n329548 );
buf ( n329550 , n324163 );
buf ( n329551 , n329550 );
buf ( n329552 , n329383 );
xor ( n329553 , n329551 , n329552 );
buf ( n329554 , n329441 );
and ( n39129 , n329553 , n329554 );
and ( n329556 , n329551 , n329552 );
or ( n329557 , n39129 , n329556 );
buf ( n329558 , n329557 );
buf ( n329559 , n329558 );
xor ( n39134 , n329537 , n329388 );
xor ( n329561 , n39134 , n329540 );
buf ( n329562 , n329561 );
or ( n39137 , n329559 , n329562 );
buf ( n39138 , n39137 );
buf ( n329565 , n39138 );
nand ( n39140 , n39123 , n329565 );
buf ( n39141 , n39140 );
buf ( n329568 , n39141 );
buf ( n329569 , n329033 );
buf ( n329570 , n329172 );
or ( n329571 , n329569 , n329570 );
buf ( n329572 , n329571 );
buf ( n329573 , n329572 );
buf ( n329574 , n329167 );
buf ( n329575 , n329298 );
or ( n39150 , n329574 , n329575 );
buf ( n39151 , n39150 );
buf ( n329578 , n39151 );
nand ( n39153 , n329573 , n329578 );
buf ( n329580 , n39153 );
buf ( n329581 , n329580 );
nor ( n39156 , n329568 , n329581 );
buf ( n329583 , n39156 );
buf ( n329584 , n329583 );
not ( n329585 , n329584 );
not ( n39160 , n33631 );
not ( n329587 , n39160 );
xor ( n329588 , n10429 , n325313 );
and ( n329589 , n329588 , n34863 );
and ( n329590 , n10429 , n325313 );
or ( n39165 , n329589 , n329590 );
xor ( n329592 , n329587 , n39165 );
buf ( n329593 , n324979 );
buf ( n39168 , n33636 );
buf ( n329595 , n39168 );
xor ( n329596 , n329593 , n329595 );
buf ( n329597 , n34594 );
xor ( n329598 , n329596 , n329597 );
buf ( n329599 , n329598 );
xnor ( n329600 , n329592 , n329599 );
buf ( n329601 , n329600 );
xor ( n39176 , n10429 , n325313 );
xor ( n329603 , n39176 , n34863 );
xor ( n329604 , n325356 , n325345 );
and ( n39179 , n329604 , n329088 );
and ( n329606 , n325356 , n325345 );
or ( n39181 , n39179 , n329606 );
nor ( n329608 , n329603 , n39181 );
buf ( n329609 , n307616 );
buf ( n39184 , n329609 );
not ( n329611 , n39184 );
or ( n329612 , n329608 , n329611 );
nand ( n39187 , n329603 , n39181 );
nand ( n329614 , n329612 , n39187 );
buf ( n329615 , n329614 );
nor ( n39190 , n329601 , n329615 );
buf ( n329617 , n39190 );
buf ( n39192 , n329617 );
not ( n39193 , n39192 );
buf ( n329620 , n39193 );
buf ( n329621 , n329620 );
not ( n39196 , n329621 );
buf ( n39197 , n39196 );
buf ( n329624 , n39197 );
buf ( n329625 , n329108 );
xor ( n329626 , n329611 , n39181 );
xnor ( n329627 , n329626 , n329603 );
buf ( n329628 , n329627 );
nor ( n329629 , n329625 , n329628 );
buf ( n329630 , n329629 );
buf ( n329631 , n329630 );
nor ( n329632 , n329624 , n329631 );
buf ( n329633 , n329632 );
buf ( n329634 , n329633 );
not ( n39209 , n329634 );
buf ( n329636 , n39209 );
buf ( n329637 , n329636 );
not ( n39212 , n329637 );
not ( n329639 , n329617 );
buf ( n329640 , n329627 );
buf ( n329641 , n329108 );
nand ( n39216 , n329640 , n329641 );
buf ( n39217 , n39216 );
not ( n329644 , n39217 );
and ( n39219 , n329639 , n329644 );
buf ( n39220 , n329600 );
buf ( n39221 , n329614 );
and ( n39222 , n39220 , n39221 );
buf ( n39223 , n39222 );
nor ( n329650 , n39219 , n39223 );
buf ( n329651 , n329650 );
not ( n329652 , n329651 );
or ( n329653 , n39212 , n329652 );
not ( n39228 , n33699 );
xor ( n329655 , n39228 , n324970 );
and ( n39230 , n329655 , n34542 );
and ( n329657 , n39228 , n324970 );
or ( n39232 , n39230 , n329657 );
xor ( n329659 , n324232 , n39232 );
not ( n329660 , n312275 );
not ( n329661 , n33807 );
nand ( n329662 , n325075 , n329661 );
not ( n39237 , n329662 );
and ( n329664 , n329660 , n39237 );
not ( n329665 , n325075 );
nand ( n39240 , n329665 , n33807 );
nor ( n329667 , n312275 , n39240 );
nor ( n39242 , n329664 , n329667 );
nand ( n39243 , n312275 , n325075 , n33807 );
nand ( n39244 , n312275 , n329665 , n329661 );
nand ( n39245 , n39242 , n39243 , n39244 );
and ( n39246 , n329659 , n39245 );
and ( n39247 , n324232 , n39232 );
or ( n39248 , n39246 , n39247 );
buf ( n329675 , n39248 );
not ( n39250 , n324116 );
xor ( n39251 , n39250 , n329399 );
nor ( n39252 , n312275 , n325075 );
or ( n39253 , n39252 , n329661 );
nand ( n39254 , n39253 , n34845 );
xor ( n39255 , n39251 , n39254 );
buf ( n329682 , n39255 );
nor ( n329683 , n329675 , n329682 );
buf ( n329684 , n329683 );
buf ( n329685 , n329684 );
xor ( n39260 , n39250 , n329399 );
and ( n329687 , n39260 , n39254 );
and ( n329688 , n39250 , n329399 );
or ( n39263 , n329687 , n329688 );
buf ( n329690 , n39263 );
buf ( n39265 , n328852 );
nor ( n39266 , n329690 , n39265 );
buf ( n39267 , n39266 );
buf ( n329694 , n39267 );
nor ( n329695 , n329685 , n329694 );
buf ( n329696 , n329695 );
xor ( n39271 , n324232 , n39232 );
xor ( n329698 , n39271 , n39245 );
not ( n329699 , n329698 );
not ( n39274 , n33706 );
buf ( n329701 , n39274 );
xor ( n39276 , n39228 , n324970 );
xor ( n39277 , n39276 , n34542 );
buf ( n329704 , n39277 );
xor ( n329705 , n329701 , n329704 );
xor ( n329706 , n329593 , n329595 );
and ( n39281 , n329706 , n329597 );
and ( n329708 , n329593 , n329595 );
or ( n39283 , n39281 , n329708 );
buf ( n329710 , n39283 );
buf ( n329711 , n329710 );
and ( n329712 , n329705 , n329711 );
and ( n39287 , n329701 , n329704 );
or ( n329714 , n329712 , n39287 );
buf ( n329715 , n329714 );
not ( n39290 , n329715 );
nand ( n329717 , n329699 , n39290 );
not ( n39292 , n329587 );
not ( n329719 , n329599 );
not ( n329720 , n329719 );
or ( n39295 , n39292 , n329720 );
nand ( n329722 , n39295 , n39165 );
nand ( n329723 , n329599 , n39160 );
nand ( n39298 , n329722 , n329723 );
buf ( n329725 , n39298 );
not ( n39300 , n329725 );
xor ( n39301 , n329701 , n329704 );
xor ( n39302 , n39301 , n329711 );
buf ( n329729 , n39302 );
buf ( n329730 , n329729 );
not ( n39305 , n329730 );
buf ( n329732 , n39305 );
buf ( n329733 , n329732 );
nand ( n329734 , n39300 , n329733 );
buf ( n329735 , n329734 );
nand ( n39310 , n329696 , n329717 , n329735 );
buf ( n39311 , n39310 );
buf ( n329738 , n328779 );
buf ( n329739 , n328857 );
nor ( n329740 , n329738 , n329739 );
buf ( n329741 , n329740 );
buf ( n329742 , n329741 );
buf ( n329743 , n328784 );
buf ( n329744 , n328729 );
nor ( n329745 , n329743 , n329744 );
buf ( n329746 , n329745 );
buf ( n329747 , n329746 );
nor ( n39322 , n329742 , n329747 );
buf ( n329749 , n39322 );
buf ( n329750 , n329749 );
xor ( n39325 , n329551 , n329552 );
xor ( n39326 , n39325 , n329554 );
buf ( n329753 , n39326 );
buf ( n329754 , n329753 );
buf ( n329755 , n34661 );
buf ( n329756 , n329484 );
xor ( n39331 , n329755 , n329756 );
buf ( n329758 , n329436 );
and ( n39333 , n39331 , n329758 );
and ( n39334 , n329755 , n329756 );
or ( n39335 , n39333 , n39334 );
buf ( n329762 , n39335 );
buf ( n329763 , n329762 );
nor ( n329764 , n329754 , n329763 );
buf ( n329765 , n329764 );
buf ( n329766 , n329765 );
buf ( n329767 , n328734 );
xor ( n39342 , n329755 , n329756 );
xor ( n39343 , n39342 , n329758 );
buf ( n329770 , n39343 );
buf ( n329771 , n329770 );
nor ( n329772 , n329767 , n329771 );
buf ( n329773 , n329772 );
buf ( n329774 , n329773 );
nor ( n329775 , n329766 , n329774 );
buf ( n329776 , n329775 );
buf ( n329777 , n329776 );
nand ( n329778 , n329750 , n329777 );
buf ( n329779 , n329778 );
buf ( n329780 , n329779 );
nor ( n329781 , n39311 , n329780 );
buf ( n329782 , n329781 );
buf ( n39357 , n329782 );
nand ( n39358 , n329653 , n39357 );
buf ( n39359 , n39358 );
buf ( n329786 , n39359 );
not ( n39361 , n329786 );
buf ( n329788 , n329219 );
buf ( n329789 , n329321 );
nor ( n329790 , n329788 , n329789 );
buf ( n329791 , n329790 );
buf ( n329792 , n329791 );
buf ( n329793 , n329316 );
buf ( n329794 , n33557 );
xor ( n39369 , n329794 , n329453 );
and ( n39370 , n39369 , n329487 );
and ( n329797 , n329794 , n329453 );
or ( n329798 , n39370 , n329797 );
buf ( n329799 , n329798 );
nor ( n39374 , n329793 , n329799 );
buf ( n39375 , n39374 );
buf ( n39376 , n39375 );
nor ( n39377 , n329792 , n39376 );
buf ( n39378 , n39377 );
buf ( n329805 , n39378 );
not ( n39380 , n329805 );
buf ( n39381 , n323640 );
not ( n329808 , n39381 );
buf ( n329809 , n329808 );
buf ( n329810 , n329448 );
xor ( n39385 , n329809 , n329810 );
buf ( n329812 , n329458 );
and ( n39387 , n39385 , n329812 );
and ( n39388 , n329809 , n329810 );
or ( n329815 , n39387 , n39388 );
buf ( n329816 , n329815 );
buf ( n39391 , n329816 );
xor ( n329818 , n329794 , n329453 );
xor ( n329819 , n329818 , n329487 );
buf ( n39394 , n329819 );
nor ( n39395 , n39391 , n39394 );
buf ( n39396 , n39395 );
buf ( n329823 , n39396 );
xor ( n39398 , n329809 , n329810 );
xor ( n329825 , n39398 , n329812 );
buf ( n329826 , n329825 );
buf ( n329827 , n329826 );
buf ( n329828 , n328660 );
nand ( n329829 , n329827 , n329828 );
buf ( n329830 , n329829 );
buf ( n329831 , n329830 );
or ( n329832 , n329823 , n329831 );
buf ( n329833 , n329816 );
buf ( n329834 , n329819 );
nand ( n329835 , n329833 , n329834 );
buf ( n329836 , n329835 );
buf ( n329837 , n329836 );
nand ( n39412 , n329832 , n329837 );
buf ( n329839 , n39412 );
buf ( n329840 , n329839 );
not ( n39415 , n329840 );
or ( n329842 , n39380 , n39415 );
buf ( n329843 , n329791 );
not ( n39418 , n329843 );
buf ( n329845 , n39418 );
buf ( n329846 , n329845 );
buf ( n329847 , n329316 );
buf ( n329848 , n329798 );
and ( n329849 , n329847 , n329848 );
buf ( n329850 , n329849 );
buf ( n329851 , n329850 );
and ( n39426 , n329846 , n329851 );
buf ( n329853 , n329219 );
buf ( n329854 , n329321 );
and ( n39429 , n329853 , n329854 );
buf ( n329856 , n39429 );
buf ( n329857 , n329856 );
nor ( n39432 , n39426 , n329857 );
buf ( n329859 , n39432 );
buf ( n329860 , n329859 );
nand ( n39435 , n329842 , n329860 );
buf ( n329862 , n39435 );
buf ( n329863 , n329862 );
not ( n329864 , n831 );
not ( n39439 , n306684 );
or ( n329866 , n329864 , n39439 );
nand ( n329867 , n329866 , n33663 );
buf ( n39442 , n329867 );
buf ( n329869 , n329425 );
xor ( n329870 , n39442 , n329869 );
xor ( n329871 , n329092 , n329093 );
xor ( n39446 , n329871 , n329095 );
buf ( n329873 , n39446 );
buf ( n329874 , n329873 );
and ( n329875 , n329870 , n329874 );
and ( n39450 , n39442 , n329869 );
or ( n329877 , n329875 , n39450 );
buf ( n329878 , n329877 );
not ( n329879 , n329878 );
not ( n329880 , n329103 );
and ( n39455 , n329879 , n329880 );
xor ( n329882 , n39442 , n329869 );
xor ( n329883 , n329882 , n329874 );
buf ( n329884 , n329883 );
buf ( n329885 , n329884 );
buf ( n329886 , n329224 );
nor ( n39461 , n329885 , n329886 );
buf ( n329888 , n39461 );
nor ( n39463 , n39455 , n329888 );
buf ( n329890 , n39463 );
and ( n329891 , n329863 , n329890 );
buf ( n329892 , n329891 );
buf ( n39467 , n329892 );
buf ( n329894 , n329884 );
buf ( n329895 , n329224 );
and ( n329896 , n329894 , n329895 );
buf ( n329897 , n329896 );
buf ( n329898 , n329897 );
not ( n329899 , n329898 );
not ( n329900 , n329103 );
buf ( n329901 , n329878 );
not ( n329902 , n329901 );
buf ( n329903 , n329902 );
nand ( n39478 , n329900 , n329903 );
buf ( n329905 , n39478 );
not ( n39480 , n329905 );
or ( n329907 , n329899 , n39480 );
buf ( n329908 , n329903 );
not ( n39483 , n329908 );
buf ( n329910 , n329103 );
nand ( n329911 , n39483 , n329910 );
buf ( n329912 , n329911 );
buf ( n329913 , n329912 );
nand ( n329914 , n329907 , n329913 );
buf ( n329915 , n329914 );
not ( n329916 , n329915 );
nand ( n39491 , n329916 , n329650 );
buf ( n329918 , n39491 );
nor ( n39493 , n39467 , n329918 );
buf ( n329920 , n39493 );
buf ( n329921 , n329920 );
not ( n329922 , n329921 );
and ( n39497 , n39361 , n329922 );
buf ( n329924 , n329717 );
not ( n39499 , n329924 );
buf ( n329926 , n39298 );
buf ( n329927 , n329729 );
nand ( n39502 , n329926 , n329927 );
buf ( n329929 , n39502 );
buf ( n329930 , n329929 );
not ( n39505 , n329930 );
buf ( n329932 , n39505 );
buf ( n329933 , n329932 );
not ( n39508 , n329933 );
or ( n329935 , n39499 , n39508 );
buf ( n329936 , n39290 );
not ( n329937 , n329936 );
buf ( n329938 , n329698 );
nand ( n329939 , n329937 , n329938 );
buf ( n329940 , n329939 );
buf ( n329941 , n329940 );
nand ( n329942 , n329935 , n329941 );
buf ( n329943 , n329942 );
buf ( n329944 , n329943 );
buf ( n329945 , n329696 );
and ( n39520 , n329944 , n329945 );
buf ( n329947 , n39248 );
buf ( n329948 , n39255 );
nand ( n329949 , n329947 , n329948 );
buf ( n329950 , n329949 );
buf ( n329951 , n329950 );
buf ( n329952 , n39267 );
or ( n329953 , n329951 , n329952 );
buf ( n329954 , n39263 );
buf ( n329955 , n328852 );
nand ( n39530 , n329954 , n329955 );
buf ( n39531 , n39530 );
buf ( n329958 , n39531 );
nand ( n39533 , n329953 , n329958 );
buf ( n329960 , n39533 );
buf ( n329961 , n329960 );
nor ( n39536 , n39520 , n329961 );
buf ( n329963 , n39536 );
buf ( n329964 , n329963 );
buf ( n329965 , n329746 );
buf ( n329966 , n328779 );
buf ( n329967 , n328857 );
nand ( n329968 , n329966 , n329967 );
buf ( n329969 , n329968 );
buf ( n329970 , n329969 );
or ( n329971 , n329965 , n329970 );
buf ( n329972 , n328784 );
buf ( n329973 , n328729 );
nand ( n329974 , n329972 , n329973 );
buf ( n329975 , n329974 );
buf ( n329976 , n329975 );
nand ( n329977 , n329971 , n329976 );
buf ( n329978 , n329977 );
buf ( n329979 , n329978 );
buf ( n329980 , n329776 );
and ( n39555 , n329979 , n329980 );
buf ( n329982 , n329765 );
buf ( n39557 , n329770 );
buf ( n39558 , n328734 );
nand ( n39559 , n39557 , n39558 );
buf ( n39560 , n39559 );
buf ( n329987 , n39560 );
or ( n39562 , n329982 , n329987 );
buf ( n329989 , n329762 );
buf ( n329990 , n329753 );
nand ( n329991 , n329989 , n329990 );
buf ( n329992 , n329991 );
buf ( n329993 , n329992 );
nand ( n39568 , n39562 , n329993 );
buf ( n329995 , n39568 );
buf ( n329996 , n329995 );
nor ( n39571 , n39555 , n329996 );
buf ( n329998 , n39571 );
buf ( n329999 , n329998 );
nand ( n39574 , n329964 , n329999 );
buf ( n330001 , n39574 );
buf ( n330002 , n330001 );
buf ( n39577 , n329998 );
buf ( n330004 , n329779 );
nand ( n39579 , n39577 , n330004 );
buf ( n330006 , n39579 );
buf ( n330007 , n330006 );
and ( n330008 , n330002 , n330007 );
nor ( n330009 , n39497 , n330008 );
buf ( n330010 , n330009 );
buf ( n330011 , n330010 );
not ( n330012 , n330011 );
buf ( n330013 , n330012 );
buf ( n330014 , n330013 );
not ( n39589 , n330014 );
or ( n39590 , n329585 , n39589 );
buf ( n39591 , n328678 );
buf ( n330018 , n328558 );
nor ( n39593 , n39591 , n330018 );
buf ( n330020 , n39593 );
buf ( n330021 , n330020 );
buf ( n39596 , n328553 );
buf ( n330023 , n323888 );
xor ( n39598 , n330023 , n329420 );
and ( n330025 , n39598 , n329466 );
and ( n39600 , n330023 , n329420 );
or ( n39601 , n330025 , n39600 );
buf ( n330028 , n39601 );
nor ( n39603 , n39596 , n330028 );
buf ( n330030 , n39603 );
buf ( n330031 , n330030 );
nor ( n39606 , n330021 , n330031 );
buf ( n330033 , n39606 );
buf ( n330034 , n330033 );
buf ( n330035 , n328655 );
xor ( n330036 , n323862 , n313441 );
xor ( n39611 , n330036 , n24026 );
xor ( n330038 , n33506 , n39611 );
and ( n39613 , n330038 , n329393 );
and ( n330040 , n33506 , n39611 );
or ( n39615 , n39613 , n330040 );
buf ( n330042 , n39615 );
nor ( n330043 , n330035 , n330042 );
buf ( n330044 , n330043 );
buf ( n330045 , n330044 );
buf ( n330046 , n328683 );
xor ( n39621 , n33506 , n39611 );
xor ( n330048 , n39621 , n329393 );
buf ( n330049 , n330048 );
nor ( n330050 , n330046 , n330049 );
buf ( n330051 , n330050 );
buf ( n330052 , n330051 );
nor ( n330053 , n330045 , n330052 );
buf ( n330054 , n330053 );
buf ( n330055 , n330054 );
nand ( n330056 , n330034 , n330055 );
buf ( n330057 , n330056 );
not ( n39632 , n330057 );
buf ( n39633 , n328756 );
buf ( n330060 , n328807 );
nor ( n39635 , n39633 , n330060 );
buf ( n39636 , n39635 );
buf ( n330063 , n39636 );
buf ( n330064 , n328802 );
buf ( n330065 , n328832 );
nand ( n39640 , n330064 , n330065 );
buf ( n330067 , n39640 );
buf ( n330068 , n330067 );
or ( n39643 , n330063 , n330068 );
buf ( n330070 , n328756 );
buf ( n330071 , n328807 );
nand ( n330072 , n330070 , n330071 );
buf ( n330073 , n330072 );
buf ( n330074 , n330073 );
nand ( n330075 , n39643 , n330074 );
buf ( n330076 , n330075 );
buf ( n330077 , n330076 );
xor ( n39652 , n330023 , n329420 );
xor ( n330079 , n39652 , n329466 );
buf ( n330080 , n330079 );
buf ( n39655 , n33469 );
xor ( n330082 , n39655 , n329415 );
and ( n330083 , n330082 , n329479 );
and ( n330084 , n39655 , n329415 );
or ( n39659 , n330083 , n330084 );
buf ( n330086 , n39659 );
nor ( n330087 , n330080 , n330086 );
buf ( n330088 , n330087 );
buf ( n330089 , n330088 );
xor ( n330090 , n39655 , n329415 );
xor ( n39665 , n330090 , n329479 );
buf ( n39666 , n39665 );
buf ( n39667 , n328761 );
nor ( n39668 , n39666 , n39667 );
buf ( n39669 , n39668 );
buf ( n330096 , n39669 );
nor ( n39671 , n330089 , n330096 );
buf ( n39672 , n39671 );
buf ( n330099 , n39672 );
nand ( n39674 , n330077 , n330099 );
buf ( n330101 , n39674 );
buf ( n330102 , n330101 );
buf ( n330103 , n330088 );
not ( n39678 , n330103 );
buf ( n330105 , n39678 );
buf ( n330106 , n330105 );
buf ( n330107 , n39665 );
buf ( n330108 , n328761 );
and ( n39683 , n330107 , n330108 );
buf ( n330110 , n39683 );
buf ( n330111 , n330110 );
and ( n330112 , n330106 , n330111 );
buf ( n330113 , n330079 );
buf ( n330114 , n39659 );
and ( n330115 , n330113 , n330114 );
buf ( n330116 , n330115 );
buf ( n330117 , n330116 );
nor ( n330118 , n330112 , n330117 );
buf ( n330119 , n330118 );
buf ( n39694 , n330119 );
and ( n39695 , n330102 , n39694 );
buf ( n39696 , n39695 );
not ( n330123 , n39696 );
and ( n39698 , n39632 , n330123 );
not ( n330125 , n330054 );
buf ( n330126 , n328553 );
buf ( n330127 , n39601 );
and ( n39702 , n330126 , n330127 );
buf ( n330129 , n39702 );
buf ( n330130 , n330129 );
not ( n39705 , n330130 );
buf ( n330132 , n330020 );
not ( n39707 , n330132 );
buf ( n330134 , n39707 );
buf ( n330135 , n330134 );
not ( n39710 , n330135 );
or ( n39711 , n39705 , n39710 );
buf ( n330138 , n328678 );
buf ( n330139 , n328558 );
nand ( n39714 , n330138 , n330139 );
buf ( n330141 , n39714 );
buf ( n330142 , n330141 );
nand ( n39717 , n39711 , n330142 );
buf ( n330144 , n39717 );
not ( n39719 , n330144 );
or ( n330146 , n330125 , n39719 );
buf ( n330147 , n330044 );
not ( n330148 , n330147 );
buf ( n39723 , n328683 );
buf ( n39724 , n330048 );
nand ( n39725 , n39723 , n39724 );
buf ( n39726 , n39725 );
buf ( n330153 , n39726 );
not ( n39728 , n330153 );
and ( n330155 , n330148 , n39728 );
buf ( n330156 , n328655 );
buf ( n330157 , n39615 );
and ( n330158 , n330156 , n330157 );
buf ( n330159 , n330158 );
buf ( n330160 , n330159 );
nor ( n330161 , n330155 , n330160 );
buf ( n330162 , n330161 );
nand ( n330163 , n330146 , n330162 );
nor ( n330164 , n39698 , n330163 );
buf ( n39739 , n330164 );
buf ( n330166 , n39672 );
buf ( n330167 , n39636 );
buf ( n330168 , n328802 );
buf ( n330169 , n328832 );
nor ( n39744 , n330168 , n330169 );
buf ( n39745 , n39744 );
buf ( n39746 , n39745 );
nor ( n39747 , n330167 , n39746 );
buf ( n330174 , n39747 );
buf ( n330175 , n330174 );
and ( n39750 , n330166 , n330175 );
buf ( n330177 , n39750 );
buf ( n330178 , n330177 );
buf ( n330179 , n328879 );
buf ( n330180 , n328924 );
nor ( n39755 , n330179 , n330180 );
buf ( n330182 , n39755 );
buf ( n330183 , n330182 );
not ( n39758 , n330183 );
buf ( n39759 , n39758 );
buf ( n330186 , n39759 );
not ( n39761 , n330186 );
buf ( n330188 , n33179 );
buf ( n330189 , n330188 );
xor ( n330190 , n320127 , n320330 );
xor ( n39765 , n330190 , n33180 );
not ( n330192 , n39765 );
not ( n330193 , n329500 );
nand ( n39768 , n330192 , n330193 );
and ( n330195 , n330189 , n39768 );
nor ( n330196 , n330192 , n330193 );
nor ( n39771 , n330195 , n330196 );
not ( n39772 , n39771 );
buf ( n39773 , n39772 );
buf ( n330200 , n328919 );
and ( n39775 , n39773 , n330200 );
buf ( n39776 , n39775 );
buf ( n330203 , n39776 );
not ( n39778 , n330203 );
or ( n39779 , n39761 , n39778 );
buf ( n330206 , n328879 );
buf ( n330207 , n328924 );
nand ( n39782 , n330206 , n330207 );
buf ( n330209 , n39782 );
buf ( n330210 , n330209 );
nand ( n39785 , n39779 , n330210 );
buf ( n330212 , n39785 );
buf ( n330213 , n330212 );
not ( n330214 , n323756 );
xor ( n330215 , n330214 , n329471 );
and ( n39790 , n330215 , n329396 );
and ( n330217 , n330214 , n329471 );
or ( n330218 , n39790 , n330217 );
nor ( n39793 , n328827 , n330218 );
buf ( n330220 , n39793 );
xor ( n330221 , n330214 , n329471 );
xor ( n39796 , n330221 , n329396 );
buf ( n330223 , n39796 );
buf ( n330224 , n328884 );
nor ( n39799 , n330223 , n330224 );
buf ( n39800 , n39799 );
buf ( n330227 , n39800 );
nor ( n39802 , n330220 , n330227 );
buf ( n39803 , n39802 );
buf ( n330230 , n39803 );
and ( n330231 , n330213 , n330230 );
nand ( n330232 , n39796 , n328884 );
or ( n39807 , n39793 , n330232 );
nand ( n330234 , n328827 , n330218 );
nand ( n330235 , n39807 , n330234 );
buf ( n330236 , n330235 );
nor ( n330237 , n330231 , n330236 );
buf ( n330238 , n330237 );
buf ( n330239 , n330238 );
xor ( n39814 , n323529 , n329409 );
xor ( n330241 , n39814 , n329474 );
buf ( n39816 , n330241 );
buf ( n39817 , n328964 );
nor ( n39818 , n39816 , n39817 );
buf ( n39819 , n39818 );
buf ( n330246 , n39819 );
buf ( n330247 , n328959 );
buf ( n330248 , n33077 );
buf ( n330249 , n329495 );
xor ( n330250 , n330248 , n330249 );
xor ( n39825 , n325728 , n292343 );
xor ( n330252 , n39825 , n325731 );
buf ( n330253 , n330252 );
and ( n39828 , n330250 , n330253 );
and ( n330255 , n330248 , n330249 );
or ( n330256 , n39828 , n330255 );
buf ( n330257 , n330256 );
buf ( n330258 , n330257 );
nand ( n39833 , n330247 , n330258 );
buf ( n330260 , n39833 );
buf ( n330261 , n330260 );
or ( n39836 , n330246 , n330261 );
buf ( n330263 , n330241 );
buf ( n330264 , n328964 );
nand ( n39839 , n330263 , n330264 );
buf ( n39840 , n39839 );
buf ( n330267 , n39840 );
nand ( n39842 , n39836 , n330267 );
buf ( n330269 , n39842 );
buf ( n330270 , n330269 );
not ( n39845 , n330270 );
and ( n39846 , n330188 , n329500 );
not ( n39847 , n330188 );
and ( n39848 , n39847 , n330193 );
nor ( n39849 , n39846 , n39848 );
and ( n39850 , n39849 , n39765 );
not ( n39851 , n39849 );
and ( n39852 , n39851 , n330192 );
nor ( n39853 , n39850 , n39852 );
buf ( n330280 , n39853 );
buf ( n330281 , n328585 );
or ( n39856 , n330280 , n330281 );
buf ( n330283 , n39856 );
buf ( n330284 , n330283 );
xor ( n39859 , n323529 , n329409 );
and ( n330286 , n39859 , n329474 );
and ( n330287 , n323529 , n329409 );
or ( n330288 , n330286 , n330287 );
or ( n330289 , n328580 , n330288 );
buf ( n330290 , n330289 );
and ( n330291 , n330284 , n330290 );
buf ( n330292 , n330291 );
buf ( n330293 , n330292 );
not ( n39868 , n330293 );
or ( n330295 , n39845 , n39868 );
buf ( n330296 , n330283 );
buf ( n330297 , n328580 );
buf ( n330298 , n330288 );
and ( n39873 , n330297 , n330298 );
buf ( n39874 , n39873 );
buf ( n39875 , n39874 );
and ( n39876 , n330296 , n39875 );
buf ( n330303 , n39853 );
buf ( n330304 , n328585 );
and ( n330305 , n330303 , n330304 );
buf ( n330306 , n330305 );
buf ( n330307 , n330306 );
nor ( n330308 , n39876 , n330307 );
buf ( n330309 , n330308 );
buf ( n330310 , n330309 );
nand ( n330311 , n330295 , n330310 );
buf ( n330312 , n330311 );
buf ( n330313 , n330312 );
buf ( n330314 , n39803 );
buf ( n330315 , n39772 );
buf ( n330316 , n328919 );
nor ( n39891 , n330315 , n330316 );
buf ( n330318 , n39891 );
buf ( n330319 , n330318 );
buf ( n330320 , n330182 );
nor ( n39895 , n330319 , n330320 );
buf ( n330322 , n39895 );
buf ( n330323 , n330322 );
and ( n39898 , n330314 , n330323 );
buf ( n330325 , n39898 );
buf ( n330326 , n330325 );
nand ( n39901 , n330313 , n330326 );
buf ( n330328 , n39901 );
buf ( n330329 , n330328 );
nand ( n330330 , n330239 , n330329 );
buf ( n330331 , n330330 );
buf ( n330332 , n330331 );
buf ( n330333 , n330057 );
not ( n39908 , n330333 );
buf ( n330335 , n39908 );
buf ( n330336 , n330335 );
nand ( n39911 , n330178 , n330332 , n330336 );
buf ( n330338 , n39911 );
buf ( n330339 , n330338 );
buf ( n330340 , n330335 );
buf ( n330341 , n330292 );
buf ( n330342 , n39819 );
buf ( n330343 , n328959 );
buf ( n330344 , n330257 );
nor ( n330345 , n330343 , n330344 );
buf ( n330346 , n330345 );
buf ( n330347 , n330346 );
nor ( n330348 , n330342 , n330347 );
buf ( n330349 , n330348 );
buf ( n330350 , n330349 );
nand ( n330351 , n330341 , n330350 );
buf ( n330352 , n330351 );
buf ( n330353 , n330352 );
not ( n330354 , n330353 );
buf ( n39929 , n330325 );
nand ( n39930 , n330354 , n39929 );
buf ( n39931 , n39930 );
buf ( n330358 , n39931 );
xor ( n39933 , n330248 , n330249 );
xor ( n330360 , n39933 , n330253 );
buf ( n330361 , n330360 );
buf ( n330362 , n330361 );
buf ( n330363 , n328990 );
nor ( n330364 , n330362 , n330363 );
buf ( n330365 , n330364 );
buf ( n330366 , n330365 );
not ( n330367 , n330366 );
buf ( n330368 , n330367 );
buf ( n39943 , n330368 );
buf ( n330370 , n329013 );
not ( n330371 , n330370 );
buf ( n330372 , n328985 );
not ( n330373 , n330372 );
buf ( n330374 , n330373 );
buf ( n330375 , n330374 );
nand ( n330376 , n330371 , n330375 );
buf ( n330377 , n330376 );
buf ( n330378 , n330377 );
nand ( n330379 , n39943 , n330378 );
buf ( n330380 , n330379 );
buf ( n330381 , n330380 );
not ( n39956 , n330381 );
buf ( n330383 , n39956 );
buf ( n330384 , n330383 );
buf ( n330385 , n329008 );
buf ( n330386 , n329061 );
nor ( n39961 , n330385 , n330386 );
buf ( n330388 , n39961 );
buf ( n330389 , n330388 );
buf ( n330390 , n329083 );
buf ( n330391 , n329056 );
nand ( n39966 , n330390 , n330391 );
buf ( n330393 , n39966 );
buf ( n330394 , n330393 );
or ( n330395 , n330389 , n330394 );
buf ( n330396 , n329008 );
buf ( n330397 , n329061 );
nand ( n330398 , n330396 , n330397 );
buf ( n330399 , n330398 );
buf ( n330400 , n330399 );
nand ( n39975 , n330395 , n330400 );
buf ( n330402 , n39975 );
buf ( n330403 , n330402 );
and ( n39978 , n330384 , n330403 );
buf ( n330405 , n328985 );
buf ( n330406 , n329013 );
nand ( n39981 , n330405 , n330406 );
buf ( n330408 , n39981 );
buf ( n330409 , n330408 );
buf ( n330410 , n330365 );
or ( n330411 , n330409 , n330410 );
buf ( n330412 , n330361 );
buf ( n330413 , n328990 );
nand ( n330414 , n330412 , n330413 );
buf ( n330415 , n330414 );
buf ( n330416 , n330415 );
nand ( n39991 , n330411 , n330416 );
buf ( n330418 , n39991 );
buf ( n39993 , n330418 );
nor ( n39994 , n39978 , n39993 );
buf ( n39995 , n39994 );
buf ( n330422 , n39995 );
buf ( n330423 , n330388 );
buf ( n330424 , n329056 );
buf ( n330425 , n329083 );
nor ( n330426 , n330424 , n330425 );
buf ( n330427 , n330426 );
buf ( n330428 , n330427 );
nor ( n330429 , n330423 , n330428 );
buf ( n330430 , n330429 );
buf ( n330431 , n330430 );
not ( n40006 , n330431 );
buf ( n330433 , n330380 );
nor ( n40008 , n40006 , n330433 );
buf ( n330435 , n40008 );
buf ( n330436 , n330435 );
buf ( n330437 , n329078 );
buf ( n330438 , n329131 );
nor ( n40013 , n330437 , n330438 );
buf ( n330440 , n40013 );
buf ( n330441 , n330440 );
buf ( n330442 , n329126 );
buf ( n330443 , n329150 );
nor ( n40018 , n330442 , n330443 );
buf ( n330445 , n40018 );
buf ( n330446 , n330445 );
nor ( n40021 , n330441 , n330446 );
buf ( n330448 , n40021 );
buf ( n40023 , n330448 );
buf ( n330450 , n329145 );
nand ( n330451 , n32793 , n32794 );
xor ( n330452 , n330451 , n329430 );
xor ( n330453 , n323395 , n323217 );
xor ( n40028 , n330453 , n32972 );
and ( n330455 , n330452 , n40028 );
and ( n330456 , n330451 , n329430 );
or ( n40031 , n330455 , n330456 );
buf ( n330458 , n40031 );
nor ( n330459 , n330450 , n330458 );
buf ( n330460 , n330459 );
buf ( n330461 , n330460 );
xor ( n330462 , n330451 , n329430 );
xor ( n40037 , n330462 , n40028 );
buf ( n330464 , n40037 );
buf ( n330465 , n329198 );
nor ( n40040 , n330464 , n330465 );
buf ( n330467 , n40040 );
buf ( n330468 , n330467 );
nor ( n330469 , n330461 , n330468 );
buf ( n330470 , n330469 );
buf ( n330471 , n330470 );
nand ( n330472 , n40023 , n330471 );
buf ( n330473 , n330472 );
buf ( n330474 , n330473 );
buf ( n330475 , n329237 );
buf ( n330476 , n329261 );
nor ( n40051 , n330475 , n330476 );
buf ( n330478 , n40051 );
buf ( n330479 , n330478 );
buf ( n330480 , n329193 );
buf ( n330481 , n329242 );
nor ( n40056 , n330480 , n330481 );
buf ( n40057 , n40056 );
buf ( n330484 , n40057 );
nor ( n40059 , n330479 , n330484 );
buf ( n40060 , n40059 );
buf ( n330487 , n40060 );
buf ( n330488 , n329256 );
buf ( n330489 , n328637 );
nor ( n330490 , n330488 , n330489 );
buf ( n330491 , n330490 );
buf ( n330492 , n330491 );
buf ( n40067 , n329340 );
buf ( n330494 , n328632 );
nand ( n330495 , n40067 , n330494 );
buf ( n330496 , n330495 );
buf ( n330497 , n330496 );
or ( n330498 , n330492 , n330497 );
buf ( n40073 , n329256 );
buf ( n40074 , n328637 );
nand ( n40075 , n40073 , n40074 );
buf ( n40076 , n40075 );
buf ( n330503 , n40076 );
nand ( n40078 , n330498 , n330503 );
buf ( n330505 , n40078 );
buf ( n330506 , n330505 );
and ( n330507 , n330487 , n330506 );
buf ( n330508 , n329261 );
buf ( n330509 , n329237 );
nand ( n40084 , n330508 , n330509 );
buf ( n330511 , n40084 );
buf ( n330512 , n330511 );
buf ( n330513 , n40057 );
or ( n330514 , n330512 , n330513 );
buf ( n40089 , n329193 );
buf ( n330516 , n329242 );
nand ( n40091 , n40089 , n330516 );
buf ( n40092 , n40091 );
buf ( n330519 , n40092 );
nand ( n330520 , n330514 , n330519 );
buf ( n330521 , n330520 );
buf ( n330522 , n330521 );
nor ( n330523 , n330507 , n330522 );
buf ( n330524 , n330523 );
buf ( n330525 , n330524 );
buf ( n330526 , n328632 );
buf ( n330527 , n329340 );
or ( n330528 , n330526 , n330527 );
buf ( n330529 , n330528 );
buf ( n330530 , n330529 );
buf ( n330531 , n329335 );
buf ( n40106 , n323001 );
not ( n40107 , n323124 );
buf ( n330534 , n40107 );
xor ( n330535 , n40106 , n330534 );
xor ( n40110 , n329322 , n329323 );
buf ( n330537 , n40110 );
buf ( n330538 , n330537 );
and ( n40113 , n330535 , n330538 );
and ( n330540 , n40106 , n330534 );
or ( n40115 , n40113 , n330540 );
buf ( n330542 , n40115 );
buf ( n330543 , n330542 );
nor ( n330544 , n330531 , n330543 );
buf ( n330545 , n330544 );
buf ( n330546 , n330545 );
xor ( n40121 , n40106 , n330534 );
xor ( n330548 , n40121 , n330538 );
buf ( n330549 , n330548 );
buf ( n330550 , n330549 );
buf ( n330551 , n329376 );
or ( n40126 , n330550 , n330551 );
buf ( n40127 , n40126 );
buf ( n40128 , n40127 );
buf ( n330555 , n323131 );
buf ( n330556 , n323039 );
not ( n330557 , n323057 );
not ( n40132 , n310283 );
or ( n330559 , n330557 , n40132 );
xor ( n330560 , n16943 , n307375 );
buf ( n330561 , n330560 );
nand ( n330562 , n831 , n330561 );
nand ( n40137 , n330559 , n330562 );
buf ( n330564 , n40137 );
and ( n40139 , n330556 , n330564 );
buf ( n330566 , n40139 );
buf ( n330567 , n330566 );
xor ( n40142 , n330555 , n330567 );
buf ( n330569 , n329371 );
and ( n40144 , n40142 , n330569 );
and ( n40145 , n330555 , n330567 );
or ( n40146 , n40144 , n40145 );
buf ( n330573 , n40146 );
buf ( n330574 , n330573 );
nand ( n40149 , n40128 , n330574 );
buf ( n330576 , n40149 );
buf ( n330577 , n330576 );
or ( n330578 , n330546 , n330577 );
buf ( n330579 , n330545 );
buf ( n330580 , n330549 );
buf ( n330581 , n329376 );
nand ( n330582 , n330580 , n330581 );
buf ( n330583 , n330582 );
buf ( n330584 , n330583 );
or ( n40159 , n330579 , n330584 );
buf ( n330586 , n329335 );
buf ( n330587 , n330542 );
nand ( n40162 , n330586 , n330587 );
buf ( n330589 , n40162 );
buf ( n330590 , n330589 );
nand ( n40165 , n330578 , n40159 , n330590 );
buf ( n330592 , n40165 );
buf ( n330593 , n330592 );
nand ( n330594 , n330530 , n330593 );
buf ( n330595 , n330594 );
buf ( n330596 , n330595 );
buf ( n330597 , n330491 );
nor ( n330598 , n330596 , n330597 );
buf ( n330599 , n330598 );
buf ( n330600 , n330599 );
buf ( n330601 , n40060 );
nand ( n330602 , n330600 , n330601 );
buf ( n330603 , n330602 );
buf ( n330604 , n330603 );
and ( n330605 , n330525 , n330604 );
buf ( n330606 , n330605 );
buf ( n330607 , n330606 );
nor ( n330608 , n330474 , n330607 );
buf ( n330609 , n330608 );
buf ( n40184 , n330609 );
nand ( n40185 , n330436 , n40184 );
buf ( n40186 , n40185 );
buf ( n330613 , n40186 );
buf ( n330614 , n330435 );
buf ( n330615 , n330460 );
buf ( n330616 , n40037 );
buf ( n330617 , n329198 );
nand ( n330618 , n330616 , n330617 );
buf ( n330619 , n330618 );
buf ( n330620 , n330619 );
or ( n330621 , n330615 , n330620 );
buf ( n330622 , n329145 );
buf ( n330623 , n40031 );
nand ( n40198 , n330622 , n330623 );
buf ( n330625 , n40198 );
buf ( n330626 , n330625 );
nand ( n330627 , n330621 , n330626 );
buf ( n330628 , n330627 );
buf ( n330629 , n330628 );
not ( n330630 , n330629 );
buf ( n330631 , n330448 );
not ( n330632 , n330631 );
or ( n330633 , n330630 , n330632 );
buf ( n330634 , n330440 );
not ( n330635 , n330634 );
buf ( n330636 , n329126 );
buf ( n330637 , n329150 );
nand ( n330638 , n330636 , n330637 );
buf ( n330639 , n330638 );
buf ( n330640 , n330639 );
not ( n330641 , n330640 );
and ( n40216 , n330635 , n330641 );
buf ( n330643 , n329078 );
buf ( n330644 , n329131 );
and ( n40219 , n330643 , n330644 );
buf ( n330646 , n40219 );
buf ( n330647 , n330646 );
nor ( n40222 , n40216 , n330647 );
buf ( n330649 , n40222 );
buf ( n330650 , n330649 );
nand ( n40225 , n330633 , n330650 );
buf ( n330652 , n40225 );
buf ( n330653 , n330652 );
nand ( n40228 , n330614 , n330653 );
buf ( n330655 , n40228 );
buf ( n330656 , n330655 );
and ( n40231 , n330422 , n330613 , n330656 );
buf ( n330658 , n40231 );
buf ( n330659 , n330658 );
nor ( n330660 , n330358 , n330659 );
buf ( n330661 , n330660 );
buf ( n330662 , n330661 );
buf ( n330663 , n330177 );
nand ( n330664 , n330340 , n330662 , n330663 );
buf ( n330665 , n330664 );
buf ( n330666 , n330665 );
nand ( n330667 , n39739 , n330339 , n330666 );
buf ( n330668 , n330667 );
buf ( n330669 , n330668 );
buf ( n330670 , n330669 );
buf ( n330671 , n330670 );
buf ( n330672 , n330671 );
buf ( n330673 , n329782 );
buf ( n330674 , n39478 );
buf ( n330675 , n329630 );
buf ( n330676 , n329888 );
nor ( n330677 , n330675 , n330676 );
buf ( n330678 , n330677 );
buf ( n330679 , n330678 );
buf ( n330680 , n329620 );
and ( n40255 , n330674 , n330679 , n330680 );
buf ( n40256 , n40255 );
buf ( n330683 , n40256 );
not ( n40258 , n330683 );
buf ( n330685 , n39378 );
buf ( n40260 , n329826 );
buf ( n330687 , n328660 );
nor ( n330688 , n40260 , n330687 );
buf ( n330689 , n330688 );
buf ( n330690 , n330689 );
buf ( n330691 , n39396 );
nor ( n330692 , n330690 , n330691 );
buf ( n330693 , n330692 );
buf ( n330694 , n330693 );
nand ( n330695 , n330685 , n330694 );
buf ( n330696 , n330695 );
buf ( n330697 , n330696 );
nor ( n330698 , n40258 , n330697 );
buf ( n330699 , n330698 );
buf ( n330700 , n330699 );
nand ( n330701 , n330673 , n330700 );
buf ( n330702 , n330701 );
buf ( n330703 , n330702 );
not ( n330704 , n330703 );
buf ( n330705 , n330704 );
buf ( n330706 , n330705 );
buf ( n330707 , n329583 );
and ( n40282 , n330672 , n330706 , n330707 );
buf ( n330709 , n329558 );
buf ( n330710 , n329561 );
nand ( n330711 , n330709 , n330710 );
buf ( n330712 , n330711 );
not ( n40287 , n330712 );
not ( n330714 , n329547 );
and ( n330715 , n40287 , n330714 );
buf ( n330716 , n329543 );
buf ( n330717 , n329293 );
and ( n330718 , n330716 , n330717 );
buf ( n330719 , n330718 );
nor ( n330720 , n330715 , n330719 );
buf ( n330721 , n330720 );
buf ( n330722 , n329580 );
or ( n330723 , n330721 , n330722 );
buf ( n330724 , n329572 );
not ( n40299 , n330724 );
buf ( n330726 , n40299 );
buf ( n330727 , n330726 );
not ( n330728 , n330727 );
buf ( n330729 , n329167 );
buf ( n330730 , n329298 );
nand ( n330731 , n330729 , n330730 );
buf ( n330732 , n330731 );
buf ( n330733 , n330732 );
not ( n40308 , n330733 );
and ( n330735 , n330728 , n40308 );
buf ( n40310 , n329172 );
buf ( n330737 , n329033 );
and ( n330738 , n40310 , n330737 );
buf ( n330739 , n330738 );
buf ( n330740 , n330739 );
nor ( n40315 , n330735 , n330740 );
buf ( n330742 , n40315 );
buf ( n330743 , n330742 );
nand ( n40318 , n330723 , n330743 );
buf ( n330745 , n40318 );
buf ( n330746 , n330745 );
buf ( n330747 , n330746 );
buf ( n330748 , n330747 );
buf ( n330749 , n330748 );
nor ( n330750 , n40282 , n330749 );
buf ( n330751 , n330750 );
buf ( n330752 , n330751 );
nand ( n40327 , n39590 , n330752 );
buf ( n330754 , n40327 );
buf ( n330755 , n330754 );
and ( n40330 , n330755 , n39109 );
not ( n330757 , n330755 );
and ( n40332 , n330757 , n39105 );
nor ( n40333 , n40330 , n40332 );
buf ( n330760 , n40333 );
buf ( n330761 , n328611 );
buf ( n330762 , n328938 );
and ( n330763 , n330761 , n330762 );
buf ( n330764 , n330763 );
buf ( n330765 , n330764 );
not ( n330766 , n330765 );
buf ( n330767 , n328611 );
buf ( n330768 , n328938 );
or ( n330769 , n330767 , n330768 );
buf ( n330770 , n330769 );
buf ( n330771 , n330770 );
nand ( n330772 , n330766 , n330771 );
buf ( n330773 , n330772 );
buf ( n330774 , n330773 );
buf ( n330775 , n330773 );
not ( n330776 , n330775 );
buf ( n330777 , n330776 );
buf ( n330778 , n330777 );
buf ( n330779 , n329583 );
buf ( n330780 , n34039 );
xor ( n40355 , n329509 , n329510 );
and ( n40356 , n40355 , n329513 );
and ( n330783 , n329509 , n329510 );
or ( n40358 , n40356 , n330783 );
buf ( n330785 , n40358 );
buf ( n330786 , n330785 );
xor ( n40361 , n330780 , n330786 );
buf ( n40362 , n33958 );
and ( n40363 , n324739 , n40362 );
not ( n40364 , n324739 );
not ( n40365 , n40362 );
and ( n40366 , n40364 , n40365 );
nor ( n40367 , n40363 , n40366 );
buf ( n330794 , n40367 );
xor ( n40369 , n40361 , n330794 );
buf ( n330796 , n40369 );
buf ( n330797 , n330796 );
xor ( n40372 , n329506 , n329507 );
and ( n40373 , n40372 , n329516 );
and ( n40374 , n329506 , n329507 );
or ( n40375 , n40373 , n40374 );
buf ( n330802 , n40375 );
buf ( n330803 , n330802 );
or ( n40378 , n330797 , n330803 );
buf ( n330805 , n40378 );
buf ( n330806 , n330805 );
buf ( n330807 , n329527 );
nand ( n40382 , n330806 , n330807 );
buf ( n330809 , n40382 );
buf ( n330810 , n330809 );
not ( n40385 , n320665 );
not ( n40386 , n40362 );
or ( n40387 , n40385 , n40386 );
or ( n40388 , n320665 , n33958 );
nand ( n40389 , n40388 , n34232 );
nand ( n40390 , n40387 , n40389 );
xor ( n40391 , n40390 , n324400 );
not ( n40392 , n34196 );
not ( n40393 , n324395 );
and ( n40394 , n40392 , n40393 );
and ( n40395 , n34196 , n324395 );
nor ( n40396 , n40394 , n40395 );
not ( n40397 , n40396 );
xor ( n40398 , n40391 , n40397 );
buf ( n40399 , n40398 );
xor ( n330826 , n330780 , n330786 );
and ( n40401 , n330826 , n330794 );
and ( n330828 , n330780 , n330786 );
or ( n330829 , n40401 , n330828 );
buf ( n330830 , n330829 );
buf ( n330831 , n330830 );
nor ( n330832 , n40399 , n330831 );
buf ( n330833 , n330832 );
buf ( n330834 , n330833 );
xor ( n330835 , n40390 , n324400 );
not ( n330836 , n40396 );
and ( n40411 , n330835 , n330836 );
and ( n330838 , n40390 , n324400 );
or ( n40413 , n40411 , n330838 );
buf ( n330840 , n40413 );
xor ( n40415 , n34159 , n324411 );
xor ( n40416 , n40415 , n34165 );
xor ( n40417 , n33979 , n40416 );
or ( n40418 , n324395 , n34107 );
nand ( n330845 , n40418 , n34086 );
nand ( n40420 , n34107 , n324395 );
nand ( n330847 , n330845 , n40420 );
xor ( n40422 , n40417 , n330847 );
buf ( n330849 , n40422 );
nor ( n330850 , n330840 , n330849 );
buf ( n330851 , n330850 );
buf ( n330852 , n330851 );
or ( n40427 , n330834 , n330852 );
buf ( n330854 , n40427 );
buf ( n330855 , n330854 );
nor ( n330856 , n330810 , n330855 );
buf ( n330857 , n330856 );
buf ( n330858 , n330857 );
and ( n40433 , n330779 , n330858 );
buf ( n40434 , n40433 );
buf ( n40435 , n40434 );
xor ( n330862 , n33979 , n40416 );
and ( n40437 , n330862 , n330847 );
and ( n330864 , n33979 , n40416 );
or ( n330865 , n40437 , n330864 );
not ( n40440 , n324411 );
not ( n40441 , n34165 );
or ( n330868 , n40440 , n40441 );
or ( n40443 , n34165 , n324411 );
nand ( n330870 , n40443 , n34159 );
nand ( n330871 , n330868 , n330870 );
xor ( n40446 , n33997 , n330871 );
xor ( n40447 , n40446 , n329490 );
nor ( n330874 , n330865 , n40447 );
buf ( n330875 , n330874 );
buf ( n330876 , n328606 );
xor ( n40451 , n33997 , n330871 );
and ( n40452 , n40451 , n329490 );
and ( n40453 , n33997 , n330871 );
or ( n40454 , n40452 , n40453 );
buf ( n330881 , n40454 );
nor ( n330882 , n330876 , n330881 );
buf ( n330883 , n330882 );
buf ( n330884 , n330883 );
nor ( n330885 , n330875 , n330884 );
buf ( n330886 , n330885 );
buf ( n330887 , n330886 );
and ( n330888 , n40435 , n330887 );
buf ( n330889 , n330888 );
buf ( n330890 , n330889 );
not ( n40465 , n330890 );
buf ( n330892 , n330013 );
not ( n40467 , n330892 );
or ( n40468 , n40465 , n40467 );
buf ( n330895 , n330671 );
buf ( n330896 , n330705 );
buf ( n330897 , n330889 );
and ( n40472 , n330895 , n330896 , n330897 );
buf ( n330899 , n330886 );
not ( n40474 , n330899 );
buf ( n330901 , n330857 );
not ( n40476 , n330901 );
buf ( n330903 , n330745 );
not ( n40478 , n330903 );
or ( n330905 , n40476 , n40478 );
buf ( n330906 , n330854 );
not ( n40481 , n330906 );
buf ( n330908 , n40481 );
buf ( n330909 , n330908 );
buf ( n330910 , n329521 );
not ( n40485 , n330910 );
buf ( n330912 , n330805 );
not ( n330913 , n330912 );
or ( n40488 , n40485 , n330913 );
buf ( n330915 , n330796 );
buf ( n330916 , n330802 );
nand ( n40491 , n330915 , n330916 );
buf ( n330918 , n40491 );
buf ( n330919 , n330918 );
nand ( n330920 , n40488 , n330919 );
buf ( n330921 , n330920 );
buf ( n330922 , n330921 );
and ( n330923 , n330909 , n330922 );
buf ( n330924 , n330830 );
buf ( n330925 , n40398 );
nand ( n330926 , n330924 , n330925 );
buf ( n330927 , n330926 );
buf ( n330928 , n330927 );
buf ( n330929 , n330851 );
or ( n40504 , n330928 , n330929 );
buf ( n330931 , n40413 );
buf ( n330932 , n40422 );
nand ( n40507 , n330931 , n330932 );
buf ( n330934 , n40507 );
buf ( n330935 , n330934 );
nand ( n40510 , n40504 , n330935 );
buf ( n330937 , n40510 );
buf ( n330938 , n330937 );
nor ( n40513 , n330923 , n330938 );
buf ( n330940 , n40513 );
buf ( n330941 , n330940 );
nand ( n40516 , n330905 , n330941 );
buf ( n330943 , n40516 );
buf ( n330944 , n330943 );
not ( n40519 , n330944 );
or ( n40520 , n40474 , n40519 );
buf ( n330947 , n330883 );
buf ( n330948 , n40447 );
buf ( n330949 , n330865 );
nand ( n40524 , n330948 , n330949 );
buf ( n330951 , n40524 );
buf ( n330952 , n330951 );
or ( n40527 , n330947 , n330952 );
buf ( n330954 , n328606 );
buf ( n330955 , n40454 );
nand ( n40530 , n330954 , n330955 );
buf ( n330957 , n40530 );
buf ( n330958 , n330957 );
nand ( n40533 , n40527 , n330958 );
buf ( n330960 , n40533 );
buf ( n330961 , n330960 );
not ( n40536 , n330961 );
buf ( n330963 , n40536 );
buf ( n330964 , n330963 );
nand ( n330965 , n40520 , n330964 );
buf ( n330966 , n330965 );
buf ( n330967 , n330966 );
nor ( n40542 , n40472 , n330967 );
buf ( n330969 , n40542 );
buf ( n330970 , n330969 );
nand ( n40545 , n40468 , n330970 );
buf ( n330972 , n40545 );
buf ( n330973 , n330972 );
and ( n40548 , n330973 , n330778 );
not ( n330975 , n330973 );
and ( n330976 , n330975 , n330774 );
nor ( n40551 , n40548 , n330976 );
buf ( n40552 , n40551 );
buf ( n330979 , n330883 );
not ( n40554 , n330979 );
buf ( n330981 , n330957 );
nand ( n40556 , n40554 , n330981 );
buf ( n40557 , n40556 );
buf ( n330984 , n40557 );
buf ( n330985 , n40557 );
not ( n40560 , n330985 );
buf ( n330987 , n40560 );
buf ( n330988 , n330987 );
buf ( n330989 , n40434 );
not ( n330990 , n330989 );
buf ( n330991 , n330990 );
buf ( n330992 , n330991 );
buf ( n330993 , n330874 );
nor ( n330994 , n330992 , n330993 );
buf ( n330995 , n330994 );
buf ( n330996 , n330995 );
not ( n40571 , n330996 );
buf ( n330998 , n330013 );
not ( n40573 , n330998 );
or ( n40574 , n40571 , n40573 );
buf ( n331001 , n330671 );
buf ( n331002 , n330705 );
buf ( n331003 , n330995 );
and ( n331004 , n331001 , n331002 , n331003 );
buf ( n331005 , n330943 );
not ( n331006 , n331005 );
buf ( n331007 , n331006 );
buf ( n331008 , n331007 );
buf ( n331009 , n330874 );
or ( n40584 , n331008 , n331009 );
buf ( n331011 , n330951 );
nand ( n40586 , n40584 , n331011 );
buf ( n331013 , n40586 );
buf ( n331014 , n331013 );
nor ( n40589 , n331004 , n331014 );
buf ( n331016 , n40589 );
buf ( n331017 , n331016 );
nand ( n40592 , n40574 , n331017 );
buf ( n331019 , n40592 );
buf ( n331020 , n331019 );
and ( n40595 , n331020 , n330988 );
not ( n40596 , n331020 );
and ( n331023 , n40596 , n330984 );
nor ( n40598 , n40595 , n331023 );
buf ( n331025 , n40598 );
buf ( n331026 , n330874 );
not ( n331027 , n331026 );
buf ( n331028 , n330951 );
nand ( n40603 , n331027 , n331028 );
buf ( n331030 , n40603 );
buf ( n331031 , n331030 );
buf ( n331032 , n331030 );
not ( n40607 , n331032 );
buf ( n331034 , n40607 );
buf ( n331035 , n331034 );
buf ( n331036 , n40434 );
not ( n331037 , n331036 );
buf ( n331038 , n330013 );
not ( n331039 , n331038 );
or ( n40614 , n331037 , n331039 );
buf ( n331041 , n330671 );
buf ( n331042 , n330705 );
buf ( n331043 , n40434 );
and ( n331044 , n331041 , n331042 , n331043 );
buf ( n331045 , n330943 );
nor ( n40620 , n331044 , n331045 );
buf ( n331047 , n40620 );
buf ( n331048 , n331047 );
nand ( n40623 , n40614 , n331048 );
buf ( n331050 , n40623 );
buf ( n331051 , n331050 );
and ( n40626 , n331051 , n331035 );
not ( n40627 , n331051 );
and ( n40628 , n40627 , n331031 );
nor ( n40629 , n40626 , n40628 );
buf ( n331056 , n40629 );
buf ( n331057 , n330851 );
not ( n40632 , n331057 );
buf ( n331059 , n330934 );
nand ( n40634 , n40632 , n331059 );
buf ( n331061 , n40634 );
buf ( n331062 , n331061 );
buf ( n331063 , n331061 );
not ( n40638 , n331063 );
buf ( n331065 , n40638 );
buf ( n331066 , n331065 );
buf ( n331067 , n329583 );
not ( n331068 , n331067 );
buf ( n331069 , n331068 );
buf ( n331070 , n331069 );
buf ( n331071 , n330809 );
not ( n40646 , n331071 );
buf ( n331073 , n330833 );
not ( n40648 , n331073 );
buf ( n331075 , n40648 );
buf ( n331076 , n331075 );
nand ( n331077 , n40646 , n331076 );
buf ( n331078 , n331077 );
buf ( n331079 , n331078 );
nor ( n331080 , n331070 , n331079 );
buf ( n331081 , n331080 );
buf ( n331082 , n331081 );
not ( n331083 , n331082 );
buf ( n331084 , n330013 );
not ( n40659 , n331084 );
or ( n331086 , n331083 , n40659 );
buf ( n331087 , n330671 );
buf ( n331088 , n330705 );
buf ( n331089 , n331081 );
and ( n40664 , n331087 , n331088 , n331089 );
buf ( n331091 , n330748 );
not ( n331092 , n331091 );
buf ( n331093 , n331092 );
buf ( n331094 , n331093 );
buf ( n331095 , n331078 );
or ( n40670 , n331094 , n331095 );
buf ( n331097 , n330921 );
buf ( n331098 , n331075 );
and ( n40673 , n331097 , n331098 );
buf ( n331100 , n330927 );
not ( n40675 , n331100 );
buf ( n331102 , n40675 );
buf ( n331103 , n331102 );
nor ( n40678 , n40673 , n331103 );
buf ( n331105 , n40678 );
buf ( n331106 , n331105 );
nand ( n40681 , n40670 , n331106 );
buf ( n331108 , n40681 );
buf ( n331109 , n331108 );
nor ( n331110 , n40664 , n331109 );
buf ( n331111 , n331110 );
buf ( n331112 , n331111 );
nand ( n40687 , n331086 , n331112 );
buf ( n331114 , n40687 );
buf ( n331115 , n331114 );
and ( n40690 , n331115 , n331066 );
not ( n40691 , n331115 );
and ( n40692 , n40691 , n331062 );
nor ( n40693 , n40690 , n40692 );
buf ( n331120 , n40693 );
buf ( n331121 , n331075 );
buf ( n331122 , n330927 );
nand ( n40697 , n331121 , n331122 );
buf ( n331124 , n40697 );
buf ( n331125 , n331124 );
buf ( n331126 , n331124 );
not ( n40701 , n331126 );
buf ( n331128 , n40701 );
buf ( n331129 , n331128 );
buf ( n331130 , n331069 );
buf ( n331131 , n330809 );
nor ( n40706 , n331130 , n331131 );
buf ( n331133 , n40706 );
buf ( n331134 , n331133 );
not ( n331135 , n331134 );
buf ( n331136 , n330013 );
not ( n40711 , n331136 );
or ( n40712 , n331135 , n40711 );
buf ( n331139 , n330671 );
buf ( n331140 , n330705 );
buf ( n331141 , n331133 );
and ( n40716 , n331139 , n331140 , n331141 );
buf ( n331143 , n331093 );
buf ( n331144 , n330809 );
or ( n40719 , n331143 , n331144 );
buf ( n331146 , n330921 );
not ( n40721 , n331146 );
buf ( n331148 , n40721 );
buf ( n331149 , n331148 );
nand ( n40724 , n40719 , n331149 );
buf ( n40725 , n40724 );
buf ( n331152 , n40725 );
nor ( n40727 , n40716 , n331152 );
buf ( n331154 , n40727 );
buf ( n331155 , n331154 );
nand ( n40730 , n40712 , n331155 );
buf ( n331157 , n40730 );
buf ( n331158 , n331157 );
and ( n40733 , n331158 , n331129 );
not ( n40734 , n331158 );
and ( n40735 , n40734 , n331125 );
nor ( n40736 , n40733 , n40735 );
buf ( n331163 , n40736 );
buf ( n331164 , n329365 );
not ( n40739 , n331164 );
xor ( n40740 , n322806 , n322878 );
xor ( n40741 , n40740 , n326869 );
and ( n40742 , n326877 , n40741 );
xor ( n40743 , n322806 , n322878 );
xor ( n40744 , n40743 , n326869 );
and ( n331171 , n329463 , n40744 );
and ( n40746 , n326877 , n329463 );
or ( n331173 , n40742 , n331171 , n40746 );
buf ( n331174 , n331173 );
not ( n40749 , n331174 );
or ( n40750 , n40739 , n40749 );
buf ( n40751 , n331173 );
buf ( n331178 , n329365 );
or ( n331179 , n40751 , n331178 );
nand ( n331180 , n40750 , n331179 );
buf ( n331181 , n331180 );
buf ( n40756 , n331181 );
buf ( n331183 , n331181 );
not ( n331184 , n331183 );
buf ( n331185 , n331184 );
buf ( n331186 , n331185 );
buf ( n331187 , n40434 );
buf ( n40762 , n330886 );
buf ( n331189 , n330770 );
buf ( n331190 , n328943 );
buf ( n331191 , n328901 );
or ( n40766 , n331190 , n331191 );
buf ( n331193 , n40766 );
buf ( n331194 , n331193 );
and ( n40769 , n331189 , n331194 );
buf ( n331196 , n40769 );
buf ( n331197 , n331196 );
nand ( n40772 , n40762 , n331197 );
buf ( n331199 , n40772 );
buf ( n331200 , n331199 );
buf ( n331201 , n328906 );
buf ( n331202 , n328527 );
nor ( n40777 , n331201 , n331202 );
buf ( n331204 , n40777 );
buf ( n331205 , n331204 );
buf ( n40780 , n38106 );
buf ( n331207 , n329275 );
nor ( n331208 , n40780 , n331207 );
buf ( n331209 , n331208 );
buf ( n331210 , n331209 );
nor ( n331211 , n331205 , n331210 );
buf ( n331212 , n331211 );
buf ( n331213 , n331212 );
buf ( n331214 , n329280 );
buf ( n331215 , n328703 );
or ( n331216 , n331214 , n331215 );
buf ( n331217 , n331216 );
buf ( n331218 , n331217 );
not ( n40793 , n331218 );
buf ( n331220 , n328708 );
xor ( n331221 , n322806 , n322878 );
xor ( n331222 , n331221 , n326869 );
xor ( n40797 , n326877 , n329463 );
xor ( n331224 , n331222 , n40797 );
buf ( n331225 , n331224 );
nor ( n331226 , n331220 , n331225 );
buf ( n331227 , n331226 );
buf ( n331228 , n331227 );
nor ( n331229 , n40793 , n331228 );
buf ( n331230 , n331229 );
buf ( n331231 , n331230 );
nand ( n331232 , n331213 , n331231 );
buf ( n331233 , n331232 );
buf ( n331234 , n331233 );
nor ( n40809 , n331200 , n331234 );
buf ( n40810 , n40809 );
buf ( n331237 , n40810 );
and ( n40812 , n331187 , n331237 );
buf ( n40813 , n40812 );
buf ( n331240 , n40813 );
not ( n40815 , n331240 );
buf ( n331242 , n330013 );
not ( n40817 , n331242 );
or ( n40818 , n40815 , n40817 );
buf ( n331245 , n330671 );
buf ( n331246 , n330705 );
buf ( n331247 , n40813 );
and ( n331248 , n331245 , n331246 , n331247 );
buf ( n331249 , n40810 );
not ( n331250 , n331249 );
buf ( n331251 , n330943 );
not ( n40826 , n331251 );
or ( n331253 , n331250 , n40826 );
buf ( n331254 , n331196 );
not ( n331255 , n331254 );
buf ( n331256 , n330960 );
not ( n40831 , n331256 );
or ( n331258 , n331255 , n40831 );
buf ( n331259 , n330764 );
buf ( n331260 , n331193 );
and ( n40835 , n331259 , n331260 );
buf ( n331262 , n328943 );
buf ( n331263 , n328901 );
and ( n40838 , n331262 , n331263 );
buf ( n40839 , n40838 );
buf ( n331266 , n40839 );
nor ( n331267 , n40835 , n331266 );
buf ( n331268 , n331267 );
buf ( n331269 , n331268 );
nand ( n331270 , n331258 , n331269 );
buf ( n331271 , n331270 );
buf ( n331272 , n331271 );
buf ( n331273 , n331233 );
not ( n40848 , n331273 );
buf ( n331275 , n40848 );
buf ( n331276 , n331275 );
and ( n40851 , n331272 , n331276 );
buf ( n331278 , n328906 );
buf ( n331279 , n328527 );
nand ( n40854 , n331278 , n331279 );
buf ( n331281 , n40854 );
buf ( n331282 , n331281 );
buf ( n331283 , n331209 );
or ( n40858 , n331282 , n331283 );
buf ( n40859 , n38106 );
buf ( n40860 , n329275 );
nand ( n40861 , n40859 , n40860 );
buf ( n40862 , n40861 );
buf ( n331289 , n40862 );
nand ( n331290 , n40858 , n331289 );
buf ( n331291 , n331290 );
buf ( n331292 , n331291 );
buf ( n331293 , n331230 );
and ( n331294 , n331292 , n331293 );
buf ( n331295 , n329280 );
buf ( n331296 , n328703 );
nand ( n331297 , n331295 , n331296 );
buf ( n331298 , n331297 );
buf ( n331299 , n331298 );
buf ( n331300 , n331227 );
or ( n331301 , n331299 , n331300 );
buf ( n331302 , n328708 );
buf ( n331303 , n331224 );
nand ( n40878 , n331302 , n331303 );
buf ( n331305 , n40878 );
buf ( n331306 , n331305 );
nand ( n40881 , n331301 , n331306 );
buf ( n331308 , n40881 );
buf ( n331309 , n331308 );
nor ( n331310 , n40851 , n331294 , n331309 );
buf ( n331311 , n331310 );
buf ( n331312 , n331311 );
nand ( n331313 , n331253 , n331312 );
buf ( n331314 , n331313 );
buf ( n331315 , n331314 );
nor ( n331316 , n331248 , n331315 );
buf ( n331317 , n331316 );
buf ( n331318 , n331317 );
nand ( n40893 , n40818 , n331318 );
buf ( n40894 , n40893 );
buf ( n331321 , n40894 );
and ( n40896 , n331321 , n331186 );
not ( n40897 , n331321 );
and ( n40898 , n40897 , n40756 );
nor ( n40899 , n40896 , n40898 );
buf ( n331326 , n40899 );
buf ( n331327 , n331217 );
buf ( n331328 , n331298 );
nand ( n331329 , n331327 , n331328 );
buf ( n331330 , n331329 );
buf ( n331331 , n331330 );
buf ( n40906 , n331330 );
not ( n331333 , n40906 );
buf ( n331334 , n331333 );
buf ( n331335 , n331334 );
buf ( n40910 , n330991 );
buf ( n331337 , n331199 );
not ( n331338 , n331337 );
buf ( n40913 , n331212 );
nand ( n40914 , n331338 , n40913 );
buf ( n40915 , n40914 );
buf ( n331342 , n40915 );
nor ( n331343 , n40910 , n331342 );
buf ( n331344 , n331343 );
buf ( n331345 , n331344 );
not ( n331346 , n331345 );
buf ( n331347 , n330013 );
not ( n331348 , n331347 );
or ( n331349 , n331346 , n331348 );
buf ( n331350 , n330671 );
buf ( n331351 , n330705 );
buf ( n331352 , n331344 );
and ( n40927 , n331350 , n331351 , n331352 );
buf ( n331354 , n331007 );
buf ( n331355 , n40915 );
or ( n40930 , n331354 , n331355 );
buf ( n331357 , n331271 );
buf ( n331358 , n331212 );
and ( n40933 , n331357 , n331358 );
buf ( n331360 , n331291 );
nor ( n331361 , n40933 , n331360 );
buf ( n331362 , n331361 );
buf ( n331363 , n331362 );
nand ( n331364 , n40930 , n331363 );
buf ( n331365 , n331364 );
buf ( n331366 , n331365 );
nor ( n40941 , n40927 , n331366 );
buf ( n40942 , n40941 );
buf ( n331369 , n40942 );
nand ( n40944 , n331349 , n331369 );
buf ( n331371 , n40944 );
buf ( n331372 , n331371 );
and ( n40947 , n331372 , n331335 );
not ( n40948 , n331372 );
and ( n40949 , n40948 , n331331 );
nor ( n40950 , n40947 , n40949 );
buf ( n331377 , n40950 );
buf ( n331378 , n39151 );
not ( n40953 , n331378 );
buf ( n331380 , n40953 );
buf ( n331381 , n331380 );
not ( n40956 , n331381 );
buf ( n331383 , n330732 );
nand ( n40958 , n40956 , n331383 );
buf ( n331385 , n40958 );
buf ( n331386 , n331385 );
buf ( n331387 , n331385 );
not ( n331388 , n331387 );
buf ( n331389 , n331388 );
buf ( n331390 , n331389 );
buf ( n331391 , n39141 );
not ( n40966 , n331391 );
buf ( n331393 , n40966 );
buf ( n331394 , n331393 );
not ( n40969 , n331394 );
buf ( n331396 , n330013 );
not ( n331397 , n331396 );
or ( n331398 , n40969 , n331397 );
buf ( n331399 , n330671 );
buf ( n331400 , n330705 );
buf ( n331401 , n331393 );
and ( n331402 , n331399 , n331400 , n331401 );
buf ( n331403 , n330720 );
not ( n331404 , n331403 );
buf ( n331405 , n331404 );
buf ( n331406 , n331405 );
nor ( n40981 , n331402 , n331406 );
buf ( n331408 , n40981 );
buf ( n331409 , n331408 );
nand ( n40984 , n331398 , n331409 );
buf ( n331411 , n40984 );
buf ( n331412 , n331411 );
and ( n40987 , n331412 , n331390 );
not ( n331414 , n331412 );
and ( n40989 , n331414 , n331386 );
nor ( n40990 , n40987 , n40989 );
buf ( n331417 , n40990 );
buf ( n331418 , n330719 );
buf ( n331419 , n329547 );
nor ( n331420 , n331418 , n331419 );
buf ( n331421 , n331420 );
buf ( n331422 , n331421 );
not ( n40997 , n331422 );
buf ( n331424 , n40997 );
buf ( n331425 , n331424 );
buf ( n331426 , n331421 );
buf ( n331427 , n39138 );
not ( n331428 , n331427 );
buf ( n331429 , n330013 );
not ( n41004 , n331429 );
or ( n331431 , n331428 , n41004 );
buf ( n331432 , n330671 );
buf ( n331433 , n330705 );
buf ( n331434 , n39138 );
and ( n331435 , n331432 , n331433 , n331434 );
buf ( n331436 , n330712 );
not ( n41011 , n331436 );
buf ( n331438 , n41011 );
buf ( n331439 , n331438 );
nor ( n41014 , n331435 , n331439 );
buf ( n41015 , n41014 );
buf ( n331442 , n41015 );
nand ( n41017 , n331431 , n331442 );
buf ( n41018 , n41017 );
buf ( n331445 , n41018 );
and ( n331446 , n331445 , n331426 );
not ( n41021 , n331445 );
and ( n331448 , n41021 , n331425 );
nor ( n331449 , n331446 , n331448 );
buf ( n331450 , n331449 );
buf ( n331451 , n331227 );
not ( n41026 , n331451 );
buf ( n331453 , n331305 );
nand ( n331454 , n41026 , n331453 );
buf ( n331455 , n331454 );
buf ( n331456 , n331455 );
buf ( n331457 , n331455 );
not ( n41032 , n331457 );
buf ( n331459 , n41032 );
buf ( n331460 , n331459 );
buf ( n331461 , n40434 );
buf ( n331462 , n331212 );
buf ( n331463 , n331217 );
and ( n41038 , n331462 , n331463 );
buf ( n331465 , n41038 );
buf ( n331466 , n331465 );
not ( n41041 , n331466 );
buf ( n331468 , n331199 );
nor ( n331469 , n41041 , n331468 );
buf ( n331470 , n331469 );
buf ( n331471 , n331470 );
and ( n331472 , n331461 , n331471 );
buf ( n331473 , n331472 );
buf ( n331474 , n331473 );
not ( n41049 , n331474 );
buf ( n331476 , n330013 );
not ( n331477 , n331476 );
or ( n41052 , n41049 , n331477 );
buf ( n331479 , n330671 );
buf ( n331480 , n330705 );
buf ( n331481 , n331473 );
and ( n331482 , n331479 , n331480 , n331481 );
buf ( n331483 , n331470 );
not ( n331484 , n331483 );
buf ( n331485 , n330943 );
not ( n41060 , n331485 );
or ( n331487 , n331484 , n41060 );
buf ( n331488 , n331271 );
buf ( n331489 , n331465 );
and ( n331490 , n331488 , n331489 );
buf ( n331491 , n331217 );
not ( n41066 , n331491 );
buf ( n331493 , n331291 );
not ( n331494 , n331493 );
or ( n331495 , n41066 , n331494 );
buf ( n331496 , n331298 );
nand ( n331497 , n331495 , n331496 );
buf ( n331498 , n331497 );
buf ( n331499 , n331498 );
nor ( n331500 , n331490 , n331499 );
buf ( n331501 , n331500 );
buf ( n331502 , n331501 );
nand ( n331503 , n331487 , n331502 );
buf ( n331504 , n331503 );
buf ( n331505 , n331504 );
nor ( n331506 , n331482 , n331505 );
buf ( n331507 , n331506 );
buf ( n331508 , n331507 );
nand ( n41083 , n41052 , n331508 );
buf ( n331510 , n41083 );
buf ( n331511 , n331510 );
and ( n41086 , n331511 , n331460 );
not ( n41087 , n331511 );
and ( n41088 , n41087 , n331456 );
nor ( n41089 , n41086 , n41088 );
buf ( n331516 , n41089 );
buf ( n41091 , n330726 );
buf ( n41092 , n330739 );
nor ( n41093 , n41091 , n41092 );
buf ( n41094 , n41093 );
buf ( n331521 , n41094 );
not ( n331522 , n331521 );
buf ( n331523 , n331522 );
buf ( n331524 , n331523 );
buf ( n331525 , n41094 );
buf ( n331526 , n39141 );
buf ( n331527 , n331380 );
nor ( n41102 , n331526 , n331527 );
buf ( n331529 , n41102 );
buf ( n331530 , n331529 );
not ( n331531 , n331530 );
buf ( n331532 , n330013 );
not ( n41107 , n331532 );
or ( n41108 , n331531 , n41107 );
buf ( n331535 , n330671 );
buf ( n331536 , n330705 );
buf ( n331537 , n331529 );
and ( n41112 , n331535 , n331536 , n331537 );
buf ( n331539 , n330720 );
buf ( n331540 , n331380 );
or ( n331541 , n331539 , n331540 );
buf ( n331542 , n330732 );
nand ( n41117 , n331541 , n331542 );
buf ( n331544 , n41117 );
buf ( n331545 , n331544 );
nor ( n41120 , n41112 , n331545 );
buf ( n331547 , n41120 );
buf ( n331548 , n331547 );
nand ( n41123 , n41108 , n331548 );
buf ( n41124 , n41123 );
buf ( n331551 , n41124 );
and ( n41126 , n331551 , n331525 );
not ( n41127 , n331551 );
and ( n331554 , n41127 , n331524 );
nor ( n41129 , n41126 , n331554 );
buf ( n331556 , n41129 );
buf ( n331557 , n331209 );
not ( n41132 , n331557 );
buf ( n331559 , n40862 );
nand ( n41134 , n41132 , n331559 );
buf ( n331561 , n41134 );
buf ( n331562 , n331561 );
buf ( n41137 , n331561 );
not ( n41138 , n41137 );
buf ( n41139 , n41138 );
buf ( n331566 , n41139 );
buf ( n331567 , n40434 );
buf ( n331568 , n331199 );
buf ( n331569 , n331204 );
nor ( n41144 , n331568 , n331569 );
buf ( n331571 , n41144 );
buf ( n331572 , n331571 );
and ( n331573 , n331567 , n331572 );
buf ( n331574 , n331573 );
buf ( n331575 , n331574 );
not ( n331576 , n331575 );
buf ( n331577 , n330013 );
not ( n331578 , n331577 );
or ( n41153 , n331576 , n331578 );
buf ( n331580 , n330671 );
buf ( n331581 , n330705 );
buf ( n331582 , n331574 );
and ( n41157 , n331580 , n331581 , n331582 );
buf ( n331584 , n331571 );
not ( n41159 , n331584 );
buf ( n331586 , n330943 );
not ( n331587 , n331586 );
or ( n331588 , n41159 , n331587 );
buf ( n331589 , n331271 );
not ( n331590 , n331589 );
buf ( n331591 , n331590 );
buf ( n331592 , n331591 );
not ( n331593 , n331592 );
buf ( n331594 , n331204 );
not ( n41169 , n331594 );
and ( n41170 , n331593 , n41169 );
buf ( n41171 , n331281 );
not ( n41172 , n41171 );
buf ( n331599 , n41172 );
buf ( n331600 , n331599 );
nor ( n41175 , n41170 , n331600 );
buf ( n331602 , n41175 );
buf ( n331603 , n331602 );
nand ( n331604 , n331588 , n331603 );
buf ( n331605 , n331604 );
buf ( n331606 , n331605 );
nor ( n331607 , n41157 , n331606 );
buf ( n331608 , n331607 );
buf ( n331609 , n331608 );
nand ( n41184 , n41153 , n331609 );
buf ( n331611 , n41184 );
buf ( n331612 , n331611 );
and ( n41187 , n331612 , n331566 );
not ( n41188 , n331612 );
and ( n41189 , n41188 , n331562 );
nor ( n41190 , n41187 , n41189 );
buf ( n331617 , n41190 );
buf ( n331618 , n331599 );
buf ( n331619 , n331204 );
nor ( n41194 , n331618 , n331619 );
buf ( n331621 , n41194 );
buf ( n331622 , n331621 );
not ( n331623 , n331622 );
buf ( n331624 , n331623 );
buf ( n331625 , n331624 );
buf ( n331626 , n331621 );
buf ( n331627 , n330991 );
buf ( n331628 , n331199 );
nor ( n41203 , n331627 , n331628 );
buf ( n331630 , n41203 );
buf ( n331631 , n331630 );
not ( n41206 , n331631 );
buf ( n331633 , n330013 );
not ( n41208 , n331633 );
or ( n41209 , n41206 , n41208 );
buf ( n331636 , n330671 );
buf ( n331637 , n330705 );
buf ( n331638 , n331630 );
and ( n41213 , n331636 , n331637 , n331638 );
buf ( n331640 , n331007 );
buf ( n331641 , n331199 );
or ( n41216 , n331640 , n331641 );
buf ( n331643 , n331591 );
nand ( n41218 , n41216 , n331643 );
buf ( n331645 , n41218 );
buf ( n331646 , n331645 );
nor ( n331647 , n41213 , n331646 );
buf ( n331648 , n331647 );
buf ( n331649 , n331648 );
nand ( n41224 , n41209 , n331649 );
buf ( n331651 , n41224 );
buf ( n331652 , n331651 );
and ( n331653 , n331652 , n331626 );
not ( n41228 , n331652 );
and ( n331655 , n41228 , n331625 );
nor ( n331656 , n331653 , n331655 );
buf ( n331657 , n331656 );
buf ( n331658 , n40839 );
not ( n41233 , n331658 );
buf ( n331660 , n331193 );
nand ( n331661 , n41233 , n331660 );
buf ( n331662 , n331661 );
buf ( n41237 , n331662 );
buf ( n331664 , n331662 );
not ( n331665 , n331664 );
buf ( n331666 , n331665 );
buf ( n331667 , n331666 );
buf ( n331668 , n330991 );
buf ( n331669 , n330886 );
buf ( n331670 , n330770 );
nand ( n331671 , n331669 , n331670 );
buf ( n331672 , n331671 );
buf ( n331673 , n331672 );
nor ( n331674 , n331668 , n331673 );
buf ( n331675 , n331674 );
buf ( n331676 , n331675 );
not ( n41251 , n331676 );
buf ( n331678 , n330013 );
not ( n41253 , n331678 );
or ( n41254 , n41251 , n41253 );
buf ( n331681 , n330671 );
buf ( n331682 , n330705 );
buf ( n331683 , n331675 );
and ( n331684 , n331681 , n331682 , n331683 );
buf ( n331685 , n331007 );
buf ( n331686 , n331672 );
or ( n331687 , n331685 , n331686 );
buf ( n331688 , n330960 );
buf ( n331689 , n330770 );
and ( n331690 , n331688 , n331689 );
buf ( n331691 , n330764 );
nor ( n331692 , n331690 , n331691 );
buf ( n331693 , n331692 );
buf ( n331694 , n331693 );
nand ( n331695 , n331687 , n331694 );
buf ( n331696 , n331695 );
buf ( n331697 , n331696 );
nor ( n331698 , n331684 , n331697 );
buf ( n331699 , n331698 );
buf ( n331700 , n331699 );
nand ( n331701 , n41254 , n331700 );
buf ( n331702 , n331701 );
buf ( n331703 , n331702 );
and ( n41278 , n331703 , n331667 );
not ( n41279 , n331703 );
and ( n41280 , n41279 , n41237 );
nor ( n41281 , n41278 , n41280 );
buf ( n331708 , n41281 );
buf ( n331709 , n329746 );
not ( n41284 , n331709 );
buf ( n331711 , n329975 );
nand ( n41286 , n41284 , n331711 );
buf ( n331713 , n41286 );
buf ( n331714 , n331713 );
buf ( n331715 , n331713 );
not ( n41290 , n331715 );
buf ( n331717 , n41290 );
buf ( n331718 , n331717 );
buf ( n331719 , n39310 );
not ( n331720 , n331719 );
buf ( n331721 , n331720 );
buf ( n331722 , n331721 );
buf ( n331723 , n329741 );
not ( n41298 , n331723 );
buf ( n41299 , n41298 );
buf ( n331726 , n41299 );
nand ( n331727 , n331722 , n331726 );
buf ( n331728 , n331727 );
buf ( n331729 , n331728 );
not ( n331730 , n330699 );
buf ( n331731 , n331730 );
nor ( n331732 , n331729 , n331731 );
buf ( n331733 , n331732 );
buf ( n331734 , n331733 );
not ( n331735 , n331734 );
buf ( n331736 , n330671 );
not ( n41311 , n331736 );
or ( n331738 , n331735 , n41311 );
buf ( n41313 , n331728 );
not ( n331740 , n41313 );
buf ( n331741 , n331740 );
buf ( n331742 , n331741 );
buf ( n41317 , n329862 );
buf ( n331744 , n40256 );
nand ( n331745 , n41317 , n331744 );
buf ( n331746 , n331745 );
buf ( n331747 , n331746 );
buf ( n331748 , n329915 );
buf ( n331749 , n329633 );
nand ( n41324 , n331748 , n331749 );
buf ( n331751 , n41324 );
buf ( n331752 , n331751 );
buf ( n331753 , n329650 );
nand ( n331754 , n331747 , n331752 , n331753 );
buf ( n331755 , n331754 );
buf ( n331756 , n331755 );
not ( n331757 , n331756 );
buf ( n331758 , n331757 );
buf ( n331759 , n331758 );
not ( n331760 , n331759 );
buf ( n331761 , n331760 );
buf ( n331762 , n331761 );
and ( n331763 , n331742 , n331762 );
buf ( n331764 , n41299 );
not ( n331765 , n331764 );
buf ( n331766 , n329963 );
not ( n331767 , n331766 );
buf ( n331768 , n331767 );
buf ( n331769 , n331768 );
not ( n331770 , n331769 );
or ( n41345 , n331765 , n331770 );
buf ( n331772 , n329969 );
nand ( n41347 , n41345 , n331772 );
buf ( n331774 , n41347 );
buf ( n331775 , n331774 );
nor ( n331776 , n331763 , n331775 );
buf ( n331777 , n331776 );
buf ( n331778 , n331777 );
nand ( n41353 , n331738 , n331778 );
buf ( n331780 , n41353 );
buf ( n331781 , n331780 );
and ( n331782 , n331781 , n331718 );
not ( n331783 , n331781 );
and ( n41358 , n331783 , n331714 );
nor ( n41359 , n331782 , n41358 );
buf ( n41360 , n41359 );
buf ( n331787 , n331438 );
not ( n41362 , n331787 );
buf ( n331789 , n39138 );
nand ( n41364 , n41362 , n331789 );
buf ( n331791 , n41364 );
buf ( n331792 , n331791 );
buf ( n331793 , n331791 );
not ( n41368 , n331793 );
buf ( n331795 , n41368 );
buf ( n331796 , n331795 );
buf ( n331797 , n330671 );
not ( n41372 , n331797 );
buf ( n331799 , n330705 );
not ( n41374 , n331799 );
or ( n331801 , n41372 , n41374 );
buf ( n331802 , n330010 );
nand ( n331803 , n331801 , n331802 );
buf ( n331804 , n331803 );
buf ( n331805 , n331804 );
and ( n331806 , n331805 , n331796 );
not ( n331807 , n331805 );
and ( n41382 , n331807 , n331792 );
nor ( n331809 , n331806 , n41382 );
buf ( n331810 , n331809 );
buf ( n331811 , n329765 );
not ( n41386 , n331811 );
buf ( n331813 , n329992 );
nand ( n41388 , n41386 , n331813 );
buf ( n331815 , n41388 );
buf ( n331816 , n331815 );
buf ( n331817 , n331815 );
not ( n41392 , n331817 );
buf ( n331819 , n41392 );
buf ( n331820 , n331819 );
buf ( n331821 , n331721 );
buf ( n331822 , n329749 );
not ( n331823 , n331822 );
buf ( n331824 , n329773 );
nor ( n41399 , n331823 , n331824 );
buf ( n331826 , n41399 );
buf ( n331827 , n331826 );
nand ( n331828 , n331821 , n331827 );
buf ( n331829 , n331828 );
buf ( n331830 , n331829 );
buf ( n331831 , n331730 );
nor ( n41406 , n331830 , n331831 );
buf ( n331833 , n41406 );
buf ( n331834 , n331833 );
not ( n41409 , n331834 );
buf ( n331836 , n330671 );
not ( n41411 , n331836 );
or ( n41412 , n41409 , n41411 );
buf ( n331839 , n331829 );
not ( n41414 , n331839 );
buf ( n331841 , n41414 );
buf ( n331842 , n331841 );
buf ( n331843 , n331761 );
and ( n41418 , n331842 , n331843 );
buf ( n41419 , n331826 );
not ( n41420 , n41419 );
buf ( n331847 , n331768 );
not ( n331848 , n331847 );
or ( n41423 , n41420 , n331848 );
buf ( n331850 , n329978 );
not ( n331851 , n331850 );
buf ( n331852 , n331851 );
buf ( n331853 , n331852 );
not ( n331854 , n331853 );
buf ( n331855 , n329773 );
not ( n41430 , n331855 );
and ( n331857 , n331854 , n41430 );
buf ( n331858 , n39560 );
not ( n41433 , n331858 );
buf ( n331860 , n41433 );
buf ( n331861 , n331860 );
nor ( n41436 , n331857 , n331861 );
buf ( n331863 , n41436 );
buf ( n331864 , n331863 );
nand ( n41439 , n41423 , n331864 );
buf ( n331866 , n41439 );
buf ( n331867 , n331866 );
nor ( n331868 , n41418 , n331867 );
buf ( n331869 , n331868 );
buf ( n331870 , n331869 );
nand ( n331871 , n41412 , n331870 );
buf ( n331872 , n331871 );
buf ( n331873 , n331872 );
and ( n331874 , n331873 , n331820 );
not ( n41449 , n331873 );
and ( n331876 , n41449 , n331816 );
nor ( n331877 , n331874 , n331876 );
buf ( n331878 , n331877 );
buf ( n331879 , n331860 );
buf ( n331880 , n329773 );
nor ( n41455 , n331879 , n331880 );
buf ( n41456 , n41455 );
buf ( n331883 , n41456 );
not ( n41458 , n331883 );
buf ( n41459 , n41458 );
buf ( n331886 , n41459 );
buf ( n331887 , n41456 );
buf ( n331888 , n330671 );
not ( n41463 , n331888 );
buf ( n41464 , n331721 );
buf ( n41465 , n329749 );
and ( n41466 , n41464 , n41465 );
buf ( n41467 , n41466 );
buf ( n331894 , n41467 );
not ( n41469 , n331894 );
buf ( n331896 , n331730 );
nor ( n41471 , n41469 , n331896 );
buf ( n331898 , n41471 );
buf ( n331899 , n331898 );
not ( n331900 , n331899 );
or ( n331901 , n41463 , n331900 );
buf ( n331902 , n331755 );
buf ( n331903 , n41467 );
and ( n41478 , n331902 , n331903 );
buf ( n331905 , n41478 );
buf ( n331906 , n331905 );
buf ( n331907 , n329749 );
not ( n41482 , n331907 );
buf ( n331909 , n331768 );
not ( n331910 , n331909 );
or ( n41485 , n41482 , n331910 );
buf ( n331912 , n331852 );
nand ( n331913 , n41485 , n331912 );
buf ( n331914 , n331913 );
buf ( n331915 , n331914 );
nor ( n41490 , n331906 , n331915 );
buf ( n331917 , n41490 );
buf ( n331918 , n331917 );
nand ( n41493 , n331901 , n331918 );
buf ( n41494 , n41493 );
buf ( n331921 , n41494 );
and ( n331922 , n331921 , n331887 );
not ( n41497 , n331921 );
and ( n331924 , n41497 , n331886 );
nor ( n41499 , n331922 , n331924 );
buf ( n331926 , n41499 );
buf ( n331927 , n330805 );
buf ( n331928 , n330918 );
nand ( n41503 , n331927 , n331928 );
buf ( n331930 , n41503 );
buf ( n331931 , n331930 );
buf ( n331932 , n331930 );
not ( n331933 , n331932 );
buf ( n331934 , n331933 );
buf ( n331935 , n331934 );
buf ( n331936 , n330705 );
buf ( n41511 , n329583 );
buf ( n331938 , n329527 );
nand ( n331939 , n41511 , n331938 );
buf ( n331940 , n331939 );
buf ( n331941 , n331940 );
not ( n331942 , n331941 );
buf ( n331943 , n331942 );
buf ( n331944 , n331943 );
and ( n331945 , n331936 , n331944 );
buf ( n331946 , n331945 );
not ( n41521 , n331946 );
not ( n331948 , n330671 );
or ( n41523 , n41521 , n331948 );
buf ( n331950 , n330001 );
not ( n41525 , n331950 );
buf ( n331952 , n41525 );
buf ( n331953 , n331952 );
not ( n41528 , n331953 );
buf ( n331955 , n331755 );
buf ( n331956 , n331721 );
nand ( n41531 , n331955 , n331956 );
buf ( n331958 , n41531 );
buf ( n331959 , n331958 );
not ( n41534 , n331959 );
or ( n41535 , n41528 , n41534 );
buf ( n331962 , n330006 );
not ( n331963 , n331962 );
buf ( n331964 , n331940 );
nor ( n331965 , n331963 , n331964 );
buf ( n331966 , n331965 );
buf ( n331967 , n331966 );
nand ( n331968 , n41535 , n331967 );
buf ( n331969 , n331968 );
buf ( n331970 , n331969 );
buf ( n331971 , n330748 );
buf ( n331972 , n329527 );
and ( n331973 , n331971 , n331972 );
buf ( n331974 , n329521 );
nor ( n331975 , n331973 , n331974 );
buf ( n331976 , n331975 );
buf ( n41551 , n331976 );
and ( n41552 , n331970 , n41551 );
buf ( n41553 , n41552 );
nand ( n331980 , n41523 , n41553 );
buf ( n331981 , n331980 );
and ( n331982 , n331981 , n331935 );
not ( n331983 , n331981 );
and ( n331984 , n331983 , n331931 );
nor ( n331985 , n331982 , n331984 );
buf ( n331986 , n331985 );
buf ( n331987 , n41299 );
buf ( n331988 , n329969 );
nand ( n41563 , n331987 , n331988 );
buf ( n41564 , n41563 );
buf ( n331991 , n41564 );
buf ( n331992 , n41564 );
not ( n41567 , n331992 );
buf ( n331994 , n41567 );
buf ( n331995 , n331994 );
buf ( n331996 , n330671 );
not ( n331997 , n331996 );
buf ( n331998 , n331730 );
buf ( n331999 , n39310 );
nor ( n41574 , n331998 , n331999 );
buf ( n332001 , n41574 );
buf ( n332002 , n332001 );
not ( n41577 , n332002 );
or ( n41578 , n331997 , n41577 );
buf ( n332005 , n331958 );
buf ( n332006 , n329963 );
and ( n41581 , n332005 , n332006 );
buf ( n332008 , n41581 );
buf ( n332009 , n332008 );
nand ( n332010 , n41578 , n332009 );
buf ( n332011 , n332010 );
buf ( n332012 , n332011 );
and ( n41587 , n332012 , n331995 );
not ( n332014 , n332012 );
and ( n41589 , n332014 , n331991 );
nor ( n41590 , n41587 , n41589 );
buf ( n332017 , n41590 );
buf ( n332018 , n39267 );
not ( n41593 , n332018 );
buf ( n332020 , n39531 );
nand ( n41595 , n41593 , n332020 );
buf ( n41596 , n41595 );
buf ( n332023 , n41596 );
buf ( n41598 , n41596 );
not ( n41599 , n41598 );
buf ( n41600 , n41599 );
buf ( n332027 , n41600 );
buf ( n332028 , n331730 );
and ( n332029 , n329717 , n329735 );
buf ( n332030 , n332029 );
buf ( n41605 , n329684 );
not ( n332032 , n41605 );
buf ( n332033 , n332032 );
buf ( n332034 , n332033 );
nand ( n332035 , n332030 , n332034 );
buf ( n332036 , n332035 );
buf ( n332037 , n332036 );
nor ( n332038 , n332028 , n332037 );
buf ( n332039 , n332038 );
buf ( n332040 , n332039 );
not ( n332041 , n332040 );
buf ( n332042 , n330671 );
not ( n41617 , n332042 );
or ( n332044 , n332041 , n41617 );
buf ( n332045 , n331761 );
buf ( n332046 , n332036 );
not ( n332047 , n332046 );
buf ( n332048 , n332047 );
buf ( n332049 , n332048 );
and ( n332050 , n332045 , n332049 );
buf ( n332051 , n332033 );
not ( n41626 , n332051 );
buf ( n332053 , n329943 );
not ( n332054 , n332053 );
or ( n41629 , n41626 , n332054 );
buf ( n332056 , n329950 );
nand ( n41631 , n41629 , n332056 );
buf ( n332058 , n41631 );
buf ( n332059 , n332058 );
nor ( n41634 , n332050 , n332059 );
buf ( n332061 , n41634 );
buf ( n332062 , n332061 );
nand ( n41637 , n332044 , n332062 );
buf ( n332064 , n41637 );
buf ( n332065 , n332064 );
and ( n332066 , n332065 , n332027 );
not ( n332067 , n332065 );
and ( n41642 , n332067 , n332023 );
nor ( n332069 , n332066 , n41642 );
buf ( n332070 , n332069 );
buf ( n332071 , n332033 );
buf ( n332072 , n329950 );
nand ( n332073 , n332071 , n332072 );
buf ( n332074 , n332073 );
buf ( n332075 , n332074 );
buf ( n332076 , n332074 );
not ( n332077 , n332076 );
buf ( n332078 , n332077 );
buf ( n332079 , n332078 );
and ( n332080 , n330699 , n332029 );
buf ( n332081 , n332080 );
not ( n41656 , n332081 );
buf ( n332083 , n330671 );
not ( n332084 , n332083 );
or ( n41659 , n41656 , n332084 );
buf ( n332086 , n331761 );
buf ( n332087 , n332029 );
and ( n41662 , n332086 , n332087 );
buf ( n332089 , n329943 );
nor ( n332090 , n41662 , n332089 );
buf ( n332091 , n332090 );
buf ( n332092 , n332091 );
nand ( n41667 , n41659 , n332092 );
buf ( n332094 , n41667 );
buf ( n332095 , n332094 );
and ( n41670 , n332095 , n332079 );
not ( n41671 , n332095 );
and ( n41672 , n41671 , n332075 );
nor ( n41673 , n41670 , n41672 );
buf ( n332100 , n41673 );
buf ( n332101 , n329630 );
not ( n41676 , n332101 );
buf ( n332103 , n41676 );
buf ( n332104 , n332103 );
buf ( n332105 , n39217 );
nand ( n41680 , n332104 , n332105 );
buf ( n332107 , n41680 );
buf ( n332108 , n332107 );
buf ( n332109 , n332107 );
not ( n41684 , n332109 );
buf ( n332111 , n41684 );
buf ( n332112 , n332111 );
buf ( n332113 , n39463 );
buf ( n332114 , n330696 );
not ( n41689 , n332114 );
buf ( n332116 , n41689 );
buf ( n332117 , n332116 );
and ( n41692 , n332113 , n332117 );
buf ( n332119 , n41692 );
buf ( n332120 , n332119 );
not ( n41695 , n332120 );
buf ( n332122 , n330671 );
not ( n41697 , n332122 );
or ( n41698 , n41695 , n41697 );
buf ( n332125 , n329892 );
buf ( n332126 , n329915 );
nor ( n41701 , n332125 , n332126 );
buf ( n332128 , n41701 );
buf ( n332129 , n332128 );
nand ( n41704 , n41698 , n332129 );
buf ( n332131 , n41704 );
buf ( n332132 , n332131 );
and ( n41707 , n332132 , n332112 );
not ( n41708 , n332132 );
and ( n41709 , n41708 , n332108 );
nor ( n332136 , n41707 , n41709 );
buf ( n332137 , n332136 );
buf ( n332138 , n329735 );
buf ( n332139 , n329929 );
nand ( n332140 , n332138 , n332139 );
buf ( n332141 , n332140 );
buf ( n332142 , n332141 );
buf ( n41717 , n332141 );
not ( n332144 , n41717 );
buf ( n332145 , n332144 );
buf ( n332146 , n332145 );
buf ( n332147 , n330671 );
not ( n332148 , n332147 );
buf ( n332149 , n330699 );
not ( n332150 , n332149 );
or ( n41725 , n332148 , n332150 );
buf ( n332152 , n331758 );
nand ( n332153 , n41725 , n332152 );
buf ( n332154 , n332153 );
buf ( n332155 , n332154 );
and ( n332156 , n332155 , n332146 );
not ( n41731 , n332155 );
and ( n41732 , n41731 , n332142 );
nor ( n332159 , n332156 , n41732 );
buf ( n332160 , n332159 );
buf ( n332161 , n39223 );
buf ( n332162 , n39197 );
nor ( n41737 , n332161 , n332162 );
buf ( n41738 , n41737 );
buf ( n41739 , n41738 );
not ( n41740 , n41739 );
buf ( n41741 , n41740 );
buf ( n332168 , n41741 );
buf ( n332169 , n41738 );
buf ( n332170 , n39463 );
buf ( n332171 , n332103 );
nand ( n41746 , n332170 , n332171 );
buf ( n332173 , n41746 );
buf ( n332174 , n332173 );
buf ( n332175 , n330696 );
nor ( n332176 , n332174 , n332175 );
buf ( n332177 , n332176 );
buf ( n332178 , n332177 );
not ( n41753 , n332178 );
buf ( n332180 , n330671 );
not ( n41755 , n332180 );
or ( n41756 , n41753 , n41755 );
buf ( n332183 , n329862 );
not ( n41758 , n332183 );
buf ( n332185 , n41758 );
buf ( n332186 , n332185 );
not ( n332187 , n332186 );
buf ( n332188 , n332173 );
not ( n41763 , n332188 );
and ( n332190 , n332187 , n41763 );
buf ( n332191 , n332103 );
not ( n332192 , n332191 );
buf ( n332193 , n329915 );
not ( n41768 , n332193 );
or ( n332195 , n332192 , n41768 );
buf ( n332196 , n39217 );
nand ( n41771 , n332195 , n332196 );
buf ( n332198 , n41771 );
buf ( n332199 , n332198 );
nor ( n41774 , n332190 , n332199 );
buf ( n41775 , n41774 );
buf ( n332202 , n41775 );
nand ( n332203 , n41756 , n332202 );
buf ( n332204 , n332203 );
buf ( n332205 , n332204 );
and ( n332206 , n332205 , n332169 );
not ( n332207 , n332205 );
and ( n332208 , n332207 , n332168 );
nor ( n332209 , n332206 , n332208 );
buf ( n332210 , n332209 );
buf ( n332211 , n39478 );
buf ( n41786 , n329912 );
nand ( n41787 , n332211 , n41786 );
buf ( n41788 , n41787 );
buf ( n332215 , n41788 );
buf ( n332216 , n41788 );
not ( n332217 , n332216 );
buf ( n332218 , n332217 );
buf ( n332219 , n332218 );
buf ( n332220 , n330696 );
buf ( n332221 , n329888 );
nor ( n332222 , n332220 , n332221 );
buf ( n332223 , n332222 );
buf ( n332224 , n332223 );
not ( n41799 , n332224 );
buf ( n332226 , n330671 );
not ( n41801 , n332226 );
or ( n41802 , n41799 , n41801 );
buf ( n332229 , n329888 );
not ( n41804 , n332229 );
buf ( n332231 , n41804 );
buf ( n332232 , n332231 );
not ( n332233 , n332232 );
buf ( n332234 , n329862 );
not ( n332235 , n332234 );
or ( n332236 , n332233 , n332235 );
buf ( n332237 , n329897 );
not ( n332238 , n332237 );
buf ( n332239 , n332238 );
buf ( n332240 , n332239 );
nand ( n332241 , n332236 , n332240 );
buf ( n332242 , n332241 );
buf ( n332243 , n332242 );
not ( n332244 , n332243 );
buf ( n332245 , n332244 );
buf ( n332246 , n332245 );
nand ( n332247 , n41802 , n332246 );
buf ( n332248 , n332247 );
buf ( n332249 , n332248 );
and ( n332250 , n332249 , n332219 );
not ( n41825 , n332249 );
and ( n332252 , n41825 , n332215 );
nor ( n332253 , n332250 , n332252 );
buf ( n332254 , n332253 );
buf ( n332255 , n332231 );
buf ( n41830 , n332239 );
nand ( n41831 , n332255 , n41830 );
buf ( n332258 , n41831 );
buf ( n41833 , n332258 );
buf ( n332260 , n332258 );
not ( n41835 , n332260 );
buf ( n41836 , n41835 );
buf ( n332263 , n41836 );
buf ( n332264 , n332116 );
not ( n332265 , n332264 );
buf ( n332266 , n330671 );
not ( n41841 , n332266 );
or ( n332268 , n332265 , n41841 );
buf ( n332269 , n332185 );
nand ( n41844 , n332268 , n332269 );
buf ( n41845 , n41844 );
buf ( n332272 , n41845 );
and ( n332273 , n332272 , n332263 );
not ( n332274 , n332272 );
and ( n41849 , n332274 , n41833 );
nor ( n332276 , n332273 , n41849 );
buf ( n332277 , n332276 );
buf ( n332278 , n329856 );
buf ( n332279 , n329791 );
nor ( n41854 , n332278 , n332279 );
buf ( n332281 , n41854 );
buf ( n332282 , n332281 );
not ( n41857 , n332282 );
buf ( n332284 , n41857 );
buf ( n332285 , n332284 );
buf ( n332286 , n332281 );
buf ( n332287 , n330693 );
buf ( n332288 , n39375 );
not ( n41863 , n332288 );
buf ( n332290 , n41863 );
buf ( n332291 , n332290 );
and ( n41866 , n332287 , n332291 );
buf ( n332293 , n41866 );
buf ( n332294 , n332293 );
not ( n332295 , n332294 );
buf ( n332296 , n330671 );
not ( n332297 , n332296 );
or ( n332298 , n332295 , n332297 );
buf ( n332299 , n329839 );
buf ( n332300 , n332290 );
and ( n332301 , n332299 , n332300 );
buf ( n332302 , n329850 );
nor ( n332303 , n332301 , n332302 );
buf ( n332304 , n332303 );
buf ( n332305 , n332304 );
nand ( n41880 , n332298 , n332305 );
buf ( n41881 , n41880 );
buf ( n41882 , n41881 );
and ( n332309 , n41882 , n332286 );
not ( n41884 , n41882 );
and ( n332311 , n41884 , n332285 );
nor ( n41886 , n332309 , n332311 );
buf ( n41887 , n41886 );
buf ( n41888 , n329850 );
buf ( n332315 , n39375 );
nor ( n332316 , n41888 , n332315 );
buf ( n332317 , n332316 );
buf ( n332318 , n332317 );
not ( n41893 , n332318 );
buf ( n332320 , n41893 );
buf ( n332321 , n332320 );
buf ( n332322 , n332317 );
buf ( n332323 , n330693 );
not ( n41898 , n332323 );
buf ( n332325 , n330671 );
not ( n332326 , n332325 );
or ( n41901 , n41898 , n332326 );
buf ( n332328 , n329839 );
not ( n41903 , n332328 );
buf ( n41904 , n41903 );
buf ( n332331 , n41904 );
nand ( n332332 , n41901 , n332331 );
buf ( n332333 , n332332 );
buf ( n332334 , n332333 );
and ( n41909 , n332334 , n332322 );
not ( n332336 , n332334 );
and ( n332337 , n332336 , n332321 );
nor ( n332338 , n41909 , n332337 );
buf ( n332339 , n332338 );
buf ( n332340 , n39396 );
not ( n332341 , n332340 );
buf ( n332342 , n329836 );
nand ( n41917 , n332341 , n332342 );
buf ( n332344 , n41917 );
buf ( n332345 , n332344 );
buf ( n332346 , n332344 );
not ( n332347 , n332346 );
buf ( n332348 , n332347 );
buf ( n332349 , n332348 );
buf ( n332350 , n330689 );
not ( n41925 , n332350 );
buf ( n332352 , n41925 );
buf ( n332353 , n332352 );
not ( n41928 , n332353 );
buf ( n332355 , n330671 );
not ( n332356 , n332355 );
or ( n41931 , n41928 , n332356 );
buf ( n332358 , n329830 );
nand ( n41933 , n41931 , n332358 );
buf ( n332360 , n41933 );
buf ( n332361 , n332360 );
and ( n41936 , n332361 , n332349 );
not ( n41937 , n332361 );
and ( n41938 , n41937 , n332345 );
nor ( n41939 , n41936 , n41938 );
buf ( n332366 , n41939 );
buf ( n332367 , n329717 );
buf ( n332368 , n329940 );
nand ( n41943 , n332367 , n332368 );
buf ( n332370 , n41943 );
buf ( n332371 , n332370 );
buf ( n332372 , n332370 );
not ( n41947 , n332372 );
buf ( n332374 , n41947 );
buf ( n332375 , n332374 );
buf ( n332376 , n329735 );
not ( n41951 , n332376 );
buf ( n332378 , n331730 );
nor ( n41953 , n41951 , n332378 );
buf ( n332380 , n41953 );
buf ( n332381 , n332380 );
not ( n332382 , n332381 );
buf ( n332383 , n330671 );
not ( n41958 , n332383 );
or ( n332385 , n332382 , n41958 );
buf ( n332386 , n329735 );
not ( n41961 , n332386 );
buf ( n332388 , n331755 );
not ( n332389 , n332388 );
or ( n332390 , n41961 , n332389 );
buf ( n332391 , n329929 );
nand ( n41966 , n332390 , n332391 );
buf ( n41967 , n41966 );
buf ( n41968 , n41967 );
not ( n41969 , n41968 );
buf ( n41970 , n41969 );
buf ( n332397 , n41970 );
nand ( n41972 , n332385 , n332397 );
buf ( n332399 , n41972 );
buf ( n332400 , n332399 );
and ( n41975 , n332400 , n332375 );
not ( n41976 , n332400 );
and ( n332403 , n41976 , n332371 );
nor ( n41978 , n41975 , n332403 );
buf ( n332405 , n41978 );
buf ( n332406 , n39636 );
not ( n41981 , n332406 );
buf ( n332408 , n330073 );
nand ( n332409 , n41981 , n332408 );
buf ( n332410 , n332409 );
buf ( n332411 , n332410 );
buf ( n332412 , n332410 );
not ( n332413 , n332412 );
buf ( n332414 , n332413 );
buf ( n332415 , n332414 );
buf ( n332416 , n39745 );
not ( n332417 , n332416 );
buf ( n41992 , n330331 );
nand ( n41993 , n332417 , n41992 );
buf ( n41994 , n41993 );
buf ( n41995 , n41994 );
buf ( n332422 , n39931 );
not ( n332423 , n332422 );
buf ( n332424 , n332423 );
buf ( n332425 , n332424 );
buf ( n332426 , n330658 );
buf ( n332427 , n39745 );
nor ( n42002 , n332426 , n332427 );
buf ( n332429 , n42002 );
buf ( n332430 , n332429 );
nand ( n42005 , n332425 , n332430 );
buf ( n332432 , n42005 );
buf ( n332433 , n332432 );
buf ( n332434 , n330067 );
nand ( n42009 , n41995 , n332433 , n332434 );
buf ( n332436 , n42009 );
buf ( n332437 , n332436 );
and ( n42012 , n332437 , n332415 );
not ( n332439 , n332437 );
and ( n42014 , n332439 , n332411 );
nor ( n42015 , n42012 , n42014 );
buf ( n332442 , n42015 );
buf ( n332443 , n330110 );
buf ( n332444 , n39669 );
nor ( n332445 , n332443 , n332444 );
buf ( n332446 , n332445 );
buf ( n332447 , n332446 );
not ( n332448 , n332447 );
buf ( n332449 , n332448 );
buf ( n332450 , n332449 );
buf ( n332451 , n332446 );
not ( n42026 , n330174 );
not ( n332453 , n330331 );
or ( n332454 , n42026 , n332453 );
buf ( n332455 , n330174 );
not ( n42030 , n332455 );
buf ( n332457 , n42030 );
buf ( n332458 , n332457 );
buf ( n332459 , n330658 );
nor ( n332460 , n332458 , n332459 );
buf ( n332461 , n332460 );
and ( n42036 , n332424 , n332461 );
nor ( n42037 , n42036 , n330076 );
nand ( n42038 , n332454 , n42037 );
buf ( n332465 , n42038 );
and ( n42040 , n332465 , n332451 );
not ( n42041 , n332465 );
and ( n332468 , n42041 , n332450 );
nor ( n332469 , n42040 , n332468 );
buf ( n332470 , n332469 );
buf ( n332471 , n330134 );
buf ( n332472 , n330141 );
nand ( n42047 , n332471 , n332472 );
buf ( n332474 , n42047 );
buf ( n332475 , n332474 );
buf ( n332476 , n332474 );
not ( n42051 , n332476 );
buf ( n332478 , n42051 );
buf ( n332479 , n332478 );
buf ( n332480 , n330177 );
not ( n42055 , n332480 );
buf ( n332482 , n42055 );
buf ( n332483 , n332482 );
buf ( n332484 , n330030 );
nor ( n42059 , n332483 , n332484 );
buf ( n332486 , n42059 );
buf ( n332487 , n332486 );
buf ( n332488 , n330331 );
nand ( n42063 , n332487 , n332488 );
buf ( n332490 , n42063 );
buf ( n332491 , n332490 );
buf ( n332492 , n332486 );
buf ( n332493 , n330661 );
nand ( n42068 , n332492 , n332493 );
buf ( n332495 , n42068 );
buf ( n332496 , n332495 );
buf ( n332497 , n39696 );
not ( n42072 , n332497 );
buf ( n332499 , n42072 );
buf ( n332500 , n332499 );
buf ( n332501 , n330030 );
not ( n42076 , n332501 );
buf ( n332503 , n42076 );
buf ( n332504 , n332503 );
nand ( n42079 , n332500 , n332504 );
buf ( n332506 , n42079 );
buf ( n332507 , n332506 );
buf ( n332508 , n330129 );
not ( n42083 , n332508 );
buf ( n332510 , n42083 );
buf ( n332511 , n332510 );
nand ( n42086 , n332491 , n332496 , n332507 , n332511 );
buf ( n332513 , n42086 );
buf ( n332514 , n332513 );
and ( n42089 , n332514 , n332479 );
not ( n42090 , n332514 );
and ( n42091 , n42090 , n332475 );
nor ( n42092 , n42089 , n42091 );
buf ( n332519 , n42092 );
buf ( n332520 , n330051 );
not ( n42095 , n332520 );
buf ( n332522 , n42095 );
buf ( n332523 , n332522 );
buf ( n332524 , n39726 );
nand ( n42099 , n332523 , n332524 );
buf ( n332526 , n42099 );
buf ( n332527 , n332526 );
buf ( n332528 , n332526 );
not ( n42103 , n332528 );
buf ( n332530 , n42103 );
buf ( n332531 , n332530 );
buf ( n332532 , n330177 );
buf ( n332533 , n330033 );
and ( n42108 , n332532 , n332533 );
buf ( n332535 , n42108 );
buf ( n332536 , n332535 );
buf ( n332537 , n330661 );
nand ( n42112 , n332536 , n332537 );
buf ( n332539 , n42112 );
buf ( n332540 , n332539 );
buf ( n332541 , n332535 );
buf ( n332542 , n330331 );
nand ( n42117 , n332541 , n332542 );
buf ( n332544 , n42117 );
buf ( n332545 , n332544 );
buf ( n332546 , n332499 );
buf ( n332547 , n330033 );
and ( n42122 , n332546 , n332547 );
buf ( n332549 , n330144 );
nor ( n42124 , n42122 , n332549 );
buf ( n332551 , n42124 );
buf ( n332552 , n332551 );
nand ( n42127 , n332540 , n332545 , n332552 );
buf ( n332554 , n42127 );
buf ( n332555 , n332554 );
and ( n42130 , n332555 , n332531 );
not ( n42131 , n332555 );
and ( n42132 , n42131 , n332527 );
nor ( n42133 , n42130 , n42132 );
buf ( n332560 , n42133 );
buf ( n332561 , n330159 );
buf ( n332562 , n330044 );
nor ( n42137 , n332561 , n332562 );
buf ( n332564 , n42137 );
buf ( n332565 , n332564 );
not ( n42140 , n332565 );
buf ( n332567 , n42140 );
buf ( n332568 , n332567 );
buf ( n332569 , n332564 );
buf ( n332570 , n330331 );
not ( n42145 , n332570 );
buf ( n332572 , n42145 );
buf ( n332573 , n332572 );
not ( n42148 , n332573 );
buf ( n332575 , n330033 );
buf ( n332576 , n332522 );
nand ( n42151 , n332575 , n332576 );
buf ( n332578 , n42151 );
buf ( n332579 , n332578 );
buf ( n332580 , n332482 );
nor ( n42155 , n332579 , n332580 );
buf ( n332582 , n42155 );
buf ( n332583 , n332582 );
nand ( n42158 , n42148 , n332583 );
buf ( n332585 , n42158 );
buf ( n332586 , n332585 );
buf ( n332587 , n332582 );
buf ( n332588 , n330661 );
nand ( n42163 , n332587 , n332588 );
buf ( n332590 , n42163 );
buf ( n332591 , n332590 );
not ( n42166 , n332578 );
not ( n42167 , n39696 );
and ( n42168 , n42166 , n42167 );
buf ( n332595 , n332522 );
not ( n42170 , n332595 );
buf ( n332597 , n330144 );
not ( n42172 , n332597 );
or ( n42173 , n42170 , n42172 );
buf ( n332600 , n39726 );
nand ( n42175 , n42173 , n332600 );
buf ( n332602 , n42175 );
nor ( n42177 , n42168 , n332602 );
buf ( n332604 , n42177 );
nand ( n42179 , n332586 , n332591 , n332604 );
buf ( n332606 , n42179 );
buf ( n332607 , n332606 );
and ( n42182 , n332607 , n332569 );
not ( n42183 , n332607 );
and ( n42184 , n42183 , n332568 );
nor ( n42185 , n42182 , n42184 );
buf ( n332612 , n42185 );
buf ( n332613 , n332352 );
buf ( n332614 , n329830 );
nand ( n42189 , n332613 , n332614 );
buf ( n332616 , n42189 );
buf ( n332617 , n332616 );
buf ( n332618 , n330671 );
buf ( n332619 , n332616 );
buf ( n332620 , n330671 );
not ( n42195 , n332617 );
not ( n42196 , n332618 );
or ( n42197 , n42195 , n42196 );
or ( n42198 , n332619 , n332620 );
nand ( n42199 , n42197 , n42198 );
buf ( n332626 , n42199 );
buf ( n332627 , n332503 );
buf ( n332628 , n332510 );
nand ( n42203 , n332627 , n332628 );
buf ( n332630 , n42203 );
buf ( n332631 , n332630 );
buf ( n332632 , n332630 );
not ( n42207 , n332632 );
buf ( n332634 , n42207 );
buf ( n332635 , n332634 );
buf ( n332636 , n330177 );
buf ( n332637 , n330331 );
nand ( n42212 , n332636 , n332637 );
buf ( n332639 , n42212 );
buf ( n332640 , n332639 );
buf ( n332641 , n332424 );
buf ( n332642 , n330177 );
buf ( n332643 , n330658 );
not ( n42218 , n332643 );
buf ( n332645 , n42218 );
buf ( n332646 , n332645 );
nand ( n42221 , n332641 , n332642 , n332646 );
buf ( n332648 , n42221 );
buf ( n332649 , n332648 );
buf ( n332650 , n39696 );
nand ( n42225 , n332640 , n332649 , n332650 );
buf ( n332652 , n42225 );
buf ( n332653 , n332652 );
and ( n42228 , n332653 , n332635 );
not ( n42229 , n332653 );
and ( n42230 , n42229 , n332631 );
nor ( n42231 , n42228 , n42230 );
buf ( n332658 , n42231 );
buf ( n332659 , n330116 );
buf ( n332660 , n330088 );
nor ( n42235 , n332659 , n332660 );
buf ( n332662 , n42235 );
buf ( n332663 , n332662 );
not ( n42238 , n332663 );
buf ( n332665 , n42238 );
buf ( n332666 , n332665 );
buf ( n332667 , n332662 );
buf ( n332668 , n330331 );
buf ( n332669 , n332457 );
buf ( n332670 , n39669 );
nor ( n42245 , n332669 , n332670 );
buf ( n332672 , n42245 );
buf ( n332673 , n332672 );
nand ( n42248 , n332668 , n332673 );
buf ( n332675 , n42248 );
buf ( n332676 , n332675 );
buf ( n332677 , n332424 );
buf ( n332678 , n332645 );
buf ( n332679 , n332672 );
nand ( n42254 , n332677 , n332678 , n332679 );
buf ( n332681 , n42254 );
buf ( n332682 , n332681 );
not ( n42257 , n330076 );
buf ( n332684 , n42257 );
not ( n42259 , n332684 );
buf ( n332686 , n39669 );
not ( n42261 , n332686 );
and ( n42262 , n42259 , n42261 );
buf ( n332689 , n330110 );
nor ( n42264 , n42262 , n332689 );
buf ( n332691 , n42264 );
buf ( n332692 , n332691 );
nand ( n42267 , n332676 , n332682 , n332692 );
buf ( n332694 , n42267 );
buf ( n332695 , n332694 );
and ( n42270 , n332695 , n332667 );
not ( n42271 , n332695 );
and ( n42272 , n42271 , n332666 );
nor ( n42273 , n42270 , n42272 );
buf ( n332700 , n42273 );
buf ( n332701 , n39745 );
not ( n42276 , n332701 );
buf ( n332703 , n330067 );
nand ( n42278 , n42276 , n332703 );
buf ( n332705 , n42278 );
buf ( n332706 , n332705 );
buf ( n332707 , n332705 );
not ( n42282 , n332707 );
buf ( n332709 , n42282 );
buf ( n332710 , n332709 );
buf ( n332711 , n330661 );
not ( n332712 , n332711 );
buf ( n332713 , n332572 );
nand ( n332714 , n332712 , n332713 );
buf ( n332715 , n332714 );
buf ( n332716 , n332715 );
and ( n332717 , n332716 , n332710 );
not ( n42292 , n332716 );
and ( n332719 , n42292 , n332706 );
nor ( n332720 , n332717 , n332719 );
buf ( n332721 , n332720 );
buf ( n332722 , n330322 );
buf ( n42297 , n39800 );
not ( n42298 , n42297 );
buf ( n42299 , n42298 );
buf ( n332726 , n42299 );
and ( n42301 , n332722 , n332726 );
buf ( n332728 , n42301 );
buf ( n42303 , n332728 );
buf ( n42304 , n330352 );
buf ( n42305 , n330658 );
nor ( n42306 , n42304 , n42305 );
buf ( n332733 , n42306 );
buf ( n42308 , n332733 );
nand ( n42309 , n42303 , n42308 );
buf ( n42310 , n42309 );
buf ( n332737 , n330349 );
buf ( n332738 , n332645 );
buf ( n332739 , n330269 );
not ( n332740 , n332739 );
buf ( n332741 , n332740 );
buf ( n332742 , n332741 );
not ( n332743 , n332737 );
not ( n42318 , n332738 );
or ( n332745 , n332743 , n42318 );
nand ( n42320 , n332745 , n332742 );
buf ( n332747 , n42320 );
buf ( n332748 , n330658 );
buf ( n332749 , n330346 );
not ( n42324 , n332749 );
buf ( n332751 , n42324 );
buf ( n332752 , n332751 );
buf ( n332753 , n330260 );
and ( n332754 , n332752 , n332753 );
buf ( n332755 , n332754 );
buf ( n332756 , n332755 );
buf ( n332757 , n332755 );
buf ( n332758 , n330658 );
not ( n42333 , n332748 );
not ( n42334 , n332756 );
or ( n332761 , n42333 , n42334 );
or ( n332762 , n332757 , n332758 );
nand ( n42337 , n332761 , n332762 );
buf ( n332764 , n42337 );
or ( n42339 , n330652 , n330609 );
and ( n332766 , n42339 , n330430 );
nor ( n332767 , n332766 , n330402 );
buf ( n332768 , n332767 );
buf ( n332769 , n330377 );
buf ( n332770 , n330408 );
and ( n42345 , n332769 , n332770 );
buf ( n42346 , n42345 );
buf ( n42347 , n42346 );
buf ( n332774 , n42346 );
buf ( n332775 , n332767 );
not ( n332776 , n332768 );
not ( n332777 , n42347 );
or ( n42352 , n332776 , n332777 );
or ( n332779 , n332774 , n332775 );
nand ( n332780 , n42352 , n332779 );
buf ( n332781 , n332780 );
buf ( n332782 , n332751 );
buf ( n332783 , n332645 );
buf ( n332784 , n330260 );
not ( n332785 , n332782 );
not ( n42360 , n332783 );
or ( n42361 , n332785 , n42360 );
nand ( n332788 , n42361 , n332784 );
buf ( n332789 , n332788 );
buf ( n42364 , n330349 );
buf ( n42365 , n330289 );
and ( n42366 , n42364 , n42365 );
buf ( n332793 , n42366 );
buf ( n332794 , n332793 );
buf ( n332795 , n332645 );
buf ( n332796 , n330269 );
buf ( n332797 , n330289 );
and ( n42372 , n332796 , n332797 );
buf ( n332799 , n39874 );
nor ( n332800 , n42372 , n332799 );
buf ( n332801 , n332800 );
buf ( n332802 , n332801 );
not ( n332803 , n332794 );
not ( n42378 , n332795 );
or ( n332805 , n332803 , n42378 );
nand ( n42380 , n332805 , n332802 );
buf ( n332807 , n42380 );
buf ( n42382 , n332645 );
buf ( n332809 , n330352 );
buf ( n332810 , n330318 );
nor ( n42385 , n332809 , n332810 );
buf ( n332812 , n42385 );
buf ( n332813 , n332812 );
nand ( n42388 , n42382 , n332813 );
buf ( n332815 , n42388 );
buf ( n332816 , n330606 );
buf ( n332817 , n330467 );
or ( n42392 , n332816 , n332817 );
buf ( n332819 , n330619 );
nand ( n42394 , n42392 , n332819 );
buf ( n332821 , n42394 );
buf ( n332822 , n332821 );
buf ( n332823 , n330460 );
not ( n42398 , n332823 );
buf ( n332825 , n330625 );
nand ( n42400 , n42398 , n332825 );
buf ( n332827 , n42400 );
buf ( n332828 , n332827 );
buf ( n332829 , n332827 );
buf ( n332830 , n332821 );
not ( n42405 , n332822 );
not ( n332832 , n332828 );
or ( n42407 , n42405 , n332832 );
or ( n42408 , n332829 , n332830 );
nand ( n42409 , n42407 , n42408 );
buf ( n332836 , n42409 );
buf ( n42411 , n330652 );
buf ( n42412 , n330427 );
not ( n332839 , n42412 );
buf ( n332840 , n332839 );
buf ( n332841 , n332840 );
nand ( n332842 , n42411 , n332841 );
buf ( n332843 , n332842 );
buf ( n332844 , n332843 );
buf ( n332845 , n330473 );
buf ( n332846 , n330427 );
nor ( n332847 , n332845 , n332846 );
buf ( n332848 , n332847 );
buf ( n332849 , n332848 );
buf ( n332850 , n330606 );
not ( n42425 , n332850 );
buf ( n332852 , n42425 );
buf ( n332853 , n332852 );
nand ( n42428 , n332849 , n332853 );
buf ( n42429 , n42428 );
buf ( n332856 , n42429 );
buf ( n332857 , n330393 );
nand ( n332858 , n332844 , n332856 , n332857 );
buf ( n332859 , n332858 );
buf ( n332860 , n332859 );
buf ( n332861 , n330388 );
not ( n332862 , n332861 );
buf ( n42437 , n330399 );
nand ( n42438 , n332862 , n42437 );
buf ( n42439 , n42438 );
buf ( n332866 , n42439 );
buf ( n332867 , n42439 );
buf ( n332868 , n332859 );
not ( n332869 , n332860 );
not ( n42444 , n332866 );
or ( n42445 , n332869 , n42444 );
or ( n42446 , n332867 , n332868 );
nand ( n42447 , n42445 , n42446 );
buf ( n332874 , n42447 );
buf ( n332875 , n332840 );
buf ( n332876 , n330393 );
nand ( n42451 , n332875 , n332876 );
buf ( n332878 , n42451 );
buf ( n332879 , n332878 );
buf ( n332880 , n330609 );
buf ( n332881 , n330652 );
or ( n42456 , n332880 , n332881 );
buf ( n332883 , n42456 );
buf ( n332884 , n332883 );
buf ( n332885 , n332878 );
buf ( n332886 , n332883 );
not ( n42461 , n332879 );
not ( n42462 , n332884 );
or ( n42463 , n42461 , n42462 );
or ( n42464 , n332885 , n332886 );
nand ( n42465 , n42463 , n42464 );
buf ( n332892 , n42465 );
buf ( n332893 , n332852 );
buf ( n332894 , n330470 );
buf ( n42469 , n330445 );
not ( n332896 , n42469 );
buf ( n332897 , n332896 );
buf ( n332898 , n332897 );
and ( n332899 , n332893 , n332894 , n332898 );
buf ( n332900 , n330628 );
not ( n332901 , n332900 );
buf ( n332902 , n332897 );
not ( n332903 , n332902 );
or ( n332904 , n332901 , n332903 );
buf ( n332905 , n330639 );
nand ( n332906 , n332904 , n332905 );
buf ( n332907 , n332906 );
buf ( n332908 , n332907 );
nor ( n42483 , n332899 , n332908 );
buf ( n332910 , n42483 );
buf ( n332911 , n332910 );
buf ( n332912 , n330646 );
buf ( n332913 , n330440 );
nor ( n332914 , n332912 , n332913 );
buf ( n332915 , n332914 );
buf ( n42490 , n332915 );
buf ( n332917 , n332915 );
buf ( n332918 , n332910 );
not ( n332919 , n332911 );
not ( n332920 , n42490 );
or ( n42495 , n332919 , n332920 );
or ( n332922 , n332917 , n332918 );
nand ( n42497 , n42495 , n332922 );
buf ( n332924 , n42497 );
buf ( n332925 , n332852 );
buf ( n332926 , n330470 );
and ( n332927 , n332925 , n332926 );
buf ( n332928 , n330628 );
nor ( n42503 , n332927 , n332928 );
buf ( n332930 , n42503 );
buf ( n332931 , n332930 );
buf ( n332932 , n332897 );
buf ( n332933 , n330639 );
and ( n42508 , n332932 , n332933 );
buf ( n42509 , n42508 );
buf ( n332936 , n42509 );
buf ( n332937 , n42509 );
buf ( n332938 , n332930 );
not ( n332939 , n332931 );
not ( n42514 , n332936 );
or ( n332941 , n332939 , n42514 );
or ( n332942 , n332937 , n332938 );
nand ( n42517 , n332941 , n332942 );
buf ( n42518 , n42517 );
buf ( n332945 , n332852 );
buf ( n332946 , n330467 );
not ( n332947 , n332946 );
buf ( n332948 , n330619 );
nand ( n42523 , n332947 , n332948 );
buf ( n332950 , n42523 );
buf ( n332951 , n332950 );
buf ( n332952 , n332950 );
buf ( n332953 , n332852 );
not ( n42528 , n332945 );
not ( n332955 , n332951 );
or ( n332956 , n42528 , n332955 );
or ( n42531 , n332952 , n332953 );
nand ( n332958 , n332956 , n42531 );
buf ( n332959 , n332958 );
buf ( n332960 , n330599 );
buf ( n332961 , n330505 );
nor ( n332962 , n332960 , n332961 );
buf ( n332963 , n332962 );
buf ( n332964 , n332963 );
buf ( n332965 , n330478 );
not ( n42540 , n332965 );
buf ( n42541 , n42540 );
buf ( n332968 , n42541 );
buf ( n332969 , n330511 );
and ( n42544 , n332968 , n332969 );
buf ( n332971 , n42544 );
buf ( n332972 , n332971 );
buf ( n332973 , n332971 );
buf ( n332974 , n332963 );
not ( n42549 , n332964 );
not ( n42550 , n332972 );
or ( n332977 , n42549 , n42550 );
or ( n42552 , n332973 , n332974 );
nand ( n42553 , n332977 , n42552 );
buf ( n332980 , n42553 );
buf ( n332981 , n330491 );
not ( n42556 , n332981 );
buf ( n332983 , n40076 );
nand ( n42558 , n42556 , n332983 );
buf ( n332985 , n42558 );
buf ( n332986 , n332985 );
buf ( n332987 , n330595 );
buf ( n332988 , n330496 );
nand ( n42563 , n332987 , n332988 );
buf ( n332990 , n42563 );
buf ( n332991 , n332990 );
buf ( n332992 , n332990 );
buf ( n332993 , n332985 );
not ( n332994 , n332986 );
not ( n332995 , n332991 );
or ( n42570 , n332994 , n332995 );
or ( n332997 , n332992 , n332993 );
nand ( n332998 , n42570 , n332997 );
buf ( n332999 , n332998 );
buf ( n333000 , n330529 );
buf ( n42575 , n330496 );
nand ( n42576 , n333000 , n42575 );
buf ( n42577 , n42576 );
buf ( n333004 , n42577 );
buf ( n333005 , n330592 );
buf ( n333006 , n42577 );
buf ( n333007 , n330592 );
not ( n333008 , n333004 );
not ( n42583 , n333005 );
or ( n333010 , n333008 , n42583 );
or ( n333011 , n333006 , n333007 );
nand ( n42586 , n333010 , n333011 );
buf ( n333013 , n42586 );
buf ( n333014 , n330545 );
not ( n42589 , n333014 );
buf ( n333016 , n330589 );
nand ( n42591 , n42589 , n333016 );
buf ( n333018 , n42591 );
buf ( n333019 , n333018 );
buf ( n333020 , n330576 );
buf ( n333021 , n330583 );
nand ( n42596 , n333020 , n333021 );
buf ( n42597 , n42596 );
buf ( n333024 , n42597 );
buf ( n333025 , n42597 );
buf ( n333026 , n333018 );
not ( n42601 , n333019 );
not ( n42602 , n333024 );
or ( n333029 , n42601 , n42602 );
or ( n333030 , n333025 , n333026 );
nand ( n42605 , n333029 , n333030 );
buf ( n333032 , n42605 );
buf ( n333033 , n40127 );
buf ( n333034 , n330583 );
nand ( n333035 , n333033 , n333034 );
buf ( n333036 , n333035 );
buf ( n333037 , n333036 );
buf ( n333038 , n330573 );
buf ( n333039 , n330573 );
buf ( n333040 , n333036 );
not ( n333041 , n333037 );
not ( n42616 , n333038 );
or ( n333043 , n333041 , n42616 );
or ( n333044 , n333039 , n333040 );
nand ( n42619 , n333043 , n333044 );
buf ( n42620 , n42619 );
xor ( n333047 , n330555 , n330567 );
xor ( n42622 , n333047 , n330569 );
buf ( n333049 , n42622 );
buf ( n333050 , n330312 );
buf ( n333051 , n330318 );
not ( n333052 , n333051 );
buf ( n333053 , n333052 );
buf ( n333054 , n333053 );
nand ( n42629 , n333050 , n333054 );
buf ( n333056 , n42629 );
buf ( n333057 , n330312 );
buf ( n333058 , n332728 );
nand ( n42633 , n333057 , n333058 );
buf ( n333060 , n42633 );
buf ( n333061 , n330212 );
buf ( n333062 , n42299 );
buf ( n333063 , n330232 );
not ( n42638 , n333063 );
buf ( n42639 , n42638 );
buf ( n333066 , n42639 );
and ( n42641 , n333061 , n333062 );
nor ( n42642 , n42641 , n333066 );
buf ( n333069 , n42642 );
xor ( n42644 , n330556 , n330564 );
buf ( n333071 , n42644 );
buf ( n42646 , n333053 );
buf ( n333073 , n39776 );
not ( n42648 , n333073 );
buf ( n42649 , n42648 );
buf ( n333076 , n42649 );
nand ( n42651 , n42646 , n333076 );
buf ( n333078 , n42651 );
buf ( n333079 , n330365 );
buf ( n333080 , n330415 );
not ( n42655 , n333079 );
nand ( n42656 , n42655 , n333080 );
buf ( n333083 , n42656 );
buf ( n333084 , n39819 );
buf ( n333085 , n39840 );
not ( n42660 , n333084 );
nand ( n42661 , n42660 , n333085 );
buf ( n333088 , n42661 );
buf ( n333089 , n330511 );
not ( n42664 , n333089 );
buf ( n333091 , n42664 );
buf ( n333092 , n332733 );
buf ( n333093 , n330312 );
or ( n42668 , n333092 , n333093 );
buf ( n333095 , n42668 );
buf ( n333096 , n333095 );
buf ( n333097 , n333078 );
xnor ( n42672 , n333096 , n333097 );
buf ( n333099 , n42672 );
buf ( n333100 , n332747 );
buf ( n333101 , n39874 );
not ( n42676 , n333101 );
buf ( n333103 , n330289 );
nand ( n42678 , n42676 , n333103 );
buf ( n333105 , n42678 );
buf ( n333106 , n333105 );
xnor ( n42681 , n333100 , n333106 );
buf ( n333108 , n42681 );
buf ( n333109 , n332789 );
buf ( n333110 , n333088 );
xnor ( n42685 , n333109 , n333110 );
buf ( n333112 , n42685 );
buf ( n333113 , n330322 );
buf ( n333114 , n330352 );
not ( n42689 , n333113 );
nor ( n42690 , n42689 , n333114 );
buf ( n333117 , n42690 );
buf ( n333118 , n332807 );
buf ( n333119 , n330283 );
not ( n42694 , n333119 );
buf ( n333121 , n330306 );
nor ( n42696 , n42694 , n333121 );
buf ( n333123 , n42696 );
buf ( n333124 , n333123 );
xor ( n42699 , n333118 , n333124 );
buf ( n333126 , n42699 );
buf ( n333127 , n323081 );
buf ( n333128 , n328621 );
not ( n42703 , n309907 );
not ( n42704 , n308644 );
or ( n42705 , n42703 , n42704 );
nand ( n42706 , n42705 , n307238 );
not ( n42707 , n16774 );
and ( n42708 , n42707 , n16812 );
and ( n42709 , n42706 , n42708 );
not ( n42710 , n42706 );
not ( n42711 , n42708 );
and ( n42712 , n42710 , n42711 );
nor ( n42713 , n42709 , n42712 );
buf ( n333140 , n42713 );
xor ( n42715 , n333127 , n333128 );
xor ( n42716 , n42715 , n333140 );
buf ( n333143 , n42716 );
xor ( n42718 , n333127 , n333128 );
and ( n42719 , n42718 , n333140 );
and ( n42720 , n333127 , n333128 );
or ( n42721 , n42719 , n42720 );
buf ( n333148 , n42721 );
buf ( n333149 , n329243 );
buf ( n333150 , n32738 );
xnor ( n42725 , n19460 , n18220 );
buf ( n333152 , n42725 );
xor ( n42727 , n333149 , n333150 );
xor ( n42728 , n42727 , n333152 );
buf ( n333155 , n42728 );
xor ( n42730 , n333149 , n333150 );
and ( n42731 , n42730 , n333152 );
and ( n42732 , n333149 , n333150 );
or ( n42733 , n42731 , n42732 );
buf ( n333160 , n42733 );
buf ( n333161 , n323181 );
buf ( n333162 , n323066 );
not ( n42737 , n309874 );
not ( n42738 , n308644 );
or ( n42739 , n42737 , n42738 );
nand ( n42740 , n42739 , n309847 );
not ( n42741 , n16820 );
nand ( n42742 , n42741 , n16769 );
not ( n42743 , n42742 );
and ( n42744 , n42740 , n42743 );
not ( n42745 , n42740 );
and ( n42746 , n42745 , n42742 );
nor ( n42747 , n42744 , n42746 );
buf ( n333174 , n42747 );
xor ( n42749 , n333161 , n333162 );
xor ( n42750 , n42749 , n333174 );
buf ( n333177 , n42750 );
xor ( n42752 , n333161 , n333162 );
and ( n42753 , n42752 , n333174 );
and ( n42754 , n333161 , n333162 );
or ( n42755 , n42753 , n42754 );
buf ( n333182 , n42755 );
buf ( n333183 , n323053 );
buf ( n333184 , n38747 );
buf ( n333185 , n307889 );
xor ( n42760 , n333183 , n333184 );
xor ( n42761 , n42760 , n333185 );
buf ( n333188 , n42761 );
xor ( n42763 , n333183 , n333184 );
and ( n42764 , n42763 , n333185 );
and ( n42765 , n333183 , n333184 );
or ( n42766 , n42764 , n42765 );
buf ( n333193 , n42766 );
buf ( n333194 , n32858 );
buf ( n333195 , n38706 );
not ( n42770 , n17049 );
nand ( n42771 , n17464 , n17467 , n307466 );
nand ( n42772 , n17464 , n307250 );
nand ( n42773 , n42770 , n42771 , n42772 );
and ( n42774 , n42773 , n309882 );
not ( n42775 , n42773 );
and ( n42776 , n42775 , n19453 );
nor ( n42777 , n42774 , n42776 );
buf ( n333204 , n42777 );
xor ( n42779 , n333194 , n333195 );
xor ( n42780 , n42779 , n333204 );
buf ( n333207 , n42780 );
xor ( n42782 , n333194 , n333195 );
and ( n42783 , n42782 , n333204 );
and ( n42784 , n333194 , n333195 );
or ( n42785 , n42783 , n42784 );
buf ( n333212 , n42785 );
buf ( n333213 , n329109 );
buf ( n333214 , n295150 );
buf ( n333215 , n307904 );
xor ( n42790 , n333213 , n333214 );
xor ( n42791 , n42790 , n333215 );
buf ( n333218 , n42791 );
xor ( n42793 , n333213 , n333214 );
and ( n42794 , n42793 , n333215 );
and ( n42795 , n333213 , n333214 );
or ( n42796 , n42794 , n42795 );
buf ( n333223 , n42796 );
buf ( n333224 , n4641 );
buf ( n333225 , n32912 );
buf ( n333226 , n307869 );
xor ( n42801 , n333224 , n333225 );
xor ( n42802 , n42801 , n333226 );
buf ( n333229 , n42802 );
xor ( n42804 , n333224 , n333225 );
and ( n42805 , n42804 , n333226 );
and ( n42806 , n333224 , n333225 );
or ( n42807 , n42805 , n42806 );
buf ( n333234 , n42807 );
buf ( n333235 , n323377 );
buf ( n333236 , n329039 );
not ( n42811 , n307864 );
not ( n42812 , n307488 );
not ( n42813 , n42812 );
or ( n42814 , n42811 , n42813 );
nand ( n42815 , n42814 , n16604 );
not ( n42816 , n307015 );
nand ( n42817 , n42816 , n307034 );
not ( n42818 , n42817 );
and ( n42819 , n42815 , n42818 );
not ( n42820 , n42815 );
and ( n42821 , n42820 , n42817 );
nor ( n42822 , n42819 , n42821 );
buf ( n333249 , n42822 );
xor ( n42824 , n333235 , n333236 );
xor ( n42825 , n42824 , n333249 );
buf ( n333252 , n42825 );
xor ( n42827 , n333235 , n333236 );
and ( n42828 , n42827 , n333249 );
and ( n42829 , n333235 , n333236 );
or ( n42830 , n42828 , n42829 );
buf ( n333257 , n42830 );
buf ( n333258 , n309969 );
buf ( n333259 , n328991 );
xnor ( n42834 , n19474 , n17434 );
buf ( n333261 , n42834 );
xor ( n42836 , n333258 , n333259 );
xor ( n42837 , n42836 , n333261 );
buf ( n333264 , n42837 );
xor ( n42839 , n333258 , n333259 );
and ( n42840 , n42839 , n333261 );
and ( n42841 , n333258 , n333259 );
or ( n42842 , n42840 , n42841 );
buf ( n333269 , n42842 );
buf ( n333270 , n33012 );
buf ( n333271 , n328965 );
buf ( n333272 , n17379 );
xor ( n42847 , n333270 , n333271 );
xor ( n42848 , n42847 , n333272 );
buf ( n333275 , n42848 );
xor ( n42850 , n333270 , n333271 );
and ( n42851 , n42850 , n333272 );
and ( n42852 , n333270 , n333271 );
or ( n42853 , n42851 , n42852 );
buf ( n333280 , n42853 );
buf ( n333281 , n323489 );
buf ( n333282 , n323481 );
buf ( n333283 , n307840 );
xor ( n42858 , n333281 , n333282 );
xor ( n42859 , n42858 , n333283 );
buf ( n333286 , n42859 );
xor ( n42861 , n333281 , n333282 );
and ( n42862 , n42861 , n333283 );
and ( n42863 , n333281 , n333282 );
or ( n42864 , n42862 , n42863 );
buf ( n333291 , n42864 );
buf ( n333292 , n323131 );
xnor ( n42867 , n309814 , n19465 );
buf ( n333294 , n42867 );
xor ( n42869 , n333292 , n333294 );
buf ( n333296 , n42869 );
and ( n42871 , n333292 , n333294 );
buf ( n333298 , n42871 );
buf ( n333299 , n324574 );
buf ( n333300 , n324569 );
xor ( n42875 , n333299 , n333300 );
buf ( n333302 , n42875 );
and ( n42877 , n333299 , n333300 );
buf ( n333304 , n42877 );
buf ( n333305 , n324522 );
buf ( n333306 , n34092 );
xor ( n42881 , n333305 , n333306 );
buf ( n333308 , n42881 );
and ( n42883 , n333305 , n333306 );
buf ( n333310 , n42883 );
buf ( n333311 , n36335 );
buf ( n333312 , n36339 );
xor ( n42887 , n333311 , n333312 );
buf ( n333314 , n42887 );
and ( n42889 , n333311 , n333312 );
buf ( n333316 , n42889 );
buf ( n333317 , n36401 );
buf ( n333318 , n36397 );
xor ( n42893 , n333317 , n333318 );
buf ( n333320 , n42893 );
and ( n42895 , n333317 , n333318 );
buf ( n333322 , n42895 );
buf ( n333323 , n326869 );
buf ( n333324 , n326877 );
xor ( n42899 , n333323 , n333324 );
buf ( n333326 , n42899 );
not ( n42901 , n19478 );
nand ( n42902 , n309807 , n309800 );
nor ( n42903 , n309815 , n42902 );
nand ( n42904 , n309928 , n42903 );
not ( n42905 , n42902 );
nand ( n42906 , n42905 , n18214 );
nand ( n42907 , n309921 , n309800 );
and ( n42908 , n42907 , n309563 );
nand ( n42909 , n42904 , n42906 , n42908 );
not ( n42910 , n42909 );
or ( n42911 , n42901 , n42910 );
not ( n42912 , n42902 );
and ( n42913 , n18214 , n42912 );
not ( n42914 , n19478 );
nand ( n42915 , n42914 , n42908 );
nor ( n42916 , n42913 , n42915 );
nand ( n42917 , n42904 , n42916 );
nand ( n42918 , n42911 , n42917 );
buf ( n42919 , n329512 );
buf ( n42920 , n42919 );
or ( n42921 , n42920 , n39079 );
and ( n42922 , n42918 , n42921 );
buf ( n42923 , n42920 );
and ( n42924 , n42923 , n39079 );
nor ( n42925 , n42922 , n42924 );
nand ( n42926 , n309928 , n309804 );
nand ( n42927 , n18214 , n19375 );
and ( n42928 , n309923 , n309802 );
nor ( n42929 , n42928 , n19138 );
nand ( n42930 , n42926 , n42927 , n42929 );
xnor ( n42931 , n33958 , n34039 );
not ( n42932 , n42931 );
not ( n42933 , n19476 );
and ( n42934 , n42932 , n42933 );
and ( n42935 , n42931 , n19476 );
nor ( n42936 , n42934 , n42935 );
xnor ( n42937 , n42930 , n42936 );
nand ( n42938 , n42925 , n42937 );
buf ( n333365 , n42938 );
or ( n42940 , n42925 , n42937 );
buf ( n333367 , n42940 );
nand ( n42942 , n333365 , n333367 );
buf ( n333369 , n42942 );
buf ( n333370 , n333369 );
buf ( n333371 , n333369 );
not ( n42946 , n333371 );
buf ( n333373 , n42946 );
buf ( n333374 , n333373 );
not ( n42949 , n308849 );
nor ( n42950 , n42949 , n18036 );
nand ( n42951 , n42950 , n308846 );
not ( n42952 , n42951 );
not ( n42953 , n17620 );
not ( n42954 , n42953 );
nand ( n42955 , n309928 , n19378 );
nand ( n42956 , n42952 , n42954 , n42955 );
not ( n42957 , n42955 );
not ( n42958 , n42950 );
nand ( n42959 , n42957 , n42958 );
nand ( n42960 , n42953 , n42958 );
or ( n42961 , n42950 , n308846 );
nand ( n42962 , n42956 , n42959 , n42960 , n42961 );
xor ( n42963 , n302980 , n328762 );
and ( n42964 , n42962 , n42963 );
not ( n42965 , n42962 );
not ( n42966 , n42963 );
and ( n42967 , n42965 , n42966 );
nor ( n42968 , n42964 , n42967 );
buf ( n333395 , n42968 );
not ( n42970 , n333395 );
buf ( n333397 , n42970 );
not ( n42972 , n309792 );
buf ( n42973 , n307500 );
not ( n42974 , n42973 );
or ( n42975 , n42972 , n42974 );
nand ( n42976 , n17577 , n17618 );
not ( n42977 , n42976 );
nand ( n42978 , n42975 , n42977 );
not ( n42979 , n12699 );
nand ( n42980 , n42979 , n328847 );
not ( n42981 , n307916 );
nand ( n42982 , n42981 , n308846 );
nand ( n42983 , n42978 , n42980 , n42982 );
not ( n42984 , n42978 );
not ( n42985 , n42980 );
nor ( n42986 , n42985 , n42982 );
and ( n42987 , n42984 , n42986 );
buf ( n42988 , n38422 );
and ( n42989 , n42988 , n12699 );
nor ( n42990 , n42987 , n42989 );
nand ( n42991 , n42983 , n42990 );
buf ( n333418 , n42991 );
not ( n42993 , n333418 );
buf ( n333420 , n42993 );
nand ( n42995 , n333397 , n333420 );
nor ( n42996 , n302980 , n328762 );
nor ( n42997 , n42996 , n42950 );
not ( n42998 , n42997 );
not ( n42999 , n42953 );
or ( n43000 , n42998 , n42999 );
or ( n43001 , n42996 , n42961 );
nand ( n43002 , n43000 , n43001 );
not ( n43003 , n43002 );
nor ( n43004 , n42996 , n42951 );
nand ( n43005 , n42955 , n42954 , n43004 );
not ( n43006 , n42955 );
nand ( n43007 , n43006 , n42997 );
nand ( n43008 , n302980 , n328762 );
nand ( n43009 , n43003 , n43005 , n43007 , n43008 );
not ( n43010 , n43009 );
not ( n43011 , n308465 );
nor ( n43012 , n43011 , n42977 );
and ( n43013 , n309792 , n308465 );
not ( n43014 , n43013 );
not ( n43015 , n307500 );
or ( n43016 , n43014 , n43015 );
not ( n43017 , n18422 );
nand ( n43018 , n43016 , n43017 );
nor ( n43019 , n43012 , n43018 );
xor ( n43020 , n17602 , n38283 );
xor ( n43021 , n43019 , n43020 );
not ( n43022 , n43021 );
and ( n43023 , n17841 , n18429 );
not ( n43024 , n43023 );
and ( n43025 , n43022 , n43024 );
and ( n43026 , n43021 , n43023 );
nor ( n43027 , n43025 , n43026 );
nand ( n43028 , n43010 , n43027 );
and ( n43029 , n42995 , n43028 );
xor ( n43030 , n34661 , n11750 );
not ( n43031 , n43030 );
nor ( n43032 , n308855 , n18432 );
not ( n43033 , n43032 );
nand ( n43034 , n307500 , n309792 , n19447 );
nand ( n43035 , n19447 , n17619 );
and ( n43036 , n18422 , n17841 );
not ( n43037 , n18429 );
nor ( n43038 , n43036 , n43037 );
nand ( n43039 , n43034 , n43035 , n43038 );
not ( n43040 , n43039 );
not ( n43041 , n43040 );
or ( n43042 , n43033 , n43041 );
not ( n43043 , n43032 );
nand ( n43044 , n43043 , n43039 );
nand ( n43045 , n43042 , n43044 );
not ( n43046 , n43045 );
or ( n43047 , n43031 , n43046 );
or ( n43048 , n43030 , n43045 );
nand ( n43049 , n43047 , n43048 );
nor ( n43050 , n17602 , n38283 );
nor ( n43051 , n43050 , n43023 );
nand ( n43052 , n43012 , n43051 );
not ( n43053 , n43050 );
nand ( n43054 , n43053 , n43023 );
or ( n43055 , n43018 , n43012 , n43054 );
nand ( n43056 , n43018 , n43051 );
nand ( n43057 , n17602 , n38283 );
and ( n43058 , n43052 , n43055 , n43056 , n43057 );
nand ( n43059 , n43049 , n43058 );
xnor ( n43060 , n329379 , n329550 );
not ( n43061 , n18039 );
not ( n43062 , n42977 );
and ( n43063 , n43061 , n43062 );
or ( n43064 , n308866 , n18211 );
nor ( n43065 , n43063 , n43064 );
not ( n43066 , n43065 );
not ( n43067 , n19393 );
not ( n43068 , n307500 );
or ( n43069 , n43067 , n43068 );
nand ( n43070 , n43069 , n19428 );
not ( n43071 , n43070 );
not ( n43072 , n43071 );
or ( n43073 , n43066 , n43072 );
nor ( n43074 , n42977 , n18039 );
or ( n43075 , n43074 , n43070 );
nand ( n43076 , n43075 , n43064 );
nand ( n43077 , n43073 , n43076 );
xor ( n43078 , n43060 , n43077 );
or ( n43079 , n11750 , n34661 );
not ( n43080 , n43079 );
not ( n43081 , n43045 );
or ( n43082 , n43080 , n43081 );
nand ( n43083 , n11750 , n34661 );
nand ( n333510 , n43082 , n43083 );
not ( n333511 , n333510 );
nand ( n333512 , n43078 , n333511 );
and ( n43087 , n43059 , n333512 );
nand ( n43088 , n43029 , n43087 );
not ( n333515 , n43088 );
xnor ( n43090 , n324232 , n33807 );
xor ( n43091 , n43090 , n309903 );
not ( n43092 , n309840 );
not ( n43093 , n307500 );
or ( n333520 , n43092 , n43093 );
not ( n333521 , n307515 );
not ( n333522 , n17288 );
or ( n333523 , n333521 , n333522 );
nand ( n43098 , n333523 , n17300 );
not ( n43099 , n19408 );
and ( n333526 , n43098 , n43099 );
not ( n43101 , n309835 );
not ( n43102 , n18229 );
or ( n43103 , n43101 , n43102 );
not ( n43104 , n17607 );
nand ( n333531 , n43103 , n43104 );
nor ( n333532 , n333526 , n333531 );
nand ( n333533 , n333520 , n333532 );
xor ( n333534 , n43091 , n333533 );
buf ( n333535 , n333534 );
not ( n43110 , n17603 );
nand ( n333537 , n43110 , n17606 );
not ( n43112 , n333537 );
not ( n43113 , n43112 );
nor ( n43114 , n43113 , n39274 );
not ( n43115 , n43114 );
nor ( n333542 , n19413 , n19411 , n309908 );
not ( n333543 , n333542 );
not ( n333544 , n307500 );
or ( n43119 , n333543 , n333544 );
not ( n333546 , n307515 );
not ( n43121 , n17288 );
or ( n43122 , n333546 , n43121 );
nand ( n333549 , n43122 , n17300 );
nor ( n43124 , n19413 , n309908 );
and ( n43125 , n333549 , n43124 );
not ( n43126 , n307969 );
not ( n43127 , n18229 );
or ( n333554 , n43126 , n43127 );
nand ( n333555 , n333554 , n308032 );
nor ( n333556 , n43125 , n333555 );
nand ( n333557 , n43119 , n333556 );
not ( n43132 , n333557 );
or ( n43133 , n43115 , n43132 );
not ( n333560 , n333557 );
not ( n43135 , n333537 );
nor ( n43136 , n43135 , n39274 );
nand ( n43137 , n333560 , n43136 );
nand ( n43138 , n43133 , n43137 );
not ( n333565 , n39228 );
or ( n333566 , n43138 , n333565 );
nand ( n333567 , n43112 , n333557 );
nand ( n333568 , n333560 , n333537 );
nand ( n43143 , n333567 , n333568 , n39274 );
nand ( n43144 , n333566 , n43143 );
buf ( n333571 , n43144 );
nor ( n43146 , n333535 , n333571 );
buf ( n333573 , n43146 );
xor ( n43148 , n333565 , n39274 );
not ( n43149 , n43148 );
not ( n333576 , n43149 );
and ( n333577 , n43112 , n333576 );
not ( n333578 , n43112 );
not ( n333579 , n43148 );
and ( n43154 , n333578 , n333579 );
or ( n43155 , n333577 , n43154 );
and ( n333582 , n333557 , n43155 );
not ( n43157 , n333557 );
not ( n43158 , n43149 );
and ( n43159 , n333537 , n43158 );
not ( n43160 , n333537 );
not ( n333587 , n43148 );
and ( n333588 , n43160 , n333587 );
or ( n333589 , n43159 , n333588 );
and ( n333590 , n43157 , n333589 );
or ( n43165 , n333582 , n333590 );
not ( n43166 , n43165 );
nand ( n333593 , n307500 , n309842 );
nand ( n43168 , n18244 , n333593 );
and ( n43169 , n307969 , n308032 );
xnor ( n43170 , n43168 , n43169 );
nor ( n43171 , n39160 , n39168 );
or ( n333598 , n43170 , n43171 );
nand ( n333599 , n39168 , n39160 );
nand ( n333600 , n333598 , n333599 );
nor ( n333601 , n43166 , n333600 );
nor ( n43176 , n333573 , n333601 );
xnor ( n43177 , n34491 , n39250 );
xor ( n333604 , n309945 , n43177 );
not ( n43179 , n309938 );
not ( n43180 , n42973 );
or ( n43181 , n43179 , n43180 );
nand ( n43182 , n43181 , n308666 );
xnor ( n333609 , n333604 , n43182 );
not ( n333610 , n309903 );
not ( n333611 , n333533 );
or ( n333612 , n333610 , n333611 );
or ( n43187 , n333533 , n309903 );
nand ( n43188 , n333612 , n43187 );
or ( n333615 , n324232 , n33807 );
and ( n43190 , n43188 , n333615 );
and ( n43191 , n324232 , n33807 );
nor ( n43192 , n43190 , n43191 );
nand ( n43193 , n333609 , n43192 );
and ( n333620 , n34491 , n39250 );
nor ( n333621 , n333620 , n309945 );
nand ( n333622 , n43182 , n333621 );
not ( n333623 , n43182 );
not ( n43198 , n309945 );
nor ( n43199 , n43198 , n333620 );
nand ( n333626 , n333623 , n43199 );
or ( n43201 , n333620 , n34491 , n39250 );
nand ( n43202 , n333622 , n333626 , n43201 );
xor ( n43203 , n12699 , n38420 );
xor ( n43204 , n42982 , n43203 );
and ( n333631 , n42978 , n43204 );
not ( n333632 , n42978 );
xnor ( n333633 , n43203 , n42982 );
and ( n333634 , n333632 , n333633 );
nor ( n43209 , n333631 , n333634 );
nand ( n43210 , n43202 , n43209 );
nand ( n333637 , n43193 , n43210 );
not ( n43212 , n333637 );
and ( n43213 , n43176 , n43212 );
nand ( n43214 , n333515 , n43213 );
not ( n43215 , n42919 );
not ( n333642 , n39079 );
or ( n333643 , n43215 , n333642 );
or ( n333644 , n39079 , n42919 );
nand ( n333645 , n333643 , n333644 );
and ( n43220 , n42918 , n333645 );
not ( n43221 , n42918 );
not ( n333648 , n333645 );
and ( n43223 , n43221 , n333648 );
nor ( n43224 , n43220 , n43223 );
not ( n43225 , n307500 );
not ( n43226 , n309828 );
or ( n333653 , n43225 , n43226 );
nand ( n333654 , n333653 , n19494 );
not ( n333655 , n309807 );
nor ( n333656 , n333655 , n42977 );
nor ( n43231 , n333654 , n333656 );
not ( n43232 , n43231 );
nor ( n333659 , n309986 , n33616 );
nand ( n43234 , n309800 , n309563 );
not ( n43235 , n43234 );
or ( n43236 , n333659 , n43235 );
not ( n43237 , n43236 );
and ( n333664 , n43232 , n43237 );
nor ( n333665 , n333659 , n43234 );
not ( n333666 , n333665 );
not ( n333667 , n43231 );
or ( n43242 , n333666 , n333667 );
nand ( n43243 , n33616 , n309986 );
nand ( n333670 , n43242 , n43243 );
nor ( n43245 , n333664 , n333670 );
nand ( n43246 , n43224 , n43245 );
not ( n43247 , n39110 );
buf ( n43248 , n43247 );
or ( n333675 , n324020 , n43248 );
not ( n333676 , n333675 );
not ( n43251 , n309901 );
not ( n333678 , n43251 );
nand ( n333679 , n307500 , n309792 , n308640 );
nand ( n43254 , n333679 , n308641 , n18451 );
not ( n43255 , n43254 );
not ( n333682 , n43255 );
or ( n43257 , n333678 , n333682 );
nand ( n43258 , n43254 , n309901 );
nand ( n43259 , n43257 , n43258 );
not ( n43260 , n43259 );
or ( n333687 , n333676 , n43260 );
nand ( n333688 , n43248 , n324020 );
nand ( n333689 , n333687 , n333688 );
not ( n333690 , n333689 );
xor ( n43265 , n33870 , n7448 );
not ( n43266 , n43265 );
not ( n333693 , n19392 );
not ( n43268 , n307500 );
or ( n43269 , n333693 , n43268 );
nand ( n43270 , n43269 , n18448 );
not ( n43271 , n43270 );
not ( n333698 , n17618 );
not ( n333699 , n17577 );
or ( n43274 , n333698 , n333699 );
not ( n333701 , n19391 );
nand ( n333702 , n43274 , n333701 );
not ( n43277 , n333702 );
not ( n43278 , n43277 );
nand ( n333705 , n43271 , n43278 );
not ( n43280 , n333705 );
or ( n43281 , n43266 , n43280 );
not ( n43282 , n43270 );
not ( n43283 , n43265 );
nand ( n333710 , n43282 , n43278 , n43283 );
nand ( n333711 , n43281 , n333710 );
not ( n43286 , n333711 );
not ( n333713 , n309728 );
and ( n333714 , n19294 , n333713 );
not ( n43289 , n333714 );
and ( n43290 , n43286 , n43289 );
not ( n333717 , n43265 );
not ( n43292 , n333705 );
or ( n43293 , n333717 , n43292 );
nand ( n43294 , n43293 , n333710 );
and ( n43295 , n43294 , n333714 );
nor ( n333722 , n43290 , n43295 );
nand ( n333723 , n333690 , n333722 );
or ( n43298 , n329379 , n329550 );
and ( n43299 , n43077 , n43298 );
and ( n333726 , n329379 , n329550 );
nor ( n333727 , n43299 , n333726 );
xor ( n43302 , n43247 , n324020 );
not ( n43303 , n43302 );
not ( n333730 , n43259 );
or ( n43305 , n43303 , n333730 );
or ( n43306 , n43302 , n43259 );
nand ( n43307 , n43305 , n43306 );
nand ( n43308 , n333727 , n43307 );
not ( n333735 , n307500 );
not ( n43310 , n309818 );
or ( n333737 , n333735 , n43310 );
nand ( n43312 , n333737 , n19303 );
not ( n333739 , n43312 );
or ( n333740 , n42977 , n309817 );
nand ( n43315 , n333739 , n333740 );
nor ( n43316 , n302388 , n33622 );
not ( n333743 , n19368 );
nor ( n43318 , n333743 , n309879 );
nor ( n43319 , n43316 , n43318 );
nand ( n43320 , n43315 , n43319 );
not ( n43321 , n43312 );
not ( n333748 , n43316 );
and ( n43323 , n43318 , n333748 );
nand ( n333750 , n43321 , n333740 , n43323 );
nand ( n333751 , n302388 , n33622 );
nand ( n333752 , n43320 , n333750 , n333751 );
not ( n43327 , n333752 );
not ( n43328 , n333659 );
nand ( n333755 , n43328 , n43243 );
and ( n43330 , n333755 , n43234 );
not ( n43331 , n333755 );
and ( n43332 , n43331 , n43235 );
or ( n43333 , n43330 , n43332 );
and ( n333760 , n43231 , n43333 );
not ( n333761 , n43231 );
and ( n43336 , n333755 , n43235 );
not ( n333763 , n333755 );
and ( n333764 , n333763 , n43234 );
or ( n43339 , n43336 , n333764 );
and ( n43340 , n333761 , n43339 );
nor ( n333767 , n333760 , n43340 );
not ( n43342 , n333767 );
nand ( n43343 , n43327 , n43342 );
and ( n43344 , n333723 , n43308 , n43343 );
nor ( n43345 , n33870 , n7448 );
not ( n333772 , n43345 );
nand ( n333773 , n333772 , n333714 );
nor ( n333774 , n43270 , n333773 );
nand ( n333775 , n333774 , n43278 );
nor ( n43350 , n43345 , n333714 );
nand ( n43351 , n43350 , n333705 );
nand ( n333778 , n33870 , n7448 );
and ( n43353 , n333775 , n43351 , n333778 );
buf ( n333780 , n43353 );
xor ( n43355 , n302388 , n33622 );
xor ( n43356 , n43318 , n43355 );
not ( n333783 , n42977 );
not ( n333784 , n309817 );
and ( n43359 , n333783 , n333784 );
nor ( n333786 , n43359 , n43312 );
xnor ( n333787 , n43356 , n333786 );
buf ( n333788 , n333787 );
not ( n43363 , n333788 );
buf ( n333790 , n43363 );
buf ( n333791 , n333790 );
nand ( n43366 , n333780 , n333791 );
buf ( n333793 , n43366 );
buf ( n43368 , n333793 );
buf ( n333795 , n43368 );
nand ( n333796 , n43246 , n43344 , n333795 );
nor ( n333797 , n43214 , n333796 );
not ( n333798 , n333797 );
not ( n43373 , n33311 );
not ( n43374 , n43373 );
or ( n333801 , n43374 , n328863 );
not ( n43376 , n333801 );
nand ( n43377 , n308673 , n17442 , n307809 );
not ( n43378 , n16434 );
nand ( n43379 , n43378 , n16437 );
not ( n333806 , n43379 );
and ( n333807 , n43377 , n333806 );
not ( n333808 , n43377 );
and ( n333809 , n333808 , n43379 );
nor ( n43384 , n333807 , n333809 );
not ( n43385 , n43384 );
or ( n333812 , n43376 , n43385 );
nand ( n43387 , n43374 , n328863 );
nand ( n43388 , n333812 , n43387 );
buf ( n333815 , n43388 );
not ( n43390 , n333815 );
buf ( n333817 , n43390 );
buf ( n43392 , n333817 );
and ( n43393 , n298380 , n328858 );
not ( n333820 , n298380 );
not ( n333821 , n328858 );
and ( n43396 , n333820 , n333821 );
nor ( n43397 , n43393 , n43396 );
not ( n333824 , n43397 );
not ( n43399 , n333824 );
and ( n43400 , n309884 , n43399 );
not ( n43401 , n309884 );
not ( n43402 , n43397 );
and ( n333829 , n43401 , n43402 );
or ( n333830 , n43400 , n333829 );
and ( n333831 , n307857 , n333830 );
not ( n333832 , n307857 );
not ( n43407 , n333824 );
and ( n43408 , n309883 , n43407 );
not ( n333835 , n309883 );
not ( n43410 , n43397 );
and ( n43411 , n333835 , n43410 );
or ( n43412 , n43408 , n43411 );
and ( n43413 , n333832 , n43412 );
or ( n333840 , n333831 , n43413 );
not ( n333841 , n333840 );
buf ( n43416 , n333841 );
nand ( n333843 , n43392 , n43416 );
buf ( n333844 , n333843 );
buf ( n333845 , n333844 );
xor ( n333846 , n43374 , n328863 );
not ( n43421 , n333846 );
not ( n43422 , n43421 );
and ( n43423 , n333806 , n43422 );
not ( n43424 , n333806 );
not ( n333851 , n333846 );
and ( n333852 , n43424 , n333851 );
or ( n333853 , n43423 , n333852 );
and ( n333854 , n43377 , n333853 );
not ( n43429 , n43377 );
not ( n43430 , n43421 );
and ( n333857 , n43379 , n43430 );
not ( n43432 , n43379 );
not ( n43433 , n333846 );
and ( n43434 , n43432 , n43433 );
or ( n43435 , n333857 , n43434 );
and ( n333862 , n43429 , n43435 );
or ( n333863 , n333854 , n333862 );
buf ( n333864 , n333863 );
not ( n43439 , n333864 );
buf ( n333866 , n43439 );
buf ( n333867 , n333866 );
or ( n333868 , n33180 , n330189 );
not ( n333869 , n333868 );
not ( n333870 , n307820 );
or ( n43445 , n333869 , n333870 );
nand ( n333872 , n33180 , n330189 );
nand ( n43447 , n43445 , n333872 );
buf ( n333874 , n43447 );
not ( n333875 , n333874 );
buf ( n333876 , n333875 );
buf ( n333877 , n333876 );
nand ( n333878 , n333867 , n333877 );
buf ( n333879 , n333878 );
buf ( n333880 , n333879 );
nand ( n333881 , n333845 , n333880 );
buf ( n333882 , n333881 );
buf ( n333883 , n333882 );
not ( n333884 , n333883 );
xor ( n43459 , n330214 , n328814 );
and ( n333886 , n43459 , n307790 );
and ( n333887 , n330214 , n328814 );
or ( n333888 , n333886 , n333887 );
not ( n43463 , n333888 );
not ( n333890 , n38382 );
and ( n333891 , n333890 , n293601 );
not ( n333892 , n333890 );
not ( n333893 , n293601 );
and ( n333894 , n333892 , n333893 );
nor ( n43469 , n333891 , n333894 );
xor ( n333896 , n307772 , n43469 );
not ( n333897 , n333896 );
and ( n43472 , n43463 , n333897 );
xor ( n333899 , n330214 , n328814 );
xor ( n333900 , n333899 , n307790 );
buf ( n333901 , n333900 );
not ( n333902 , n298380 );
nand ( n333903 , n333902 , n333821 );
not ( n43478 , n333903 );
and ( n333905 , n307857 , n309884 );
not ( n333906 , n307857 );
and ( n43481 , n333906 , n309883 );
nor ( n333908 , n333905 , n43481 );
not ( n333909 , n333908 );
or ( n43484 , n43478 , n333909 );
nand ( n333911 , n298380 , n328858 );
nand ( n43486 , n43484 , n333911 );
buf ( n333913 , n43486 );
nor ( n333914 , n333901 , n333913 );
buf ( n333915 , n333914 );
nor ( n43490 , n43472 , n333915 );
buf ( n333917 , n43490 );
nand ( n43492 , n333884 , n333917 );
buf ( n333919 , n43492 );
buf ( n333920 , n333919 );
not ( n43495 , n333920 );
buf ( n43496 , n43495 );
buf ( n43497 , n333286 );
not ( n43498 , n43497 );
buf ( n333925 , n43498 );
buf ( n333926 , n33077 );
buf ( n333927 , n1916 );
xor ( n333928 , n333926 , n333927 );
buf ( n333929 , n307852 );
and ( n333930 , n333928 , n333929 );
and ( n43505 , n333926 , n333927 );
or ( n333932 , n333930 , n43505 );
buf ( n333933 , n333932 );
buf ( n333934 , n333933 );
not ( n333935 , n333934 );
buf ( n333936 , n333935 );
nand ( n333937 , n333925 , n333936 );
buf ( n333938 , n333291 );
not ( n43513 , n333938 );
buf ( n333940 , n43513 );
buf ( n333941 , n333940 );
xor ( n43516 , n323529 , n10720 );
and ( n43517 , n307877 , n307107 );
not ( n333944 , n17448 );
not ( n43519 , n16626 );
or ( n333946 , n333944 , n43519 );
nand ( n333947 , n333946 , n309877 );
not ( n43522 , n333947 );
not ( n43523 , n307823 );
nand ( n43524 , n43523 , n17448 , n307746 );
nand ( n43525 , n43522 , n43524 );
xor ( n43526 , n43517 , n43525 );
xor ( n43527 , n43516 , n43526 );
buf ( n333954 , n43527 );
not ( n43529 , n333954 );
buf ( n333956 , n43529 );
buf ( n43531 , n333956 );
nand ( n43532 , n333941 , n43531 );
buf ( n43533 , n43532 );
and ( n333960 , n333937 , n43533 );
xor ( n43535 , n33180 , n330188 );
and ( n333962 , n307820 , n43535 );
not ( n333963 , n307820 );
not ( n333964 , n43535 );
and ( n43539 , n333963 , n333964 );
nor ( n333966 , n333962 , n43539 );
not ( n43541 , n333966 );
or ( n333968 , n38133 , n328573 );
not ( n43543 , n333968 );
not ( n333970 , n16681 );
nor ( n43545 , n333970 , n16683 );
and ( n333972 , n16626 , n17450 );
not ( n333973 , n307877 );
not ( n43548 , n307103 );
or ( n333975 , n333973 , n43548 );
nand ( n333976 , n333975 , n307107 );
nor ( n333977 , n333972 , n333976 );
nand ( n43552 , n333977 , n17451 );
xor ( n43553 , n43545 , n43552 );
not ( n43554 , n43553 );
or ( n43555 , n43543 , n43554 );
nand ( n333982 , n38133 , n328573 );
nand ( n333983 , n43555 , n333982 );
not ( n43558 , n333983 );
nand ( n333985 , n43541 , n43558 );
xor ( n333986 , n38133 , n328573 );
and ( n43561 , n43553 , n333986 );
not ( n333988 , n43553 );
not ( n333989 , n333986 );
and ( n333990 , n333988 , n333989 );
or ( n333991 , n43561 , n333990 );
buf ( n333992 , n333991 );
xor ( n333993 , n323529 , n10720 );
and ( n333994 , n333993 , n43526 );
and ( n333995 , n323529 , n10720 );
or ( n333996 , n333994 , n333995 );
buf ( n333997 , n333996 );
not ( n333998 , n333997 );
buf ( n333999 , n333998 );
buf ( n334000 , n333999 );
nand ( n334001 , n333992 , n334000 );
buf ( n334002 , n334001 );
and ( n43577 , n333985 , n334002 );
nand ( n334004 , n333960 , n43577 );
not ( n334005 , n334004 );
nand ( n43580 , n43496 , n334005 );
not ( n334007 , n43580 );
buf ( n334008 , n333257 );
buf ( n334009 , n333264 );
nor ( n334010 , n334008 , n334009 );
buf ( n334011 , n334010 );
buf ( n334012 , n334011 );
not ( n334013 , n334012 );
buf ( n334014 , n334013 );
not ( n334015 , n334014 );
buf ( n334016 , n333252 );
buf ( n43591 , n333234 );
and ( n43592 , n334016 , n43591 );
buf ( n334019 , n43592 );
not ( n43594 , n334019 );
or ( n43595 , n334015 , n43594 );
buf ( n334022 , n333257 );
buf ( n334023 , n333264 );
nand ( n334024 , n334022 , n334023 );
buf ( n334025 , n334024 );
nand ( n43600 , n43595 , n334025 );
buf ( n334027 , n333269 );
buf ( n43602 , n333275 );
nor ( n43603 , n334027 , n43602 );
buf ( n43604 , n43603 );
xor ( n334031 , n323498 , n1916 );
xnor ( n334032 , n334031 , n307852 );
nor ( n43607 , n334032 , n333280 );
nor ( n43608 , n43604 , n43607 );
nand ( n43609 , n43600 , n43608 );
buf ( n334036 , n43607 );
not ( n43611 , n334036 );
buf ( n334038 , n43611 );
buf ( n43613 , n333275 );
buf ( n334040 , n333269 );
and ( n334041 , n43613 , n334040 );
buf ( n334042 , n334041 );
and ( n43617 , n334038 , n334042 );
buf ( n334044 , n333280 );
xor ( n334045 , n333926 , n333927 );
xor ( n43620 , n334045 , n333929 );
buf ( n334047 , n43620 );
buf ( n334048 , n334047 );
nand ( n43623 , n334044 , n334048 );
buf ( n334050 , n43623 );
buf ( n334051 , n334050 );
not ( n334052 , n334051 );
buf ( n334053 , n334052 );
nor ( n43628 , n43617 , n334053 );
nand ( n334055 , n43609 , n43628 );
not ( n334056 , n334055 );
buf ( n334057 , n333229 );
buf ( n334058 , n333223 );
nor ( n334059 , n334057 , n334058 );
buf ( n334060 , n334059 );
buf ( n334061 , n334060 );
buf ( n334062 , n333218 );
buf ( n334063 , n333212 );
nor ( n334064 , n334062 , n334063 );
buf ( n334065 , n334064 );
buf ( n334066 , n334065 );
nor ( n43641 , n334061 , n334066 );
buf ( n334068 , n43641 );
buf ( n334069 , n334068 );
not ( n43644 , n334069 );
buf ( n334071 , n333193 );
xor ( n334072 , n330451 , n323217 );
xor ( n43647 , n334072 , n307913 );
buf ( n334074 , n43647 );
nand ( n334075 , n334071 , n334074 );
buf ( n334076 , n334075 );
not ( n334077 , n334076 );
not ( n334078 , n334077 );
xor ( n334079 , n330451 , n323217 );
and ( n43654 , n334079 , n307913 );
and ( n334081 , n330451 , n323217 );
or ( n43656 , n43654 , n334081 );
or ( n43657 , n43656 , n333207 );
not ( n43658 , n43657 );
or ( n334085 , n334078 , n43658 );
nand ( n334086 , n333207 , n43656 );
nand ( n43661 , n334085 , n334086 );
buf ( n334088 , n43661 );
not ( n334089 , n334088 );
or ( n43664 , n43644 , n334089 );
buf ( n334091 , n334060 );
not ( n43666 , n334091 );
buf ( n334093 , n333218 );
buf ( n334094 , n333212 );
nand ( n334095 , n334093 , n334094 );
buf ( n334096 , n334095 );
buf ( n334097 , n334096 );
not ( n334098 , n334097 );
and ( n43673 , n43666 , n334098 );
buf ( n334100 , n333229 );
buf ( n334101 , n333223 );
and ( n43676 , n334100 , n334101 );
buf ( n334103 , n43676 );
buf ( n334104 , n334103 );
nor ( n43679 , n43673 , n334104 );
buf ( n334106 , n43679 );
buf ( n334107 , n334106 );
nand ( n43682 , n43664 , n334107 );
buf ( n334109 , n43682 );
buf ( n334110 , n43657 );
buf ( n334111 , n333193 );
buf ( n334112 , n43647 );
or ( n43687 , n334111 , n334112 );
buf ( n334114 , n43687 );
buf ( n334115 , n334114 );
and ( n43690 , n334110 , n334115 );
buf ( n334117 , n43690 );
buf ( n334118 , n334117 );
buf ( n334119 , n334068 );
nand ( n334120 , n334118 , n334119 );
buf ( n334121 , n334120 );
buf ( n334122 , n334121 );
or ( n43697 , n329327 , n323104 );
not ( n334124 , n43697 );
and ( n334125 , n309907 , n307238 );
not ( n43700 , n334125 );
not ( n334127 , n307465 );
or ( n334128 , n43700 , n334127 );
not ( n43703 , n307238 );
not ( n43704 , n309907 );
or ( n334131 , n43703 , n43704 );
nand ( n43706 , n334131 , n308644 );
nand ( n334133 , n334128 , n43706 );
not ( n334134 , n334133 );
or ( n43709 , n334124 , n334134 );
nand ( n334136 , n329327 , n323104 );
nand ( n334137 , n43709 , n334136 );
buf ( n334138 , n334137 );
buf ( n334139 , n333143 );
nand ( n43714 , n334138 , n334139 );
buf ( n43715 , n43714 );
buf ( n334142 , n43715 );
buf ( n334143 , n333155 );
buf ( n334144 , n333148 );
nor ( n334145 , n334143 , n334144 );
buf ( n334146 , n334145 );
buf ( n334147 , n334146 );
or ( n334148 , n334142 , n334147 );
buf ( n334149 , n333148 );
buf ( n334150 , n333155 );
nand ( n334151 , n334149 , n334150 );
buf ( n334152 , n334151 );
buf ( n334153 , n334152 );
nand ( n43728 , n334148 , n334153 );
buf ( n334155 , n43728 );
buf ( n334156 , n334155 );
buf ( n334157 , n333188 );
buf ( n334158 , n333182 );
nor ( n334159 , n334157 , n334158 );
buf ( n334160 , n334159 );
buf ( n334161 , n334160 );
nor ( n334162 , n333177 , n333160 );
buf ( n334163 , n334162 );
nor ( n334164 , n334161 , n334163 );
buf ( n334165 , n334164 );
buf ( n334166 , n334165 );
nand ( n43741 , n334156 , n334166 );
buf ( n334168 , n43741 );
buf ( n334169 , n334168 );
buf ( n334170 , n334146 );
buf ( n43745 , n333143 );
buf ( n334172 , n334137 );
nor ( n334173 , n43745 , n334172 );
buf ( n334174 , n334173 );
buf ( n334175 , n334174 );
nor ( n334176 , n334170 , n334175 );
buf ( n334177 , n334176 );
buf ( n334178 , n334177 );
xnor ( n334179 , n329327 , n323104 );
not ( n334180 , n334179 );
not ( n43755 , n334133 );
or ( n334182 , n334180 , n43755 );
or ( n334183 , n334133 , n334179 );
nand ( n43758 , n334182 , n334183 );
buf ( n334185 , n43758 );
not ( n334186 , n323118 );
not ( n334187 , n40107 );
or ( n43762 , n334186 , n334187 );
or ( n334189 , n40107 , n323118 );
and ( n334190 , n309947 , n309789 );
not ( n43765 , n309947 );
not ( n334192 , n309789 );
and ( n334193 , n43765 , n334192 );
nor ( n43768 , n334190 , n334193 );
nand ( n334195 , n334189 , n43768 );
nand ( n334196 , n43762 , n334195 );
buf ( n334197 , n334196 );
nor ( n43772 , n334185 , n334197 );
buf ( n334199 , n43772 );
buf ( n334200 , n334199 );
buf ( n334201 , n18256 );
buf ( n334202 , n40137 );
or ( n334203 , n334201 , n334202 );
buf ( n334204 , n334203 );
buf ( n43779 , n334204 );
buf ( n43780 , n32707 );
xor ( n43781 , n43779 , n43780 );
buf ( n43782 , n333296 );
and ( n43783 , n43781 , n43782 );
and ( n43784 , n43779 , n43780 );
or ( n43785 , n43783 , n43784 );
buf ( n43786 , n43785 );
buf ( n334213 , n43786 );
xor ( n43788 , n40107 , n323118 );
xor ( n334215 , n43788 , n309947 );
xnor ( n334216 , n334215 , n334192 );
buf ( n334217 , n334216 );
buf ( n334218 , n333298 );
or ( n334219 , n334217 , n334218 );
buf ( n334220 , n334219 );
buf ( n43795 , n334220 );
nand ( n43796 , n334213 , n43795 );
buf ( n43797 , n43796 );
buf ( n334224 , n43797 );
or ( n43799 , n334200 , n334224 );
buf ( n334226 , n334199 );
buf ( n43801 , n334216 );
buf ( n334228 , n333298 );
nand ( n43803 , n43801 , n334228 );
buf ( n334230 , n43803 );
buf ( n334231 , n334230 );
or ( n334232 , n334226 , n334231 );
buf ( n334233 , n334196 );
buf ( n43808 , n43758 );
nand ( n334235 , n334233 , n43808 );
buf ( n334236 , n334235 );
buf ( n334237 , n334236 );
nand ( n43812 , n43799 , n334232 , n334237 );
buf ( n334239 , n43812 );
buf ( n334240 , n334239 );
and ( n334241 , n334178 , n334240 );
buf ( n334242 , n334241 );
buf ( n334243 , n334242 );
buf ( n334244 , n334165 );
nand ( n334245 , n334243 , n334244 );
buf ( n334246 , n334245 );
buf ( n334247 , n334246 );
buf ( n334248 , n333160 );
buf ( n334249 , n333177 );
nand ( n334250 , n334248 , n334249 );
buf ( n334251 , n334250 );
buf ( n334252 , n334251 );
not ( n334253 , n334252 );
buf ( n334254 , n334160 );
not ( n43829 , n334254 );
and ( n334256 , n334253 , n43829 );
buf ( n334257 , n333188 );
buf ( n334258 , n333182 );
and ( n334259 , n334257 , n334258 );
buf ( n334260 , n334259 );
buf ( n334261 , n334260 );
nor ( n334262 , n334256 , n334261 );
buf ( n334263 , n334262 );
buf ( n334264 , n334263 );
and ( n334265 , n334169 , n334247 , n334264 );
buf ( n334266 , n334265 );
buf ( n334267 , n334266 );
nor ( n334268 , n334122 , n334267 );
buf ( n334269 , n334268 );
or ( n334270 , n334109 , n334269 );
nor ( n334271 , n43607 , n43604 );
buf ( n334272 , n334271 );
buf ( n334273 , n333252 );
buf ( n334274 , n333234 );
nor ( n43849 , n334273 , n334274 );
buf ( n334276 , n43849 );
buf ( n43851 , n334276 );
buf ( n43852 , n334011 );
nor ( n43853 , n43851 , n43852 );
buf ( n43854 , n43853 );
buf ( n334281 , n43854 );
and ( n43856 , n334272 , n334281 );
buf ( n43857 , n43856 );
nand ( n334284 , n334270 , n43857 );
nand ( n43859 , n334056 , n334284 );
nand ( n334286 , n334007 , n43859 );
buf ( n334287 , n334286 );
nand ( n43862 , n333985 , n334002 );
buf ( n334289 , n43533 );
buf ( n334290 , n333936 );
buf ( n334291 , n333925 );
nor ( n334292 , n334290 , n334291 );
buf ( n334293 , n334292 );
buf ( n334294 , n334293 );
and ( n334295 , n334289 , n334294 );
buf ( n43870 , n333940 );
buf ( n334297 , n333956 );
nor ( n334298 , n43870 , n334297 );
buf ( n334299 , n334298 );
buf ( n334300 , n334299 );
nor ( n43875 , n334295 , n334300 );
buf ( n334302 , n43875 );
nor ( n334303 , n43862 , n334302 );
buf ( n334304 , n334303 );
nor ( n334305 , n333991 , n333999 );
not ( n334306 , n334305 );
not ( n43881 , n333985 );
or ( n334308 , n334306 , n43881 );
nand ( n334309 , n333966 , n333983 );
nand ( n43884 , n334308 , n334309 );
buf ( n334311 , n43884 );
nor ( n334312 , n334304 , n334311 );
buf ( n334313 , n334312 );
buf ( n334314 , n334313 );
not ( n334315 , n334314 );
buf ( n334316 , n333919 );
not ( n43891 , n334316 );
and ( n43892 , n334315 , n43891 );
buf ( n334319 , n43490 );
not ( n334320 , n334319 );
buf ( n334321 , n333863 );
buf ( n334322 , n43447 );
and ( n334323 , n334321 , n334322 );
buf ( n334324 , n334323 );
buf ( n334325 , n334324 );
not ( n334326 , n334325 );
buf ( n334327 , n333844 );
not ( n334328 , n334327 );
or ( n43903 , n334326 , n334328 );
buf ( n334330 , n43388 );
not ( n43905 , n333841 );
buf ( n334332 , n43905 );
nand ( n334333 , n334330 , n334332 );
buf ( n334334 , n334333 );
buf ( n334335 , n334334 );
nand ( n334336 , n43903 , n334335 );
buf ( n334337 , n334336 );
buf ( n334338 , n334337 );
not ( n334339 , n334338 );
or ( n334340 , n334320 , n334339 );
buf ( n334341 , n333900 );
buf ( n334342 , n43486 );
nand ( n334343 , n334341 , n334342 );
buf ( n334344 , n334343 );
buf ( n334345 , n334344 );
not ( n43920 , n334345 );
buf ( n43921 , n43920 );
buf ( n334348 , n43921 );
or ( n43923 , n333896 , n333888 );
buf ( n334350 , n43923 );
and ( n334351 , n334348 , n334350 );
buf ( n334352 , n333888 );
buf ( n334353 , n333896 );
and ( n334354 , n334352 , n334353 );
buf ( n334355 , n334354 );
buf ( n334356 , n334355 );
nor ( n334357 , n334351 , n334356 );
buf ( n334358 , n334357 );
buf ( n334359 , n334358 );
nand ( n334360 , n334340 , n334359 );
buf ( n334361 , n334360 );
buf ( n334362 , n334361 );
nor ( n334363 , n43892 , n334362 );
buf ( n334364 , n334363 );
buf ( n334365 , n334364 );
nand ( n334366 , n334287 , n334365 );
buf ( n334367 , n334366 );
buf ( n334368 , n334367 );
or ( n334369 , n38359 , n296411 );
not ( n334370 , n334369 );
not ( n43945 , n307758 );
or ( n334372 , n334370 , n43945 );
nand ( n334373 , n38359 , n296411 );
nand ( n43948 , n334372 , n334373 );
not ( n43949 , n43948 );
xor ( n334376 , n38309 , n328740 );
and ( n334377 , n17332 , n17444 );
not ( n43952 , n334377 );
nand ( n334379 , n307745 , n17319 );
nand ( n334380 , n334379 , n17387 );
not ( n43955 , n334380 );
or ( n334382 , n43952 , n43955 );
and ( n334383 , n307738 , n17444 );
nor ( n43958 , n334383 , n306989 );
nand ( n334385 , n334382 , n43958 );
nand ( n334386 , n16565 , n306975 );
not ( n43961 , n334386 );
and ( n334388 , n334385 , n43961 );
not ( n334389 , n334385 );
and ( n334390 , n334389 , n334386 );
nor ( n43965 , n334388 , n334390 );
and ( n334392 , n334376 , n43965 );
not ( n43967 , n334376 );
not ( n43968 , n43965 );
and ( n43969 , n43967 , n43968 );
nor ( n334396 , n334392 , n43969 );
not ( n334397 , n334396 );
nand ( n43972 , n43949 , n334397 );
buf ( n334399 , n43972 );
xnor ( n43974 , n38359 , n296411 );
xor ( n334401 , n43974 , n307758 );
buf ( n334402 , n333890 );
not ( n334403 , n334402 );
nand ( n43978 , n334403 , n333893 );
not ( n334405 , n43978 );
not ( n334406 , n307772 );
or ( n43981 , n334405 , n334406 );
nand ( n43982 , n293601 , n334402 );
nand ( n43983 , n43981 , n43982 );
not ( n43984 , n43983 );
nand ( n43985 , n334401 , n43984 );
buf ( n334412 , n43985 );
nand ( n334413 , n334399 , n334412 );
buf ( n334414 , n334413 );
buf ( n43989 , n334414 );
not ( n334416 , n43989 );
buf ( n334417 , n334416 );
or ( n334418 , n4309 , n39655 );
not ( n334419 , n334418 );
nand ( n43994 , n17447 , n308674 , n19482 );
not ( n334421 , n16563 );
and ( n334422 , n306995 , n334421 );
xor ( n334423 , n43994 , n334422 );
not ( n43998 , n334423 );
or ( n334425 , n334419 , n43998 );
nand ( n334426 , n4309 , n39655 );
nand ( n44001 , n334425 , n334426 );
or ( n334428 , n323889 , n330023 );
nand ( n44003 , n323889 , n330023 );
nand ( n44004 , n334428 , n44003 );
not ( n334431 , n19471 );
not ( n44006 , n309928 );
or ( n334433 , n334431 , n44006 );
or ( n334434 , n309928 , n19471 );
nand ( n44009 , n334433 , n334434 );
xnor ( n334436 , n44004 , n44009 );
nor ( n334437 , n44001 , n334436 );
and ( n334438 , n334418 , n334426 );
and ( n334439 , n334438 , n334423 );
not ( n44014 , n334438 );
not ( n334441 , n334423 );
and ( n334442 , n44014 , n334441 );
nor ( n44017 , n334439 , n334442 );
not ( n334444 , n328740 );
not ( n334445 , n38309 );
or ( n44020 , n334444 , n334445 );
or ( n44021 , n38309 , n328740 );
nand ( n334448 , n44021 , n43965 );
nand ( n44023 , n44020 , n334448 );
nor ( n334450 , n44017 , n44023 );
nor ( n334451 , n334437 , n334450 );
and ( n44026 , n334417 , n334451 );
buf ( n334453 , n44026 );
nand ( n334454 , n334368 , n334453 );
buf ( n334455 , n334454 );
nor ( n334456 , n334436 , n44001 );
not ( n334457 , n334456 );
nor ( n44032 , n334401 , n43984 );
not ( n334459 , n44032 );
not ( n334460 , n43972 );
or ( n44035 , n334459 , n334460 );
nand ( n334462 , n334396 , n43948 );
nand ( n334463 , n44035 , n334462 );
or ( n44038 , n44017 , n44023 );
nand ( n44039 , n334457 , n334463 , n44038 );
not ( n44040 , n334437 );
nand ( n334467 , n44017 , n44023 );
not ( n334468 , n334467 );
and ( n44043 , n44040 , n334468 );
and ( n44044 , n334436 , n44001 );
nor ( n44045 , n44043 , n44044 );
nand ( n334472 , n44039 , n44045 );
buf ( n334473 , n334472 );
not ( n44048 , n334473 );
buf ( n334475 , n44048 );
buf ( n44050 , n328661 );
or ( n334477 , n296368 , n44050 );
not ( n334478 , n334477 );
not ( n44053 , n309872 );
not ( n44054 , n307500 );
or ( n44055 , n44053 , n44054 );
nand ( n334482 , n44055 , n309876 );
and ( n334483 , n334482 , n309897 );
not ( n44058 , n334482 );
and ( n44059 , n44058 , n19468 );
nor ( n44060 , n334483 , n44059 );
not ( n334487 , n44060 );
or ( n334488 , n334478 , n334487 );
nand ( n334489 , n296368 , n44050 );
nand ( n334490 , n334488 , n334489 );
not ( n334491 , n334490 );
not ( n334492 , n334491 );
nand ( n44067 , n307503 , n17079 );
not ( n334494 , n44067 );
not ( n334495 , n309873 );
not ( n44070 , n307500 );
or ( n334497 , n334495 , n44070 );
nand ( n334498 , n334497 , n309855 );
not ( n334499 , n334498 );
or ( n44074 , n334494 , n334499 );
or ( n334501 , n44067 , n334498 );
nand ( n334502 , n44074 , n334501 );
not ( n44077 , n334502 );
or ( n334504 , n323862 , n33506 );
nand ( n334505 , n323862 , n33506 );
nand ( n44080 , n334504 , n334505 );
not ( n334507 , n44080 );
nand ( n334508 , n44077 , n334507 );
nand ( n334509 , n334502 , n44080 );
nand ( n334510 , n334508 , n334509 );
not ( n44085 , n334510 );
not ( n334512 , n44085 );
or ( n334513 , n334492 , n334512 );
not ( n44088 , n328638 );
and ( n334515 , n44088 , n328648 );
not ( n334516 , n328648 );
and ( n334517 , n328638 , n334516 );
nor ( n44092 , n334515 , n334517 );
not ( n334519 , n44092 );
not ( n334520 , n334519 );
not ( n334521 , n17094 );
not ( n334522 , n334521 );
or ( n44097 , n334520 , n334522 );
nand ( n334524 , n17094 , n44092 );
nand ( n334525 , n44097 , n334524 );
not ( n44100 , n334525 );
nand ( n334527 , n334504 , n334502 );
nand ( n334528 , n44100 , n334527 , n334505 );
nand ( n44103 , n334513 , n334528 );
not ( n334530 , n44103 );
not ( n334531 , n334428 );
not ( n334532 , n44009 );
or ( n44107 , n334531 , n334532 );
nand ( n44108 , n44107 , n44003 );
xor ( n44109 , n328533 , n12778 );
not ( n44110 , n44109 );
not ( n44111 , n16405 );
nand ( n44112 , n44111 , n307512 );
not ( n44113 , n44112 );
and ( n44114 , n44110 , n44113 );
and ( n44115 , n44112 , n44109 );
nor ( n334542 , n44114 , n44115 );
not ( n44117 , n306801 );
not ( n334544 , n307500 );
or ( n334545 , n44117 , n334544 );
nand ( n44120 , n334545 , n309898 );
xnor ( n44121 , n334542 , n44120 );
nand ( n44122 , n44108 , n44121 );
buf ( n334549 , n44122 );
not ( n44124 , n334549 );
or ( n334551 , n328533 , n12778 );
not ( n334552 , n334551 );
not ( n334553 , n44112 );
not ( n334554 , n44120 );
or ( n44129 , n334553 , n334554 );
or ( n334556 , n44120 , n44112 );
nand ( n44131 , n44129 , n334556 );
not ( n334558 , n44131 );
or ( n334559 , n334552 , n334558 );
nand ( n44134 , n328533 , n12778 );
nand ( n334561 , n334559 , n44134 );
buf ( n334562 , n334561 );
xor ( n44137 , n44050 , n296368 );
not ( n44138 , n44137 );
not ( n44139 , n44138 );
and ( n44140 , n309897 , n44139 );
not ( n44141 , n309897 );
not ( n44142 , n44137 );
and ( n44143 , n44141 , n44142 );
or ( n44144 , n44140 , n44143 );
and ( n44145 , n334482 , n44144 );
not ( n44146 , n334482 );
not ( n44147 , n44138 );
and ( n44148 , n19468 , n44147 );
not ( n44149 , n19468 );
not ( n334576 , n44137 );
and ( n44151 , n44149 , n334576 );
or ( n44152 , n44148 , n44151 );
and ( n44153 , n44146 , n44152 );
or ( n44154 , n44145 , n44153 );
buf ( n334581 , n44154 );
nand ( n334582 , n334562 , n334581 );
buf ( n334583 , n334582 );
buf ( n334584 , n334583 );
not ( n334585 , n334584 );
or ( n44160 , n44124 , n334585 );
buf ( n334587 , n334561 );
buf ( n334588 , n44154 );
or ( n44163 , n334587 , n334588 );
buf ( n44164 , n44163 );
buf ( n334591 , n44164 );
nand ( n44166 , n44160 , n334591 );
buf ( n44167 , n44166 );
not ( n334594 , n44167 );
and ( n44169 , n334530 , n334594 );
not ( n334596 , n334525 );
nand ( n334597 , n334504 , n334502 );
and ( n44172 , n334597 , n334505 );
and ( n334599 , n334596 , n44172 );
not ( n334600 , n334509 );
not ( n334601 , n334508 );
or ( n334602 , n334600 , n334601 );
nand ( n44177 , n334602 , n334490 );
or ( n44178 , n334599 , n44177 );
or ( n334605 , n44172 , n334596 );
nand ( n334606 , n44178 , n334605 );
nor ( n44181 , n44169 , n334606 );
nand ( n334608 , n334455 , n334475 , n44181 );
buf ( n334609 , n334608 );
not ( n44184 , n17307 );
xor ( n334611 , n38777 , n16425 );
or ( n334612 , n44184 , n334611 );
not ( n44187 , n334611 );
or ( n334614 , n44187 , n17307 );
nand ( n44189 , n334612 , n334614 );
not ( n334616 , n44189 );
not ( n334617 , n334616 );
or ( n44192 , n38873 , n16421 );
not ( n44193 , n44192 );
not ( n334620 , n19443 );
not ( n334621 , n307500 );
or ( n44196 , n334620 , n334621 );
nand ( n334623 , n44196 , n309782 );
xnor ( n334624 , n334623 , n309895 );
not ( n44199 , n334624 );
or ( n334626 , n44193 , n44199 );
nand ( n334627 , n38873 , n16421 );
nand ( n44202 , n334626 , n334627 );
not ( n44203 , n44202 );
not ( n334630 , n44203 );
or ( n334631 , n334617 , n334630 );
xor ( n44206 , n38873 , n16421 );
and ( n334633 , n44206 , n334624 );
not ( n334634 , n44206 );
not ( n44209 , n334624 );
and ( n334636 , n334634 , n44209 );
nor ( n334637 , n334633 , n334636 );
not ( n44212 , n334637 );
not ( n334639 , n329794 );
not ( n334640 , n33553 );
not ( n44215 , n334640 );
or ( n334642 , n334639 , n44215 );
or ( n334643 , n334640 , n329794 );
nand ( n334644 , n17197 , n334643 );
nand ( n44219 , n334642 , n334644 );
not ( n334646 , n44219 );
nand ( n334647 , n44212 , n334646 );
nand ( n44222 , n334631 , n334647 );
nand ( n334649 , n44088 , n334516 );
not ( n334650 , n334649 );
not ( n44225 , n17094 );
or ( n334652 , n334650 , n44225 );
nand ( n334653 , n328638 , n328648 );
nand ( n44228 , n334652 , n334653 );
not ( n334655 , n329444 );
not ( n334656 , n39381 );
not ( n44231 , n307537 );
nand ( n44232 , n44231 , n17111 );
not ( n44233 , n44232 );
and ( n334660 , n334656 , n44233 );
and ( n44235 , n39381 , n44232 );
nor ( n334662 , n334660 , n44235 );
xor ( n334663 , n334655 , n334662 );
nor ( n334664 , n16429 , n306685 );
not ( n44239 , n334664 );
not ( n334666 , n307500 );
or ( n334667 , n44239 , n334666 );
and ( n334668 , n17088 , n16258 );
not ( n44243 , n16259 );
nor ( n334670 , n334668 , n44243 );
nand ( n44245 , n334667 , n334670 );
xnor ( n334672 , n334663 , n44245 );
or ( n44247 , n44228 , n334672 );
not ( n334674 , n329808 );
not ( n44249 , n329444 );
or ( n44250 , n334674 , n44249 );
not ( n44251 , n44232 );
or ( n44252 , n44245 , n44251 );
nand ( n44253 , n44245 , n44251 );
nand ( n44254 , n334655 , n39381 );
nand ( n44255 , n44252 , n44253 , n44254 );
nand ( n334682 , n44250 , n44255 );
not ( n44257 , n334682 );
xor ( n334684 , n334640 , n329794 );
and ( n334685 , n334684 , n17197 );
not ( n44260 , n334684 );
not ( n44261 , n17197 );
and ( n44262 , n44260 , n44261 );
nor ( n334689 , n334685 , n44262 );
not ( n334690 , n334689 );
nand ( n44265 , n44257 , n334690 );
nand ( n334692 , n44247 , n44265 );
nor ( n334693 , n44222 , n334692 );
not ( n44268 , n329091 );
not ( n334695 , n329867 );
nand ( n334696 , n44268 , n334695 );
not ( n44271 , n334696 );
not ( n334698 , n17263 );
nor ( n334699 , n19411 , n334698 );
not ( n44274 , n334699 );
not ( n334701 , n307500 );
or ( n334702 , n44274 , n334701 );
not ( n334703 , n334698 );
and ( n44278 , n334703 , n43098 );
not ( n44279 , n307690 );
nor ( n44280 , n44278 , n44279 );
nand ( n44281 , n334702 , n44280 );
nand ( n334708 , n308014 , n308009 );
not ( n334709 , n334708 );
and ( n44284 , n44281 , n334709 );
not ( n334711 , n44281 );
and ( n334712 , n334711 , n334708 );
nor ( n44287 , n44284 , n334712 );
not ( n334714 , n44287 );
or ( n334715 , n44271 , n334714 );
nand ( n44290 , n329867 , n329091 );
nand ( n334717 , n334715 , n44290 );
xor ( n334718 , n329088 , n329084 );
and ( n44293 , n334718 , n309900 );
not ( n334720 , n334718 );
not ( n334721 , n309900 );
and ( n44296 , n334720 , n334721 );
or ( n334723 , n44293 , n44296 );
nor ( n334724 , n19411 , n309939 );
not ( n44299 , n334724 );
not ( n334726 , n307500 );
or ( n44301 , n44299 , n334726 );
not ( n334728 , n43098 );
nor ( n334729 , n334728 , n309939 );
nor ( n334730 , n334729 , n309862 );
nand ( n44305 , n44301 , n334730 );
buf ( n334732 , n44305 );
and ( n334733 , n334723 , n334732 );
not ( n44308 , n334723 );
not ( n334735 , n334732 );
and ( n334736 , n44308 , n334735 );
nor ( n44311 , n334733 , n334736 );
nor ( n334738 , n334717 , n44311 );
not ( n334739 , n334738 );
or ( n44314 , n38777 , n16425 );
not ( n334741 , n44314 );
not ( n334742 , n17307 );
or ( n44317 , n334741 , n334742 );
nand ( n44318 , n38777 , n16425 );
nand ( n334745 , n44317 , n44318 );
not ( n334746 , n334745 );
and ( n44321 , n329091 , n334695 );
not ( n334748 , n329091 );
and ( n334749 , n334748 , n329867 );
or ( n44324 , n44321 , n334749 );
and ( n334751 , n44287 , n44324 );
not ( n334752 , n44287 );
not ( n44327 , n44324 );
and ( n334754 , n334752 , n44327 );
nor ( n44329 , n334751 , n334754 );
not ( n44330 , n44329 );
nand ( n334757 , n334746 , n44330 );
nand ( n44332 , n334739 , n334757 );
not ( n334759 , n309949 );
not ( n44334 , n334759 );
not ( n334761 , n19515 );
not ( n334762 , n307500 );
or ( n44337 , n334761 , n334762 );
and ( n334764 , n19513 , n307729 );
nor ( n334765 , n334764 , n309866 );
nand ( n44340 , n44337 , n334765 );
not ( n334767 , n44340 );
not ( n334768 , n334767 );
or ( n44343 , n44334 , n334768 );
nand ( n44344 , n44340 , n309949 );
nand ( n334771 , n44343 , n44344 );
not ( n44346 , n10429 );
not ( n334773 , n44346 );
nand ( n44348 , n334773 , n39184 );
or ( n334775 , n10429 , n39184 );
and ( n334776 , n44348 , n334775 );
not ( n44351 , n334776 );
and ( n334778 , n334771 , n44351 );
not ( n334779 , n334771 );
and ( n334780 , n334779 , n334776 );
nor ( n44355 , n334778 , n334780 );
not ( n44356 , n334721 );
xnor ( n334783 , n44305 , n44356 );
or ( n44358 , n329088 , n329084 );
and ( n334785 , n334783 , n44358 );
and ( n44360 , n329088 , n329084 );
nor ( n334787 , n334785 , n44360 );
nand ( n44362 , n44355 , n334787 );
nand ( n44363 , n44346 , n329611 );
not ( n44364 , n44363 );
not ( n334791 , n334771 );
or ( n334792 , n44364 , n334791 );
nand ( n44367 , n334792 , n44348 );
not ( n334794 , n44367 );
not ( n334795 , n43169 );
xnor ( n44370 , n39160 , n39168 );
not ( n334797 , n44370 );
not ( n334798 , n43168 );
or ( n334799 , n334797 , n334798 );
not ( n44374 , n44370 );
nand ( n44375 , n44374 , n18244 , n333593 );
nand ( n334802 , n334799 , n44375 );
not ( n334803 , n334802 );
or ( n44378 , n334795 , n334803 );
or ( n334805 , n43169 , n334802 );
nand ( n334806 , n44378 , n334805 );
nand ( n44381 , n334794 , n334806 );
nand ( n334808 , n44362 , n44381 );
nor ( n334809 , n44332 , n334808 );
nand ( n44384 , n334693 , n334809 );
not ( n334811 , n44384 );
buf ( n44386 , n334811 );
buf ( n334813 , n44121 );
buf ( n334814 , n44108 );
nor ( n334815 , n334813 , n334814 );
buf ( n334816 , n334815 );
buf ( n334817 , n334816 );
not ( n334818 , n334817 );
buf ( n334819 , n334818 );
nand ( n334820 , n44164 , n334819 );
nor ( n334821 , n44103 , n334820 );
not ( n334822 , n334821 );
nand ( n44397 , n334822 , n44181 );
buf ( n334824 , n44397 );
nand ( n334825 , n334609 , n44386 , n334824 );
buf ( n334826 , n334825 );
and ( n334827 , n44228 , n334672 );
nand ( n334828 , n44265 , n334827 );
nand ( n44403 , n334689 , n334682 );
nand ( n334830 , n334828 , n44403 );
not ( n334831 , n334830 );
not ( n44406 , n334616 );
not ( n334833 , n44203 );
or ( n334834 , n44406 , n334833 );
nand ( n44409 , n334834 , n334647 );
not ( n334836 , n44409 );
not ( n334837 , n334836 );
or ( n44412 , n334831 , n334837 );
and ( n334839 , n44219 , n334637 );
nand ( n334840 , n44203 , n334616 );
and ( n44415 , n334839 , n334840 );
buf ( n44416 , n44202 );
buf ( n44417 , n44189 );
and ( n44418 , n44416 , n44417 );
buf ( n44419 , n44418 );
nor ( n334846 , n44415 , n44419 );
nand ( n44421 , n44412 , n334846 );
nand ( n334848 , n44421 , n334809 );
buf ( n334849 , n334848 );
buf ( n334850 , n334808 );
not ( n334851 , n334850 );
buf ( n334852 , n334851 );
not ( n334853 , n334852 );
nand ( n44428 , n44329 , n334745 );
nor ( n334855 , n334717 , n44311 );
or ( n334856 , n44428 , n334855 );
nand ( n44431 , n334717 , n44311 );
nand ( n334858 , n334856 , n44431 );
not ( n334859 , n334858 );
or ( n44434 , n334853 , n334859 );
nor ( n334861 , n334787 , n44355 );
and ( n334862 , n334861 , n44381 );
not ( n44437 , n44367 );
nor ( n334864 , n334806 , n44437 );
nor ( n334865 , n334862 , n334864 );
nand ( n334866 , n44434 , n334865 );
buf ( n44441 , n334866 );
not ( n44442 , n44441 );
buf ( n334869 , n44442 );
buf ( n334870 , n334869 );
and ( n334871 , n334849 , n334870 );
buf ( n334872 , n334871 );
nand ( n44447 , n334826 , n334872 );
not ( n44448 , n44447 );
or ( n334875 , n333798 , n44448 );
buf ( n334876 , n43088 );
not ( n44451 , n334876 );
buf ( n44452 , n44451 );
buf ( n334879 , n44452 );
not ( n334880 , n334879 );
not ( n44455 , n43212 );
nand ( n44456 , n43166 , n333600 );
or ( n334883 , n333573 , n44456 );
buf ( n334884 , n43144 );
buf ( n334885 , n333534 );
nand ( n334886 , n334884 , n334885 );
buf ( n334887 , n334886 );
nand ( n334888 , n334883 , n334887 );
not ( n334889 , n334888 );
or ( n334890 , n44455 , n334889 );
nor ( n44465 , n333609 , n43192 );
and ( n44466 , n44465 , n43210 );
nor ( n44467 , n43202 , n43209 );
nor ( n44468 , n44466 , n44467 );
nand ( n44469 , n334890 , n44468 );
buf ( n334896 , n44469 );
buf ( n334897 , n334896 );
not ( n334898 , n334897 );
or ( n334899 , n334880 , n334898 );
buf ( n334900 , n43087 );
not ( n44475 , n334900 );
not ( n334902 , n43028 );
buf ( n44477 , n42968 );
buf ( n44478 , n42991 );
and ( n44479 , n44477 , n44478 );
buf ( n44480 , n44479 );
not ( n334907 , n44480 );
or ( n44482 , n334902 , n334907 );
not ( n334909 , n43027 );
nand ( n334910 , n334909 , n43009 );
nand ( n44485 , n44482 , n334910 );
buf ( n334912 , n44485 );
not ( n334913 , n334912 );
or ( n334914 , n44475 , n334913 );
nor ( n334915 , n43049 , n43058 );
nand ( n44490 , n333511 , n43078 );
and ( n334917 , n334915 , n44490 );
not ( n44492 , n43078 );
nand ( n44493 , n44492 , n333510 );
not ( n44494 , n44493 );
nor ( n334921 , n334917 , n44494 );
buf ( n334922 , n334921 );
nand ( n44497 , n334914 , n334922 );
buf ( n334924 , n44497 );
buf ( n334925 , n334924 );
not ( n334926 , n334925 );
buf ( n334927 , n334926 );
buf ( n334928 , n334927 );
nand ( n334929 , n334899 , n334928 );
buf ( n334930 , n334929 );
buf ( n334931 , n333796 );
not ( n334932 , n334931 );
buf ( n334933 , n334932 );
and ( n334934 , n334930 , n334933 );
buf ( n334935 , n43246 );
not ( n334936 , n334935 );
and ( n334937 , n333793 , n43343 );
not ( n44512 , n334937 );
not ( n334939 , n333723 );
nor ( n334940 , n333727 , n43307 );
not ( n334941 , n334940 );
or ( n334942 , n334939 , n334941 );
not ( n44517 , n333722 );
nand ( n334944 , n44517 , n333689 );
nand ( n44519 , n334942 , n334944 );
not ( n334946 , n44519 );
or ( n334947 , n44512 , n334946 );
buf ( n334948 , n43343 );
nor ( n44523 , n43353 , n333790 );
and ( n334950 , n334948 , n44523 );
and ( n334951 , n333752 , n333767 );
nor ( n44526 , n334950 , n334951 );
nand ( n44527 , n334947 , n44526 );
buf ( n334954 , n44527 );
buf ( n44529 , n334954 );
buf ( n334956 , n44529 );
buf ( n334957 , n334956 );
not ( n334958 , n334957 );
or ( n44533 , n334936 , n334958 );
nor ( n334960 , n43224 , n43245 );
buf ( n334961 , n334960 );
not ( n44536 , n334961 );
buf ( n44537 , n44536 );
buf ( n334964 , n44537 );
nand ( n44539 , n44533 , n334964 );
buf ( n44540 , n44539 );
nor ( n334967 , n334934 , n44540 );
nand ( n44542 , n334875 , n334967 );
buf ( n334969 , n44542 );
and ( n334970 , n334969 , n333374 );
not ( n44545 , n334969 );
and ( n334972 , n44545 , n333370 );
nor ( n334973 , n334970 , n334972 );
buf ( n334974 , n334973 );
buf ( n334975 , n334944 );
buf ( n44550 , n333723 );
nand ( n334977 , n334975 , n44550 );
buf ( n334978 , n334977 );
buf ( n334979 , n334977 );
not ( n334980 , n334979 );
buf ( n334981 , n334980 );
buf ( n334982 , n334981 );
buf ( n334983 , n43308 );
not ( n334984 , n334983 );
buf ( n44559 , n43214 );
nor ( n44560 , n334984 , n44559 );
buf ( n44561 , n44560 );
buf ( n334988 , n44561 );
not ( n44563 , n334988 );
buf ( n334990 , n44447 );
not ( n334991 , n334990 );
or ( n44566 , n44563 , n334991 );
buf ( n334993 , n334930 );
buf ( n334994 , n43308 );
and ( n334995 , n334993 , n334994 );
buf ( n334996 , n334940 );
nor ( n334997 , n334995 , n334996 );
buf ( n334998 , n334997 );
buf ( n334999 , n334998 );
nand ( n335000 , n44566 , n334999 );
buf ( n335001 , n335000 );
buf ( n335002 , n335001 );
and ( n335003 , n335002 , n334982 );
not ( n335004 , n335002 );
and ( n44579 , n335004 , n334978 );
nor ( n335006 , n335003 , n44579 );
buf ( n335007 , n335006 );
not ( n44582 , n33986 );
not ( n335009 , n309886 );
not ( n335010 , n19504 );
or ( n44585 , n335009 , n335010 );
or ( n335012 , n19504 , n309886 );
nand ( n335013 , n44585 , n335012 );
not ( n44588 , n335013 );
or ( n335015 , n44582 , n44588 );
nand ( n335016 , n33979 , n324411 );
nand ( n335017 , n335015 , n335016 );
xor ( n44592 , n34002 , n33997 );
not ( n335019 , n309890 );
not ( n335020 , n335019 );
nor ( n335021 , n309808 , n19213 );
nand ( n44596 , n309807 , n335021 );
not ( n335023 , n44596 );
nand ( n335024 , n335023 , n18214 );
and ( n335025 , n309921 , n335021 );
nor ( n44600 , n335025 , n19277 );
buf ( n335027 , n44600 );
not ( n335028 , n309822 );
not ( n44603 , n44596 );
nand ( n335030 , n307500 , n335028 , n44603 );
nand ( n335031 , n335024 , n335027 , n335030 );
not ( n44606 , n335031 );
or ( n335033 , n335020 , n44606 );
and ( n335034 , n335030 , n309890 );
nand ( n44609 , n335034 , n335024 , n335027 );
nand ( n335036 , n335033 , n44609 );
xnor ( n335037 , n44592 , n335036 );
and ( n44612 , n335017 , n335037 );
buf ( n335039 , n44612 );
not ( n335040 , n335039 );
buf ( n335041 , n335040 );
not ( n335042 , n335017 );
not ( n44617 , n335037 );
nand ( n335044 , n335042 , n44617 );
buf ( n335045 , n335044 );
nand ( n44620 , n335041 , n335045 );
buf ( n335047 , n44620 );
buf ( n44622 , n44620 );
not ( n335049 , n44622 );
buf ( n335050 , n335049 );
buf ( n335051 , n335050 );
nand ( n335052 , n43344 , n43368 );
not ( n335053 , n335052 );
xor ( n335054 , n33979 , n324411 );
not ( n44629 , n335054 );
not ( n335056 , n44629 );
and ( n335057 , n19459 , n335056 );
not ( n44632 , n19459 );
not ( n335059 , n335054 );
and ( n335060 , n44632 , n335059 );
or ( n44635 , n335057 , n335060 );
and ( n335062 , n19504 , n44635 );
not ( n335063 , n19504 );
not ( n44638 , n44629 );
and ( n335065 , n309886 , n44638 );
not ( n335066 , n309886 );
not ( n44641 , n335054 );
and ( n44642 , n335066 , n44641 );
or ( n335069 , n335065 , n44642 );
and ( n44644 , n335063 , n335069 );
or ( n335071 , n335062 , n44644 );
not ( n44646 , n335071 );
not ( n335073 , n33975 );
not ( n335074 , n309892 );
nand ( n44649 , n42973 , n309826 );
and ( n335076 , n309923 , n19396 );
nor ( n335077 , n335076 , n309860 );
nand ( n335078 , n44649 , n335077 , n19506 );
not ( n44653 , n335078 );
or ( n335080 , n335074 , n44653 );
not ( n335081 , n309892 );
nand ( n44656 , n335081 , n44649 , n335077 , n19506 );
nand ( n335083 , n335080 , n44656 );
not ( n335084 , n335083 );
or ( n44659 , n335073 , n335084 );
nand ( n335086 , n44659 , n34037 );
not ( n335087 , n335086 );
nand ( n44662 , n44646 , n335087 );
or ( n44663 , n34039 , n33958 );
nand ( n335090 , n44663 , n19476 );
not ( n44665 , n335090 );
not ( n335092 , n44665 );
not ( n44667 , n42929 );
not ( n335094 , n44667 );
or ( n335095 , n335092 , n335094 );
nand ( n44670 , n335095 , n34040 );
not ( n335097 , n44670 );
not ( n335098 , n44667 );
not ( n44673 , n44663 );
nor ( n44674 , n44673 , n19476 );
nand ( n335101 , n335098 , n42927 , n42926 , n44674 );
not ( n335102 , n42927 );
nand ( n44677 , n335102 , n44665 );
or ( n335104 , n42926 , n335090 );
nand ( n335105 , n335097 , n335101 , n44677 , n335104 );
not ( n44680 , n335105 );
xnor ( n335107 , n324395 , n324400 );
not ( n335108 , n335107 );
not ( n44683 , n309892 );
and ( n335110 , n335108 , n44683 );
and ( n44685 , n335107 , n309892 );
nor ( n335112 , n335110 , n44685 );
and ( n44687 , n335078 , n335112 );
not ( n335114 , n335078 );
not ( n335115 , n335112 );
and ( n44690 , n335114 , n335115 );
nor ( n335117 , n44687 , n44690 );
not ( n335118 , n335117 );
nand ( n335119 , n44680 , n335118 );
and ( n44694 , n43246 , n44662 , n335119 , n42938 );
nand ( n335121 , n335053 , n44694 );
buf ( n335122 , n335121 );
not ( n44697 , n335122 );
buf ( n335124 , n44697 );
not ( n335125 , n335124 );
nor ( n44700 , n334866 , n44469 );
nand ( n335127 , n334848 , n44700 );
not ( n335128 , n335127 );
nor ( n44703 , n44469 , n43213 );
nor ( n335130 , n44703 , n43088 );
not ( n335131 , n335130 );
or ( n44706 , n335128 , n335131 );
nand ( n44707 , n44706 , n334927 );
buf ( n335134 , n44707 );
buf ( n335135 , n335134 );
not ( n44710 , n335135 );
or ( n335137 , n335125 , n44710 );
and ( n335138 , n43859 , n334417 , n334451 );
or ( n44713 , n333919 , n334004 );
nor ( n335140 , n44713 , n44103 );
not ( n335141 , n334820 );
nand ( n44716 , n335138 , n335140 , n335141 );
buf ( n335143 , n334364 );
not ( n44718 , n335143 );
buf ( n335145 , n44718 );
nand ( n335146 , n44026 , n335145 , n334821 );
not ( n44721 , n44045 );
not ( n335148 , n44039 );
or ( n44723 , n44721 , n335148 );
nand ( n335150 , n44723 , n334821 );
nand ( n44725 , n44716 , n335146 , n44181 , n335150 );
buf ( n335152 , n44725 );
buf ( n335153 , n335152 );
buf ( n335154 , n43176 );
buf ( n335155 , n43212 );
nand ( n44730 , n43087 , n335154 , n43029 , n335155 );
nor ( n335157 , n44384 , n44730 );
buf ( n335158 , n335157 );
buf ( n335159 , n335158 );
buf ( n335160 , n44697 );
and ( n335161 , n335153 , n335159 , n335160 );
not ( n335162 , n44694 );
not ( n44737 , n44527 );
or ( n335164 , n335162 , n44737 );
buf ( n335165 , n334960 );
not ( n335166 , n335165 );
buf ( n335167 , n42938 );
not ( n44742 , n335167 );
or ( n335169 , n335166 , n44742 );
buf ( n335170 , n42940 );
nand ( n335171 , n335169 , n335170 );
buf ( n335172 , n335171 );
and ( n335173 , n44662 , n335119 );
and ( n44748 , n335172 , n335173 );
buf ( n335175 , n44662 );
not ( n335176 , n335175 );
buf ( n335177 , n335176 );
nand ( n335178 , n335117 , n335105 );
or ( n335179 , n335177 , n335178 );
nand ( n44754 , n335071 , n335086 );
nand ( n335181 , n335179 , n44754 );
nor ( n44756 , n44748 , n335181 );
nand ( n335183 , n335164 , n44756 );
buf ( n335184 , n335183 );
buf ( n335185 , n335184 );
nor ( n335186 , n335161 , n335185 );
buf ( n335187 , n335186 );
buf ( n335188 , n335187 );
nand ( n44763 , n335137 , n335188 );
buf ( n335190 , n44763 );
buf ( n335191 , n335190 );
and ( n335192 , n335191 , n335051 );
not ( n44767 , n335191 );
and ( n335194 , n44767 , n335047 );
nor ( n335195 , n335192 , n335194 );
buf ( n335196 , n335195 );
buf ( n335197 , n44662 );
buf ( n335198 , n44754 );
nand ( n335199 , n335197 , n335198 );
buf ( n335200 , n335199 );
buf ( n335201 , n335200 );
buf ( n335202 , n335200 );
not ( n44777 , n335202 );
buf ( n335204 , n44777 );
buf ( n335205 , n335204 );
buf ( n335206 , n335119 );
not ( n44781 , n335206 );
nand ( n335208 , n43246 , n42938 );
buf ( n44783 , n335208 );
nor ( n44784 , n44781 , n44783 );
buf ( n44785 , n44784 );
buf ( n335212 , n44785 );
not ( n44787 , n335212 );
not ( n335214 , n335052 );
not ( n44789 , n335214 );
buf ( n335216 , n44789 );
nor ( n335217 , n44787 , n335216 );
buf ( n335218 , n335217 );
buf ( n335219 , n335218 );
not ( n335220 , n335219 );
buf ( n335221 , n335134 );
not ( n44796 , n335221 );
or ( n335223 , n335220 , n44796 );
buf ( n335224 , n44725 );
buf ( n335225 , n335224 );
buf ( n335226 , n335158 );
buf ( n335227 , n335218 );
and ( n44802 , n335225 , n335226 , n335227 );
buf ( n335229 , n44785 );
not ( n335230 , n335229 );
buf ( n335231 , n334956 );
not ( n44806 , n335231 );
or ( n44807 , n335230 , n44806 );
not ( n44808 , n335119 );
not ( n335235 , n335172 );
or ( n335236 , n44808 , n335235 );
nand ( n44811 , n335236 , n335178 );
buf ( n335238 , n44811 );
not ( n44813 , n335238 );
buf ( n44814 , n44813 );
buf ( n335241 , n44814 );
nand ( n335242 , n44807 , n335241 );
buf ( n335243 , n335242 );
buf ( n335244 , n335243 );
nor ( n335245 , n44802 , n335244 );
buf ( n335246 , n335245 );
buf ( n335247 , n335246 );
nand ( n44822 , n335223 , n335247 );
buf ( n335249 , n44822 );
buf ( n335250 , n335249 );
and ( n335251 , n335250 , n335205 );
not ( n44826 , n335250 );
and ( n44827 , n44826 , n335201 );
nor ( n335254 , n335251 , n44827 );
buf ( n335255 , n335254 );
nand ( n335256 , n335119 , n335178 );
buf ( n335257 , n335256 );
buf ( n335258 , n335256 );
not ( n44833 , n335258 );
buf ( n335260 , n44833 );
buf ( n335261 , n335260 );
not ( n335262 , n335208 );
not ( n335263 , n335262 );
nor ( n335264 , n335263 , n44789 );
buf ( n335265 , n335264 );
not ( n335266 , n335265 );
buf ( n335267 , n335134 );
not ( n335268 , n335267 );
or ( n335269 , n335266 , n335268 );
buf ( n335270 , n335224 );
buf ( n335271 , n335158 );
buf ( n335272 , n335264 );
and ( n335273 , n335270 , n335271 , n335272 );
buf ( n335274 , n335262 );
not ( n44849 , n335274 );
buf ( n335276 , n334956 );
not ( n44851 , n335276 );
or ( n335278 , n44849 , n44851 );
buf ( n335279 , n335172 );
not ( n44854 , n335279 );
buf ( n44855 , n44854 );
buf ( n335282 , n44855 );
nand ( n44857 , n335278 , n335282 );
buf ( n335284 , n44857 );
buf ( n335285 , n335284 );
nor ( n44860 , n335273 , n335285 );
buf ( n44861 , n44860 );
buf ( n44862 , n44861 );
nand ( n44863 , n335269 , n44862 );
buf ( n44864 , n44863 );
buf ( n335291 , n44864 );
and ( n44866 , n335291 , n335261 );
not ( n44867 , n335291 );
and ( n335294 , n44867 , n335257 );
nor ( n44869 , n44866 , n335294 );
buf ( n44870 , n44869 );
buf ( n335297 , n43246 );
buf ( n335298 , n44537 );
nand ( n335299 , n335297 , n335298 );
buf ( n335300 , n335299 );
buf ( n335301 , n335300 );
buf ( n335302 , n335300 );
not ( n44877 , n335302 );
buf ( n335304 , n44877 );
buf ( n335305 , n335304 );
not ( n335306 , n335214 );
not ( n335307 , n335134 );
or ( n44882 , n335306 , n335307 );
and ( n44883 , n335152 , n335158 , n335214 );
nor ( n44884 , n44883 , n334956 );
nand ( n44885 , n44882 , n44884 );
buf ( n335312 , n44885 );
and ( n44887 , n335312 , n335305 );
not ( n335314 , n335312 );
and ( n44889 , n335314 , n335301 );
nor ( n335316 , n44887 , n44889 );
buf ( n335317 , n335316 );
buf ( n335318 , n334951 );
not ( n44893 , n335318 );
buf ( n335320 , n334948 );
nand ( n44895 , n44893 , n335320 );
buf ( n44896 , n44895 );
buf ( n44897 , n44896 );
buf ( n335324 , n44896 );
not ( n335325 , n335324 );
buf ( n335326 , n335325 );
buf ( n335327 , n335326 );
not ( n44902 , n333795 );
buf ( n335329 , n44902 );
nand ( n335330 , n43308 , n333723 );
buf ( n335331 , n335330 );
nor ( n335332 , n335329 , n335331 );
buf ( n335333 , n335332 );
buf ( n335334 , n335333 );
not ( n335335 , n335334 );
buf ( n335336 , n335134 );
not ( n335337 , n335336 );
or ( n335338 , n335335 , n335337 );
buf ( n335339 , n335152 );
buf ( n335340 , n335158 );
buf ( n335341 , n335333 );
and ( n335342 , n335339 , n335340 , n335341 );
buf ( n335343 , n44519 );
not ( n44918 , n335343 );
buf ( n335345 , n44918 );
buf ( n335346 , n335345 );
buf ( n335347 , n44902 );
or ( n335348 , n335346 , n335347 );
buf ( n335349 , n44523 );
not ( n335350 , n335349 );
buf ( n335351 , n335350 );
buf ( n335352 , n335351 );
nand ( n335353 , n335348 , n335352 );
buf ( n335354 , n335353 );
buf ( n335355 , n335354 );
nor ( n335356 , n335342 , n335355 );
buf ( n335357 , n335356 );
buf ( n335358 , n335357 );
nand ( n44933 , n335338 , n335358 );
buf ( n335360 , n44933 );
buf ( n335361 , n335360 );
and ( n335362 , n335361 , n335327 );
not ( n335363 , n335361 );
and ( n335364 , n335363 , n44897 );
nor ( n44939 , n335362 , n335364 );
buf ( n44940 , n44939 );
buf ( n335367 , n44902 );
buf ( n44942 , n44523 );
buf ( n335369 , n44942 );
nor ( n44944 , n335367 , n335369 );
buf ( n335371 , n44944 );
buf ( n335372 , n335371 );
not ( n335373 , n335372 );
buf ( n335374 , n335373 );
buf ( n335375 , n335374 );
buf ( n335376 , n335371 );
buf ( n335377 , n335330 );
not ( n44952 , n335377 );
buf ( n335379 , n44952 );
buf ( n335380 , n335379 );
not ( n335381 , n335380 );
buf ( n335382 , n335134 );
not ( n44957 , n335382 );
or ( n335384 , n335381 , n44957 );
buf ( n335385 , n335152 );
buf ( n335386 , n335158 );
buf ( n335387 , n335379 );
and ( n44962 , n335385 , n335386 , n335387 );
buf ( n335389 , n335345 );
not ( n44964 , n335389 );
buf ( n44965 , n44964 );
buf ( n335392 , n44965 );
nor ( n335393 , n44962 , n335392 );
buf ( n335394 , n335393 );
buf ( n335395 , n335394 );
nand ( n44970 , n335384 , n335395 );
buf ( n335397 , n44970 );
buf ( n335398 , n335397 );
and ( n335399 , n335398 , n335376 );
not ( n335400 , n335398 );
and ( n44975 , n335400 , n335375 );
nor ( n44976 , n335399 , n44975 );
buf ( n335403 , n44976 );
not ( n44978 , n44465 );
buf ( n335405 , n43193 );
buf ( n335406 , n335405 );
buf ( n335407 , n335406 );
nand ( n335408 , n44978 , n335407 );
buf ( n335409 , n335408 );
buf ( n335410 , n335408 );
not ( n44985 , n335410 );
buf ( n335412 , n44985 );
buf ( n335413 , n335412 );
not ( n44988 , n334811 );
buf ( n335415 , n44988 );
nor ( n335416 , n333573 , n333601 );
buf ( n335417 , n335416 );
not ( n335418 , n335417 );
buf ( n335419 , n335418 );
buf ( n335420 , n335419 );
nor ( n335421 , n335415 , n335420 );
buf ( n335422 , n335421 );
buf ( n335423 , n335422 );
not ( n44998 , n335423 );
buf ( n335425 , n335224 );
not ( n335426 , n335425 );
or ( n335427 , n44998 , n335426 );
not ( n45002 , n334872 );
and ( n335429 , n45002 , n335416 );
buf ( n335430 , n334888 );
nor ( n335431 , n335429 , n335430 );
buf ( n45006 , n335431 );
nand ( n45007 , n335427 , n45006 );
buf ( n335434 , n45007 );
buf ( n335435 , n335434 );
and ( n45010 , n335435 , n335413 );
not ( n335437 , n335435 );
and ( n335438 , n335437 , n335409 );
nor ( n335439 , n45010 , n335438 );
buf ( n335440 , n335439 );
buf ( n335441 , n44467 );
not ( n45016 , n335441 );
buf ( n335443 , n43210 );
nand ( n45018 , n45016 , n335443 );
buf ( n335445 , n45018 );
buf ( n335446 , n335445 );
buf ( n335447 , n335445 );
not ( n335448 , n335447 );
buf ( n335449 , n335448 );
buf ( n335450 , n335449 );
buf ( n335451 , n335407 );
not ( n45026 , n335451 );
buf ( n335453 , n335419 );
nor ( n45028 , n45026 , n335453 );
buf ( n335455 , n45028 );
buf ( n335456 , n335455 );
not ( n335457 , n335456 );
buf ( n335458 , n44384 );
nor ( n45033 , n335457 , n335458 );
buf ( n335460 , n45033 );
buf ( n335461 , n335460 );
not ( n45036 , n335461 );
buf ( n335463 , n335224 );
not ( n335464 , n335463 );
or ( n335465 , n45036 , n335464 );
buf ( n335466 , n335455 );
buf ( n335467 , n45002 );
and ( n335468 , n335466 , n335467 );
not ( n335469 , n44465 );
nand ( n45044 , n335407 , n335430 );
nand ( n335471 , n335469 , n45044 );
buf ( n335472 , n335471 );
nor ( n335473 , n335468 , n335472 );
buf ( n335474 , n335473 );
buf ( n335475 , n335474 );
nand ( n335476 , n335465 , n335475 );
buf ( n335477 , n335476 );
buf ( n335478 , n335477 );
and ( n45053 , n335478 , n335450 );
not ( n335480 , n335478 );
and ( n335481 , n335480 , n335446 );
nor ( n45056 , n45053 , n335481 );
buf ( n335483 , n45056 );
buf ( n335484 , n43308 );
not ( n45059 , n335484 );
buf ( n335486 , n334940 );
nor ( n335487 , n45059 , n335486 );
buf ( n335488 , n335487 );
buf ( n45063 , n335488 );
not ( n45064 , n45063 );
buf ( n45065 , n45064 );
buf ( n335492 , n45065 );
buf ( n335493 , n335488 );
not ( n45068 , n335158 );
not ( n45069 , n335224 );
or ( n45070 , n45068 , n45069 );
not ( n335497 , n335134 );
nand ( n335498 , n45070 , n335497 );
buf ( n335499 , n335498 );
and ( n335500 , n335499 , n335493 );
not ( n335501 , n335499 );
and ( n335502 , n335501 , n335492 );
nor ( n335503 , n335500 , n335502 );
buf ( n335504 , n335503 );
nand ( n45079 , n44493 , n44490 );
buf ( n335506 , n45079 );
buf ( n335507 , n45079 );
not ( n335508 , n335507 );
buf ( n335509 , n335508 );
buf ( n45084 , n335509 );
and ( n45085 , n42995 , n43028 );
buf ( n335512 , n45085 );
buf ( n335513 , n43059 );
and ( n335514 , n335512 , n335513 );
buf ( n335515 , n335514 );
buf ( n335516 , n335515 );
buf ( n335517 , n43213 );
buf ( n45092 , n335517 );
buf ( n335519 , n45092 );
buf ( n335520 , n335519 );
nand ( n45095 , n335516 , n335520 );
buf ( n45096 , n45095 );
buf ( n335523 , n45096 );
buf ( n335524 , n44988 );
nor ( n45099 , n335523 , n335524 );
buf ( n45100 , n45099 );
buf ( n45101 , n45100 );
not ( n45102 , n45101 );
buf ( n45103 , n335224 );
not ( n45104 , n45103 );
or ( n45105 , n45102 , n45104 );
buf ( n335532 , n45002 );
buf ( n335533 , n45096 );
not ( n335534 , n335533 );
buf ( n335535 , n335534 );
buf ( n335536 , n335535 );
and ( n335537 , n335532 , n335536 );
buf ( n335538 , n335515 );
not ( n335539 , n335538 );
buf ( n335540 , n334896 );
not ( n45115 , n335540 );
or ( n45116 , n335539 , n45115 );
buf ( n335543 , n43059 );
not ( n335544 , n335543 );
buf ( n335545 , n44485 );
not ( n335546 , n335545 );
or ( n335547 , n335544 , n335546 );
buf ( n335548 , n334915 );
not ( n45123 , n335548 );
buf ( n335550 , n45123 );
buf ( n335551 , n335550 );
nand ( n335552 , n335547 , n335551 );
buf ( n335553 , n335552 );
buf ( n335554 , n335553 );
not ( n45129 , n335554 );
buf ( n45130 , n45129 );
buf ( n335557 , n45130 );
nand ( n335558 , n45116 , n335557 );
buf ( n335559 , n335558 );
buf ( n335560 , n335559 );
nor ( n45135 , n335537 , n335560 );
buf ( n335562 , n45135 );
buf ( n335563 , n335562 );
nand ( n45138 , n45105 , n335563 );
buf ( n335565 , n45138 );
buf ( n335566 , n335565 );
and ( n335567 , n335566 , n45084 );
not ( n45142 , n335566 );
and ( n335569 , n45142 , n335506 );
nor ( n335570 , n335567 , n335569 );
buf ( n335571 , n335570 );
nand ( n335572 , n334910 , n43028 );
buf ( n335573 , n335572 );
buf ( n335574 , n335572 );
not ( n45149 , n335574 );
buf ( n335576 , n45149 );
buf ( n335577 , n335576 );
buf ( n335578 , n44988 );
buf ( n335579 , n335519 );
buf ( n45154 , n42995 );
buf ( n335581 , n45154 );
buf ( n335582 , n335581 );
buf ( n335583 , n335582 );
nand ( n335584 , n335579 , n335583 );
buf ( n335585 , n335584 );
buf ( n335586 , n335585 );
nor ( n45161 , n335578 , n335586 );
buf ( n335588 , n45161 );
buf ( n335589 , n335588 );
not ( n45164 , n335589 );
buf ( n335591 , n335224 );
not ( n335592 , n335591 );
or ( n335593 , n45164 , n335592 );
buf ( n335594 , n335585 );
not ( n335595 , n335594 );
buf ( n335596 , n335595 );
buf ( n335597 , n335596 );
buf ( n335598 , n45002 );
and ( n45173 , n335597 , n335598 );
buf ( n335600 , n335582 );
not ( n335601 , n335600 );
buf ( n335602 , n334896 );
not ( n45177 , n335602 );
or ( n45178 , n335601 , n45177 );
buf ( n335605 , n44480 );
not ( n45180 , n335605 );
buf ( n45181 , n45180 );
buf ( n335608 , n45181 );
nand ( n335609 , n45178 , n335608 );
buf ( n335610 , n335609 );
buf ( n335611 , n335610 );
nor ( n335612 , n45173 , n335611 );
buf ( n335613 , n335612 );
buf ( n45188 , n335613 );
nand ( n335615 , n335593 , n45188 );
buf ( n335616 , n335615 );
buf ( n335617 , n335616 );
and ( n45192 , n335617 , n335577 );
not ( n45193 , n335617 );
and ( n45194 , n45193 , n335573 );
nor ( n335621 , n45192 , n45194 );
buf ( n335622 , n335621 );
buf ( n335623 , n335582 );
buf ( n45198 , n45181 );
nand ( n45199 , n335623 , n45198 );
buf ( n45200 , n45199 );
buf ( n335627 , n45200 );
buf ( n335628 , n45200 );
not ( n45203 , n335628 );
buf ( n335630 , n45203 );
buf ( n335631 , n335630 );
buf ( n335632 , n335519 );
not ( n335633 , n335632 );
buf ( n335634 , n44384 );
nor ( n335635 , n335633 , n335634 );
buf ( n335636 , n335635 );
buf ( n335637 , n335636 );
not ( n45212 , n335637 );
buf ( n335639 , n335224 );
not ( n45214 , n335639 );
or ( n335641 , n45212 , n45214 );
buf ( n335642 , n45002 );
buf ( n335643 , n335519 );
and ( n45218 , n335642 , n335643 );
buf ( n335645 , n334896 );
nor ( n335646 , n45218 , n335645 );
buf ( n335647 , n335646 );
buf ( n335648 , n335647 );
nand ( n45223 , n335641 , n335648 );
buf ( n45224 , n45223 );
buf ( n335651 , n45224 );
and ( n45226 , n335651 , n335631 );
not ( n335653 , n335651 );
and ( n335654 , n335653 , n335627 );
nor ( n45229 , n45226 , n335654 );
buf ( n335656 , n45229 );
buf ( n45231 , n44403 );
nand ( n335658 , n44265 , n45231 );
buf ( n335659 , n335658 );
buf ( n335660 , n335658 );
not ( n335661 , n335660 );
buf ( n335662 , n335661 );
buf ( n335663 , n335662 );
buf ( n335664 , n44247 );
not ( n45239 , n335664 );
buf ( n335666 , n335224 );
not ( n335667 , n335666 );
or ( n335668 , n45239 , n335667 );
buf ( n335669 , n44228 );
buf ( n45244 , n334672 );
nand ( n45245 , n335669 , n45244 );
buf ( n45246 , n45245 );
buf ( n335673 , n45246 );
nand ( n335674 , n335668 , n335673 );
buf ( n335675 , n335674 );
buf ( n335676 , n335675 );
and ( n45251 , n335676 , n335663 );
not ( n45252 , n335676 );
and ( n45253 , n45252 , n335659 );
nor ( n45254 , n45251 , n45253 );
buf ( n335681 , n45254 );
buf ( n335682 , n44456 );
not ( n335683 , n333601 );
buf ( n335684 , n335683 );
nand ( n335685 , n335682 , n335684 );
buf ( n335686 , n335685 );
buf ( n335687 , n335686 );
buf ( n45262 , n44447 );
buf ( n45263 , n335686 );
buf ( n45264 , n44447 );
not ( n45265 , n335687 );
not ( n45266 , n45262 );
or ( n45267 , n45265 , n45266 );
or ( n45268 , n45263 , n45264 );
nand ( n45269 , n45267 , n45268 );
buf ( n45270 , n45269 );
not ( n335697 , n334864 );
nand ( n335698 , n335697 , n44381 );
buf ( n335699 , n335698 );
buf ( n335700 , n335698 );
not ( n335701 , n335700 );
buf ( n335702 , n335701 );
buf ( n335703 , n335702 );
buf ( n335704 , n334693 );
buf ( n45279 , n335704 );
buf ( n45280 , n45279 );
buf ( n335707 , n45280 );
not ( n335708 , n335707 );
buf ( n335709 , n44332 );
not ( n45284 , n335709 );
buf ( n335711 , n45284 );
buf ( n335712 , n335711 );
buf ( n45287 , n44362 );
buf ( n335714 , n45287 );
nand ( n335715 , n335712 , n335714 );
buf ( n335716 , n335715 );
buf ( n45291 , n335716 );
nor ( n45292 , n335708 , n45291 );
buf ( n45293 , n45292 );
buf ( n45294 , n45293 );
not ( n335721 , n45294 );
buf ( n335722 , n335224 );
not ( n45297 , n335722 );
or ( n335724 , n335721 , n45297 );
buf ( n335725 , n335716 );
not ( n335726 , n335725 );
buf ( n335727 , n335726 );
buf ( n335728 , n44421 );
and ( n45303 , n335727 , n335728 );
buf ( n335730 , n45287 );
not ( n335731 , n335730 );
buf ( n335732 , n334858 );
not ( n335733 , n335732 );
or ( n45308 , n335731 , n335733 );
buf ( n335735 , n334861 );
not ( n335736 , n335735 );
buf ( n335737 , n335736 );
buf ( n335738 , n335737 );
nand ( n45313 , n45308 , n335738 );
buf ( n335740 , n45313 );
nor ( n45315 , n45303 , n335740 );
buf ( n335742 , n45315 );
nand ( n45317 , n335724 , n335742 );
buf ( n45318 , n45317 );
buf ( n335745 , n45318 );
and ( n335746 , n335745 , n335703 );
not ( n45321 , n335745 );
and ( n335748 , n45321 , n335699 );
nor ( n335749 , n335746 , n335748 );
buf ( n335750 , n335749 );
buf ( n335751 , n45287 );
buf ( n335752 , n335737 );
nand ( n45327 , n335751 , n335752 );
buf ( n335754 , n45327 );
buf ( n335755 , n335754 );
buf ( n335756 , n335754 );
not ( n45331 , n335756 );
buf ( n45332 , n45331 );
buf ( n335759 , n45332 );
buf ( n45334 , n45280 );
buf ( n45335 , n335711 );
and ( n45336 , n45334 , n45335 );
buf ( n45337 , n45336 );
buf ( n335764 , n45337 );
not ( n335765 , n335764 );
buf ( n335766 , n335224 );
not ( n45341 , n335766 );
or ( n45342 , n335765 , n45341 );
and ( n45343 , n335728 , n335711 );
nor ( n45344 , n45343 , n334858 );
buf ( n335771 , n45344 );
nand ( n335772 , n45342 , n335771 );
buf ( n335773 , n335772 );
buf ( n335774 , n335773 );
and ( n335775 , n335774 , n335759 );
not ( n45350 , n335774 );
and ( n335777 , n45350 , n335755 );
nor ( n335778 , n335775 , n335777 );
buf ( n335779 , n335778 );
not ( n45354 , n334738 );
nand ( n335781 , n45354 , n44431 );
buf ( n335782 , n335781 );
buf ( n335783 , n335781 );
not ( n335784 , n335783 );
buf ( n335785 , n335784 );
buf ( n335786 , n335785 );
buf ( n335787 , n45280 );
buf ( n335788 , n334757 );
and ( n335789 , n335787 , n335788 );
buf ( n335790 , n335789 );
buf ( n335791 , n335790 );
not ( n335792 , n335791 );
buf ( n335793 , n335224 );
not ( n45368 , n335793 );
or ( n45369 , n335792 , n45368 );
and ( n45370 , n335728 , n334757 );
not ( n45371 , n44428 );
nor ( n335798 , n45370 , n45371 );
buf ( n335799 , n335798 );
nand ( n335800 , n45369 , n335799 );
buf ( n335801 , n335800 );
buf ( n335802 , n335801 );
and ( n335803 , n335802 , n335786 );
not ( n335804 , n335802 );
and ( n335805 , n335804 , n335782 );
nor ( n335806 , n335803 , n335805 );
buf ( n335807 , n335806 );
not ( n45382 , n45371 );
nand ( n45383 , n45382 , n334757 );
buf ( n335810 , n45383 );
buf ( n335811 , n45383 );
not ( n335812 , n335811 );
buf ( n335813 , n335812 );
buf ( n335814 , n335813 );
buf ( n335815 , n45280 );
not ( n45390 , n335815 );
buf ( n335817 , n335224 );
not ( n335818 , n335817 );
or ( n45393 , n45390 , n335818 );
not ( n45394 , n335728 );
buf ( n335821 , n45394 );
nand ( n45396 , n45393 , n335821 );
buf ( n335823 , n45396 );
buf ( n335824 , n335823 );
and ( n45399 , n335824 , n335814 );
not ( n45400 , n335824 );
and ( n335827 , n45400 , n335810 );
nor ( n335828 , n45399 , n335827 );
buf ( n335829 , n335828 );
not ( n335830 , n44419 );
nand ( n45405 , n335830 , n334840 );
buf ( n335832 , n45405 );
buf ( n335833 , n45405 );
not ( n335834 , n335833 );
buf ( n335835 , n335834 );
buf ( n335836 , n335835 );
buf ( n45411 , n334647 );
not ( n45412 , n45411 );
nor ( n45413 , n45412 , n334692 );
buf ( n335840 , n45413 );
not ( n45415 , n335840 );
buf ( n335842 , n335224 );
not ( n335843 , n335842 );
or ( n45418 , n45415 , n335843 );
not ( n335845 , n45411 );
buf ( n335846 , n334830 );
not ( n335847 , n335846 );
or ( n335848 , n335845 , n335847 );
buf ( n335849 , n334839 );
not ( n335850 , n335849 );
buf ( n335851 , n335850 );
nand ( n335852 , n335848 , n335851 );
buf ( n45427 , n335852 );
not ( n45428 , n45427 );
buf ( n45429 , n45428 );
buf ( n335856 , n45429 );
nand ( n335857 , n45418 , n335856 );
buf ( n335858 , n335857 );
buf ( n335859 , n335858 );
and ( n45434 , n335859 , n335836 );
not ( n45435 , n335859 );
and ( n45436 , n45435 , n335832 );
nor ( n45437 , n45434 , n45436 );
buf ( n45438 , n45437 );
nand ( n335865 , n335851 , n45411 );
buf ( n335866 , n335865 );
buf ( n335867 , n335865 );
not ( n335868 , n335867 );
buf ( n335869 , n335868 );
buf ( n335870 , n335869 );
buf ( n335871 , n334692 );
not ( n335872 , n335871 );
buf ( n335873 , n335872 );
buf ( n335874 , n335873 );
not ( n335875 , n335874 );
buf ( n335876 , n335224 );
not ( n335877 , n335876 );
or ( n45452 , n335875 , n335877 );
not ( n335879 , n335846 );
buf ( n335880 , n335879 );
nand ( n335881 , n45452 , n335880 );
buf ( n335882 , n335881 );
buf ( n335883 , n335882 );
and ( n335884 , n335883 , n335870 );
not ( n335885 , n335883 );
and ( n45460 , n335885 , n335866 );
nor ( n335887 , n335884 , n45460 );
buf ( n335888 , n335887 );
nand ( n335889 , n334605 , n334528 );
buf ( n335890 , n335889 );
buf ( n335891 , n335889 );
not ( n335892 , n335891 );
buf ( n335893 , n335892 );
buf ( n45468 , n335893 );
nand ( n45469 , n44085 , n334491 );
buf ( n335896 , n45469 );
not ( n335897 , n335896 );
buf ( n335898 , n335897 );
buf ( n335899 , n335898 );
buf ( n335900 , n334820 );
nor ( n335901 , n335899 , n335900 );
buf ( n335902 , n335901 );
buf ( n335903 , n335902 );
buf ( n335904 , n44026 );
and ( n335905 , n335903 , n335904 );
buf ( n335906 , n335905 );
buf ( n335907 , n335906 );
not ( n335908 , n334286 );
buf ( n335909 , n335908 );
nand ( n335910 , n335907 , n335909 );
buf ( n335911 , n335910 );
buf ( n335912 , n335911 );
buf ( n45487 , n335906 );
buf ( n335914 , n335145 );
buf ( n335915 , n335914 );
nand ( n335916 , n45487 , n335915 );
buf ( n335917 , n335916 );
buf ( n45492 , n335917 );
buf ( n335919 , n334472 );
buf ( n335920 , n335902 );
and ( n335921 , n335919 , n335920 );
buf ( n335922 , n44167 );
buf ( n335923 , n335898 );
nor ( n335924 , n335922 , n335923 );
buf ( n335925 , n335924 );
buf ( n335926 , n335925 );
buf ( n335927 , n44177 );
not ( n335928 , n335927 );
buf ( n335929 , n335928 );
buf ( n335930 , n335929 );
nor ( n45505 , n335921 , n335926 , n335930 );
buf ( n45506 , n45505 );
buf ( n335933 , n45506 );
nand ( n335934 , n335912 , n45492 , n335933 );
buf ( n335935 , n335934 );
buf ( n335936 , n335935 );
and ( n335937 , n335936 , n45468 );
not ( n335938 , n335936 );
and ( n45513 , n335938 , n335890 );
nor ( n45514 , n335937 , n45513 );
buf ( n45515 , n45514 );
buf ( n45516 , n43972 );
buf ( n45517 , n334462 );
nand ( n45518 , n45516 , n45517 );
buf ( n45519 , n45518 );
buf ( n45520 , n45519 );
buf ( n335947 , n45519 );
not ( n45522 , n335947 );
buf ( n45523 , n45522 );
buf ( n335950 , n45523 );
nand ( n335951 , n43985 , n335914 );
buf ( n45526 , n43859 );
not ( n335953 , n43580 );
and ( n335954 , n45526 , n335953 , n43985 );
nor ( n335955 , n335954 , n44032 );
nand ( n45530 , n335951 , n335955 );
buf ( n335957 , n45530 );
and ( n335958 , n335957 , n335950 );
not ( n335959 , n335957 );
and ( n45534 , n335959 , n45520 );
nor ( n335961 , n335958 , n45534 );
buf ( n335962 , n335961 );
buf ( n335963 , n44038 );
buf ( n335964 , n334467 );
nand ( n335965 , n335963 , n335964 );
buf ( n335966 , n335965 );
buf ( n335967 , n335966 );
buf ( n335968 , n335966 );
not ( n335969 , n335968 );
buf ( n335970 , n335969 );
buf ( n45545 , n335970 );
buf ( n335972 , n334417 );
buf ( n45547 , n335972 );
buf ( n45548 , n45547 );
nand ( n335975 , n45548 , n335914 );
and ( n335976 , n45526 , n45548 , n335953 );
nor ( n45551 , n335976 , n334463 );
nand ( n335978 , n335975 , n45551 );
buf ( n335979 , n335978 );
and ( n335980 , n335979 , n45545 );
not ( n45555 , n335979 );
and ( n335982 , n45555 , n335967 );
nor ( n335983 , n335980 , n335982 );
buf ( n335984 , n335983 );
not ( n45559 , n44032 );
nand ( n335986 , n45559 , n43985 );
buf ( n45561 , n335986 );
buf ( n335988 , n335986 );
not ( n45563 , n335988 );
buf ( n45564 , n45563 );
buf ( n335991 , n45564 );
buf ( n335992 , n334367 );
and ( n45567 , n335992 , n335991 );
not ( n45568 , n335992 );
and ( n335995 , n45568 , n45561 );
nor ( n335996 , n45567 , n335995 );
buf ( n335997 , n335996 );
buf ( n335998 , n43923 );
not ( n335999 , n335998 );
buf ( n336000 , n334355 );
nor ( n336001 , n335999 , n336000 );
buf ( n336002 , n336001 );
buf ( n336003 , n336002 );
buf ( n336004 , n336002 );
not ( n336005 , n336004 );
buf ( n336006 , n336005 );
buf ( n336007 , n336006 );
buf ( n336008 , n333882 );
buf ( n45583 , n336008 );
buf ( n336010 , n45583 );
buf ( n336011 , n336010 );
buf ( n336012 , n333915 );
nor ( n336013 , n336011 , n336012 );
buf ( n336014 , n336013 );
and ( n336015 , n45526 , n336014 , n334005 );
buf ( n336016 , n336015 );
buf ( n336017 , n336014 );
buf ( n336018 , n334313 );
not ( n336019 , n336018 );
buf ( n336020 , n336019 );
buf ( n336021 , n336020 );
nand ( n336022 , n336017 , n336021 );
buf ( n336023 , n336022 );
buf ( n336024 , n336023 );
buf ( n336025 , n334337 );
buf ( n336026 , n333915 );
not ( n336027 , n336026 );
buf ( n336028 , n336027 );
buf ( n336029 , n336028 );
nand ( n336030 , n336025 , n336029 );
buf ( n336031 , n336030 );
buf ( n45606 , n336031 );
buf ( n336033 , n334344 );
nand ( n336034 , n336024 , n45606 , n336033 );
buf ( n336035 , n336034 );
buf ( n45610 , n336035 );
nor ( n45611 , n336016 , n45610 );
buf ( n45612 , n45611 );
buf ( n336039 , n45612 );
and ( n336040 , n336039 , n336007 );
not ( n45615 , n336039 );
and ( n336042 , n45615 , n336003 );
nor ( n336043 , n336040 , n336042 );
buf ( n336044 , n336043 );
buf ( n336045 , n333844 );
buf ( n336046 , n334334 );
nand ( n336047 , n336045 , n336046 );
buf ( n336048 , n336047 );
buf ( n336049 , n336048 );
buf ( n336050 , n336048 );
not ( n336051 , n336050 );
buf ( n336052 , n336051 );
buf ( n336053 , n336052 );
nand ( n336054 , n333960 , n43577 );
buf ( n45629 , n336054 );
buf ( n336056 , n333879 );
not ( n45631 , n336056 );
buf ( n45632 , n45631 );
buf ( n336059 , n45632 );
nor ( n336060 , n45629 , n336059 );
buf ( n336061 , n336060 );
buf ( n336062 , n336061 );
not ( n45637 , n336062 );
buf ( n336064 , n45526 );
not ( n45639 , n336064 );
or ( n45640 , n45637 , n45639 );
buf ( n336067 , n336020 );
buf ( n336068 , n333879 );
and ( n45643 , n336067 , n336068 );
buf ( n336070 , n334324 );
nor ( n336071 , n45643 , n336070 );
buf ( n336072 , n336071 );
buf ( n336073 , n336072 );
nand ( n336074 , n45640 , n336073 );
buf ( n336075 , n336074 );
buf ( n336076 , n336075 );
and ( n45651 , n336076 , n336053 );
not ( n336078 , n336076 );
and ( n336079 , n336078 , n336049 );
nor ( n336080 , n45651 , n336079 );
buf ( n336081 , n336080 );
buf ( n336082 , n334324 );
buf ( n336083 , n45632 );
nor ( n336084 , n336082 , n336083 );
buf ( n336085 , n336084 );
buf ( n336086 , n336085 );
not ( n336087 , n336086 );
buf ( n336088 , n336087 );
buf ( n336089 , n336088 );
buf ( n336090 , n336085 );
nand ( n336091 , n334005 , n45526 );
nand ( n336092 , n336091 , n334313 );
buf ( n336093 , n336092 );
and ( n336094 , n336093 , n336090 );
not ( n336095 , n336093 );
and ( n336096 , n336095 , n336089 );
nor ( n45671 , n336094 , n336096 );
buf ( n45672 , n45671 );
buf ( n45673 , n333985 );
buf ( n45674 , n334309 );
nand ( n45675 , n45673 , n45674 );
buf ( n45676 , n45675 );
buf ( n45677 , n45676 );
buf ( n336104 , n45676 );
not ( n45679 , n336104 );
buf ( n45680 , n45679 );
buf ( n336107 , n45680 );
and ( n336108 , n333960 , n334002 );
buf ( n336109 , n336108 );
not ( n336110 , n336109 );
buf ( n336111 , n45526 );
not ( n336112 , n336111 );
or ( n45687 , n336110 , n336112 );
buf ( n336114 , n334002 );
not ( n336115 , n336114 );
buf ( n336116 , n334302 );
not ( n45691 , n336116 );
buf ( n45692 , n45691 );
buf ( n336119 , n45692 );
not ( n45694 , n336119 );
or ( n45695 , n336115 , n45694 );
buf ( n336122 , n334305 );
not ( n336123 , n336122 );
buf ( n336124 , n336123 );
buf ( n336125 , n336124 );
nand ( n336126 , n45695 , n336125 );
buf ( n336127 , n336126 );
buf ( n336128 , n336127 );
not ( n45703 , n336128 );
buf ( n45704 , n45703 );
buf ( n336131 , n45704 );
nand ( n336132 , n45687 , n336131 );
buf ( n336133 , n336132 );
buf ( n336134 , n336133 );
and ( n336135 , n336134 , n336107 );
not ( n336136 , n336134 );
and ( n45711 , n336136 , n45677 );
nor ( n336138 , n336135 , n45711 );
buf ( n336139 , n336138 );
buf ( n336140 , n334002 );
buf ( n336141 , n336124 );
nand ( n336142 , n336140 , n336141 );
buf ( n336143 , n336142 );
buf ( n336144 , n336143 );
buf ( n336145 , n336143 );
not ( n336146 , n336145 );
buf ( n336147 , n336146 );
buf ( n45722 , n336147 );
not ( n45723 , n333960 );
not ( n336150 , n43859 );
or ( n45725 , n45723 , n336150 );
nand ( n45726 , n45725 , n334302 );
buf ( n336153 , n45726 );
and ( n45728 , n336153 , n45722 );
not ( n45729 , n336153 );
and ( n45730 , n45729 , n336144 );
nor ( n45731 , n45728 , n45730 );
buf ( n336158 , n45731 );
buf ( n336159 , n334299 );
not ( n45734 , n336159 );
buf ( n336161 , n43533 );
nand ( n45736 , n45734 , n336161 );
buf ( n336163 , n45736 );
buf ( n336164 , n336163 );
buf ( n336165 , n336163 );
not ( n45740 , n336165 );
buf ( n336167 , n45740 );
buf ( n336168 , n336167 );
not ( n45743 , n333937 );
not ( n45744 , n43859 );
or ( n45745 , n45743 , n45744 );
not ( n45746 , n334293 );
nand ( n45747 , n45745 , n45746 );
buf ( n336174 , n45747 );
and ( n45749 , n336174 , n336168 );
not ( n45750 , n336174 );
and ( n45751 , n45750 , n336164 );
nor ( n45752 , n45749 , n45751 );
buf ( n336179 , n45752 );
buf ( n336180 , n336028 );
buf ( n336181 , n334344 );
nand ( n45756 , n336180 , n336181 );
buf ( n336183 , n45756 );
buf ( n336184 , n336183 );
buf ( n336185 , n336183 );
not ( n45760 , n336185 );
buf ( n336187 , n45760 );
buf ( n336188 , n336187 );
buf ( n336189 , n336010 );
buf ( n336190 , n336054 );
nor ( n45765 , n336189 , n336190 );
buf ( n336192 , n45765 );
buf ( n336193 , n336192 );
not ( n45768 , n336193 );
buf ( n336195 , n45526 );
not ( n45770 , n336195 );
or ( n45771 , n45768 , n45770 );
buf ( n336198 , n336020 );
buf ( n336199 , n336010 );
not ( n45774 , n336199 );
buf ( n336201 , n45774 );
buf ( n336202 , n336201 );
and ( n45777 , n336198 , n336202 );
buf ( n336204 , n334337 );
nor ( n45779 , n45777 , n336204 );
buf ( n336206 , n45779 );
buf ( n336207 , n336206 );
nand ( n45782 , n45771 , n336207 );
buf ( n336209 , n45782 );
buf ( n336210 , n336209 );
and ( n45785 , n336210 , n336188 );
not ( n45786 , n336210 );
and ( n45787 , n45786 , n336184 );
nor ( n45788 , n45785 , n45787 );
buf ( n336215 , n45788 );
nand ( n45790 , n334451 , n334417 );
buf ( n336217 , n45790 );
buf ( n336218 , n334816 );
nor ( n45793 , n336217 , n336218 );
buf ( n336220 , n45793 );
buf ( n336221 , n336220 );
buf ( n336222 , n335908 );
nand ( n45797 , n336221 , n336222 );
buf ( n336224 , n45797 );
buf ( n336225 , n336224 );
buf ( n336226 , n336220 );
buf ( n336227 , n335145 );
nand ( n45802 , n336226 , n336227 );
buf ( n336229 , n45802 );
buf ( n336230 , n336229 );
buf ( n336231 , n334819 );
buf ( n336232 , n334472 );
nand ( n45807 , n336231 , n336232 );
buf ( n336234 , n45807 );
buf ( n336235 , n336234 );
buf ( n336236 , n44122 );
and ( n45811 , n336225 , n336230 , n336235 , n336236 );
buf ( n336238 , n45811 );
buf ( n336239 , n335908 );
buf ( n45814 , n334820 );
buf ( n336241 , n45814 );
buf ( n336242 , n45790 );
nor ( n45817 , n336241 , n336242 );
buf ( n336244 , n45817 );
buf ( n336245 , n336244 );
nand ( n45820 , n336239 , n336245 );
buf ( n336247 , n45820 );
buf ( n336248 , n334065 );
not ( n45823 , n336248 );
buf ( n336250 , n45823 );
buf ( n336251 , n336250 );
buf ( n336252 , n334096 );
nand ( n45827 , n336251 , n336252 );
buf ( n336254 , n45827 );
buf ( n336255 , n336254 );
buf ( n336256 , n336254 );
not ( n45831 , n336256 );
buf ( n336258 , n45831 );
buf ( n336259 , n336258 );
buf ( n336260 , n334117 );
not ( n45835 , n336260 );
buf ( n336262 , n334266 );
not ( n45837 , n336262 );
buf ( n336264 , n45837 );
buf ( n336265 , n336264 );
not ( n45840 , n336265 );
or ( n45841 , n45835 , n45840 );
buf ( n336268 , n43661 );
not ( n45843 , n336268 );
buf ( n336270 , n45843 );
buf ( n336271 , n336270 );
nand ( n45846 , n45841 , n336271 );
buf ( n336273 , n45846 );
buf ( n336274 , n336273 );
and ( n45849 , n336274 , n336259 );
not ( n45850 , n336274 );
and ( n45851 , n45850 , n336255 );
nor ( n45852 , n45849 , n45851 );
buf ( n336279 , n45852 );
buf ( n336280 , n43657 );
buf ( n336281 , n334086 );
nand ( n45856 , n336280 , n336281 );
buf ( n336283 , n45856 );
buf ( n336284 , n336283 );
buf ( n336285 , n336283 );
not ( n45860 , n336285 );
buf ( n336287 , n45860 );
buf ( n336288 , n336287 );
buf ( n336289 , n334114 );
not ( n45864 , n336289 );
buf ( n336291 , n336264 );
not ( n45866 , n336291 );
or ( n45867 , n45864 , n45866 );
buf ( n336294 , n334076 );
nand ( n45869 , n45867 , n336294 );
buf ( n336296 , n45869 );
buf ( n336297 , n336296 );
and ( n45872 , n336297 , n336288 );
not ( n45873 , n336297 );
and ( n45874 , n45873 , n336284 );
nor ( n45875 , n45872 , n45874 );
buf ( n336302 , n45875 );
buf ( n336303 , n334114 );
buf ( n336304 , n334076 );
nand ( n45879 , n336303 , n336304 );
buf ( n336306 , n45879 );
buf ( n336307 , n336306 );
buf ( n336308 , n336306 );
not ( n45883 , n336308 );
buf ( n336310 , n45883 );
buf ( n336311 , n336310 );
buf ( n336312 , n336264 );
and ( n45887 , n336312 , n336311 );
not ( n45888 , n336312 );
and ( n45889 , n45888 , n336307 );
nor ( n45890 , n45887 , n45889 );
buf ( n336317 , n45890 );
buf ( n336318 , n334121 );
not ( n45893 , n336318 );
buf ( n336320 , n45893 );
buf ( n336321 , n336320 );
buf ( n336322 , n334276 );
not ( n45897 , n336322 );
buf ( n336324 , n45897 );
buf ( n336325 , n336324 );
buf ( n336326 , n336264 );
nand ( n45901 , n336321 , n336325 , n336326 );
buf ( n336328 , n45901 );
buf ( n336329 , n336320 );
buf ( n336330 , n43854 );
buf ( n336331 , n336264 );
nand ( n45906 , n336329 , n336330 , n336331 );
buf ( n336333 , n45906 );
not ( n45908 , n334162 );
buf ( n336335 , n45908 );
buf ( n336336 , n334155 );
nand ( n45911 , n336335 , n336336 );
buf ( n336338 , n45911 );
buf ( n336339 , n336338 );
buf ( n336340 , n45908 );
buf ( n336341 , n334177 );
buf ( n336342 , n334239 );
nand ( n45917 , n336340 , n336341 , n336342 );
buf ( n336344 , n45917 );
buf ( n336345 , n336344 );
buf ( n336346 , n334251 );
and ( n45921 , n336339 , n336345 , n336346 );
buf ( n336348 , n45921 );
buf ( n336349 , n336348 );
buf ( n336350 , n334160 );
buf ( n336351 , n334260 );
nor ( n45926 , n336350 , n336351 );
buf ( n336353 , n45926 );
buf ( n336354 , n336353 );
buf ( n336355 , n336353 );
buf ( n336356 , n336348 );
not ( n45931 , n336349 );
not ( n45932 , n336354 );
or ( n45933 , n45931 , n45932 );
or ( n45934 , n336355 , n336356 );
nand ( n45935 , n45933 , n45934 );
buf ( n336362 , n45935 );
buf ( n336363 , n45908 );
buf ( n336364 , n334251 );
nand ( n45939 , n336363 , n336364 );
buf ( n336366 , n45939 );
buf ( n336367 , n336366 );
buf ( n336368 , n334242 );
buf ( n336369 , n334155 );
or ( n45944 , n336368 , n336369 );
buf ( n336371 , n45944 );
buf ( n336372 , n336371 );
buf ( n336373 , n336371 );
buf ( n336374 , n336366 );
not ( n45949 , n336367 );
not ( n45950 , n336372 );
or ( n45951 , n45949 , n45950 );
or ( n45952 , n336373 , n336374 );
nand ( n45953 , n45951 , n45952 );
buf ( n336380 , n45953 );
buf ( n336381 , n334174 );
not ( n45956 , n336381 );
buf ( n336383 , n45956 );
buf ( n336384 , n336383 );
buf ( n336385 , n43715 );
nand ( n45960 , n336384 , n336385 );
buf ( n336387 , n45960 );
buf ( n336388 , n336387 );
buf ( n336389 , n334239 );
buf ( n336390 , n334239 );
buf ( n336391 , n336387 );
not ( n45966 , n336388 );
not ( n45967 , n336389 );
or ( n45968 , n45966 , n45967 );
or ( n45969 , n336390 , n336391 );
nand ( n45970 , n45968 , n45969 );
buf ( n336397 , n45970 );
buf ( n336398 , n45002 );
buf ( n336399 , n335519 );
buf ( n336400 , n45085 );
nand ( n45975 , n336399 , n336400 );
buf ( n336402 , n45975 );
buf ( n336403 , n336402 );
not ( n45978 , n336403 );
buf ( n336405 , n45978 );
buf ( n336406 , n336405 );
buf ( n336407 , n45085 );
not ( n45982 , n336407 );
buf ( n336409 , n334896 );
not ( n45984 , n336409 );
or ( n45985 , n45982 , n45984 );
buf ( n336412 , n44485 );
not ( n45987 , n336412 );
buf ( n336414 , n45987 );
buf ( n336415 , n336414 );
nand ( n45990 , n45985 , n336415 );
buf ( n336417 , n45990 );
buf ( n336418 , n336417 );
and ( n45993 , n336398 , n336406 );
nor ( n45994 , n45993 , n336418 );
buf ( n336421 , n45994 );
buf ( n336422 , n334220 );
buf ( n336423 , n334230 );
nand ( n45998 , n336422 , n336423 );
buf ( n336425 , n45998 );
buf ( n336426 , n336425 );
buf ( n336427 , n43786 );
buf ( n336428 , n43786 );
buf ( n336429 , n336425 );
not ( n46004 , n336426 );
not ( n46005 , n336427 );
or ( n46006 , n46004 , n46005 );
or ( n46007 , n336428 , n336429 );
nand ( n46008 , n46006 , n46007 );
buf ( n336435 , n46008 );
xor ( n46010 , n43779 , n43780 );
xor ( n46011 , n46010 , n43782 );
buf ( n336438 , n46011 );
buf ( n336439 , n334109 );
buf ( n336440 , n336324 );
nand ( n46015 , n336439 , n336440 );
buf ( n336442 , n46015 );
buf ( n336443 , n334109 );
buf ( n336444 , n43854 );
nand ( n46019 , n336443 , n336444 );
buf ( n336446 , n46019 );
buf ( n336447 , n335122 );
not ( n46022 , n33997 );
nand ( n46023 , n46022 , n335036 );
not ( n46024 , n46023 );
not ( n46025 , n34002 );
or ( n46026 , n46024 , n46025 );
not ( n46027 , n335036 );
nand ( n46028 , n46027 , n33997 );
nand ( n46029 , n46026 , n46028 );
not ( n46030 , n46029 );
and ( n46031 , n309831 , n309928 );
not ( n46032 , n309829 );
not ( n46033 , n309923 );
or ( n46034 , n46032 , n46033 );
nand ( n46035 , n46034 , n19275 );
nor ( n46036 , n46031 , n46035 );
not ( n46037 , n309830 );
nand ( n46038 , n46037 , n18214 );
nand ( n46039 , n46036 , n46038 );
not ( n46040 , n19344 );
nand ( n46041 , n46040 , n309766 );
not ( n46042 , n46041 );
and ( n46043 , n46039 , n46042 );
not ( n46044 , n46039 );
and ( n46045 , n46044 , n46041 );
nor ( n46046 , n46043 , n46045 );
buf ( n46047 , n328586 );
xor ( n46048 , n46047 , n33989 );
xor ( n46049 , n46046 , n46048 );
not ( n46050 , n46049 );
nand ( n46051 , n46030 , n46050 );
buf ( n46052 , n46047 );
or ( n46053 , n46052 , n33989 );
not ( n46054 , n46053 );
not ( n46055 , n46046 );
or ( n46056 , n46054 , n46055 );
nand ( n46057 , n46052 , n33989 );
nand ( n46058 , n46056 , n46057 );
buf ( n336485 , n46058 );
not ( n46060 , n336485 );
buf ( n336487 , n46060 );
xnor ( n46062 , n34015 , n34010 );
not ( n46063 , n46062 );
not ( n46064 , n310321 );
xnor ( n46065 , n310014 , n310008 );
not ( n46066 , n46065 );
and ( n46067 , n46064 , n46066 );
and ( n46068 , n310321 , n46065 );
nor ( n46069 , n46067 , n46068 );
not ( n46070 , n46069 );
nand ( n46071 , n309812 , n309928 );
and ( n46072 , n309921 , n19382 );
nor ( n46073 , n46072 , n309774 );
nand ( n46074 , n309936 , n46071 , n46073 );
not ( n46075 , n46074 );
or ( n46076 , n46070 , n46075 );
xor ( n46077 , n310321 , n326872 );
and ( n46078 , n46073 , n46077 );
nand ( n46079 , n46071 , n46078 , n309936 );
nand ( n46080 , n46076 , n46079 );
not ( n46081 , n46080 );
or ( n46082 , n46063 , n46081 );
or ( n46083 , n46062 , n46080 );
nand ( n46084 , n46082 , n46083 );
not ( n46085 , n46084 );
and ( n46086 , n336487 , n46085 );
or ( n46087 , n34015 , n34010 );
not ( n46088 , n46087 );
not ( n46089 , n46080 );
or ( n46090 , n46088 , n46089 );
nand ( n46091 , n34015 , n34010 );
nand ( n46092 , n46090 , n46091 );
buf ( n336519 , n46092 );
not ( n46094 , n336519 );
buf ( n336521 , n46094 );
buf ( n336522 , n333308 );
not ( n46097 , n336522 );
buf ( n336524 , n46097 );
and ( n46099 , n336521 , n336524 );
nor ( n46100 , n46086 , n46099 );
nand ( n46101 , n335044 , n46051 , n46100 );
not ( n46102 , n46101 );
buf ( n336529 , n46102 );
buf ( n336530 , n333304 );
buf ( n336531 , n333314 );
nor ( n46106 , n336530 , n336531 );
buf ( n336533 , n46106 );
not ( n46108 , n336533 );
or ( n46109 , n333310 , n333302 );
and ( n46110 , n46108 , n46109 );
buf ( n336537 , n46110 );
buf ( n336538 , n333316 );
buf ( n336539 , n333320 );
or ( n46114 , n336538 , n336539 );
buf ( n336541 , n46114 );
buf ( n336542 , n336541 );
and ( n46117 , n336537 , n336542 );
buf ( n336544 , n46117 );
buf ( n336545 , n336544 );
nand ( n46120 , n336529 , n336545 );
buf ( n336547 , n46120 );
buf ( n336548 , n336547 );
nor ( n46123 , n336447 , n336548 );
buf ( n336550 , n46123 );
buf ( n336551 , n335122 );
buf ( n336552 , n46102 );
buf ( n336553 , n46110 );
nand ( n46128 , n336552 , n336553 );
buf ( n336555 , n46128 );
buf ( n336556 , n336555 );
nor ( n46131 , n336551 , n336556 );
buf ( n336558 , n46131 );
buf ( n336559 , n335122 );
nand ( n46134 , n46102 , n46109 );
buf ( n336561 , n46134 );
nor ( n46136 , n336559 , n336561 );
buf ( n336563 , n46136 );
nand ( n46138 , n46085 , n336487 );
buf ( n336565 , n46138 );
not ( n46140 , n336565 );
not ( n46141 , n44612 );
buf ( n336568 , n46029 );
not ( n46143 , n336568 );
buf ( n336570 , n46050 );
nand ( n46145 , n46143 , n336570 );
buf ( n336572 , n46145 );
not ( n46147 , n336572 );
or ( n46148 , n46141 , n46147 );
buf ( n336575 , n46029 );
buf ( n336576 , n46049 );
nand ( n46151 , n336575 , n336576 );
buf ( n336578 , n46151 );
nand ( n46153 , n46148 , n336578 );
buf ( n336580 , n46153 );
not ( n46155 , n336580 );
or ( n46156 , n46140 , n46155 );
buf ( n336583 , n46084 );
buf ( n336584 , n336487 );
not ( n46159 , n336584 );
and ( n46160 , n336583 , n46159 );
buf ( n336587 , n46160 );
buf ( n336588 , n336587 );
not ( n46163 , n336588 );
buf ( n336590 , n46163 );
buf ( n336591 , n336590 );
nand ( n46166 , n46156 , n336591 );
buf ( n336593 , n46166 );
buf ( n336594 , n336593 );
not ( n46169 , n336594 );
buf ( n336596 , n46169 );
buf ( n336597 , n336541 );
nand ( n46172 , n333310 , n333302 );
or ( n46173 , n336533 , n46172 );
buf ( n336600 , n333304 );
buf ( n336601 , n333314 );
nand ( n46176 , n336600 , n336601 );
buf ( n336603 , n46176 );
nand ( n46178 , n46173 , n336603 );
buf ( n336605 , n46178 );
buf ( n336606 , n333316 );
buf ( n336607 , n333320 );
nand ( n46182 , n336606 , n336607 );
buf ( n336609 , n46182 );
buf ( n336610 , n336609 );
not ( n46185 , n336597 );
not ( n46186 , n336605 );
or ( n46187 , n46185 , n46186 );
nand ( n46188 , n46187 , n336610 );
buf ( n336615 , n46188 );
buf ( n336616 , n336555 );
not ( n46191 , n336616 );
buf ( n336618 , n46191 );
buf ( n336619 , n336547 );
not ( n46194 , n336619 );
buf ( n336621 , n46194 );
buf ( n336622 , n46134 );
not ( n46197 , n336622 );
buf ( n336624 , n46197 );
buf ( n336625 , n43661 );
buf ( n336626 , n336250 );
nand ( n46201 , n336625 , n336626 );
buf ( n336628 , n46201 );
buf ( n336629 , n334417 );
buf ( n336630 , n44038 );
and ( n46205 , n336629 , n336630 );
buf ( n336632 , n46205 );
buf ( n336633 , n46153 );
not ( n46208 , n336633 );
buf ( n336635 , n46208 );
buf ( n336636 , n336324 );
buf ( n336637 , n334019 );
not ( n46212 , n336637 );
buf ( n336639 , n46212 );
buf ( n336640 , n336639 );
nand ( n46215 , n336636 , n336640 );
buf ( n336642 , n46215 );
buf ( n336643 , n333937 );
buf ( n336644 , n45746 );
and ( n46219 , n336643 , n336644 );
buf ( n336646 , n46219 );
buf ( n336647 , n334038 );
buf ( n336648 , n334050 );
nand ( n46223 , n336647 , n336648 );
buf ( n336650 , n46223 );
buf ( n336651 , n40137 );
buf ( n336652 , n18256 );
buf ( n336653 , n334204 );
not ( n46228 , n336651 );
not ( n46229 , n336652 );
or ( n46230 , n46228 , n46229 );
nand ( n46231 , n46230 , n336653 );
buf ( n336658 , n46231 );
buf ( n336659 , n44164 );
buf ( n336660 , n334583 );
nand ( n46235 , n336659 , n336660 );
buf ( n336662 , n46235 );
buf ( n336663 , n336521 );
buf ( n336664 , n336524 );
nor ( n46239 , n336663 , n336664 );
buf ( n336666 , n46239 );
buf ( n336667 , n43604 );
not ( n46242 , n336667 );
buf ( n336669 , n46242 );
buf ( n336670 , n334109 );
buf ( n336671 , n334269 );
or ( n46246 , n336670 , n336671 );
buf ( n336673 , n46246 );
buf ( n336674 , n336673 );
buf ( n336675 , n336642 );
xnor ( n46250 , n336674 , n336675 );
buf ( n336677 , n46250 );
and ( n46252 , n43600 , n336669 );
nor ( n46253 , n46252 , n334042 );
or ( n46254 , n334109 , n334269 );
buf ( n336681 , n43854 );
not ( n46256 , n336681 );
buf ( n336683 , n43604 );
nor ( n46258 , n46256 , n336683 );
buf ( n336685 , n46258 );
nand ( n46260 , n46254 , n336685 );
nand ( n46261 , n46253 , n46260 );
buf ( n336688 , n46261 );
buf ( n336689 , n336650 );
xnor ( n46264 , n336688 , n336689 );
buf ( n336691 , n46264 );
buf ( n336692 , n336238 );
buf ( n336693 , n336662 );
xor ( n46268 , n336692 , n336693 );
buf ( n336695 , n46268 );
buf ( n336696 , n325721 );
buf ( n46272 , n36664 );
buf ( n336698 , n46272 );
nand ( n46274 , n336696 , n336698 );
buf ( n336700 , n46274 );
buf ( n336701 , n34449 );
buf ( n336702 , n36120 );
buf ( n336703 , n36259 );
not ( n46279 , n336701 );
nand ( n46280 , n46279 , n336702 , n336703 );
buf ( n336706 , n46280 );
buf ( n336707 , n36120 );
buf ( n336708 , n328264 );
buf ( n336709 , n36145 );
nand ( n46285 , n336707 , n336708 , n336709 );
buf ( n336711 , n46285 );
buf ( n336712 , n36120 );
buf ( n336713 , n328279 );
buf ( n336714 , n36259 );
nand ( n46290 , n336712 , n336713 , n336714 );
buf ( n336716 , n46290 );
buf ( n336717 , n328493 );
buf ( n336718 , n36120 );
buf ( n336719 , n328493 );
buf ( n336720 , n36120 );
not ( n46296 , n336717 );
not ( n46297 , n336718 );
or ( n46298 , n46296 , n46297 );
or ( n46299 , n336719 , n336720 );
nand ( n46300 , n46298 , n46299 );
buf ( n336726 , n46300 );
buf ( n336727 , n328329 );
buf ( n336728 , n36120 );
buf ( n336729 , n36145 );
nand ( n46305 , n336727 , n336728 , n336729 );
buf ( n336731 , n46305 );
buf ( n336732 , n36120 );
buf ( n336733 , n328288 );
buf ( n336734 , n36145 );
nand ( n46310 , n336732 , n336733 , n336734 );
buf ( n336736 , n46310 );
buf ( n336737 , n327709 );
buf ( n336738 , n36078 );
buf ( n336739 , n326515 );
not ( n46315 , n336737 );
not ( n46316 , n336738 );
or ( n46317 , n46315 , n46316 );
nand ( n46318 , n46317 , n336739 );
buf ( n336744 , n46318 );
buf ( n336745 , n36120 );
buf ( n336746 , n36259 );
buf ( n336747 , n36260 );
nand ( n46323 , n336745 , n336746 , n336747 );
buf ( n336749 , n46323 );
buf ( n336750 , n335224 );
buf ( n336751 , n335158 );
not ( n46327 , n46102 );
nor ( n46328 , n335122 , n46327 );
buf ( n336754 , n46328 );
buf ( n336755 , n46102 );
not ( n46331 , n336755 );
buf ( n336757 , n335183 );
not ( n46333 , n336757 );
or ( n46334 , n46331 , n46333 );
nand ( n46335 , n336521 , n336524 );
and ( n46336 , n46138 , n46335 );
not ( n46337 , n46336 );
not ( n46338 , n46153 );
or ( n46339 , n46337 , n46338 );
not ( n46340 , n46335 );
not ( n46341 , n336587 );
or ( n46342 , n46340 , n46341 );
not ( n46343 , n336666 );
nand ( n46344 , n46342 , n46343 );
not ( n46345 , n46344 );
nand ( n46346 , n46339 , n46345 );
not ( n46347 , n46346 );
buf ( n336773 , n46347 );
nand ( n46349 , n46334 , n336773 );
buf ( n336775 , n46349 );
buf ( n336776 , n336775 );
and ( n46352 , n336750 , n336751 , n336754 );
nor ( n46353 , n46352 , n336776 );
buf ( n336779 , n46353 );
buf ( n336780 , n335224 );
buf ( n336781 , n335158 );
buf ( n336782 , n336550 );
buf ( n336783 , n336621 );
not ( n46359 , n336783 );
not ( n46360 , n44694 );
not ( n46361 , n44527 );
or ( n46362 , n46360 , n46361 );
nand ( n46363 , n46362 , n44756 );
buf ( n336789 , n46363 );
not ( n46365 , n336789 );
or ( n46366 , n46359 , n46365 );
not ( n46367 , n46336 );
not ( n46368 , n46153 );
or ( n46369 , n46367 , n46368 );
nand ( n46370 , n46369 , n46345 );
and ( n46371 , n46370 , n336544 );
nor ( n46372 , n46371 , n336615 );
buf ( n336798 , n46372 );
nand ( n46374 , n46366 , n336798 );
buf ( n336800 , n46374 );
buf ( n336801 , n336800 );
and ( n46377 , n336780 , n336781 , n336782 );
nor ( n46378 , n46377 , n336801 );
buf ( n336804 , n46378 );
buf ( n336805 , n335152 );
buf ( n336806 , n335158 );
buf ( n336807 , n336558 );
buf ( n336808 , n336618 );
not ( n46384 , n336808 );
buf ( n336810 , n46363 );
not ( n46386 , n336810 );
or ( n46387 , n46384 , n46386 );
and ( n46388 , n46346 , n46110 );
nor ( n46389 , n46388 , n46178 );
buf ( n336815 , n46389 );
nand ( n46391 , n46387 , n336815 );
buf ( n336817 , n46391 );
buf ( n336818 , n336817 );
and ( n46394 , n336805 , n336806 , n336807 );
nor ( n46395 , n46394 , n336818 );
buf ( n336821 , n46395 );
buf ( n336822 , n335152 );
buf ( n336823 , n335158 );
nand ( n46399 , n335042 , n44617 );
nand ( n46400 , n46138 , n46051 , n46399 );
nor ( n46401 , n335122 , n46400 );
buf ( n336827 , n46401 );
not ( n46403 , n46400 );
not ( n46404 , n46403 );
not ( n46405 , n46363 );
or ( n46406 , n46404 , n46405 );
nand ( n46407 , n46406 , n336596 );
buf ( n336833 , n46407 );
and ( n46409 , n336822 , n336823 , n336827 );
nor ( n46410 , n46409 , n336833 );
buf ( n336836 , n46410 );
buf ( n336837 , n335152 );
buf ( n336838 , n335158 );
not ( n46414 , n335045 );
nor ( n46415 , n46414 , n335122 );
buf ( n336841 , n46415 );
not ( n46417 , n335045 );
not ( n46418 , n335183 );
or ( n46419 , n46417 , n46418 );
nand ( n46420 , n46419 , n335041 );
buf ( n336846 , n46420 );
and ( n46422 , n336837 , n336838 , n336841 );
nor ( n46423 , n46422 , n336846 );
buf ( n336849 , n46423 );
buf ( n336850 , n335152 );
buf ( n336851 , n335158 );
buf ( n336852 , n336563 );
not ( n46428 , n336624 );
not ( n46429 , n46363 );
or ( n46430 , n46428 , n46429 );
and ( n46431 , n46370 , n46109 );
not ( n46432 , n46172 );
nor ( n46433 , n46431 , n46432 );
nand ( n46434 , n46430 , n46433 );
buf ( n336860 , n46434 );
and ( n46436 , n336850 , n336851 , n336852 );
nor ( n46437 , n46436 , n336860 );
buf ( n336863 , n46437 );
buf ( n336864 , n335224 );
buf ( n336865 , n335158 );
nand ( n46441 , n335044 , n46051 );
nor ( n46442 , n335122 , n46441 );
buf ( n336868 , n46442 );
not ( n46444 , n46441 );
buf ( n336870 , n46444 );
not ( n46446 , n336870 );
buf ( n336872 , n335183 );
not ( n46448 , n336872 );
or ( n46449 , n46446 , n46448 );
buf ( n336875 , n336635 );
nand ( n46451 , n46449 , n336875 );
buf ( n336877 , n46451 );
buf ( n336878 , n336877 );
and ( n46454 , n336864 , n336865 , n336868 );
nor ( n46455 , n46454 , n336878 );
buf ( n336881 , n46455 );
buf ( n336882 , n37475 );
buf ( n336883 , n326456 );
nand ( n46459 , n336882 , n336883 );
buf ( n336885 , n46459 );
nand ( n46461 , n327748 , n36118 , n336885 );
not ( n46462 , n36098 );
and ( n46463 , n326532 , n326487 );
nor ( n46464 , n46463 , n36117 );
nand ( n46465 , n46462 , n46464 );
buf ( n336891 , n37225 );
buf ( n336892 , n325653 );
nor ( n46468 , n336891 , n336892 );
buf ( n336894 , n46468 );
nand ( n46470 , n46461 , n46465 , n336894 );
not ( n46471 , n36170 );
nand ( n46472 , n336706 , n328341 , n46471 );
nand ( n46473 , n328374 , n328354 );
not ( n46474 , n46473 );
and ( n46475 , n46472 , n46474 );
not ( n46476 , n46472 );
and ( n46477 , n46476 , n46473 );
nor ( n46478 , n46475 , n46477 );
buf ( n336904 , n328328 );
not ( n46480 , n336904 );
buf ( n336906 , n36530 );
not ( n46482 , n336906 );
or ( n46483 , n46480 , n46482 );
buf ( n336909 , n328459 );
nand ( n46485 , n46483 , n336909 );
buf ( n336911 , n46485 );
not ( n46487 , n336911 );
nand ( n46488 , n46487 , n328333 , n336731 );
not ( n46489 , n324378 );
not ( n46490 , n324374 );
or ( n46491 , n46489 , n46490 );
or ( n46492 , n324374 , n324378 );
nand ( n46493 , n46491 , n46492 );
not ( n46494 , n46493 );
and ( n46495 , n46488 , n46494 );
not ( n46496 , n46488 );
and ( n46497 , n46496 , n46493 );
nor ( n46498 , n46495 , n46497 );
buf ( n336924 , n328295 );
not ( n46500 , n336924 );
buf ( n336926 , n36530 );
not ( n46502 , n336926 );
or ( n46503 , n46500 , n46502 );
buf ( n336929 , n38039 );
nand ( n46505 , n46503 , n336929 );
buf ( n336931 , n46505 );
not ( n46507 , n336931 );
nand ( n46508 , n36120 , n37870 , n36145 );
nand ( n46509 , n46507 , n328299 , n46508 );
nand ( n46510 , n326929 , n327006 );
not ( n46511 , n46510 );
and ( n46512 , n46509 , n46511 );
not ( n46513 , n46509 );
and ( n46514 , n46513 , n46510 );
nor ( n46515 , n46512 , n46514 );
buf ( n336941 , n328261 );
not ( n46517 , n336941 );
buf ( n336943 , n36530 );
not ( n46519 , n336943 );
or ( n46520 , n46517 , n46519 );
buf ( n336946 , n328499 );
nand ( n46522 , n46520 , n336946 );
buf ( n336948 , n46522 );
not ( n46524 , n336948 );
nand ( n46525 , n46524 , n328267 , n336711 );
nand ( n46526 , n328274 , n328408 );
not ( n46527 , n46526 );
and ( n46528 , n46525 , n46527 );
not ( n46529 , n46525 );
and ( n46530 , n46529 , n46526 );
nor ( n46531 , n46528 , n46530 );
buf ( n336957 , n37859 );
not ( n46533 , n336957 );
buf ( n336959 , n36530 );
not ( n46535 , n336959 );
or ( n46536 , n46533 , n46535 );
buf ( n336962 , n328496 );
nand ( n46538 , n46536 , n336962 );
buf ( n336964 , n46538 );
not ( n46540 , n336964 );
nand ( n46541 , n46540 , n328291 , n336736 );
nand ( n46542 , n326975 , n36542 );
not ( n46543 , n46542 );
and ( n46544 , n46541 , n46543 );
not ( n46545 , n46541 );
and ( n46546 , n46545 , n46542 );
nor ( n46547 , n46544 , n46546 );
nand ( n46548 , n36120 , n36145 , n46272 );
not ( n46549 , n36530 );
nand ( n46550 , n336700 , n46548 , n46549 );
nand ( n46551 , n37859 , n328496 );
not ( n46552 , n46551 );
and ( n46553 , n46550 , n46552 );
not ( n46554 , n46550 );
and ( n46555 , n46554 , n46551 );
nor ( n46556 , n46553 , n46555 );
not ( n46557 , n335134 );
not ( n46558 , n46328 );
or ( n46559 , n46557 , n46558 );
nand ( n46560 , n46559 , n336779 );
nand ( n46561 , n46109 , n46172 );
not ( n46562 , n46561 );
and ( n46563 , n46560 , n46562 );
not ( n46564 , n46560 );
and ( n46565 , n46564 , n46561 );
nor ( n46566 , n46563 , n46565 );
not ( n46567 , n335134 );
not ( n46568 , n46415 );
or ( n46569 , n46567 , n46568 );
nand ( n46570 , n46569 , n336849 );
nand ( n46571 , n336572 , n336578 );
not ( n46572 , n46571 );
and ( n46573 , n46570 , n46572 );
not ( n46574 , n46570 );
and ( n46575 , n46574 , n46571 );
nor ( n46576 , n46573 , n46575 );
not ( n46577 , n46442 );
not ( n46578 , n335134 );
or ( n46579 , n46577 , n46578 );
nand ( n46580 , n46579 , n336881 );
nand ( n46581 , n336590 , n46138 );
not ( n46582 , n46581 );
and ( n46583 , n46580 , n46582 );
not ( n46584 , n46580 );
and ( n46585 , n46584 , n46581 );
nor ( n46586 , n46583 , n46585 );
not ( n46587 , n46401 );
not ( n46588 , n335134 );
or ( n46589 , n46587 , n46588 );
nand ( n46590 , n46589 , n336836 );
not ( n46591 , n336666 );
nand ( n46592 , n46591 , n46335 );
not ( n46593 , n46592 );
and ( n46594 , n46590 , n46593 );
not ( n46595 , n46590 );
and ( n46596 , n46595 , n46592 );
nor ( n46597 , n46594 , n46596 );
not ( n46598 , n336550 );
not ( n46599 , n335134 );
or ( n46600 , n46598 , n46599 );
nand ( n46601 , n46600 , n336804 );
xor ( n46602 , n333326 , n333322 );
and ( n46603 , n46601 , n46602 );
not ( n46604 , n46601 );
not ( n46605 , n46602 );
and ( n46606 , n46604 , n46605 );
nor ( n46607 , n46603 , n46606 );
not ( n46608 , n336558 );
not ( n46609 , n335134 );
or ( n46610 , n46608 , n46609 );
nand ( n46611 , n46610 , n336821 );
nand ( n46612 , n336541 , n336609 );
not ( n46613 , n46612 );
and ( n46614 , n46611 , n46613 );
not ( n46615 , n46611 );
and ( n46616 , n46615 , n46612 );
nor ( n46617 , n46614 , n46616 );
not ( n46618 , n336563 );
not ( n46619 , n335134 );
or ( n46620 , n46618 , n46619 );
nand ( n46621 , n46620 , n336863 );
not ( n46622 , n336533 );
nand ( n46623 , n46622 , n336603 );
not ( n46624 , n46623 );
and ( n46625 , n46621 , n46624 );
not ( n46626 , n46621 );
and ( n46627 , n46626 , n46623 );
nor ( n46628 , n46625 , n46627 );
not ( n46629 , n36297 );
nand ( n46630 , n328350 , n336749 , n46629 );
nand ( n46631 , n36301 , n36261 );
not ( n46632 , n46631 );
and ( n46633 , n46630 , n46632 );
not ( n46634 , n46630 );
and ( n46635 , n46634 , n46631 );
nor ( n46636 , n46633 , n46635 );
not ( n46637 , n327319 );
not ( n46638 , n46470 );
or ( n46639 , n46637 , n46638 );
nor ( n46640 , n34714 , n325275 );
buf ( n337066 , n46640 );
buf ( n337067 , n327216 );
and ( n46643 , n337066 , n337067 );
buf ( n337069 , n46643 );
nand ( n46645 , n46639 , n337069 );
nand ( n46646 , n46645 , n328419 , n327220 );
nand ( n46647 , n36158 , n36151 );
not ( n46648 , n46647 );
and ( n46649 , n46646 , n46648 );
not ( n46650 , n46646 );
and ( n46651 , n46650 , n46647 );
nor ( n46652 , n46649 , n46651 );
not ( n46653 , n328386 );
not ( n46654 , n327319 );
not ( n46655 , n46470 );
or ( n46656 , n46654 , n46655 );
buf ( n337082 , n46640 );
not ( n46658 , n337082 );
buf ( n337084 , n328355 );
nor ( n46660 , n46658 , n337084 );
buf ( n337086 , n46660 );
nand ( n46662 , n46656 , n337086 );
not ( n46663 , n46662 );
or ( n46664 , n46653 , n46663 );
and ( n46665 , n326626 , n324765 );
not ( n46666 , n46665 );
nand ( n46667 , n46664 , n46666 );
nand ( n46668 , n46662 , n328386 , n46665 );
nand ( n46669 , n46667 , n46668 );
buf ( n337095 , n43144 );
buf ( n337096 , n333534 );
nor ( n46672 , n337095 , n337096 );
buf ( n337098 , n46672 );
buf ( n337099 , n44988 );
buf ( n337100 , n336402 );
nor ( n46676 , n337099 , n337100 );
buf ( n337102 , n46676 );
buf ( n337103 , n35567 );
buf ( n337104 , n38063 );
xnor ( n46680 , n337103 , n337104 );
buf ( n337106 , n46680 );
nand ( n46682 , n46470 , n327319 );
nand ( n46683 , n36271 , n35254 );
not ( n46684 , n46683 );
and ( n46685 , n46682 , n46684 );
not ( n46686 , n46682 );
and ( n46687 , n46686 , n46683 );
nor ( n46688 , n46685 , n46687 );
not ( n46689 , n327692 );
not ( n46690 , n326454 );
nor ( n46691 , n46690 , n37282 );
not ( n46692 , n44038 );
not ( n46693 , n334463 );
or ( n46694 , n46692 , n46693 );
nand ( n46695 , n46694 , n334467 );
and ( n46696 , n46689 , n46691 , n37264 );
nor ( n46697 , n46696 , n336744 );
nand ( n46698 , n328282 , n336716 , n37989 );
not ( n46699 , n326995 );
nand ( n46700 , n46699 , n326920 );
not ( n46701 , n46700 );
and ( n46702 , n46698 , n46701 );
not ( n46703 , n46698 );
and ( n46704 , n46703 , n46700 );
nor ( n46705 , n46702 , n46704 );
buf ( n337131 , n335914 );
buf ( n337132 , n336244 );
nand ( n46708 , n337131 , n337132 );
buf ( n337134 , n46708 );
buf ( n337135 , n45814 );
not ( n46711 , n337135 );
buf ( n337137 , n334472 );
nand ( n46713 , n46711 , n337137 );
buf ( n337139 , n46713 );
nand ( n46715 , n336247 , n337134 , n337139 , n44167 );
nand ( n46716 , n44177 , n45469 );
not ( n46717 , n46716 );
and ( n46718 , n46715 , n46717 );
not ( n46719 , n46715 );
and ( n46720 , n46719 , n46716 );
nor ( n46721 , n46718 , n46720 );
not ( n46722 , n46691 );
not ( n46723 , n37258 );
or ( n46724 , n46722 , n46723 );
nand ( n46725 , n46724 , n46697 );
nor ( n46726 , n326521 , n326510 );
and ( n46727 , n46725 , n46726 );
not ( n46728 , n46725 );
not ( n46729 , n46726 );
and ( n46730 , n46728 , n46729 );
nor ( n46731 , n46727 , n46730 );
buf ( n337157 , n37258 );
buf ( n337158 , n326456 );
nand ( n46734 , n337157 , n337158 );
buf ( n337160 , n46734 );
buf ( n337161 , n326456 );
buf ( n337162 , n37264 );
buf ( n337163 , n46689 );
nand ( n46739 , n337161 , n337162 , n337163 );
buf ( n337165 , n46739 );
nand ( n46741 , n337160 , n327748 , n337165 );
not ( n46742 , n326528 );
nand ( n46743 , n46742 , n35930 );
not ( n46744 , n46743 );
and ( n46745 , n46741 , n46744 );
not ( n46746 , n46741 );
and ( n46747 , n46746 , n46743 );
nor ( n46748 , n46745 , n46747 );
nand ( n46749 , n335908 , n44026 );
buf ( n337175 , n44026 );
buf ( n337176 , n335914 );
nand ( n46752 , n337175 , n337176 );
buf ( n337178 , n46752 );
nand ( n46754 , n46749 , n337178 , n334475 );
nand ( n46755 , n334819 , n44122 );
not ( n46756 , n46755 );
and ( n46757 , n46754 , n46756 );
not ( n46758 , n46754 );
and ( n46759 , n46758 , n46755 );
nor ( n46760 , n46757 , n46759 );
nand ( n46761 , n336632 , n335914 );
and ( n46762 , n336632 , n45526 , n335953 );
nor ( n46763 , n46762 , n46695 );
nand ( n46764 , n46761 , n46763 );
nor ( n46765 , n44044 , n334456 );
and ( n46766 , n46764 , n46765 );
not ( n46767 , n46764 );
not ( n46768 , n46765 );
and ( n46769 , n46767 , n46768 );
nor ( n46770 , n46766 , n46769 );
nand ( n46771 , n326061 , n326033 );
not ( n46772 , n46771 );
buf ( n337198 , n35567 );
buf ( n337199 , n325870 );
buf ( n337200 , n326046 );
nand ( n46776 , n337198 , n337199 , n337200 );
buf ( n337202 , n46776 );
nand ( n46778 , n337202 , n328469 , n328162 );
not ( n46779 , n46778 );
or ( n46780 , n46772 , n46779 );
or ( n46781 , n46771 , n46778 );
nand ( n46782 , n46780 , n46781 );
nand ( n46783 , n42299 , n330232 );
not ( n46784 , n334042 );
nand ( n46785 , n46784 , n336669 );
not ( n46786 , n46785 );
not ( n46787 , n43600 );
nand ( n46788 , n46787 , n336446 , n336333 );
not ( n46789 , n46788 );
or ( n46790 , n46786 , n46789 );
or ( n46791 , n46785 , n46788 );
nand ( n46792 , n46790 , n46791 );
nand ( n46793 , n39759 , n330209 );
not ( n46794 , n46793 );
nand ( n46795 , n333056 , n332815 , n42649 );
not ( n46796 , n46795 );
or ( n46797 , n46794 , n46796 );
or ( n46798 , n46793 , n46795 );
nand ( n46799 , n46797 , n46798 );
not ( n46800 , n39793 );
nand ( n46801 , n46800 , n330234 );
not ( n46802 , n46801 );
nand ( n46803 , n42310 , n333060 , n333069 );
not ( n46804 , n46803 );
or ( n46805 , n46802 , n46804 );
or ( n46806 , n46801 , n46803 );
nand ( n46807 , n46805 , n46806 );
nand ( n46808 , n334014 , n334025 );
not ( n46809 , n46808 );
nand ( n46810 , n336442 , n336328 , n336639 );
not ( n46811 , n46810 );
or ( n46812 , n46809 , n46811 );
or ( n46813 , n46808 , n46810 );
nand ( n46814 , n46812 , n46813 );
not ( n46815 , n334199 );
nand ( n46816 , n46815 , n334236 );
not ( n46817 , n46816 );
nand ( n46818 , n334230 , n43797 );
not ( n46819 , n46818 );
or ( n46820 , n46817 , n46819 );
or ( n46821 , n46818 , n46816 );
nand ( n46822 , n46820 , n46821 );
not ( n46823 , n334239 );
not ( n46824 , n336383 );
or ( n46825 , n46823 , n46824 );
nand ( n46826 , n46825 , n43715 );
not ( n46827 , n46826 );
not ( n46828 , n334146 );
nand ( n46829 , n46828 , n334152 );
not ( n46830 , n46829 );
or ( n46831 , n46827 , n46830 );
or ( n46832 , n46829 , n46826 );
nand ( n46833 , n46831 , n46832 );
not ( n46834 , n40057 );
nand ( n46835 , n46834 , n40092 );
not ( n46836 , n46835 );
not ( n46837 , n333091 );
or ( n46838 , n330599 , n330505 );
nand ( n46839 , n46838 , n42541 );
nand ( n46840 , n46837 , n46839 );
not ( n46841 , n46840 );
or ( n46842 , n46836 , n46841 );
or ( n46843 , n46835 , n46840 );
nand ( n46844 , n46842 , n46843 );
not ( n46845 , n35528 );
nand ( n46846 , n325959 , n325898 );
not ( n46847 , n46846 );
or ( n46848 , n46845 , n46847 );
or ( n46849 , n46846 , n35528 );
nand ( n46850 , n46848 , n46849 );
not ( n46851 , n335224 );
nor ( n46852 , n44988 , n333601 );
not ( n46853 , n46852 );
or ( n46854 , n46851 , n46853 );
and ( n46855 , n335683 , n45002 );
not ( n46856 , n44456 );
nor ( n46857 , n46855 , n46856 );
nand ( n46858 , n46854 , n46857 );
not ( n46859 , n334887 );
nor ( n46860 , n46859 , n337098 );
and ( n46861 , n46858 , n46860 );
not ( n46862 , n46858 );
not ( n46863 , n46860 );
and ( n46864 , n46862 , n46863 );
nor ( n46865 , n46861 , n46864 );
not ( n46866 , n337102 );
not ( n46867 , n335224 );
or ( n46868 , n46866 , n46867 );
nand ( n46869 , n46868 , n336421 );
nand ( n46870 , n335550 , n43059 );
not ( n46871 , n46870 );
and ( n46872 , n46869 , n46871 );
not ( n46873 , n46869 );
and ( n46874 , n46873 , n46870 );
nor ( n46875 , n46872 , n46874 );
not ( n46876 , n35046 );
nor ( n46877 , n46876 , n327123 );
not ( n46878 , n46877 );
not ( n46879 , n36120 );
or ( n46880 , n46878 , n46879 );
nand ( n46881 , n46880 , n328440 );
nand ( n46882 , n327143 , n34991 );
not ( n46883 , n46882 );
and ( n46884 , n46881 , n46883 );
not ( n46885 , n46881 );
and ( n46886 , n46885 , n46882 );
nor ( n46887 , n46884 , n46886 );
and ( n46888 , n37655 , n328485 );
nor ( n46889 , n46888 , n35700 );
nand ( n46890 , n328485 , n37660 );
nand ( n46891 , n46889 , n46890 );
nand ( n46892 , n328064 , n326089 );
not ( n46893 , n46892 );
and ( n46894 , n46891 , n46893 );
not ( n46895 , n46891 );
and ( n46896 , n46895 , n46892 );
nor ( n46897 , n46894 , n46896 );
or ( n46898 , n334103 , n334060 );
not ( n46899 , n46898 );
nand ( n46900 , n336250 , n334117 , n336264 );
nand ( n46901 , n46900 , n336628 , n334096 );
not ( n46902 , n46901 );
or ( n46903 , n46899 , n46902 );
or ( n46904 , n46898 , n46901 );
nand ( n46905 , n46903 , n46904 );
nand ( n46906 , n44247 , n45246 );
not ( n46907 , n46906 );
and ( n46908 , n335224 , n46907 );
not ( n46909 , n335224 );
and ( n46910 , n46909 , n46906 );
nor ( n46911 , n46908 , n46910 );
buf ( n337337 , n328475 );
buf ( n337338 , n328478 );
nand ( n46914 , n37297 , n35432 );
nand ( n46915 , n46914 , n35862 );
buf ( n337341 , n46915 );
and ( n46917 , n337341 , n337338 );
not ( n46918 , n337341 );
and ( n46919 , n46918 , n337337 );
nor ( n46920 , n46917 , n46919 );
buf ( n337346 , n46920 );
nand ( n46922 , n325772 , n326265 );
xor ( n46923 , n336646 , n45526 );
buf ( n337349 , n333083 );
buf ( n337350 , n330430 );
buf ( n337351 , n330377 );
and ( n46927 , n337350 , n337351 );
buf ( n337353 , n46927 );
buf ( n337354 , n337353 );
buf ( n337355 , n330609 );
nand ( n46931 , n337354 , n337355 );
buf ( n337357 , n46931 );
buf ( n337358 , n337357 );
buf ( n337359 , n337353 );
buf ( n337360 , n330652 );
nand ( n46936 , n337359 , n337360 );
buf ( n337362 , n46936 );
buf ( n337363 , n337362 );
buf ( n337364 , n330377 );
buf ( n337365 , n330402 );
nand ( n46941 , n337364 , n337365 );
buf ( n337367 , n46941 );
buf ( n337368 , n337367 );
buf ( n337369 , n330408 );
nand ( n46945 , n337358 , n337363 , n337368 , n337369 );
buf ( n337371 , n46945 );
buf ( n337372 , n337371 );
buf ( n337373 , n333083 );
buf ( n337374 , n337371 );
not ( n46950 , n337349 );
not ( n46951 , n337372 );
or ( n46952 , n46950 , n46951 );
or ( n46953 , n337373 , n337374 );
nand ( n46954 , n46952 , n46953 );
buf ( n337380 , n46954 );
and ( n46956 , n46922 , n327692 );
not ( n46957 , n46922 );
and ( n46958 , n46957 , n37297 );
nor ( n46959 , n46956 , n46958 );
not ( n46960 , n46783 );
buf ( n337386 , n330312 );
buf ( n337387 , n330322 );
nand ( n46963 , n337386 , n337387 );
buf ( n337389 , n46963 );
not ( n46965 , n330212 );
buf ( n337391 , n332645 );
buf ( n337392 , n333117 );
nand ( n46968 , n337391 , n337392 );
buf ( n337394 , n46968 );
nand ( n46970 , n337389 , n46965 , n337394 );
not ( n46971 , n46970 );
or ( n46972 , n46960 , n46971 );
or ( n46973 , n46783 , n46970 );
nand ( n46974 , n46972 , n46973 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
