// IWLS benchmark module "i6" printed on Wed May 29 17:26:47 2002
module i6(\V138(0) , \V138(2) , \V32(27) , \V32(26) , \V32(25) , \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V96(27) , \V138(4) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V131(27) , \V131(26) , \V131(25) , \V131(24) , \V131(23) , \V131(22) , \V131(21) , \V131(20) , \V131(19) , \V131(18) , \V131(17) , \V131(16) , \V131(15) , \V131(14) , \V131(13) , \V131(12) , \V131(11) , \V131(10) , \V131(9) , \V131(8) , \V131(7) , \V131(6) , \V131(5) , \V131(4) , \V131(3) , \V131(2) , \V131(1) , \V131(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V99(0) , \V138(3) , \V98(0) , \V97(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V134(0) , \V133(1) , \V133(0) , \V131(31) , \V131(30) , \V131(29) , \V131(28) , \V166(27) , \V166(26) , \V166(25) , \V166(24) , \V166(23) , \V166(22) , \V166(21) , \V166(20) , \V166(19) , \V166(18) , \V166(17) , \V166(16) , \V166(15) , \V166(14) , \V166(13) , \V166(12) , \V166(11) , \V166(10) , \V166(9) , \V166(8) , \V166(7) , \V166(6) , \V166(5) , \V166(4) , \V166(3) , \V166(2) , \V166(1) , \V166(0) , \V198(31) , \V198(30) , \V198(29) , \V198(28) , \V198(27) , \V198(26) , \V198(25) , \V198(24) , \V198(23) , \V198(22) , \V198(21) , \V198(20) , \V198(19) , \V198(18) , \V198(17) , \V198(16) , \V198(15) , \V198(14) , \V198(13) , \V198(12) , \V198(11) , \V198(10) , \V198(9) , \V198(8) , \V198(7) , \V198(6) , \V198(5) , \V198(4) , \V198(3) , \V198(2) , \V198(1) , \V198(0) , \V205(6) , \V205(5) , \V205(4) , \V205(3) , \V205(2) , \V205(1) , \V205(0) );
input
  \V138(0) ,
  \V96(0) ,
  \V96(1) ,
  \V64(13) ,
  \V96(2) ,
  \V64(12) ,
  \V96(3) ,
  \V64(15) ,
  \V96(4) ,
  \V64(14) ,
  \V96(5) ,
  \V96(6) ,
  \V96(7) ,
  \V64(11) ,
  \V96(8) ,
  \V64(10) ,
  \V96(9) ,
  \V97(0) ,
  \V64(17) ,
  \V64(16) ,
  \V64(19) ,
  \V64(18) ,
  \V64(23) ,
  \V64(22) ,
  \V64(25) ,
  \V64(24) ,
  \V98(0) ,
  \V64(21) ,
  \V64(20) ,
  \V64(27) ,
  \V64(26) ,
  \V64(29) ,
  \V64(28) ,
  \V99(0) ,
  \V64(31) ,
  \V64(30) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(13) ,
  \V32(4) ,
  \V32(12) ,
  \V32(5) ,
  \V32(15) ,
  \V32(6) ,
  \V32(14) ,
  \V32(7) ,
  \V32(8) ,
  \V32(9) ,
  \V32(11) ,
  \V32(10) ,
  \V32(17) ,
  \V32(16) ,
  \V32(19) ,
  \V32(18) ,
  \V32(23) ,
  \V32(22) ,
  \V32(25) ,
  \V32(24) ,
  \V32(21) ,
  \V32(20) ,
  \V131(27) ,
  \V131(26) ,
  \V32(27) ,
  \V131(29) ,
  \V96(13) ,
  \V32(26) ,
  \V131(28) ,
  \V96(12) ,
  \V32(29) ,
  \V96(15) ,
  \V32(28) ,
  \V96(14) ,
  \V96(11) ,
  \V96(10) ,
  \V131(21) ,
  \V131(20) ,
  \V32(31) ,
  \V131(23) ,
  \V131(3) ,
  \V32(30) ,
  \V131(22) ,
  \V131(2) ,
  \V131(25) ,
  \V131(5) ,
  \V96(17) ,
  \V131(24) ,
  \V131(4) ,
  \V96(16) ,
  \V131(17) ,
  \V96(19) ,
  \V131(16) ,
  \V96(18) ,
  \V131(19) ,
  \V131(1) ,
  \V96(23) ,
  \V131(18) ,
  \V131(0) ,
  \V96(22) ,
  \V96(25) ,
  \V96(24) ,
  \V131(7) ,
  \V96(21) ,
  \V131(6) ,
  \V96(20) ,
  \V131(11) ,
  \V131(9) ,
  \V131(10) ,
  \V131(8) ,
  \V131(13) ,
  \V131(12) ,
  \V131(15) ,
  \V96(27) ,
  \V131(14) ,
  \V96(26) ,
  \V96(29) ,
  \V96(28) ,
  \V64(0) ,
  \V96(31) ,
  \V133(1) ,
  \V64(1) ,
  \V96(30) ,
  \V133(0) ,
  \V64(2) ,
  \V64(3) ,
  \V64(4) ,
  \V64(5) ,
  \V64(6) ,
  \V64(7) ,
  \V64(8) ,
  \V64(9) ,
  \V134(0) ,
  \V131(31) ,
  \V131(30) ,
  \V138(3) ,
  \V138(2) ,
  \V138(4) ;
output
  \V198(11) ,
  \V198(10) ,
  \V198(13) ,
  \V198(12) ,
  \V198(15) ,
  \V198(14) ,
  \V166(3) ,
  \V166(2) ,
  \V166(5) ,
  \V166(4) ,
  \V166(1) ,
  \V166(0) ,
  \V166(7) ,
  \V166(6) ,
  \V166(9) ,
  \V166(8) ,
  \V198(31) ,
  \V198(30) ,
  \V205(3) ,
  \V205(2) ,
  \V205(5) ,
  \V205(4) ,
  \V166(27) ,
  \V166(26) ,
  \V198(3) ,
  \V198(2) ,
  \V205(1) ,
  \V198(5) ,
  \V205(0) ,
  \V198(4) ,
  \V198(1) ,
  \V198(0) ,
  \V205(6) ,
  \V166(21) ,
  \V166(20) ,
  \V166(23) ,
  \V166(22) ,
  \V198(7) ,
  \V166(25) ,
  \V198(6) ,
  \V166(24) ,
  \V198(9) ,
  \V166(17) ,
  \V198(8) ,
  \V166(16) ,
  \V166(19) ,
  \V166(18) ,
  \V166(11) ,
  \V166(10) ,
  \V166(13) ,
  \V166(12) ,
  \V166(15) ,
  \V166(14) ,
  \V198(27) ,
  \V198(26) ,
  \V198(29) ,
  \V198(28) ,
  \V198(21) ,
  \V198(20) ,
  \V198(23) ,
  \V198(22) ,
  \V198(25) ,
  \V198(24) ,
  \V198(17) ,
  \V198(16) ,
  \V198(19) ,
  \V198(18) ;
wire
  \V291(21) ,
  \V291(20) ,
  \V291(23) ,
  \V291(22) ,
  \V291(25) ,
  \V291(24) ,
  \V291(17) ,
  \V291(16) ,
  \V291(19) ,
  \V291(18) ,
  \V389(3) ,
  \V389(2) ,
  \V291(11) ,
  \V291(10) ,
  \V291(13) ,
  \V291(12) ,
  \V389(1) ,
  \V291(15) ,
  \V389(0) ,
  \V291(14) ,
  \V417(27) ,
  \V417(26) ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \V417(21) ,
  \[4] ,
  \V417(20) ,
  \[5] ,
  \V417(23) ,
  \[6] ,
  \V417(22) ,
  \[7] ,
  \V417(25) ,
  \[8] ,
  \V417(24) ,
  \[9] ,
  \V417(17) ,
  \V417(16) ,
  \V417(19) ,
  \V417(18) ,
  \V417(11) ,
  \V417(10) ,
  \V417(13) ,
  \V417(12) ,
  \V417(15) ,
  \V417(14) ,
  V206,
  V207,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V214,
  V215,
  V216,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V223,
  V224,
  V225,
  V226,
  V227,
  V228,
  V229,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V242,
  V243,
  V244,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V257,
  V258,
  V259,
  V260,
  V261,
  V262,
  V263,
  V292,
  V293,
  V294,
  V295,
  V296,
  V297,
  V298,
  V299,
  V300,
  V301,
  V302,
  V303,
  V304,
  V305,
  V306,
  V307,
  V308,
  V309,
  V310,
  V311,
  V312,
  V313,
  V314,
  V315,
  V316,
  V317,
  V318,
  V319,
  V320,
  V321,
  V322,
  V323,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  V330,
  V331,
  V332,
  V333,
  V334,
  V335,
  V336,
  V337,
  V338,
  V339,
  V340,
  V341,
  V342,
  V343,
  V344,
  V345,
  V346,
  V347,
  V348,
  V349,
  V350,
  V351,
  V352,
  V353,
  V354,
  V355,
  V356,
  V357,
  V358,
  V359,
  V360,
  V361,
  V362,
  V363,
  V364,
  V365,
  V366,
  V367,
  V368,
  V369,
  V370,
  V371,
  V372,
  V373,
  V374,
  V375,
  V376,
  V377,
  V378,
  V379,
  V380,
  V381,
  V382,
  V383,
  V384,
  V385,
  V418,
  V419,
  V420,
  V421,
  V422,
  V423,
  V424,
  V425,
  V426,
  V427,
  V428,
  V429,
  V430,
  V431,
  V432,
  V433,
  V434,
  V435,
  V436,
  V437,
  V438,
  V439,
  V440,
  V441,
  V442,
  V443,
  V444,
  V445,
  V446,
  V447,
  V448,
  V449,
  V450,
  V451,
  V452,
  V453,
  V454,
  V455,
  V456,
  V457,
  V458,
  V459,
  V460,
  V461,
  V462,
  V463,
  V464,
  V465,
  V466,
  V467,
  V474,
  V475,
  V476,
  V477,
  V478,
  V479,
  \V417(3) ,
  V480,
  V481,
  V482,
  \V417(2) ,
  \V417(5) ,
  \V417(4) ,
  \[10] ,
  \[11] ,
  \[12] ,
  \V417(1) ,
  \[13] ,
  \V417(0) ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \V417(7) ,
  \[19] ,
  \V417(6) ,
  \V417(9) ,
  \V417(8) ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \V471(3) ,
  \[29] ,
  \V471(2) ,
  \V471(1) ,
  \V471(0) ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \V291(3) ,
  \[39] ,
  \V291(2) ,
  \V291(5) ,
  \V291(4) ,
  \V291(1) ,
  \V291(0) ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \V291(7) ,
  \V473(1) ,
  \[45] ,
  \V291(6) ,
  \V473(0) ,
  \[46] ,
  \V291(9) ,
  \[47] ,
  \V291(8) ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \V291(27) ,
  \V291(26) ;
assign
  \V291(21)  = ~\V64(21) ,
  \V198(11)  = \[48] ,
  \V291(20)  = ~\V64(20) ,
  \V198(10)  = \[49] ,
  \V291(23)  = ~\V64(23) ,
  \V198(13)  = \[46] ,
  \V291(22)  = ~\V64(22) ,
  \V198(12)  = \[47] ,
  \V291(25)  = ~\V64(25) ,
  \V198(15)  = \[44] ,
  \V291(24)  = ~\V64(24) ,
  \V198(14)  = \[45] ,
  \V291(17)  = ~\V64(17) ,
  \V291(16)  = ~\V64(16) ,
  \V291(19)  = ~\V64(19) ,
  \V291(18)  = ~\V64(18) ,
  \V389(3)  = ~\V64(31) ,
  \V166(3)  = \[24] ,
  \V389(2)  = ~\V64(30) ,
  \V166(2)  = \[25] ,
  \V291(11)  = ~\V64(11) ,
  \V166(5)  = \[22] ,
  \V291(10)  = ~\V64(10) ,
  \V166(4)  = \[23] ,
  \V291(13)  = ~\V64(13) ,
  \V291(12)  = ~\V64(12) ,
  \V389(1)  = ~\V64(29) ,
  \V291(15)  = ~\V64(15) ,
  \V166(1)  = \[26] ,
  \V389(0)  = ~\V64(28) ,
  \V291(14)  = ~\V64(14) ,
  \V166(0)  = \[27] ,
  \V166(7)  = \[20] ,
  \V166(6)  = \[21] ,
  \V166(9)  = \[18] ,
  \V417(27)  = ~\V131(27) ,
  \V166(8)  = \[19] ,
  \V417(26)  = ~\V131(26) ,
  \V198(31)  = \[28] ,
  \V198(30)  = \[29] ,
  \[0]  = V292 | (V236 | V208),
  \[1]  = V293 | (V237 | V209),
  \[2]  = V294 | (V238 | V210),
  \[3]  = V295 | (V239 | V211),
  \V417(21)  = ~\V131(21) ,
  \[4]  = V296 | (V240 | V212),
  \V417(20)  = ~\V131(20) ,
  \[5]  = V297 | (V241 | V213),
  \V417(23)  = ~\V131(23) ,
  \[6]  = V298 | (V242 | V214),
  \V417(22)  = ~\V131(22) ,
  \[7]  = V299 | (V243 | V215),
  \V417(25)  = ~\V131(25) ,
  \[8]  = V300 | (V244 | V216),
  \V417(24)  = ~\V131(24) ,
  \[9]  = V301 | (V245 | V217),
  \V417(17)  = ~\V131(17) ,
  \V417(16)  = ~\V131(16) ,
  \V417(19)  = ~\V131(19) ,
  \V417(18)  = ~\V131(18) ,
  \V417(11)  = ~\V131(11) ,
  \V417(10)  = ~\V131(10) ,
  \V417(13)  = ~\V131(13) ,
  \V417(12)  = ~\V131(12) ,
  \V417(15)  = ~\V131(15) ,
  \V417(14)  = ~\V131(14) ,
  \V205(3)  = \[63] ,
  \V205(2)  = \[64] ,
  \V205(5)  = \[61] ,
  \V205(4)  = \[62] ,
  \V166(27)  = \[0] ,
  \V166(26)  = \[1] ,
  \V198(3)  = \[56] ,
  \V198(2)  = \[57] ,
  \V205(1)  = \[65] ,
  \V198(5)  = \[54] ,
  \V205(0)  = \[66] ,
  \V198(4)  = \[55] ,
  \V198(1)  = \[58] ,
  \V198(0)  = \[59] ,
  \V205(6)  = \[60] ,
  \V166(21)  = \[6] ,
  V206 = ~\V138(0) ,
  V207 = ~\V138(2) ,
  \V166(20)  = \[7] ,
  V208 = V206 & (V207 & \V32(27) ),
  V209 = V206 & (V207 & \V32(26) ),
  V210 = V206 & (V207 & \V32(25) ),
  V211 = V206 & (V207 & \V32(24) ),
  V212 = V206 & (V207 & \V32(23) ),
  V213 = V206 & (V207 & \V32(22) ),
  V214 = V206 & (V207 & \V32(21) ),
  V215 = V206 & (V207 & \V32(20) ),
  V216 = V206 & (V207 & \V32(19) ),
  V217 = V206 & (V207 & \V32(18) ),
  \V166(23)  = \[4] ,
  V218 = V206 & (V207 & \V32(17) ),
  V219 = V206 & (V207 & \V32(16) ),
  V220 = V206 & (V207 & \V32(15) ),
  V221 = V206 & (V207 & \V32(14) ),
  V222 = V206 & (V207 & \V32(13) ),
  V223 = V206 & (V207 & \V32(12) ),
  V224 = V206 & (V207 & \V32(11) ),
  V225 = V206 & (V207 & \V32(10) ),
  V226 = V206 & (V207 & \V32(9) ),
  V227 = V206 & (V207 & \V32(8) ),
  \V166(22)  = \[5] ,
  \V198(7)  = \[52] ,
  V228 = V206 & (V207 & \V32(7) ),
  V229 = V206 & (V207 & \V32(6) ),
  V230 = V206 & (V207 & \V32(5) ),
  V231 = V206 & (V207 & \V32(4) ),
  V232 = V206 & (V207 & \V32(3) ),
  V233 = V206 & (V207 & \V32(2) ),
  V234 = V206 & (V207 & \V32(1) ),
  V235 = V206 & (V207 & \V32(0) ),
  V236 = \V138(0)  & (V207 & \V64(27) ),
  V237 = \V138(0)  & (V207 & \V64(26) ),
  \V166(25)  = \[2] ,
  \V198(6)  = \[53] ,
  V238 = \V138(0)  & (V207 & \V64(25) ),
  V239 = \V138(0)  & (V207 & \V64(24) ),
  V240 = \V138(0)  & (V207 & \V64(23) ),
  V241 = \V138(0)  & (V207 & \V64(22) ),
  V242 = \V138(0)  & (V207 & \V64(21) ),
  V243 = \V138(0)  & (V207 & \V64(20) ),
  V244 = \V138(0)  & (V207 & \V64(19) ),
  V245 = \V138(0)  & (V207 & \V64(18) ),
  V246 = \V138(0)  & (V207 & \V64(17) ),
  V247 = \V138(0)  & (V207 & \V64(16) ),
  \V166(24)  = \[3] ,
  \V198(9)  = \[50] ,
  V248 = \V138(0)  & (V207 & \V64(15) ),
  V249 = \V138(0)  & (V207 & \V64(14) ),
  V250 = \V138(0)  & (V207 & \V64(13) ),
  V251 = \V138(0)  & (V207 & \V64(12) ),
  V252 = \V138(0)  & (V207 & \V64(11) ),
  V253 = \V138(0)  & (V207 & \V64(10) ),
  V254 = \V138(0)  & (V207 & \V64(9) ),
  V255 = \V138(0)  & (V207 & \V64(8) ),
  V256 = \V138(0)  & (V207 & \V64(7) ),
  V257 = \V138(0)  & (V207 & \V64(6) ),
  \V166(17)  = \[10] ,
  \V198(8)  = \[51] ,
  V258 = \V138(0)  & (V207 & \V64(5) ),
  V259 = \V138(0)  & (V207 & \V64(4) ),
  V260 = \V138(0)  & (V207 & \V64(3) ),
  V261 = \V138(0)  & (V207 & \V64(2) ),
  V262 = \V138(0)  & (V207 & \V64(1) ),
  V263 = \V138(0)  & (V207 & \V64(0) ),
  \V166(16)  = \[11] ,
  \V166(19)  = \[8] ,
  \V166(18)  = \[9] ,
  V292 = \V138(0)  & (\V138(2)  & \V291(27) ),
  V293 = \V138(0)  & (\V138(2)  & \V291(26) ),
  V294 = \V138(0)  & (\V138(2)  & \V291(25) ),
  V295 = \V138(0)  & (\V138(2)  & \V291(24) ),
  V296 = \V138(0)  & (\V138(2)  & \V291(23) ),
  V297 = \V138(0)  & (\V138(2)  & \V291(22) ),
  V298 = \V138(0)  & (\V138(2)  & \V291(21) ),
  V299 = \V138(0)  & (\V138(2)  & \V291(20) ),
  \V166(11)  = \[16] ,
  V300 = \V138(0)  & (\V138(2)  & \V291(19) ),
  V301 = \V138(0)  & (\V138(2)  & \V291(18) ),
  V302 = \V138(0)  & (\V138(2)  & \V291(17) ),
  V303 = \V138(0)  & (\V138(2)  & \V291(16) ),
  V304 = \V138(0)  & (\V138(2)  & \V291(15) ),
  V305 = \V138(0)  & (\V138(2)  & \V291(14) ),
  V306 = \V138(0)  & (\V138(2)  & \V291(13) ),
  V307 = \V138(0)  & (\V138(2)  & \V291(12) ),
  \V166(10)  = \[17] ,
  V308 = \V138(0)  & (\V138(2)  & \V291(11) ),
  V309 = \V138(0)  & (\V138(2)  & \V291(10) ),
  V310 = \V138(0)  & (\V138(2)  & \V291(9) ),
  V311 = \V138(0)  & (\V138(2)  & \V291(8) ),
  V312 = \V138(0)  & (\V138(2)  & \V291(7) ),
  V313 = \V138(0)  & (\V138(2)  & \V291(6) ),
  V314 = \V138(0)  & (\V138(2)  & \V291(5) ),
  V315 = \V138(0)  & (\V138(2)  & \V291(4) ),
  V316 = \V138(0)  & (\V138(2)  & \V291(3) ),
  V317 = \V138(0)  & (\V138(2)  & \V291(2) ),
  \V166(13)  = \[14] ,
  V318 = \V138(0)  & (\V138(2)  & \V291(1) ),
  V319 = \V138(0)  & (\V138(2)  & \V291(0) ),
  V320 = ~\V138(0) ,
  V321 = ~\V138(2) ,
  V322 = \V138(4)  & (V321 & (V320 & \V96(27) )),
  V323 = \V138(4)  & (V321 & (V320 & \V96(26) )),
  V324 = \V138(4)  & (V321 & (V320 & \V96(25) )),
  V325 = \V138(4)  & (V321 & (V320 & \V96(24) )),
  V326 = \V138(4)  & (V321 & (V320 & \V96(23) )),
  V327 = \V138(4)  & (V321 & (V320 & \V96(22) )),
  \V166(12)  = \[15] ,
  V328 = \V138(4)  & (V321 & (V320 & \V96(21) )),
  V329 = \V138(4)  & (V321 & (V320 & \V96(20) )),
  V330 = \V138(4)  & (V321 & (V320 & \V96(19) )),
  V331 = \V138(4)  & (V321 & (V320 & \V96(18) )),
  V332 = \V138(4)  & (V321 & (V320 & \V96(17) )),
  V333 = \V138(4)  & (V321 & (V320 & \V96(16) )),
  V334 = \V138(4)  & (V321 & (V320 & \V96(15) )),
  V335 = \V138(4)  & (V321 & (V320 & \V96(14) )),
  V336 = \V138(4)  & (V321 & (V320 & \V96(13) )),
  V337 = \V138(4)  & (V321 & (V320 & \V96(12) )),
  \V166(15)  = \[12] ,
  V338 = \V138(4)  & (V321 & (V320 & \V96(11) )),
  V339 = \V138(4)  & (V321 & (V320 & \V96(10) )),
  V340 = \V138(4)  & (V321 & (V320 & \V96(9) )),
  V341 = \V138(4)  & (V321 & (V320 & \V96(8) )),
  V342 = \V138(4)  & (V321 & (V320 & \V96(7) )),
  V343 = \V138(4)  & (V321 & (V320 & \V96(6) )),
  V344 = \V138(4)  & (V321 & (V320 & \V96(5) )),
  V345 = \V138(4)  & (V321 & (V320 & \V96(4) )),
  V346 = \V138(4)  & (V321 & (V320 & \V96(3) )),
  V347 = \V138(4)  & (V321 & (V320 & \V96(2) )),
  \V166(14)  = \[13] ,
  V348 = \V138(4)  & (V321 & (V320 & \V96(1) )),
  V349 = \V138(4)  & (V321 & (V320 & \V96(0) )),
  V350 = \V138(4)  & (V321 & (V320 & \V32(31) )),
  V351 = \V138(4)  & (V321 & (V320 & \V32(30) )),
  V352 = \V138(4)  & (V321 & (V320 & \V32(29) )),
  V353 = \V138(4)  & (V321 & (V320 & \V32(28) )),
  V354 = \V138(4)  & (V321 & (\V138(0)  & \V131(27) )),
  V355 = \V138(4)  & (V321 & (\V138(0)  & \V131(26) )),
  V356 = \V138(4)  & (V321 & (\V138(0)  & \V131(25) )),
  V357 = \V138(4)  & (V321 & (\V138(0)  & \V131(24) )),
  V358 = \V138(4)  & (V321 & (\V138(0)  & \V131(23) )),
  V359 = \V138(4)  & (V321 & (\V138(0)  & \V131(22) )),
  V360 = \V138(4)  & (V321 & (\V138(0)  & \V131(21) )),
  V361 = \V138(4)  & (V321 & (\V138(0)  & \V131(20) )),
  V362 = \V138(4)  & (V321 & (\V138(0)  & \V131(19) )),
  V363 = \V138(4)  & (V321 & (\V138(0)  & \V131(18) )),
  V364 = \V138(4)  & (V321 & (\V138(0)  & \V131(17) )),
  V365 = \V138(4)  & (V321 & (\V138(0)  & \V131(16) )),
  V366 = \V138(4)  & (V321 & (\V138(0)  & \V131(15) )),
  V367 = \V138(4)  & (V321 & (\V138(0)  & \V131(14) )),
  V368 = \V138(4)  & (V321 & (\V138(0)  & \V131(13) )),
  V369 = \V138(4)  & (V321 & (\V138(0)  & \V131(12) )),
  V370 = \V138(4)  & (V321 & (\V138(0)  & \V131(11) )),
  V371 = \V138(4)  & (V321 & (\V138(0)  & \V131(10) )),
  V372 = \V138(4)  & (V321 & (\V138(0)  & \V131(9) )),
  V373 = \V138(4)  & (V321 & (\V138(0)  & \V131(8) )),
  V374 = \V138(4)  & (V321 & (\V138(0)  & \V131(7) )),
  V375 = \V138(4)  & (V321 & (\V138(0)  & \V131(6) )),
  V376 = \V138(4)  & (V321 & (\V138(0)  & \V131(5) )),
  V377 = \V138(4)  & (V321 & (\V138(0)  & \V131(4) )),
  V378 = \V138(4)  & (V321 & (\V138(0)  & \V131(3) )),
  V379 = \V138(4)  & (V321 & (\V138(0)  & \V131(2) )),
  V380 = \V138(4)  & (V321 & (\V138(0)  & \V131(1) )),
  V381 = \V138(4)  & (V321 & (\V138(0)  & \V131(0) )),
  V382 = \V138(4)  & (V321 & (\V138(0)  & \V64(31) )),
  V383 = \V138(4)  & (V321 & (\V138(0)  & \V64(30) )),
  V384 = \V138(4)  & (V321 & (\V138(0)  & \V64(29) )),
  V385 = \V138(4)  & (V321 & (\V138(0)  & \V64(28) )),
  V418 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(27) )),
  V419 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(26) )),
  V420 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(25) )),
  V421 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(24) )),
  V422 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(23) )),
  V423 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(22) )),
  V424 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(21) )),
  V425 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(20) )),
  V426 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(19) )),
  V427 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(18) )),
  V428 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(17) )),
  V429 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(16) )),
  V430 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(15) )),
  V431 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(14) )),
  V432 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(13) )),
  V433 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(12) )),
  V434 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(11) )),
  V435 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(10) )),
  V436 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(9) )),
  V437 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(8) )),
  V438 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(7) )),
  V439 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(6) )),
  V440 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(5) )),
  V441 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(4) )),
  V442 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(3) )),
  V443 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(2) )),
  V444 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(1) )),
  V445 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V417(0) )),
  V446 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V389(3) )),
  V447 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V389(2) )),
  V448 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V389(1) )),
  V449 = \V138(4)  & (\V138(2)  & (\V138(0)  & \V389(0) )),
  V450 = ~\V138(4) ,
  V451 = V450 & \V138(2) ,
  V452 = ~\V138(0) ,
  V453 = ~\V138(2) ,
  V454 = \V138(3)  & (V453 & (V452 & \V99(0) )),
  V455 = \V138(3)  & (V453 & (V452 & \V98(0) )),
  V456 = \V138(3)  & (V453 & (V452 & \V97(0) )),
  V457 = \V138(3)  & (V453 & (V452 & \V96(31) )),
  V458 = \V138(3)  & (V453 & (V452 & \V96(30) )),
  V459 = \V138(3)  & (V453 & (V452 & \V96(29) )),
  V460 = \V138(3)  & (V453 & (V452 & \V96(28) )),
  V461 = \V138(3)  & (V453 & (\V138(0)  & \V134(0) )),
  V462 = \V138(3)  & (V453 & (\V138(0)  & \V133(1) )),
  V463 = \V138(3)  & (V453 & (\V138(0)  & \V133(0) )),
  V464 = \V138(3)  & (V453 & (\V138(0)  & \V131(31) )),
  V465 = \V138(3)  & (V453 & (\V138(0)  & \V131(30) )),
  V466 = \V138(3)  & (V453 & (\V138(0)  & \V131(29) )),
  V467 = \V138(3)  & (V453 & (\V138(0)  & \V131(28) )),
  V474 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V134(0) )),
  V475 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V473(1) )),
  V476 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V473(0) )),
  V477 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V471(3) )),
  V478 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V471(2) )),
  V479 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V471(1) )),
  \V417(3)  = ~\V131(3) ,
  V480 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V471(0) )),
  V481 = ~\V138(3) ,
  V482 = V481 & \V138(2) ,
  \V417(2)  = ~\V131(2) ,
  \V417(5)  = ~\V131(5) ,
  \V417(4)  = ~\V131(4) ,
  \[10]  = V302 | (V246 | V218),
  \[11]  = V303 | (V247 | V219),
  \[12]  = V304 | (V248 | V220),
  \V417(1)  = ~\V131(1) ,
  \[13]  = V305 | (V249 | V221),
  \V417(0)  = ~\V131(0) ,
  \[14]  = V306 | (V250 | V222),
  \[15]  = V307 | (V251 | V223),
  \[16]  = V308 | (V252 | V224),
  \[17]  = V309 | (V253 | V225),
  \[18]  = V310 | (V254 | V226),
  \V417(7)  = ~\V131(7) ,
  \[19]  = V311 | (V255 | V227),
  \V417(6)  = ~\V131(6) ,
  \V417(9)  = ~\V131(9) ,
  \V417(8)  = ~\V131(8) ,
  \[20]  = V312 | (V256 | V228),
  \[21]  = V313 | (V257 | V229),
  \[22]  = V314 | (V258 | V230),
  \[23]  = V315 | (V259 | V231),
  \[24]  = V316 | (V260 | V232),
  \[25]  = V317 | (V261 | V233),
  \[26]  = V318 | (V262 | V234),
  \[27]  = V319 | (V263 | V235),
  \[28]  = V451 | (V418 | (V354 | V322)),
  \V471(3)  = ~\V131(31) ,
  \[29]  = V451 | (V419 | (V355 | V323)),
  \V471(2)  = ~\V131(30) ,
  \V471(1)  = ~\V131(29) ,
  \V471(0)  = ~\V131(28) ,
  \[30]  = V451 | (V420 | (V356 | V324)),
  \[31]  = V451 | (V421 | (V357 | V325)),
  \[32]  = V451 | (V422 | (V358 | V326)),
  \[33]  = V451 | (V423 | (V359 | V327)),
  \[34]  = V451 | (V424 | (V360 | V328)),
  \[35]  = V451 | (V425 | (V361 | V329)),
  \[36]  = V451 | (V426 | (V362 | V330)),
  \[37]  = V451 | (V427 | (V363 | V331)),
  \[38]  = V451 | (V428 | (V364 | V332)),
  \V291(3)  = ~\V64(3) ,
  \[39]  = V451 | (V429 | (V365 | V333)),
  \V291(2)  = ~\V64(2) ,
  \V291(5)  = ~\V64(5) ,
  \V291(4)  = ~\V64(4) ,
  \V291(1)  = ~\V64(1) ,
  \V291(0)  = ~\V64(0) ,
  \[40]  = V451 | (V430 | (V366 | V334)),
  \[41]  = V451 | (V431 | (V367 | V335)),
  \[42]  = V451 | (V432 | (V368 | V336)),
  \[43]  = V451 | (V433 | (V369 | V337)),
  \[44]  = V451 | (V434 | (V370 | V338)),
  \V291(7)  = ~\V64(7) ,
  \V473(1)  = ~\V133(1) ,
  \[45]  = V451 | (V435 | (V371 | V339)),
  \V291(6)  = ~\V64(6) ,
  \V473(0)  = ~\V133(0) ,
  \[46]  = V451 | (V436 | (V372 | V340)),
  \V291(9)  = ~\V64(9) ,
  \[47]  = V451 | (V437 | (V373 | V341)),
  \V291(8)  = ~\V64(8) ,
  \[48]  = V451 | (V438 | (V374 | V342)),
  \[49]  = V451 | (V439 | (V375 | V343)),
  \[50]  = V451 | (V440 | (V376 | V344)),
  \[51]  = V451 | (V441 | (V377 | V345)),
  \[52]  = V451 | (V442 | (V378 | V346)),
  \[53]  = V451 | (V443 | (V379 | V347)),
  \[54]  = V451 | (V444 | (V380 | V348)),
  \[55]  = V451 | (V445 | (V381 | V349)),
  \[56]  = V451 | (V446 | (V382 | V350)),
  \[57]  = V451 | (V447 | (V383 | V351)),
  \[58]  = V451 | (V448 | (V384 | V352)),
  \[59]  = V451 | (V449 | (V385 | V353)),
  \[60]  = V474 | (V461 | V454),
  \[61]  = V482 | (V475 | (V462 | V455)),
  \[62]  = V482 | (V476 | (V463 | V456)),
  \[63]  = V482 | (V477 | (V464 | V457)),
  \V198(27)  = \[32] ,
  \[64]  = V482 | (V478 | (V465 | V458)),
  \V198(26)  = \[33] ,
  \[65]  = V482 | (V479 | (V466 | V459)),
  \V198(29)  = \[30] ,
  \[66]  = V482 | (V480 | (V467 | V460)),
  \V198(28)  = \[31] ,
  \V198(21)  = \[38] ,
  \V198(20)  = \[39] ,
  \V198(23)  = \[36] ,
  \V198(22)  = \[37] ,
  \V198(25)  = \[34] ,
  \V198(24)  = \[35] ,
  \V291(27)  = ~\V64(27) ,
  \V198(17)  = \[42] ,
  \V291(26)  = ~\V64(26) ,
  \V198(16)  = \[43] ,
  \V198(19)  = \[40] ,
  \V198(18)  = \[41] ;
endmodule

