module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 ;
output g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
     n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , 
     n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , 
     n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , 
     n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
     n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
     n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
     n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
     n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , 
     n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , 
     n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , 
     n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , 
     n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , 
     n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , 
     n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , 
     n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , 
     n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , 
     n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
     n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
     n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
     n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
     n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
     n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , 
     n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
     n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
     n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
     n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
     n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
     n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
     n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
     n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
     n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
     n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
     n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
     n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
     n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
     n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
     n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
     n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
     n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
     n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
     n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
     n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
     n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
     n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
     n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
     n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
     n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
     n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
     n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , 
     n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , 
     n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , 
     n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , 
     n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , 
     n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , 
     n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , 
     n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , 
     n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , 
     n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , 
     n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , 
     n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , 
     n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , 
     n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , 
     n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , 
     n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , 
     n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , 
     n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , 
     n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , 
     n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , 
     n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , 
     n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , 
     n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , 
     n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , 
     n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , 
     n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , 
     n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , 
     n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , 
     n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , 
     n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , 
     n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , 
     n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , 
     n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , 
     n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , 
     n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , 
     n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , 
     n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , 
     n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , 
     n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , 
     n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , 
     n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , 
     n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , 
     n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , 
     n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , 
     n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , 
     n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , 
     n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , 
     n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , 
     n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , 
     n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , 
     n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , 
     n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , 
     n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , 
     n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , 
     n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , 
     n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , 
     n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , 
     n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , 
     n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , 
     n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , 
     n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , 
     n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , 
     n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , 
     n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , 
     n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , 
     n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , 
     n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , 
     n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
     n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
     n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , 
     n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , 
     n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , 
     n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , 
     n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , 
     n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , 
     n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , 
     n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , 
     n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , 
     n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , 
     n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , 
     n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , 
     n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , 
     n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , 
     n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , 
     n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , 
     n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , 
     n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , 
     n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , 
     n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , 
     n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , 
     n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , 
     n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , 
     n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , 
     n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , 
     n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , 
     n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , 
     n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , 
     n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , 
     n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , 
     n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , 
     n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , 
     n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , 
     n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , 
     n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , 
     n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , 
     n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , 
     n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , 
     n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , 
     n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , 
     n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , 
     n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , 
     n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , 
     n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , 
     n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , 
     n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , 
     n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , 
     n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , 
     n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , 
     n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , 
     n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , 
     n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , 
     n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , 
     n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , 
     n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , 
     n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , 
     n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , 
     n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , 
     n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , 
     n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , 
     n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , 
     n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , 
     n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , 
     n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , 
     n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , 
     n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , 
     n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , 
     n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , 
     n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , 
     n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , 
     n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , 
     n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , 
     n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , 
     n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , 
     n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , 
     n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , 
     n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , 
     n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , 
     n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , 
     n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , 
     n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , 
     n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , 
     n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , 
     n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , 
     n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , 
     n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , 
     n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , 
     n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , 
     n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , 
     n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , 
     n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , 
     n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , 
     n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , 
     n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , 
     n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , 
     n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , 
     n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , 
     n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , 
     n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , 
     n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , 
     n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , 
     n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , 
     n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , 
     n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , 
     n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , 
     n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , 
     n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , 
     n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , 
     n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , 
     n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , 
     n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , 
     n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , 
     n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , 
     n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , 
     n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , 
     n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , 
     n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , 
     n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , 
     n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , 
     n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , 
     n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , 
     n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , 
     n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , 
     n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , 
     n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , 
     n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , 
     n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , 
     n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , 
     n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , 
     n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , 
     n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , 
     n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , 
     n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , 
     n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , 
     n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , 
     n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , 
     n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , 
     n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , 
     n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , 
     n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , 
     n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , 
     n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , 
     n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , 
     n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , 
     n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , 
     n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , 
     n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , 
     n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , 
     n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , 
     n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , 
     n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , 
     n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , 
     n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , 
     n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , 
     n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , 
     n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , 
     n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , 
     n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , 
     n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , 
     n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , 
     n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , 
     n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , 
     n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , 
     n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , 
     n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , 
     n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , 
     n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , 
     n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , 
     n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , 
     n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , 
     n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , 
     n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , 
     n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , 
     n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , 
     n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , 
     n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , 
     n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , 
     n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , 
     n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , 
     n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , 
     n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , 
     n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , 
     n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , 
     n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , 
     n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , 
     n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , 
     n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , 
     n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , 
     n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , 
     n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , 
     n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , 
     n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , 
     n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , 
     n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , 
     n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , 
     n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , 
     n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , 
     n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , 
     n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , 
     n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , 
     n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , 
     n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , 
     n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , 
     n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , 
     n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , 
     n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , 
     n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , 
     n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , 
     n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , 
     n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , 
     n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , 
     n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , 
     n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , 
     n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , 
     n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , 
     n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , 
     n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , 
     n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , 
     n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , 
     n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , 
     n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , 
     n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , 
     n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , 
     n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , 
     n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , 
     n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , 
     n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , 
     n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , 
     n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , 
     n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , 
     n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , 
     n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , 
     n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , 
     n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , 
     n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , 
     n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , 
     n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , 
     n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , 
     n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , 
     n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , 
     n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , 
     n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , 
     n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , 
     n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , 
     n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , 
     n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , 
     n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , 
     n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , 
     n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , 
     n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , 
     n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , 
     n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , 
     n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , 
     n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , 
     n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , 
     n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , 
     n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , 
     n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , 
     n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , 
     n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , 
     n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , 
     n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , 
     n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , 
     n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , 
     n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , 
     n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , 
     n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , 
     n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , 
     n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , 
     n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , 
     n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , 
     n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , 
     n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , 
     n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , 
     n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , 
     n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , 
     n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , 
     n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , 
     n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , 
     n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , 
     n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , 
     n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , 
     n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , 
     n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , 
     n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , 
     n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , 
     n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , 
     n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , 
     n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , 
     n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , 
     n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , 
     n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , 
     n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , 
     n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , 
     n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , 
     n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , 
     n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , 
     n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , 
     n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , 
     n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , 
     n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , 
     n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , 
     n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , 
     n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , 
     n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , 
     n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , 
     n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , 
     n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , 
     n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , 
     n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , 
     n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , 
     n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , 
     n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , 
     n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , 
     n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , 
     n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , 
     n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , 
     n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , 
     n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , 
     n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , 
     n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , 
     n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , 
     n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , 
     n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , 
     n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , 
     n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , 
     n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , 
     n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , 
     n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , 
     n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , 
     n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , 
     n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , 
     n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , 
     n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , 
     n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , 
     n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , 
     n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , 
     n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , 
     n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , 
     n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , 
     n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , 
     n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , 
     n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , 
     n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , 
     n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , 
     n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , 
     n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , 
     n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , 
     n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , 
     n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , 
     n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , 
     n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , 
     n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , 
     n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , 
     n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , 
     n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , 
     n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , 
     n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , 
     n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , 
     n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , 
     n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , 
     n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , 
     n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , 
     n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , 
     n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , 
     n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , 
     n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , 
     n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , 
     n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , 
     n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , 
     n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , 
     n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , 
     n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , 
     n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , 
     n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , 
     n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , 
     n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , 
     n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , 
     n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , 
     n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , 
     n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , 
     n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , 
     n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , 
     n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , 
     n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , 
     n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , 
     n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , 
     n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , 
     n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , 
     n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , 
     n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , 
     n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , 
     n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , 
     n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , 
     n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , 
     n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , 
     n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , 
     n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , 
     n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , 
     n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , 
     n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , 
     n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , 
     n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , 
     n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , 
     n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , 
     n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , 
     n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , 
     n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , 
     n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , 
     n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , 
     n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , 
     n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , 
     n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , 
     n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , 
     n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , 
     n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , 
     n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , 
     n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , 
     n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , 
     n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , 
     n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , 
     n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , 
     n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , 
     n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , 
     n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , 
     n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , 
     n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , 
     n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , 
     n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , 
     n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , 
     n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , 
     n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , 
     n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , 
     n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , 
     n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , 
     n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , 
     n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , 
     n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , 
     n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , 
     n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , 
     n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , 
     n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , 
     n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , 
     n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , 
     n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , 
     n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , 
     n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , 
     n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , 
     n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , 
     n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , 
     n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , 
     n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , 
     n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , 
     n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , 
     n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , 
     n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , 
     n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , 
     n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , 
     n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , 
     n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , 
     n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , 
     n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , 
     n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , 
     n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , 
     n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , 
     n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , 
     n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , 
     n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , 
     n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , 
     n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , 
     n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , 
     n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , 
     n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , 
     n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , 
     n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , 
     n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , 
     n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , 
     n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , 
     n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , 
     n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , 
     n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , 
     n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , 
     n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , 
     n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , 
     n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , 
     n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , 
     n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , 
     n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , 
     n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , 
     n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , 
     n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , 
     n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , 
     n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , 
     n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , 
     n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , 
     n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , 
     n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , 
     n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
     n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
     n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , 
     n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , 
     n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , 
     n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , 
     n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , 
     n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , 
     n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , 
     n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , 
     n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , 
     n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , 
     n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , 
     n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , 
     n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , 
     n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , 
     n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , 
     n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , 
     n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , 
     n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , 
     n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , 
     n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , 
     n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , 
     n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , 
     n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , 
     n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , 
     n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , 
     n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , 
     n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , 
     n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , 
     n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , 
     n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , 
     n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , 
     n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , 
     n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , 
     n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , 
     n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , 
     n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , 
     n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , 
     n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , 
     n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , 
     n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , 
     n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , 
     n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , 
     n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , 
     n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , 
     n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , 
     n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , 
     n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , 
     n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , 
     n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , 
     n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , 
     n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , 
     n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , 
     n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , 
     n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , 
     n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , 
     n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , 
     n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , 
     n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , 
     n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , 
     n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , 
     n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , 
     n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , 
     n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , 
     n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , 
     n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , 
     n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , 
     n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , 
     n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , 
     n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , 
     n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , 
     n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , 
     n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , 
     n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , 
     n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , 
     n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , 
     n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , 
     n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , 
     n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , 
     n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , 
     n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , 
     n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , 
     n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , 
     n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , 
     n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , 
     n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , 
     n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , 
     n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , 
     n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , 
     n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , 
     n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , 
     n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , 
     n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , 
     n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , 
     n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , 
     n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , 
     n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , 
     n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , 
     n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , 
     n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , 
     n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , 
     n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , 
     n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , 
     n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , 
     n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , 
     n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , 
     n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , 
     n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , 
     n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , 
     n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , 
     n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , 
     n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , 
     n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , 
     n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , 
     n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , 
     n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , 
     n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , 
     n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , 
     n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , 
     n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , 
     n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , 
     n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , 
     n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , 
     n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , 
     n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , 
     n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , 
     n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , 
     n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , 
     n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , 
     n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , 
     n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , 
     n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , 
     n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , 
     n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , 
     n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , 
     n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , 
     n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , 
     n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , 
     n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , 
     n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , 
     n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , 
     n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , 
     n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , 
     n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , 
     n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , 
     n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , 
     n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , 
     n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , 
     n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , 
     n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , 
     n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , 
     n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , 
     n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , 
     n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , 
     n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , 
     n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , 
     n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , 
     n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , 
     n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , 
     n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , 
     n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , 
     n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , 
     n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , 
     n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , 
     n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , 
     n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , 
     n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , 
     n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , 
     n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , 
     n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , 
     n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , 
     n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , 
     n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , 
     n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , 
     n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , 
     n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , 
     n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , 
     n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , 
     n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , 
     n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , 
     n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , 
     n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , 
     n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , 
     n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , 
     n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , 
     n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , 
     n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , 
     n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , 
     n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , 
     n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , 
     n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , 
     n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , 
     n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , 
     n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , 
     n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , 
     n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , 
     n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , 
     n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , 
     n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , 
     n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , 
     n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , 
     n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , 
     n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , 
     n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , 
     n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , 
     n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , 
     n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , 
     n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , 
     n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , 
     n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , 
     n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , 
     n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , 
     n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , 
     n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , 
     n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , 
     n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , 
     n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , 
     n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , 
     n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , 
     n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , 
     n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , 
     n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , 
     n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , 
     n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , 
     n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , 
     n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , 
     n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , 
     n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , 
     n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , 
     n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , 
     n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , 
     n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , 
     n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , 
     n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , 
     n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , 
     n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , 
     n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , 
     n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , 
     n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , 
     n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , 
     n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , 
     n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , 
     n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , 
     n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , 
     n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , 
     n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , 
     n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , 
     n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , 
     n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , 
     n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , 
     n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , 
     n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , 
     n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , 
     n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , 
     n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , 
     n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , 
     n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , 
     n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , 
     n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , 
     n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , 
     n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , 
     n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , 
     n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , 
     n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , 
     n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , 
     n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , 
     n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , 
     n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , 
     n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , 
     n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , 
     n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , 
     n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , 
     n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , 
     n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , 
     n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , 
     n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , 
     n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , 
     n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , 
     n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , 
     n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , 
     n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , 
     n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , 
     n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , 
     n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , 
     n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , 
     n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , 
     n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , 
     n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , 
     n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , 
     n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , 
     n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , 
     n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , 
     n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , 
     n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , 
     n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , 
     n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , 
     n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , 
     n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , 
     n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , 
     n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , 
     n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , 
     n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , 
     n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , 
     n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , 
     n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , 
     n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , 
     n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , 
     n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , 
     n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , 
     n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , 
     n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , 
     n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , 
     n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , 
     n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , 
     n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , 
     n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , 
     n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , 
     n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , 
     n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , 
     n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , 
     n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , 
     n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , 
     n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , 
     n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , 
     n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , 
     n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , 
     n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , 
     n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , 
     n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , 
     n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , 
     n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , 
     n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , 
     n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , 
     n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , 
     n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , 
     n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , 
     n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , 
     n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , 
     n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , 
     n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , 
     n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , 
     n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , 
     n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , 
     n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , 
     n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , 
     n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , 
     n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , 
     n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , 
     n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , 
     n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , 
     n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , 
     n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , 
     n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , 
     n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , 
     n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , 
     n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , 
     n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , 
     n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , 
     n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , 
     n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , 
     n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , 
     n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , 
     n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , 
     n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , 
     n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , 
     n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , 
     n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , 
     n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , 
     n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , 
     n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , 
     n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , 
     n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , 
     n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , 
     n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , 
     n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , 
     n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , 
     n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , 
     n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , 
     n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , 
     n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , 
     n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , 
     n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , 
     n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , 
     n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , 
     n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , 
     n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , 
     n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , 
     n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , 
     n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , 
     n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , 
     n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , 
     n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , 
     n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , 
     n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , 
     n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , 
     n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , 
     n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , 
     n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , 
     n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , 
     n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , 
     n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , 
     n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , 
     n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , 
     n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , 
     n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , 
     n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , 
     n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , 
     n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , 
     n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , 
     n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , 
     n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , 
     n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , 
     n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , 
     n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , 
     n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , 
     n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , 
     n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , 
     n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , 
     n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , 
     n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , 
     n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , 
     n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , 
     n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , 
     n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , 
     n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , 
     n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , 
     n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , 
     n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , 
     n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , 
     n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , 
     n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , 
     n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , 
     n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , 
     n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , 
     n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , 
     n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , 
     n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , 
     n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , 
     n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , 
     n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , 
     n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , 
     n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , 
     n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , 
     n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , 
     n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , 
     n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , 
     n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , 
     n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , 
     n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , 
     n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , 
     n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , 
     n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , 
     n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , 
     n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , 
     n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , 
     n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , 
     n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , 
     n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , 
     n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , 
     n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , 
     n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , 
     n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , 
     n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , 
     n24070 , n24071 , n24072 , n24073 , n24074 , n24075 ;
wire t_0 , t_1 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( n246 , g245 );
buf ( n247 , g246 );
buf ( n248 , g247 );
buf ( n249 , g248 );
buf ( n250 , g249 );
buf ( n251 , g250 );
buf ( n252 , g251 );
buf ( n253 , g252 );
buf ( n254 , g253 );
buf ( n255 , g254 );
buf ( n256 , g255 );
buf ( n257 , g256 );
buf ( n258 , g257 );
buf ( n259 , g258 );
buf ( n260 , g259 );
buf ( n261 , g260 );
buf ( n262 , g261 );
buf ( n263 , g262 );
buf ( n264 , g263 );
buf ( n265 , g264 );
buf ( n266 , g265 );
buf ( n267 , g266 );
buf ( n268 , g267 );
buf ( n269 , g268 );
buf ( n270 , g269 );
buf ( n271 , g270 );
buf ( n272 , g271 );
buf ( n273 , g272 );
buf ( n274 , g273 );
buf ( n275 , g274 );
buf ( n276 , g275 );
buf ( n277 , g276 );
buf ( n278 , g277 );
buf ( n279 , g278 );
buf ( n280 , g279 );
buf ( n281 , g280 );
buf ( n282 , g281 );
buf ( n283 , g282 );
buf ( n284 , g283 );
buf ( n285 , g284 );
buf ( n286 , g285 );
buf ( n287 , g286 );
buf ( n288 , g287 );
buf ( n289 , g288 );
buf ( n290 , g289 );
buf ( n291 , g290 );
buf ( n292 , g291 );
buf ( n293 , g292 );
buf ( n294 , g293 );
buf ( n295 , g294 );
buf ( n296 , g295 );
buf ( n297 , g296 );
buf ( n298 , g297 );
buf ( n299 , g298 );
buf ( n300 , g299 );
buf ( n301 , g300 );
buf ( n302 , g301 );
buf ( n303 , g302 );
buf ( n304 , g303 );
buf ( n305 , g304 );
buf ( n306 , g305 );
buf ( n307 , g306 );
buf ( n308 , g307 );
buf ( n309 , g308 );
buf ( n310 , g309 );
buf ( n311 , g310 );
buf ( n312 , g311 );
buf ( n313 , g312 );
buf ( n314 , g313 );
buf ( n315 , g314 );
buf ( n316 , g315 );
buf ( n317 , g316 );
buf ( n318 , g317 );
buf ( n319 , g318 );
buf ( n320 , g319 );
buf ( n321 , g320 );
buf ( n322 , g321 );
buf ( n323 , g322 );
buf ( n324 , g323 );
buf ( n325 , g324 );
buf ( n326 , g325 );
buf ( n327 , g326 );
buf ( n328 , g327 );
buf ( n329 , g328 );
buf ( n330 , g329 );
buf ( n331 , g330 );
buf ( n332 , g331 );
buf ( n333 , g332 );
buf ( n334 , g333 );
buf ( n335 , g334 );
buf ( n336 , g335 );
buf ( n337 , g336 );
buf ( n338 , g337 );
buf ( n339 , g338 );
buf ( n340 , g339 );
buf ( n341 , g340 );
buf ( n342 , g341 );
buf ( n343 , g342 );
buf ( n344 , g343 );
buf ( n345 , g344 );
buf ( n346 , g345 );
buf ( n347 , g346 );
buf ( n348 , g347 );
buf ( n349 , g348 );
buf ( n350 , g349 );
buf ( n351 , g350 );
buf ( n352 , g351 );
buf ( n353 , g352 );
buf ( n354 , g353 );
buf ( n355 , g354 );
buf ( n356 , g355 );
buf ( n357 , g356 );
buf ( n358 , g357 );
buf ( n359 , g358 );
buf ( n360 , g359 );
buf ( n361 , g360 );
buf ( n362 , g361 );
buf ( n363 , g362 );
buf ( n364 , g363 );
buf ( n365 , g364 );
buf ( n366 , g365 );
buf ( n367 , g366 );
buf ( n368 , g367 );
buf ( n369 , g368 );
buf ( n370 , g369 );
buf ( n371 , g370 );
buf ( n372 , g371 );
buf ( n373 , g372 );
buf ( n374 , g373 );
buf ( n375 , g374 );
buf ( n376 , g375 );
buf ( n377 , g376 );
buf ( n378 , g377 );
buf ( n379 , g378 );
buf ( n380 , g379 );
buf ( n381 , g380 );
buf ( n382 , g381 );
buf ( n383 , g382 );
buf ( n384 , g383 );
buf ( n385 , g384 );
buf ( n386 , g385 );
buf ( n387 , g386 );
buf ( n388 , g387 );
buf ( n389 , g388 );
buf ( n390 , g389 );
buf ( n391 , g390 );
buf ( n392 , g391 );
buf ( n393 , g392 );
buf ( n394 , g393 );
buf ( n395 , g394 );
buf ( n396 , g395 );
buf ( n397 , g396 );
buf ( n398 , g397 );
buf ( n399 , g398 );
buf ( n400 , g399 );
buf ( n401 , g400 );
buf ( n402 , g401 );
buf ( n403 , g402 );
buf ( n404 , g403 );
buf ( n405 , g404 );
buf ( n406 , g405 );
buf ( n407 , g406 );
buf ( n408 , g407 );
buf ( n409 , g408 );
buf ( n410 , g409 );
buf ( n411 , g410 );
buf ( n412 , g411 );
buf ( n413 , g412 );
buf ( n414 , g413 );
buf ( n415 , g414 );
buf ( n416 , g415 );
buf ( n417 , g416 );
buf ( n418 , g417 );
buf ( n419 , g418 );
buf ( n420 , g419 );
buf ( n421 , g420 );
buf ( n422 , g421 );
buf ( n423 , g422 );
buf ( n424 , g423 );
buf ( n425 , g424 );
buf ( n426 , g425 );
buf ( n427 , g426 );
buf ( n428 , g427 );
buf ( n429 , g428 );
buf ( n430 , g429 );
buf ( n431 , g430 );
buf ( n432 , g431 );
buf ( n433 , g432 );
buf ( n434 , g433 );
buf ( n435 , g434 );
buf ( n436 , g435 );
buf ( n437 , g436 );
buf ( n438 , g437 );
buf ( n439 , g438 );
buf ( n440 , g439 );
buf ( n441 , g440 );
buf ( n442 , g441 );
buf ( n443 , g442 );
buf ( n444 , g443 );
buf ( n445 , g444 );
buf ( n446 , g445 );
buf ( n447 , g446 );
buf ( n448 , g447 );
buf ( n449 , g448 );
buf ( n450 , g449 );
buf ( g450 , n451 );
buf ( g451 , n452 );
buf ( g452 , n453 );
buf ( g453 , n454 );
buf ( g454 , n455 );
buf ( g455 , n456 );
buf ( g456 , n457 );
buf ( g457 , n458 );
buf ( g458 , n459 );
buf ( g459 , n460 );
buf ( g460 , n461 );
buf ( g461 , n462 );
buf ( g462 , n463 );
buf ( g463 , n464 );
buf ( g464 , n465 );
buf ( g465 , n466 );
buf ( g466 , n467 );
buf ( g467 , n468 );
buf ( g468 , n469 );
buf ( g469 , n470 );
buf ( g470 , n471 );
buf ( g471 , n472 );
buf ( g472 , n473 );
buf ( g473 , n474 );
buf ( g474 , n475 );
buf ( g475 , n476 );
buf ( g476 , n477 );
buf ( g477 , n478 );
buf ( g478 , n479 );
buf ( g479 , n480 );
buf ( g480 , n481 );
buf ( g481 , n482 );
buf ( g482 , n483 );
buf ( g483 , n484 );
buf ( g484 , n485 );
buf ( g485 , n486 );
buf ( g486 , n487 );
buf ( g487 , n488 );
buf ( g488 , n489 );
buf ( g489 , n490 );
buf ( g490 , n491 );
buf ( g491 , n492 );
buf ( g492 , n493 );
buf ( g493 , n494 );
buf ( g494 , n495 );
buf ( g495 , n496 );
buf ( g496 , n497 );
buf ( g497 , n498 );
buf ( g498 , n499 );
buf ( g499 , n500 );
buf ( g500 , n501 );
buf ( g501 , n502 );
buf ( g502 , n503 );
buf ( g503 , n504 );
buf ( g504 , n505 );
buf ( g505 , n506 );
buf ( g506 , n507 );
buf ( g507 , n508 );
buf ( g508 , n509 );
buf ( g509 , n510 );
buf ( g510 , n511 );
buf ( g511 , n512 );
buf ( g512 , n513 );
buf ( g513 , n514 );
buf ( g514 , n515 );
buf ( g515 , n516 );
buf ( g516 , n517 );
buf ( g517 , n518 );
buf ( g518 , n519 );
buf ( g519 , n520 );
buf ( g520 , n521 );
buf ( g521 , n522 );
buf ( g522 , n523 );
buf ( g523 , n524 );
buf ( g524 , n525 );
buf ( g525 , n526 );
buf ( g526 , n527 );
buf ( g527 , n528 );
buf ( g528 , n529 );
buf ( g529 , n530 );
buf ( g530 , n531 );
buf ( g531 , n532 );
buf ( g532 , n533 );
buf ( g533 , n534 );
buf ( g534 , n535 );
buf ( g535 , n536 );
buf ( g536 , n537 );
buf ( g537 , n538 );
buf ( g538 , n539 );
buf ( g539 , n540 );
buf ( g540 , n541 );
buf ( g541 , n542 );
buf ( g542 , n543 );
buf ( g543 , n544 );
buf ( g544 , n545 );
buf ( g545 , n546 );
buf ( g546 , n547 );
buf ( g547 , n548 );
buf ( g548 , n549 );
buf ( g549 , n550 );
buf ( g550 , n551 );
buf ( g551 , n552 );
buf ( g552 , n553 );
buf ( g553 , n554 );
buf ( g554 , n555 );
buf ( g555 , n556 );
buf ( g556 , n557 );
buf ( g557 , n558 );
buf ( g558 , n559 );
buf ( g559 , n560 );
buf ( g560 , n561 );
buf ( g561 , n562 );
buf ( g562 , n563 );
buf ( g563 , n564 );
buf ( g564 , n565 );
buf ( g565 , n566 );
buf ( g566 , n567 );
buf ( g567 , n568 );
buf ( g568 , n569 );
buf ( g569 , n570 );
buf ( g570 , n571 );
buf ( g571 , n572 );
buf ( g572 , n573 );
buf ( g573 , n574 );
buf ( g574 , n575 );
buf ( g575 , n576 );
buf ( g576 , n577 );
buf ( g577 , n578 );
buf ( g578 , n579 );
buf ( g579 , n580 );
buf ( g580 , n581 );
buf ( g581 , n582 );
buf ( g582 , n583 );
buf ( g583 , n584 );
buf ( g584 , n585 );
buf ( g585 , n586 );
buf ( g586 , n587 );
buf ( g587 , n588 );
buf ( g588 , n589 );
buf ( g589 , n590 );
buf ( g590 , n591 );
buf ( g591 , n592 );
buf ( g592 , n593 );
buf ( g593 , n594 );
buf ( g594 , n595 );
buf ( g595 , n596 );
buf ( g596 , n597 );
buf ( g597 , n598 );
buf ( g598 , n599 );
buf ( g599 , n600 );
buf ( g600 , n601 );
buf ( g601 , n602 );
buf ( g602 , n603 );
buf ( g603 , n604 );
buf ( g604 , n605 );
buf ( g605 , n606 );
buf ( g606 , n607 );
buf ( g607 , n608 );
buf ( g608 , n609 );
buf ( g609 , n610 );
buf ( g610 , n611 );
buf ( g611 , n612 );
buf ( g612 , n613 );
buf ( g613 , n614 );
buf ( g614 , n615 );
buf ( g615 , n616 );
buf ( g616 , n617 );
buf ( g617 , n618 );
buf ( g618 , n619 );
buf ( g619 , n620 );
buf ( g620 , n621 );
buf ( g621 , n622 );
buf ( g622 , n623 );
buf ( g623 , n624 );
buf ( g624 , n625 );
buf ( g625 , n626 );
buf ( g626 , n627 );
buf ( g627 , n628 );
buf ( g628 , n629 );
buf ( g629 , n630 );
buf ( g630 , n631 );
buf ( g631 , n632 );
buf ( g632 , n633 );
buf ( g633 , n634 );
buf ( g634 , n635 );
buf ( g635 , n636 );
buf ( g636 , n637 );
buf ( g637 , n638 );
buf ( g638 , n639 );
buf ( g639 , n640 );
buf ( g640 , n641 );
buf ( g641 , n642 );
buf ( g642 , n643 );
buf ( g643 , n644 );
buf ( g644 , n645 );
buf ( g645 , n646 );
buf ( g646 , n647 );
buf ( g647 , n648 );
buf ( g648 , n649 );
buf ( g649 , n650 );
buf ( g650 , n651 );
buf ( g651 , n652 );
buf ( g652 , n653 );
buf ( g653 , n654 );
buf ( g654 , n655 );
buf ( g655 , n656 );
buf ( g656 , n657 );
buf ( g657 , n658 );
buf ( g658 , n659 );
buf ( g659 , n660 );
buf ( g660 , n661 );
buf ( g661 , n662 );
buf ( g662 , n663 );
buf ( g663 , n664 );
buf ( g664 , n665 );
buf ( g665 , n666 );
buf ( g666 , n667 );
buf ( g667 , n668 );
buf ( g668 , n669 );
buf ( g669 , n670 );
buf ( g670 , n671 );
buf ( g671 , n672 );
buf ( g672 , n673 );
buf ( g673 , n674 );
buf ( g674 , n675 );
buf ( g675 , n676 );
buf ( g676 , n677 );
buf ( g677 , n678 );
buf ( g678 , n679 );
buf ( g679 , n680 );
buf ( g680 , n681 );
buf ( g681 , n682 );
buf ( g682 , n683 );
buf ( g683 , n684 );
buf ( g684 , n685 );
buf ( g685 , n686 );
buf ( g686 , n687 );
buf ( g687 , n688 );
buf ( g688 , n689 );
buf ( g689 , n690 );
buf ( g690 , n691 );
buf ( g691 , n692 );
buf ( g692 , n693 );
buf ( g693 , n694 );
buf ( g694 , n695 );
buf ( g695 , n696 );
buf ( g696 , n697 );
buf ( g697 , n698 );
buf ( g698 , n699 );
buf ( g699 , n700 );
buf ( g700 , n701 );
buf ( g701 , n702 );
buf ( g702 , n703 );
buf ( g703 , n704 );
buf ( g704 , n705 );
buf ( g705 , n706 );
buf ( g706 , n707 );
buf ( g707 , n708 );
buf ( g708 , n709 );
buf ( g709 , n710 );
buf ( g710 , n711 );
buf ( g711 , n712 );
buf ( g712 , n713 );
buf ( g713 , n714 );
buf ( g714 , n715 );
buf ( g715 , n716 );
buf ( g716 , n717 );
buf ( g717 , n718 );
buf ( g718 , n719 );
buf ( g719 , n720 );
buf ( g720 , n721 );
buf ( g721 , n722 );
buf ( g722 , n723 );
buf ( g723 , n724 );
buf ( g724 , n725 );
buf ( g725 , n726 );
buf ( g726 , n727 );
buf ( g727 , n728 );
buf ( g728 , n729 );
buf ( g729 , n730 );
buf ( g730 , n731 );
buf ( g731 , n732 );
buf ( n451 , n21374 );
buf ( n452 , n21613 );
buf ( n453 , n21773 );
buf ( n454 , n23489 );
buf ( n455 , n23508 );
buf ( n456 , n18510 );
buf ( n457 , n21802 );
buf ( n458 , n21819 );
buf ( n459 , n23493 );
buf ( n460 , n21835 );
buf ( n461 , n23824 );
buf ( n462 , n22761 );
buf ( n463 , n21859 );
buf ( n464 , n22790 );
buf ( n465 , n21881 );
buf ( n466 , n23721 );
buf ( n467 , n22818 );
buf ( n468 , n23724 );
buf ( n469 , n23728 );
buf ( n470 , n22843 );
buf ( n471 , n22870 );
buf ( n472 , n21044 );
buf ( n473 , n6496 );
buf ( n474 , n6531 );
buf ( n475 , n23733 );
buf ( n476 , n21907 );
buf ( n477 , n14623 );
buf ( n478 , n21943 );
buf ( n479 , n13729 );
buf ( n480 , n23468 );
buf ( n481 , n23738 );
buf ( n482 , n23807 );
buf ( n483 , n23473 );
buf ( n484 , n23829 );
buf ( n485 , n23484 );
buf ( n486 , n23743 );
buf ( n487 , n18537 );
buf ( n488 , n22898 );
buf ( n489 , n18254 );
buf ( n490 , n14090 );
buf ( n491 , n18285 );
buf ( n492 , n2354 );
buf ( n493 , n21970 );
buf ( n494 , n14247 );
buf ( n495 , n14650 );
buf ( n496 , n9119 );
buf ( n497 , n14689 );
buf ( n498 , n23792 );
buf ( n499 , n23503 );
buf ( n500 , n23479 );
buf ( n501 , n23748 );
buf ( n502 , n23834 );
buf ( n503 , n23839 );
buf ( n504 , n23513 );
buf ( n505 , n23498 );
buf ( n506 , n23844 );
buf ( n507 , n23518 );
buf ( n508 , n23797 );
buf ( n509 , n23522 );
buf ( n510 , n23527 );
buf ( n511 , n23819 );
buf ( n512 , n23803 );
buf ( n513 , n23753 );
buf ( n514 , n23531 );
buf ( n515 , n23814 );
buf ( n516 , n23768 );
buf ( n517 , n23716 );
buf ( n518 , n19919 );
buf ( n519 , n22922 );
buf ( n520 , n22944 );
buf ( n521 , n22984 );
buf ( n522 , n19104 );
buf ( n523 , n19464 );
buf ( n524 , n22097 );
buf ( n525 , n22222 );
buf ( n526 , n23011 );
buf ( n527 , n19781 );
buf ( n528 , n22247 );
buf ( n529 , n23786 );
buf ( n530 , n8260 );
buf ( n531 , n23407 );
buf ( n532 , n14725 );
buf ( n533 , n23039 );
buf ( n534 , n22279 );
buf ( n535 , n23066 );
buf ( n536 , n19946 );
buf ( n537 , n15033 );
buf ( n538 , n23422 );
buf ( n539 , n22737 );
buf ( n540 , n23088 );
buf ( n541 , n15748 );
buf ( n542 , n20203 );
buf ( n543 , n22310 );
buf ( n544 , n23113 );
buf ( n545 , n16255 );
buf ( n546 , n20233 );
buf ( n547 , n23148 );
buf ( n548 , n23180 );
buf ( n549 , n20270 );
buf ( n550 , n4026 );
buf ( n551 , n22331 );
buf ( n552 , n20307 );
buf ( n553 , n9078 );
buf ( n554 , n22352 );
buf ( n555 , n23208 );
buf ( n556 , n20446 );
buf ( n557 , n22388 );
buf ( n558 , n23238 );
buf ( n559 , n20461 );
buf ( n560 , n22419 );
buf ( n561 , n16299 );
buf ( n562 , n20595 );
buf ( n563 , n13094 );
buf ( n564 , n22711 );
buf ( n565 , n20634 );
buf ( n566 , n23257 );
buf ( n567 , n22445 );
buf ( n568 , n23435 );
buf ( n569 , n17452 );
buf ( n570 , n17884 );
buf ( n571 , n23276 );
buf ( n572 , n20676 );
buf ( n573 , n18023 );
buf ( n574 , n22468 );
buf ( n575 , n20803 );
buf ( n576 , n17013 );
buf ( n577 , n20840 );
buf ( n578 , n20884 );
buf ( n579 , n17169 );
buf ( n580 , n9800 );
buf ( n581 , n22507 );
buf ( n582 , n18043 );
buf ( n583 , n20907 );
buf ( n584 , n22531 );
buf ( n585 , n17666 );
buf ( n586 , n17705 );
buf ( n587 , n20928 );
buf ( n588 , n10951 );
buf ( n589 , n16747 );
buf ( n590 , n12691 );
buf ( n591 , n18079 );
buf ( n592 , n23300 );
buf ( n593 , n24006 );
buf ( n594 , n23331 );
buf ( n595 , n23463 );
buf ( n596 , n22593 );
buf ( n597 , n22667 );
buf ( n598 , n22560 );
buf ( n599 , n11225 );
buf ( n600 , n22633 );
buf ( n601 , n20943 );
buf ( n602 , n23360 );
buf ( n603 , n18109 );
buf ( n604 , n20976 );
buf ( n605 , n12035 );
buf ( n606 , n22682 );
buf ( n607 , n18145 );
buf ( n608 , n18184 );
buf ( n609 , n23379 );
buf ( n610 , n21008 );
buf ( n611 , n12176 );
buf ( n612 , n12317 );
buf ( n613 , n5681 );
buf ( n614 , n18203 );
buf ( n615 , n10671 );
buf ( n616 , n106 );
buf ( n617 , n392 );
buf ( n618 , n24026 );
buf ( n619 , n392 );
buf ( n620 , n23866 );
buf ( n621 , n392 );
buf ( n622 , n24058 );
buf ( n623 , n392 );
buf ( n624 , n23922 );
buf ( n625 , n392 );
buf ( n626 , n23938 );
buf ( n627 , n392 );
buf ( n628 , n23942 );
buf ( n629 , n392 );
buf ( n630 , n23934 );
buf ( n631 , n392 );
buf ( n632 , n23990 );
buf ( n633 , n392 );
buf ( n634 , n24075 );
buf ( n635 , n392 );
buf ( n636 , n23926 );
buf ( n637 , n392 );
buf ( n638 , n23998 );
buf ( n639 , n392 );
buf ( n640 , n23862 );
buf ( n641 , n392 );
buf ( n642 , n23930 );
buf ( n643 , n392 );
buf ( n644 , n23886 );
buf ( n645 , n392 );
buf ( n646 , n23894 );
buf ( n647 , n392 );
buf ( n648 , n24010 );
buf ( n649 , n392 );
buf ( n650 , n24018 );
buf ( n651 , n392 );
buf ( n652 , n24014 );
buf ( n653 , n392 );
buf ( n654 , n24022 );
buf ( n655 , n392 );
buf ( n656 , n23950 );
buf ( n657 , n392 );
buf ( n658 , n23870 );
buf ( n659 , n392 );
buf ( n660 , n23962 );
buf ( n661 , n392 );
buf ( n662 , n23910 );
buf ( n663 , n392 );
buf ( n664 , n23914 );
buf ( n665 , n392 );
buf ( n666 , n24042 );
buf ( n667 , n392 );
buf ( n668 , n23902 );
buf ( n669 , n392 );
buf ( n670 , n24002 );
buf ( n671 , n392 );
buf ( n672 , n24050 );
buf ( n673 , n392 );
buf ( n674 , n24066 );
buf ( n675 , n392 );
buf ( n676 , n24062 );
buf ( n677 , n392 );
buf ( n678 , n23854 );
buf ( n679 , n392 );
buf ( n680 , n23954 );
buf ( n681 , n392 );
buf ( n682 , n23982 );
buf ( n683 , n392 );
buf ( n684 , n23978 );
buf ( n685 , n392 );
buf ( n686 , n23946 );
buf ( n687 , n392 );
buf ( n688 , n23858 );
buf ( n689 , n392 );
buf ( n690 , n23898 );
buf ( n691 , n392 );
buf ( n692 , n24054 );
buf ( n693 , n392 );
buf ( n694 , n23874 );
buf ( n695 , n392 );
buf ( n696 , n23958 );
buf ( n697 , n392 );
buf ( n698 , n24034 );
buf ( n699 , n392 );
buf ( n700 , n23849 );
buf ( n701 , n392 );
buf ( n702 , n23966 );
buf ( n703 , n392 );
buf ( n704 , n23994 );
buf ( n705 , n392 );
buf ( n706 , n23970 );
buf ( n707 , n392 );
buf ( n708 , n24046 );
buf ( n709 , n392 );
buf ( n710 , n23847 );
buf ( n711 , n392 );
buf ( n712 , n23882 );
buf ( n713 , n392 );
buf ( n714 , n24030 );
buf ( n715 , n392 );
buf ( n716 , n23986 );
buf ( n717 , n392 );
buf ( n718 , n23974 );
buf ( n719 , n392 );
buf ( n720 , n23890 );
buf ( n721 , n392 );
buf ( n722 , n23906 );
buf ( n723 , n392 );
buf ( n724 , n23918 );
buf ( n725 , n392 );
buf ( n726 , n24070 );
buf ( n727 , n392 );
buf ( n728 , n24038 );
buf ( n729 , n392 );
buf ( n730 , n24074 );
buf ( n731 , n392 );
buf ( n732 , n23878 );
not ( n735 , n1 );
and ( n736 , n89 , n79 );
not ( n737 , n89 );
not ( n738 , n79 );
and ( n739 , n737 , n738 );
nor ( n740 , n736 , n739 );
not ( n741 , n740 );
or ( n742 , n735 , n741 );
nor ( n743 , n13 , n16 );
buf ( n744 , n743 );
nor ( n745 , n14 , n15 );
not ( n746 , n745 );
not ( n747 , n746 );
nand ( n748 , n747 , n12 );
not ( n749 , n12 );
not ( n750 , n11 );
nand ( n751 , n750 , n14 );
not ( n752 , n751 );
and ( n753 , n749 , n752 );
not ( n754 , n753 );
not ( n755 , n11 );
nor ( n756 , n755 , n14 );
nand ( n757 , n15 , n756 );
not ( n758 , n757 );
not ( n759 , n12 );
nand ( n760 , n758 , n759 );
nand ( n761 , n748 , n754 , n760 );
and ( n762 , n744 , n761 );
nand ( n763 , n14 , n15 );
not ( n764 , n763 );
not ( n765 , n764 );
not ( n766 , n12 );
nand ( n767 , n766 , n13 );
or ( n768 , n765 , n767 );
nand ( n769 , n11 , n14 );
nor ( n770 , n15 , n769 );
nand ( n771 , n13 , n770 );
nand ( n772 , n768 , n771 );
and ( n773 , n16 , n772 );
nor ( n774 , n762 , n773 );
not ( n775 , n12 );
not ( n776 , n757 );
not ( n777 , n776 );
nor ( n778 , n775 , n777 );
nand ( n779 , n16 , n778 );
not ( n780 , n16 );
nand ( n781 , n13 , n780 );
not ( n782 , n781 );
not ( n783 , n15 );
not ( n784 , n11 );
nor ( n785 , n784 , n14 );
nand ( n786 , n783 , n785 );
not ( n787 , n786 );
not ( n788 , n12 );
nand ( n789 , n787 , n788 );
not ( n790 , n789 );
nand ( n791 , n782 , n790 );
and ( n792 , n774 , n779 , n791 );
not ( n793 , n17 );
nor ( n794 , n792 , n793 );
nand ( n795 , n12 , n13 );
not ( n796 , n795 );
not ( n797 , n751 );
not ( n798 , n15 );
nand ( n799 , n797 , n798 );
not ( n800 , n799 );
not ( n801 , n800 );
not ( n802 , n801 );
nand ( n803 , n796 , n802 );
not ( n804 , n786 );
nand ( n805 , n804 , n796 );
not ( n806 , n805 );
nand ( n807 , n16 , n806 );
and ( n808 , n803 , n807 );
nand ( n809 , n13 , n16 );
not ( n810 , n809 );
nand ( n811 , n11 , n14 );
not ( n812 , n811 );
and ( n813 , n798 , n812 );
not ( n814 , n813 );
nor ( n815 , n814 , n12 );
not ( n816 , n815 );
not ( n817 , n816 );
nand ( n818 , n810 , n817 );
nor ( n819 , n769 , n12 );
nand ( n820 , n13 , n819 );
not ( n821 , n820 );
not ( n822 , n16 );
nand ( n823 , n821 , n793 , n822 );
not ( n824 , n16 );
not ( n825 , n13 );
not ( n826 , n12 );
and ( n827 , n755 , n745 );
not ( n828 , n827 );
nor ( n829 , n826 , n828 );
nand ( n830 , n825 , n829 );
or ( n831 , n824 , n830 );
not ( n832 , n16 );
nor ( n833 , n832 , n13 );
nor ( n834 , n12 , n15 );
and ( n835 , n752 , n834 );
nand ( n836 , n833 , n835 );
nand ( n837 , n831 , n836 );
nand ( n838 , n793 , n837 );
nand ( n839 , n808 , n818 , n823 , n838 );
nor ( n840 , n794 , n839 );
not ( n841 , n10 );
not ( n842 , n760 );
not ( n843 , n786 );
nand ( n844 , n843 , n13 );
nor ( n845 , n12 , n13 );
buf ( n846 , n845 );
not ( n847 , n811 );
nand ( n848 , n15 , n847 );
not ( n849 , n848 );
nand ( n850 , n846 , n849 );
not ( n851 , n848 );
nand ( n852 , n12 , n851 );
not ( n853 , n852 );
nand ( n854 , n13 , n853 );
and ( n855 , n755 , n834 );
not ( n856 , n855 );
not ( n857 , n13 );
nand ( n858 , n857 , n12 );
not ( n859 , n858 );
not ( n860 , n751 );
nand ( n861 , n860 , n15 );
not ( n862 , n861 );
nand ( n863 , n859 , n862 );
not ( n864 , n829 );
nor ( n865 , n11 , n14 );
buf ( n866 , n865 );
and ( n867 , n16 , n12 , n866 );
nand ( n868 , n11 , n15 );
nand ( n869 , n769 , n868 );
and ( n870 , n833 , n869 );
nor ( n871 , n867 , n870 );
and ( n872 , n864 , n871 );
not ( n873 , n13 );
not ( n874 , n12 );
not ( n875 , n15 );
nand ( n876 , n875 , n11 );
not ( n877 , n876 );
nand ( n878 , n874 , n877 );
not ( n879 , n878 );
nand ( n880 , n873 , n879 );
nand ( n881 , n782 , n778 );
nand ( n882 , n872 , n880 , n881 );
nand ( n883 , n793 , n882 );
not ( n884 , n835 );
or ( n885 , n13 , n884 );
or ( n886 , n809 , n856 );
nand ( n887 , n885 , n886 );
not ( n888 , n16 );
not ( n889 , n888 );
and ( n890 , n12 , n752 );
not ( n891 , n890 );
not ( n892 , n13 );
nor ( n893 , n891 , n892 );
nor ( n894 , n852 , n13 );
nor ( n895 , n893 , n894 );
not ( n896 , n895 );
not ( n897 , n896 );
or ( n898 , n889 , n897 );
not ( n899 , n16 );
not ( n900 , n848 );
not ( n901 , n12 );
nand ( n902 , n900 , n901 );
or ( n903 , n899 , n902 );
nand ( n904 , n898 , n903 );
nor ( n905 , n887 , n904 );
nand ( n906 , t_1 , n883 , n905 );
and ( n907 , n841 , n906 );
not ( n908 , n841 );
not ( n909 , n12 );
not ( n910 , n800 );
and ( n911 , n910 , n786 );
or ( n912 , n909 , n911 );
not ( n913 , n12 );
buf ( n914 , n785 );
nand ( n915 , n13 , n914 );
nor ( n916 , n913 , n915 );
not ( n917 , n916 );
nand ( n918 , n912 , n917 );
nand ( n919 , n16 , n918 );
not ( n920 , n16 );
nand ( n921 , n13 , n849 );
not ( n922 , n757 );
nand ( n923 , n922 , n12 );
not ( n924 , n923 );
not ( n925 , n13 );
nand ( n926 , n924 , n925 );
nand ( n927 , n880 , n921 , n926 );
nand ( n928 , n920 , n927 );
not ( n929 , n767 );
nand ( n930 , n929 , n862 );
nand ( n931 , n16 , n862 );
nand ( n932 , n764 , n845 );
nand ( n933 , n931 , n932 );
not ( n934 , n933 );
buf ( n935 , n786 );
nor ( n936 , n809 , n935 );
not ( n937 , n13 );
not ( n938 , n12 );
nand ( n939 , n938 , n866 );
not ( n940 , n939 );
nand ( n941 , n937 , n940 );
nand ( n942 , n743 , n813 );
nand ( n943 , n941 , n942 );
nor ( n944 , n936 , n943 );
not ( n945 , n11 );
nand ( n946 , n945 , n15 );
nor ( n947 , n12 , n946 );
nand ( n948 , n16 , n947 );
nor ( n949 , n781 , n801 );
nor ( n950 , n806 , n949 );
nand ( n951 , n934 , n944 , n948 , n950 );
and ( n952 , n793 , n951 );
not ( n953 , n793 );
not ( n954 , n16 );
not ( n955 , n13 );
not ( n956 , n14 );
nand ( n957 , n956 , n15 );
not ( n958 , n957 );
nand ( n959 , n955 , n958 );
not ( n960 , n776 );
nand ( n961 , n12 , n877 );
nand ( n962 , n959 , n960 , n961 );
not ( n963 , n962 );
or ( n964 , n954 , n963 );
nand ( n965 , n964 , n771 );
not ( n966 , n965 );
not ( n967 , n13 );
not ( n968 , n12 );
nor ( n969 , n968 , n868 );
nand ( n970 , n967 , n969 );
not ( n971 , n970 );
nor ( n972 , n971 , n778 );
not ( n973 , n13 );
nand ( n974 , n973 , n752 );
nor ( n975 , n16 , n974 );
not ( n976 , n16 );
buf ( n977 , n827 );
and ( n978 , n976 , n977 );
nor ( n979 , n975 , n978 );
nand ( n980 , n966 , n972 , n979 );
and ( n981 , n953 , n980 );
nor ( n982 , n952 , n981 );
nand ( n983 , n919 , n928 , n930 , n982 );
and ( n984 , n908 , n983 );
nor ( n985 , n907 , n984 );
nand ( n986 , n840 , n985 );
not ( n987 , n986 );
and ( n988 , n987 , n738 );
not ( n989 , n987 );
and ( n990 , n989 , n79 );
nor ( n991 , n988 , n990 );
not ( n992 , n8 );
not ( n993 , n992 );
nor ( n994 , n3 , n4 );
nor ( n995 , n2 , n5 );
and ( n996 , n994 , n995 );
not ( n997 , n996 );
not ( n998 , n2 );
nand ( n999 , n998 , n6 );
nor ( n1000 , n4 , n999 );
not ( n1001 , n1000 );
not ( n1002 , n1001 );
nand ( n1003 , n1002 , n7 );
not ( n1004 , n5 );
nand ( n1005 , n1004 , n2 );
not ( n1006 , n1005 );
not ( n1007 , n6 );
nand ( n1008 , n1006 , n1007 );
not ( n1009 , n1008 );
nand ( n1010 , n1009 , n3 );
not ( n1011 , n1010 );
nand ( n1012 , n7 , n1011 );
and ( n1013 , n997 , n1003 , n1012 );
not ( n1014 , n5 );
nor ( n1015 , n1014 , n2 );
nand ( n1016 , n6 , n1015 );
not ( n1017 , n1016 );
nand ( n1018 , n7 , n1017 );
not ( n1019 , n3 );
nand ( n1020 , n2 , n5 );
not ( n1021 , n1020 );
not ( n1022 , n6 );
nand ( n1023 , n1021 , n1022 );
not ( n1024 , n1023 );
nand ( n1025 , n1019 , n1024 );
not ( n1026 , n1025 );
not ( n1027 , n6 );
nand ( n1028 , n1027 , n1015 );
not ( n1029 , n1028 );
nand ( n1030 , n1029 , n3 );
not ( n1031 , n1030 );
or ( n1032 , n1026 , n1031 );
not ( n1033 , n7 );
nand ( n1034 , n1032 , n1033 );
nand ( n1035 , n1018 , n1034 );
not ( n1036 , n1035 );
nand ( n1037 , n5 , n6 );
not ( n1038 , n1037 );
nor ( n1039 , n3 , n4 );
nand ( n1040 , n1038 , n1039 );
not ( n1041 , n1008 );
nand ( n1042 , n1041 , n4 );
not ( n1043 , n1042 );
nand ( n1044 , n1043 , n3 );
nand ( n1045 , n1013 , n1036 , n1040 , n1044 );
not ( n1046 , n1045 );
or ( n1047 , n993 , n1046 );
not ( n1048 , n4 );
nand ( n1049 , n1048 , n3 );
not ( n1050 , n1049 );
not ( n1051 , n1016 );
nand ( n1052 , n1050 , n1051 );
nand ( n1053 , n1047 , n1052 );
not ( n1054 , n1053 );
not ( n1055 , n4 );
not ( n1056 , n1028 );
not ( n1057 , n1056 );
not ( n1058 , n1008 );
not ( n1059 , n1058 );
nand ( n1060 , n1057 , n1059 );
not ( n1061 , n1060 );
or ( n1062 , n1055 , n1061 );
not ( n1063 , n1005 );
nand ( n1064 , n3 , n1063 );
not ( n1065 , n1064 );
nand ( n1066 , n1065 , n4 );
nand ( n1067 , n1062 , n1066 );
nand ( n1068 , n7 , n1067 );
not ( n1069 , n7 );
not ( n1070 , n3 );
not ( n1071 , n6 );
nand ( n1072 , n1071 , n2 );
nor ( n1073 , n4 , n1072 );
nand ( n1074 , n1070 , n1073 );
nand ( n1075 , n2 , n5 );
not ( n1076 , n1075 );
nand ( n1077 , n1076 , n6 );
not ( n1078 , n1077 );
nand ( n1079 , n3 , n1078 );
not ( n1080 , n1005 );
nand ( n1081 , n1080 , n6 );
not ( n1082 , n1081 );
nand ( n1083 , n1082 , n4 );
not ( n1084 , n1083 );
not ( n1085 , n3 );
nand ( n1086 , n1084 , n1085 );
nand ( n1087 , n1074 , n1079 , n1086 );
nand ( n1088 , n1069 , n1087 );
not ( n1089 , n7 );
not ( n1090 , n5 );
nand ( n1091 , n1090 , n6 );
not ( n1092 , n1091 );
not ( n1093 , n3 );
nand ( n1094 , n1092 , n1093 );
not ( n1095 , n1081 );
not ( n1096 , n1095 );
not ( n1097 , n1072 );
nand ( n1098 , n4 , n1097 );
nand ( n1099 , n1094 , n1096 , n1098 );
not ( n1100 , n1099 );
or ( n1101 , n1089 , n1100 );
not ( n1102 , n1024 );
not ( n1103 , n3 );
nor ( n1104 , n1102 , n1103 );
not ( n1105 , n1104 );
nand ( n1106 , n1101 , n1105 );
not ( n1107 , n7 );
not ( n1108 , n5 );
nor ( n1109 , n1108 , n2 );
not ( n1110 , n1109 );
nor ( n1111 , n3 , n1110 );
nand ( n1112 , n1107 , n1111 );
not ( n1113 , n7 );
not ( n1114 , n2 );
nor ( n1115 , n5 , n6 );
nand ( n1116 , n1113 , n1114 , n1115 );
and ( n1117 , n1112 , n1116 );
not ( n1118 , n3 );
not ( n1119 , n4 );
nand ( n1120 , n2 , n6 );
nor ( n1121 , n1119 , n1120 );
nand ( n1122 , n1118 , n1121 );
not ( n1123 , n1122 );
not ( n1124 , n1123 );
not ( n1125 , n1083 );
not ( n1126 , n1125 );
nand ( n1127 , n1117 , n1124 , n1126 );
or ( n1128 , n1106 , n1127 );
nand ( n1129 , n1128 , n8 );
nand ( n1130 , n1068 , n1088 , n1129 );
not ( n1131 , n1130 );
and ( n1132 , n1054 , n1131 );
not ( n1133 , n9 );
nor ( n1134 , n1132 , n1133 );
not ( n1135 , n1134 );
not ( n1136 , n4 );
nand ( n1137 , n1136 , n1056 );
buf ( n1138 , n1137 );
nor ( n1139 , n3 , n1138 );
not ( n1140 , n1139 );
not ( n1141 , n1077 );
nand ( n1142 , n1141 , n1136 );
not ( n1143 , n1142 );
nand ( n1144 , n7 , n1143 );
not ( n1145 , n6 );
nor ( n1146 , n2 , n5 );
nand ( n1147 , n1145 , n1146 );
not ( n1148 , n1147 );
nand ( n1149 , n4 , n1148 );
not ( n1150 , n1149 );
not ( n1151 , n7 );
and ( n1152 , n4 , n995 );
not ( n1153 , n1152 );
or ( n1154 , n1151 , n1153 );
not ( n1155 , n1075 );
not ( n1156 , n1120 );
or ( n1157 , n1155 , n1156 );
not ( n1158 , n7 );
nor ( n1159 , n1158 , n3 );
nand ( n1160 , n1157 , n1159 );
nand ( n1161 , n1154 , n1160 );
nor ( n1162 , n1150 , n1161 );
not ( n1163 , n3 );
nor ( n1164 , n1163 , n7 );
nand ( n1165 , n1164 , n1125 );
nand ( n1166 , n1162 , n1074 , n1165 );
nand ( n1167 , n992 , n1166 );
nand ( n1168 , n1140 , n1144 , n1167 );
nand ( n1169 , n3 , n7 );
not ( n1170 , n1169 );
not ( n1171 , n4 );
nor ( n1172 , n2 , n6 );
nand ( n1173 , n1171 , n1172 );
not ( n1174 , n1173 );
nand ( n1175 , n1170 , n1174 );
and ( n1176 , n4 , n1109 );
not ( n1177 , n1176 );
not ( n1178 , n1177 );
nand ( n1179 , n1178 , n3 );
not ( n1180 , n1179 );
nand ( n1181 , n1078 , n4 );
nor ( n1182 , n3 , n1181 );
not ( n1183 , n1182 );
not ( n1184 , n1183 );
or ( n1185 , n1180 , n1184 );
not ( n1186 , n7 );
nand ( n1187 , n1185 , n1186 );
not ( n1188 , n7 );
not ( n1189 , n1188 );
not ( n1190 , n1095 );
nor ( n1191 , n1190 , n4 );
not ( n1192 , n1191 );
or ( n1193 , n1189 , n1192 );
not ( n1194 , n1010 );
not ( n1195 , n3 );
nor ( n1196 , n1181 , n1195 );
nor ( n1197 , n1194 , n1196 );
nand ( n1198 , n1193 , n1197 );
not ( n1199 , n1142 );
not ( n1200 , n3 );
nand ( n1201 , n1199 , n1200 );
not ( n1202 , n1173 );
not ( n1203 , n3 );
nor ( n1204 , n1016 , n1136 );
nand ( n1205 , n1203 , n1204 );
not ( n1206 , n1205 );
or ( n1207 , n1202 , n1206 );
nand ( n1208 , n1207 , n7 );
nand ( n1209 , n1201 , n1208 );
or ( n1210 , n1198 , n1209 );
nand ( n1211 , n1210 , n8 );
nand ( n1212 , n1175 , n1187 , n1211 );
nor ( n1213 , n1168 , n1212 );
or ( n1214 , n9 , n1213 );
not ( n1215 , n1125 );
not ( n1216 , n1215 );
nand ( n1217 , n7 , n1216 );
not ( n1218 , n1008 );
not ( n1219 , n1218 );
nor ( n1220 , n1219 , n4 );
not ( n1221 , n1220 );
not ( n1222 , n1221 );
nand ( n1223 , n1164 , n1222 );
and ( n1224 , n1217 , n1223 );
not ( n1225 , n1050 );
or ( n1226 , n1037 , n1225 );
nand ( n1227 , n1226 , n1105 );
nand ( n1228 , n7 , n1227 );
nor ( n1229 , n3 , n7 );
nor ( n1230 , n4 , n1110 );
not ( n1231 , n1230 );
nor ( n1232 , n5 , n6 );
nand ( n1233 , n4 , n1232 );
buf ( n1234 , n1233 );
not ( n1235 , n1234 );
not ( n1236 , n1235 );
not ( n1237 , n1191 );
nand ( n1238 , n1231 , n1236 , n1237 );
nand ( n1239 , n1229 , n1238 );
nand ( n1240 , n1224 , n1228 , n1239 );
nand ( n1241 , n1240 , n8 );
nand ( n1242 , n1214 , n1241 );
not ( n1243 , n1242 );
nor ( n1244 , n7 , n8 );
nor ( n1245 , n4 , n1075 );
not ( n1246 , n1245 );
not ( n1247 , n3 );
nor ( n1248 , n1246 , n1247 );
nand ( n1249 , n1244 , n1248 );
not ( n1250 , n3 );
not ( n1251 , n1028 );
nand ( n1252 , n1251 , n4 );
nor ( n1253 , n1250 , n1252 );
not ( n1254 , n1253 );
not ( n1255 , n1044 );
nand ( n1256 , n7 , n1255 );
nand ( n1257 , n1254 , n1256 );
not ( n1258 , n992 );
not ( n1259 , n7 );
not ( n1260 , n1149 );
not ( n1261 , n3 );
nand ( n1262 , n1260 , n1261 );
or ( n1263 , n1259 , n1262 );
not ( n1264 , n1138 );
nand ( n1265 , n1159 , n1264 );
nand ( n1266 , n1263 , n1265 );
not ( n1267 , n1266 );
or ( n1268 , n1258 , n1267 );
not ( n1269 , n1023 );
nand ( n1270 , n1269 , n1136 );
not ( n1271 , n1270 );
nand ( n1272 , n1170 , n1271 );
nand ( n1273 , n1268 , n1272 );
nor ( n1274 , n1257 , n1273 );
nand ( n1275 , n1135 , n1243 , n1249 , n1274 );
not ( n1276 , n1275 );
buf ( n1277 , n1039 );
nand ( n1278 , n1277 , n1051 );
not ( n1279 , n1278 );
nand ( n1280 , n3 , n1150 );
not ( n1281 , n1280 );
or ( n1282 , n1279 , n1281 );
not ( n1283 , n7 );
nand ( n1284 , n1282 , n1283 );
and ( n1285 , n7 , n992 );
not ( n1286 , n3 );
not ( n1287 , n4 );
nor ( n1288 , n1287 , n1037 );
nand ( n1289 , n1286 , n1288 );
buf ( n1290 , n1148 );
nand ( n1291 , n3 , n1290 );
not ( n1292 , n1023 );
nand ( n1293 , n1292 , n4 );
not ( n1294 , n1293 );
nand ( n1295 , n3 , n1294 );
nand ( n1296 , n1289 , n1291 , n1295 );
nand ( n1297 , n1285 , n1296 );
nand ( n1298 , n3 , n1073 );
not ( n1299 , n1298 );
not ( n1300 , n7 );
nand ( n1301 , n1299 , n1300 );
not ( n1302 , n3 );
nand ( n1303 , n1302 , n1078 );
not ( n1304 , n1303 );
not ( n1305 , n3 );
nand ( n1306 , n1305 , n1000 );
not ( n1307 , n1306 );
or ( n1308 , n1304 , n1307 );
not ( n1309 , n7 );
nand ( n1310 , n1308 , n1309 );
nand ( n1311 , n1301 , n1124 , n1310 );
nand ( n1312 , n992 , n1311 );
nand ( n1313 , n1284 , n1297 , n1312 );
not ( n1314 , n1313 );
not ( n1315 , n3 );
nand ( n1316 , n6 , n1146 );
not ( n1317 , n1316 );
not ( n1318 , n1317 );
nor ( n1319 , n1315 , n1318 );
not ( n1320 , n1319 );
not ( n1321 , n1320 );
not ( n1322 , n4 );
nor ( n1323 , n1322 , n1091 );
not ( n1324 , n1323 );
not ( n1325 , n1324 );
nand ( n1326 , n1142 , n1137 );
not ( n1327 , n1326 );
not ( n1328 , n1327 );
or ( n1329 , n1325 , n1328 );
nand ( n1330 , n1329 , n3 );
not ( n1331 , n1330 );
or ( n1332 , n1321 , n1331 );
not ( n1333 , n7 );
nand ( n1334 , n1332 , n1333 );
not ( n1335 , n1334 );
not ( n1336 , n3 );
not ( n1337 , n1336 );
not ( n1338 , n1245 );
nand ( n1339 , n1136 , n1317 );
nand ( n1340 , n1338 , n1042 , n1339 );
not ( n1341 , n1340 );
or ( n1342 , n1337 , n1341 );
nand ( n1343 , n3 , n1017 );
and ( n1344 , n1343 , n1270 );
nand ( n1345 , n1342 , n1344 );
nand ( n1346 , n7 , n1345 );
not ( n1347 , n1346 );
or ( n1348 , n1335 , n1347 );
nand ( n1349 , n1348 , n8 );
nor ( n1350 , n2 , n4 );
and ( n1351 , n1350 , n1232 );
nand ( n1352 , n1170 , n1351 );
not ( n1353 , n7 );
not ( n1354 , n2 );
nor ( n1355 , n1354 , n4 );
nand ( n1356 , n1353 , n1355 );
not ( n1357 , n1356 );
nor ( n1358 , n4 , n1120 );
nand ( n1359 , n3 , n1358 );
not ( n1360 , n1359 );
or ( n1361 , n1357 , n1360 );
nand ( n1362 , n1361 , n992 );
and ( n1363 , n1352 , n1362 );
not ( n1364 , n1181 );
nand ( n1365 , n4 , n1317 );
not ( n1366 , n1365 );
or ( n1367 , n1364 , n1366 );
nand ( n1368 , n1367 , n1170 );
nand ( n1369 , n1363 , n1310 , n1368 );
not ( n1370 , n1369 );
not ( n1371 , n1150 );
not ( n1372 , n1371 );
not ( n1373 , n1204 );
not ( n1374 , n1373 );
nand ( n1375 , n3 , n1374 );
not ( n1376 , n1375 );
or ( n1377 , n1372 , n1376 );
not ( n1378 , n7 );
nand ( n1379 , n1377 , n1378 );
not ( n1380 , n1170 );
not ( n1381 , n1098 );
not ( n1382 , n1381 );
or ( n1383 , n1380 , n1382 );
nand ( n1384 , n7 , n1290 );
nand ( n1385 , n1383 , n1384 );
and ( n1386 , n992 , n1385 );
not ( n1387 , n992 );
not ( n1388 , n1024 );
not ( n1389 , n3 );
nand ( n1390 , n1389 , n4 );
not ( n1391 , n1390 );
not ( n1392 , n1391 );
nor ( n1393 , n1388 , n1392 );
not ( n1394 , n1393 );
not ( n1395 , n5 );
nor ( n1396 , n1395 , n6 );
nand ( n1397 , n4 , n1396 );
not ( n1398 , n1397 );
nand ( n1399 , n1159 , n1398 );
not ( n1400 , n3 );
nor ( n1401 , n1400 , n5 );
nand ( n1402 , n4 , n1401 );
not ( n1403 , n1402 );
not ( n1404 , n1030 );
or ( n1405 , n1403 , n1404 );
not ( n1406 , n7 );
nand ( n1407 , n1405 , n1406 );
not ( n1408 , n1096 );
nand ( n1409 , n1408 , n3 );
nand ( n1410 , n1394 , n1399 , n1407 , n1409 );
and ( n1411 , n1387 , n1410 );
nor ( n1412 , n1386 , n1411 );
nand ( n1413 , n1370 , n1379 , n1412 );
nand ( n1414 , n1133 , n1413 );
not ( n1415 , n3 );
nand ( n1416 , n1415 , n1176 );
not ( n1417 , n1416 );
not ( n1418 , n7 );
nand ( n1419 , n1417 , n1418 );
not ( n1420 , n1295 );
nand ( n1421 , n1229 , n1058 );
not ( n1422 , n1421 );
or ( n1423 , n1420 , n1422 );
nand ( n1424 , n1423 , n8 );
and ( n1425 , n7 , n8 );
not ( n1426 , n1108 );
not ( n1427 , n4 );
and ( n1428 , n1426 , n1427 );
not ( n1429 , n1110 );
and ( n1430 , n3 , n1429 );
nor ( n1431 , n1428 , n1430 );
not ( n1432 , n3 );
nand ( n1433 , n1432 , n995 );
nand ( n1434 , n1431 , n1234 , n1433 );
nand ( n1435 , n1425 , n1434 );
nand ( n1436 , n1419 , n1424 , n1435 );
not ( n1437 , n1436 );
not ( n1438 , n7 );
not ( n1439 , n3 );
nand ( n1440 , n1439 , n1245 );
not ( n1441 , n3 );
nand ( n1442 , n1441 , n1323 );
nand ( n1443 , n1440 , n1373 , n1442 );
not ( n1444 , n1443 );
or ( n1445 , n1438 , n1444 );
not ( n1446 , n6 );
nand ( n1447 , n1446 , n5 );
nor ( n1448 , n4 , n1447 );
nand ( n1449 , n1170 , n1448 );
nand ( n1450 , n1445 , n1449 );
not ( n1451 , n1450 );
not ( n1452 , n999 );
nand ( n1453 , n1452 , n1391 );
not ( n1454 , n7 );
or ( n1455 , n1454 , n1074 );
nor ( n1456 , n1091 , n4 );
nand ( n1457 , n3 , n1456 );
nand ( n1458 , n1455 , n1457 );
not ( n1459 , n1458 );
not ( n1460 , n7 );
not ( n1461 , n1288 );
nand ( n1462 , n1234 , n1461 , n1177 );
nand ( n1463 , n1460 , n1462 );
not ( n1464 , n7 );
nand ( n1465 , n1464 , n1051 );
and ( n1466 , n1416 , n1112 );
nand ( n1467 , n1459 , n1463 , n1465 , n1466 );
nand ( n1468 , n992 , n1467 );
nand ( n1469 , n1437 , n1451 , n1453 , n1468 );
nand ( n1470 , n9 , n1469 );
nand ( n1471 , n1314 , n1349 , n1414 , n1470 );
buf ( n1472 , n1471 );
not ( n1473 , n1472 );
and ( n1474 , n1276 , n1473 );
not ( n1475 , n1276 );
and ( n1476 , n1475 , n1472 );
nor ( n1477 , n1474 , n1476 );
and ( n1478 , n991 , n1477 );
not ( n1479 , n991 );
not ( n1480 , n1477 );
and ( n1481 , n1479 , n1480 );
nor ( n1482 , n1478 , n1481 );
not ( n1483 , n34 );
not ( n1484 , n33 );
not ( n1485 , n32 );
not ( n1486 , n31 );
not ( n1487 , n27 );
not ( n1488 , n29 );
nand ( n1489 , n1488 , n28 );
not ( n1490 , n1489 );
nand ( n1491 , n30 , n1490 );
not ( n1492 , n1491 );
nand ( n1493 , n1487 , n1492 );
nor ( n1494 , n1486 , n1493 );
nand ( n1495 , n1485 , n1494 );
not ( n1496 , n27 );
nor ( n1497 , n28 , n29 );
and ( n1498 , n1496 , n1497 );
and ( n1499 , n32 , n1498 );
not ( n1500 , n32 );
not ( n1501 , n28 );
not ( n1502 , n27 );
nor ( n1503 , n1502 , n31 );
not ( n1504 , n1503 );
or ( n1505 , n1501 , n1504 );
nor ( n1506 , n28 , n30 );
nand ( n1507 , n27 , n1506 );
nand ( n1508 , n1505 , n1507 );
and ( n1509 , n1500 , n1508 );
nor ( n1510 , n1499 , n1509 );
nand ( n1511 , n1495 , n1510 );
not ( n1512 , n1511 );
or ( n1513 , n1484 , n1512 );
nand ( n1514 , n31 , n32 );
not ( n1515 , n1514 );
nor ( n1516 , n28 , n29 );
nand ( n1517 , n30 , n1516 );
not ( n1518 , n1517 );
not ( n1519 , n1518 );
not ( n1520 , n27 );
nor ( n1521 , n1519 , n1520 );
not ( n1522 , n1521 );
nand ( n1523 , n28 , n29 );
not ( n1524 , n1523 );
nand ( n1525 , n1524 , n30 );
not ( n1526 , n1525 );
not ( n1527 , n1526 );
not ( n1528 , n30 );
buf ( n1529 , n1489 );
not ( n1530 , n1529 );
nand ( n1531 , n1528 , n1530 );
buf ( n1532 , n1531 );
not ( n1533 , n1532 );
nand ( n1534 , n1533 , n27 );
nand ( n1535 , n1522 , n1527 , n1534 );
nand ( n1536 , n1515 , n1535 );
nand ( n1537 , n1513 , n1536 );
not ( n1538 , n1537 );
nor ( n1539 , n27 , n31 );
not ( n1540 , n30 );
not ( n1541 , n28 );
nand ( n1542 , n1541 , n29 );
not ( n1543 , n1542 );
nand ( n1544 , n1540 , n1543 );
not ( n1545 , n1544 );
nand ( n1546 , n1539 , n1545 );
not ( n1547 , n1519 );
nand ( n1548 , n1539 , n1547 );
and ( n1549 , n1546 , n1548 );
not ( n1550 , n32 );
not ( n1551 , n1491 );
not ( n1552 , n31 );
nand ( n1553 , n1551 , n1552 );
or ( n1554 , n1550 , n1553 );
not ( n1555 , n1529 );
not ( n1556 , n1555 );
nor ( n1557 , n31 , n1556 );
not ( n1558 , n1557 );
and ( n1559 , n32 , n1558 );
not ( n1560 , n32 );
not ( n1561 , n31 );
nand ( n1562 , n1561 , n1498 );
and ( n1563 , n1560 , n1562 );
nor ( n1564 , n1559 , n1563 );
nand ( n1565 , n28 , n29 );
not ( n1566 , n1565 );
not ( n1567 , n1566 );
nor ( n1568 , n27 , n1567 );
nand ( n1569 , n31 , n1568 );
not ( n1570 , n31 );
not ( n1571 , n29 );
nand ( n1572 , n1571 , n30 );
nor ( n1573 , n27 , n1572 );
nand ( n1574 , n1570 , n1573 );
not ( n1575 , n31 );
nand ( n1576 , n1575 , n1547 );
nand ( n1577 , n1569 , n1574 , n1576 );
not ( n1578 , n1577 );
not ( n1579 , n32 );
nand ( n1580 , n1540 , n1566 );
not ( n1581 , n1580 );
nand ( n1582 , n1581 , n27 );
not ( n1583 , n1582 );
not ( n1584 , n1583 );
not ( n1585 , n1584 );
nand ( n1586 , n1579 , n1585 );
not ( n1587 , n1542 );
not ( n1588 , n1587 );
nor ( n1589 , n27 , n1588 );
nand ( n1590 , n32 , n1589 );
not ( n1591 , n1590 );
nand ( n1592 , n32 , n1492 );
not ( n1593 , n1592 );
nor ( n1594 , n1591 , n1593 );
nand ( n1595 , n1578 , n1586 , n1594 );
or ( n1596 , n1564 , n1595 );
not ( n1597 , n33 );
nand ( n1598 , n1596 , n1597 );
nand ( n1599 , n1538 , n1549 , n1554 , n1598 );
not ( n1600 , n1599 );
or ( n1601 , n1483 , n1600 );
not ( n1602 , n33 );
not ( n1603 , n1602 );
not ( n1604 , n1507 );
nand ( n1605 , n31 , n1604 );
nor ( n1606 , n27 , n1544 );
not ( n1607 , n1606 );
nor ( n1608 , n31 , n32 );
nand ( n1609 , n1608 , n1547 );
and ( n1610 , n1605 , n1607 , n1609 );
nor ( n1611 , n28 , n30 );
nand ( n1612 , n31 , n1611 );
not ( n1613 , n31 );
not ( n1614 , n27 );
nand ( n1615 , n29 , n30 );
nor ( n1616 , n1614 , n1615 );
nand ( n1617 , n1613 , n1616 );
not ( n1618 , n1617 );
not ( n1619 , n1618 );
not ( n1620 , n1525 );
not ( n1621 , n27 );
nand ( n1622 , n1620 , n1621 );
not ( n1623 , n1622 );
nand ( n1624 , n31 , n1623 );
nand ( n1625 , n1612 , n1619 , n1624 );
nand ( n1626 , n32 , n1625 );
not ( n1627 , n1491 );
nand ( n1628 , n27 , n31 );
not ( n1629 , n1628 );
nand ( n1630 , n1627 , n1629 );
not ( n1631 , n1630 );
not ( n1632 , n31 );
not ( n1633 , n1587 );
nor ( n1634 , n1632 , n1633 );
nand ( n1635 , n27 , n1634 );
not ( n1636 , n1635 );
not ( n1637 , n27 );
nand ( n1638 , n1637 , n1518 );
not ( n1639 , n1638 );
nor ( n1640 , n1636 , n1639 );
not ( n1641 , n1640 );
or ( n1642 , n1631 , n1641 );
not ( n1643 , n32 );
nand ( n1644 , n1642 , n1643 );
nand ( n1645 , n1610 , n1626 , n1644 );
not ( n1646 , n1645 );
or ( n1647 , n1603 , n1646 );
not ( n1648 , n1525 );
not ( n1649 , n1648 );
not ( n1650 , n27 );
nor ( n1651 , n1649 , n1650 );
not ( n1652 , n1651 );
not ( n1653 , n1652 );
nand ( n1654 , n31 , n1653 );
or ( n1655 , n32 , n1654 );
not ( n1656 , n1588 );
nand ( n1657 , n1656 , n1503 );
not ( n1658 , n1657 );
nor ( n1659 , n30 , n1523 );
not ( n1660 , n1659 );
nor ( n1661 , n1660 , n27 );
not ( n1662 , n1661 );
not ( n1663 , n1662 );
or ( n1664 , n1658 , n1663 );
not ( n1665 , n32 );
nand ( n1666 , n1664 , n1665 );
not ( n1667 , n31 );
nand ( n1668 , n1667 , n1659 );
buf ( n1669 , n1668 );
nand ( n1670 , n1655 , n1666 , n1669 );
nand ( n1671 , n33 , n1670 );
nand ( n1672 , n1647 , n1671 );
not ( n1673 , n34 );
not ( n1674 , n1673 );
not ( n1675 , n32 );
not ( n1676 , n31 );
nor ( n1677 , n1676 , n1638 );
nand ( n1678 , n1675 , n1677 );
not ( n1679 , n1678 );
nor ( n1680 , n1514 , n1584 );
nand ( n1681 , n29 , n30 );
nor ( n1682 , n28 , n1681 );
not ( n1683 , n1682 );
not ( n1684 , n27 );
nor ( n1685 , n1683 , n1684 );
buf ( n1686 , n1685 );
not ( n1687 , n1686 );
not ( n1688 , n1687 );
nor ( n1689 , n1679 , n1680 , n1688 );
not ( n1690 , n33 );
not ( n1691 , n32 );
nand ( n1692 , n1691 , n31 );
or ( n1693 , n1572 , n1692 );
nand ( n1694 , n1693 , n1617 );
nand ( n1695 , n1690 , n1694 );
not ( n1696 , n32 );
not ( n1697 , n30 );
nand ( n1698 , n1697 , n28 );
not ( n1699 , n1698 );
nand ( n1700 , n31 , n1699 );
not ( n1701 , n1567 );
nand ( n1702 , n31 , n1701 );
not ( n1703 , n27 );
nor ( n1704 , n29 , n30 );
and ( n1705 , n1703 , n1704 );
not ( n1706 , n1705 );
nand ( n1707 , n1700 , n1702 , n1706 );
nand ( n1708 , n1696 , n1707 );
nor ( n1709 , n28 , n1681 );
not ( n1710 , n1709 );
not ( n1711 , n1710 );
nand ( n1712 , n1711 , n31 );
not ( n1713 , n31 );
nand ( n1714 , n1713 , n1497 );
not ( n1715 , n1714 );
nor ( n1716 , n27 , n1529 );
nand ( n1717 , n31 , n1716 );
not ( n1718 , n1717 );
or ( n1719 , n1715 , n1718 );
nand ( n1720 , n1719 , n32 );
nand ( n1721 , n1708 , n1712 , n1720 );
nand ( n1722 , n33 , n1721 );
nand ( n1723 , n1689 , n1695 , n1722 );
not ( n1724 , n1723 );
or ( n1725 , n1674 , n1724 );
not ( n1726 , n32 );
nand ( n1727 , n31 , n1606 );
not ( n1728 , n1727 );
nand ( n1729 , n1726 , n1728 );
not ( n1730 , n29 );
nor ( n1731 , n1730 , n30 );
not ( n1732 , n1731 );
not ( n1733 , n1732 );
not ( n1734 , n1733 );
not ( n1735 , n1547 );
nand ( n1736 , n1734 , n1735 );
nand ( n1737 , n1736 , n32 , n1539 );
nand ( n1738 , n1729 , n1737 );
and ( n1739 , n32 , n33 );
not ( n1740 , n1739 );
not ( n1741 , n27 );
nand ( n1742 , n1741 , n29 );
or ( n1743 , n31 , n1742 );
nand ( n1744 , n1743 , n1584 );
not ( n1745 , n1744 );
or ( n1746 , n1740 , n1745 );
not ( n1747 , n1531 );
not ( n1748 , n27 );
nand ( n1749 , n1747 , n1748 );
not ( n1750 , n1749 );
and ( n1751 , n31 , n33 );
nand ( n1752 , n1750 , n32 , n1751 );
nand ( n1753 , n1746 , n1752 );
nor ( n1754 , n1738 , n1753 );
nand ( n1755 , n1725 , n1754 );
nor ( n1756 , n1672 , n1755 );
nand ( n1757 , n1601 , n1756 );
not ( n1758 , n1757 );
not ( n1759 , n20 );
nand ( n1760 , n1759 , n21 );
not ( n1761 , n1760 );
nand ( n1762 , n24 , n1761 );
not ( n1763 , n1762 );
nand ( n1764 , n1763 , n22 );
not ( n1765 , n1764 );
not ( n1766 , n1765 );
not ( n1767 , n25 );
and ( n1768 , n23 , n1767 );
not ( n1769 , n1768 );
nor ( n1770 , n1766 , n1769 );
nor ( n1771 , n20 , n21 );
not ( n1772 , n1771 );
not ( n1773 , n1772 );
nand ( n1774 , n22 , n1773 );
not ( n1775 , n1774 );
nand ( n1776 , n25 , n1775 );
not ( n1777 , n23 );
not ( n1778 , n24 );
nand ( n1779 , n1778 , n21 );
nor ( n1780 , n22 , n1779 );
nand ( n1781 , n1777 , n1780 );
and ( n1782 , n1776 , n1781 );
not ( n1783 , n24 );
nand ( n1784 , n1771 , n1783 );
not ( n1785 , n1784 );
nand ( n1786 , n22 , n1785 );
nand ( n1787 , n20 , n21 );
not ( n1788 , n1787 );
nand ( n1789 , n21 , n24 );
not ( n1790 , n1789 );
or ( n1791 , n1788 , n1790 );
not ( n1792 , n23 );
nand ( n1793 , n1792 , n25 );
not ( n1794 , n1793 );
nand ( n1795 , n1791 , n1794 );
nand ( n1796 , n1782 , n1786 , n1795 );
nor ( n1797 , n1770 , n1796 );
or ( n1798 , n26 , n1797 );
nand ( n1799 , n23 , n25 );
not ( n1800 , n1799 );
not ( n1801 , n22 );
nor ( n1802 , n21 , n24 );
nand ( n1803 , n1801 , n1802 );
not ( n1804 , n1803 );
nand ( n1805 , n1800 , n1804 );
not ( n1806 , n23 );
not ( n1807 , n21 );
nand ( n1808 , n1807 , n20 );
not ( n1809 , n1808 );
nand ( n1810 , n1783 , n1809 );
not ( n1811 , n1810 );
not ( n1812 , n22 );
nand ( n1813 , n1811 , n1812 );
not ( n1814 , n1813 );
nand ( n1815 , n1806 , n1814 );
nand ( n1816 , n1798 , n1805 , n1815 );
not ( n1817 , n1808 );
nand ( n1818 , n1817 , n24 );
not ( n1819 , n1818 );
nand ( n1820 , n1819 , n22 );
nand ( n1821 , n20 , n21 );
not ( n1822 , n1821 );
nand ( n1823 , n1822 , n24 );
not ( n1824 , n1823 );
nand ( n1825 , n1824 , n22 );
not ( n1826 , n1825 );
nand ( n1827 , n23 , n1826 );
not ( n1828 , n1762 );
and ( n1829 , n1828 , n1812 );
nand ( n1830 , n1783 , n1761 );
not ( n1831 , n1830 );
nand ( n1832 , n23 , n1831 );
not ( n1833 , n1832 );
not ( n1834 , n1833 );
not ( n1835 , n1823 );
nand ( n1836 , n1835 , n1812 );
not ( n1837 , n1836 );
not ( n1838 , n23 );
nand ( n1839 , n1837 , n1838 );
not ( n1840 , n26 );
or ( n1841 , t_0 , n1840 );
not ( n1842 , n23 );
nand ( n1843 , n22 , n1809 );
nor ( n1844 , n1842 , n1843 );
nor ( n1845 , n23 , n1825 );
nor ( n1846 , n1844 , n1845 );
or ( n1847 , n25 , n1846 );
not ( n1848 , n25 );
not ( n1849 , n1837 );
or ( n1850 , n1848 , n1849 );
nand ( n1851 , n1841 , n1847 , n1850 );
or ( n1852 , n1816 , n1851 );
not ( n1853 , n19 );
nand ( n1854 , n1852 , n1853 );
nor ( n1855 , n23 , n25 );
not ( n1856 , n1809 );
nor ( n1857 , n1856 , n22 );
not ( n1858 , n1857 );
nor ( n1859 , n20 , n24 );
nand ( n1860 , n22 , n1859 );
not ( n1861 , n1829 );
nand ( n1862 , n1858 , n1860 , n1861 );
nand ( n1863 , n1855 , n1862 );
not ( n1864 , n1764 );
nand ( n1865 , n25 , n1864 );
not ( n1866 , n1831 );
nor ( n1867 , n1866 , n22 );
nand ( n1868 , n23 , n1867 );
nor ( n1869 , n25 , n1868 );
not ( n1870 , n1869 );
nand ( n1871 , n1863 , n1865 , n1870 );
nand ( n1872 , n26 , n1871 );
not ( n1873 , n25 );
nor ( n1874 , n24 , n1821 );
nand ( n1875 , n1812 , n1874 );
not ( n1876 , n1875 );
nand ( n1877 , n23 , n1876 );
or ( n1878 , n1873 , n1877 );
nand ( n1879 , n1854 , n1872 , n1878 );
not ( n1880 , n19 );
not ( n1881 , n25 );
not ( n1882 , n23 );
not ( n1883 , n20 );
nand ( n1884 , n1883 , n24 );
not ( n1885 , n1884 );
nand ( n1886 , n1882 , n1885 );
not ( n1887 , n1828 );
not ( n1888 , n1779 );
nand ( n1889 , n22 , n1888 );
nand ( n1890 , n1886 , n1887 , n1889 );
not ( n1891 , n1890 );
or ( n1892 , n1881 , n1891 );
nor ( n1893 , n24 , n1787 );
nand ( n1894 , n23 , n1893 );
nand ( n1895 , n1892 , n1894 );
not ( n1896 , n1895 );
not ( n1897 , n23 );
not ( n1898 , n22 );
nor ( n1899 , n1898 , n1789 );
nand ( n1900 , n1897 , n1899 );
not ( n1901 , n1900 );
nor ( n1902 , n1901 , n1864 );
not ( n1903 , n23 );
nand ( n1904 , n1903 , n1809 );
nor ( n1905 , n25 , n1904 );
not ( n1906 , n1785 );
nor ( n1907 , n1906 , n25 );
nor ( n1908 , n1905 , n1907 );
nand ( n1909 , n1896 , n1902 , n1908 );
and ( n1910 , n26 , n1909 );
not ( n1911 , n26 );
not ( n1912 , n25 );
not ( n1913 , n1818 );
not ( n1914 , n1913 );
nor ( n1915 , n1912 , n1914 );
nand ( n1916 , n20 , n24 );
not ( n1917 , n23 );
nand ( n1918 , n1812 , n1917 );
nor ( n1919 , n1916 , n1918 );
not ( n1920 , n1772 );
nand ( n1921 , n1812 , n1920 );
nor ( n1922 , n23 , n1921 );
nor ( n1923 , n1915 , n1919 , n1922 );
not ( n1924 , n21 );
nand ( n1925 , n1924 , n24 );
nor ( n1926 , n22 , n1925 );
not ( n1927 , n1926 );
not ( n1928 , n1927 );
nand ( n1929 , n1928 , n25 );
not ( n1930 , n23 );
nand ( n1931 , n1930 , n1893 );
not ( n1932 , n1931 );
not ( n1933 , n1810 );
nand ( n1934 , n23 , n1933 );
not ( n1935 , n1934 );
or ( n1936 , n1932 , n1935 );
not ( n1937 , n25 );
nand ( n1938 , n1936 , n1937 );
nand ( n1939 , n22 , n23 );
not ( n1940 , n1939 );
nand ( n1941 , n1940 , n1831 );
not ( n1942 , n1941 );
not ( n1943 , n25 );
nor ( n1944 , n1943 , n1832 );
nor ( n1945 , n1942 , n1944 );
nand ( n1946 , n1923 , n1929 , n1938 , n1945 );
and ( n1947 , n1911 , n1946 );
nor ( n1948 , n1910 , n1947 );
not ( n1949 , n25 );
not ( n1950 , n1781 );
not ( n1951 , n1950 );
not ( n1952 , n1823 );
nand ( n1953 , n23 , n1952 );
not ( n1954 , n1764 );
not ( n1955 , n23 );
nand ( n1956 , n1954 , n1955 );
nand ( n1957 , n1951 , n1953 , n1956 );
nand ( n1958 , n1949 , n1957 );
not ( n1959 , n23 );
nor ( n1960 , n1959 , n22 );
not ( n1961 , n1914 );
nand ( n1962 , n1960 , n1961 );
not ( n1963 , n1831 );
and ( n1964 , n1963 , n1810 );
or ( n1965 , n1964 , n1812 );
not ( n1966 , n23 );
not ( n1967 , n1761 );
nor ( n1968 , n1966 , n1967 );
nand ( n1969 , n22 , n1968 );
nand ( n1970 , n1965 , n1969 );
nand ( n1971 , n25 , n1970 );
nand ( n1972 , n1948 , n1958 , n1962 , n1971 );
not ( n1973 , n1972 );
or ( n1974 , n1880 , n1973 );
nor ( n1975 , n25 , n26 );
not ( n1976 , n23 );
nor ( n1977 , n22 , n1787 );
not ( n1978 , n1977 );
or ( n1979 , n1976 , n1978 );
not ( n1980 , n1979 );
and ( n1981 , n1975 , n1980 );
and ( n1982 , n1940 , n1933 );
not ( n1983 , n1830 );
nand ( n1984 , n1983 , n22 );
nor ( n1985 , n1799 , n1984 );
nor ( n1986 , n1981 , n1982 , n1985 );
and ( n1987 , n25 , n26 );
not ( n1988 , n1960 );
or ( n1989 , n1916 , n1988 );
nand ( n1990 , n1989 , n1894 );
nand ( n1991 , n1987 , n1990 );
not ( n1992 , n26 );
not ( n1993 , n25 );
not ( n1994 , n1784 );
not ( n1995 , n23 );
nand ( n1996 , n1995 , n22 );
not ( n1997 , n1996 );
nand ( n1998 , n1994 , n1997 );
or ( n1999 , n1993 , n1998 );
nand ( n2000 , n1794 , n1814 );
nand ( n2001 , n1999 , n2000 );
nand ( n2002 , n1992 , n2001 );
and ( n2003 , n1986 , n1991 , n2002 );
nand ( n2004 , n1974 , n2003 );
nor ( n2005 , n1879 , n2004 );
not ( n2006 , n2005 );
not ( n2007 , n2006 );
and ( n2008 , n1758 , n2007 );
not ( n2009 , n1758 );
and ( n2010 , n2009 , n2006 );
nor ( n2011 , n2008 , n2010 );
not ( n2012 , n31 );
nand ( n2013 , n2012 , n1526 );
not ( n2014 , n2013 );
not ( n2015 , n1574 );
or ( n2016 , n2014 , n2015 );
not ( n2017 , n32 );
nand ( n2018 , n2016 , n2017 );
not ( n2019 , n1652 );
not ( n2020 , n1521 );
not ( n2021 , n2020 );
or ( n2022 , n2019 , n2021 );
nand ( n2023 , n2022 , n1515 );
not ( n2024 , n33 );
not ( n2025 , n1515 );
nand ( n2026 , n27 , n1731 );
not ( n2027 , n2026 );
not ( n2028 , n2027 );
or ( n2029 , n2025 , n2028 );
not ( n2030 , n1516 );
nor ( n2031 , n2030 , n30 );
not ( n2032 , n2031 );
not ( n2033 , n2032 );
nand ( n2034 , n32 , n2033 );
nand ( n2035 , n2029 , n2034 );
nand ( n2036 , n2024 , n2035 );
and ( n2037 , n2018 , n2023 , n2036 );
not ( n2038 , n27 );
and ( n2039 , n2038 , n2031 );
nand ( n2040 , n1515 , n2039 );
not ( n2041 , n2032 );
nand ( n2042 , n2041 , n27 );
not ( n2043 , n2042 );
not ( n2044 , n1630 );
or ( n2045 , n2043 , n2044 );
not ( n2046 , n32 );
nand ( n2047 , n2045 , n2046 );
and ( n2048 , n2040 , n2047 );
not ( n2049 , n33 );
not ( n2050 , n32 );
not ( n2051 , n2050 );
not ( n2052 , n1742 );
not ( n2053 , n2052 );
or ( n2054 , n2051 , n2053 );
nor ( n2055 , n27 , n1615 );
nand ( n2056 , n31 , n2055 );
nand ( n2057 , n2054 , n2056 );
nand ( n2058 , n2049 , n2057 );
not ( n2059 , n31 );
nand ( n2060 , n2059 , n1583 );
nand ( n2061 , n1712 , n2060 );
not ( n2062 , n32 );
not ( n2063 , n2062 );
not ( n2064 , n28 );
not ( n2065 , n2064 );
not ( n2066 , n1629 );
or ( n2067 , n2065 , n2066 );
not ( n2068 , n1531 );
nand ( n2069 , n2068 , n31 );
nand ( n2070 , n2067 , n2069 );
not ( n2071 , n2070 );
or ( n2072 , n2063 , n2071 );
not ( n2073 , n32 );
nor ( n2074 , n2073 , n31 );
not ( n2075 , n2074 );
not ( n2076 , n1698 );
nand ( n2077 , n2076 , n27 );
or ( n2078 , n2075 , n2077 );
nand ( n2079 , n2072 , n2078 );
or ( n2080 , n2061 , n2079 );
nand ( n2081 , n2080 , n33 );
nand ( n2082 , n2037 , n2048 , n2058 , n2081 );
and ( n2083 , n1673 , n2082 );
not ( n2084 , n1739 );
not ( n2085 , n2084 );
not ( n2086 , n32 );
not ( n2087 , n2086 );
nand ( n2088 , n1555 , n27 );
nand ( n2089 , n28 , n30 );
not ( n2090 , n2089 );
nand ( n2091 , n2090 , n27 );
nand ( n2092 , n2088 , n2091 , n1507 );
not ( n2093 , n2092 );
or ( n2094 , n2087 , n2093 );
not ( n2095 , n32 );
nand ( n2096 , n2095 , n1557 );
nand ( n2097 , n2094 , n2096 );
not ( n2098 , n27 );
not ( n2099 , n29 );
nor ( n2100 , n2099 , n30 );
nand ( n2101 , n2098 , n2100 );
nor ( n2102 , n31 , n2101 );
nand ( n2103 , n32 , n2102 );
not ( n2104 , n32 );
nand ( n2105 , n2104 , n1492 );
not ( n2106 , n28 );
nand ( n2107 , n2106 , n30 );
nor ( n2108 , n27 , n2107 );
nand ( n2109 , n31 , n2108 );
nand ( n2110 , n2103 , n2105 , n2109 );
nor ( n2111 , n2097 , n2110 );
or ( n2112 , n2111 , n33 );
not ( n2113 , n31 );
not ( n2114 , n2088 );
nand ( n2115 , n2113 , n2114 );
nand ( n2116 , n2112 , n2115 );
not ( n2117 , n2116 );
or ( n2118 , n2085 , n2117 );
not ( n2119 , n27 );
nand ( n2120 , n2119 , n28 );
nand ( n2121 , n31 , n1555 );
nand ( n2122 , n2120 , n2121 , n1507 , n1714 );
and ( n2123 , n2122 , n1739 );
not ( n2124 , n31 );
nand ( n2125 , n2124 , n27 );
nor ( n2126 , n1572 , n2125 );
nor ( n2127 , n2123 , n2126 );
not ( n2128 , n27 );
nand ( n2129 , n2128 , n1699 );
not ( n2130 , n2129 );
nand ( n2131 , n1515 , n2130 );
not ( n2132 , n1582 );
nand ( n2133 , n31 , n2132 );
not ( n2134 , n2133 );
nand ( n2135 , n1608 , n1545 );
not ( n2136 , n2135 );
or ( n2137 , n2134 , n2136 );
nand ( n2138 , n2137 , n33 );
not ( n2139 , n31 );
nand ( n2140 , n2139 , n1568 );
not ( n2141 , n1491 );
nand ( n2142 , n2141 , n27 );
not ( n2143 , n31 );
not ( n2144 , n27 );
nor ( n2145 , n2144 , n2107 );
nand ( n2146 , n2143 , n2145 );
nand ( n2147 , n2140 , n2142 , n2146 );
nand ( n2148 , n32 , n2147 );
and ( n2149 , n2127 , n2131 , n2138 , n2148 );
nand ( n2150 , n2118 , n2149 );
nand ( n2151 , n2150 , n34 );
not ( n2152 , n2151 );
nor ( n2153 , n2083 , n2152 );
not ( n2154 , n33 );
not ( n2155 , n1692 );
not ( n2156 , n2155 );
not ( n2157 , n2145 );
not ( n2158 , n1623 );
nand ( n2159 , n1735 , n2157 , n2158 , n1749 );
not ( n2160 , n2159 );
or ( n2161 , n2156 , n2160 );
not ( n2162 , n31 );
not ( n2163 , n2162 );
not ( n2164 , n1568 );
not ( n2165 , n1544 );
nand ( n2166 , n27 , n2165 );
nand ( n2167 , n2164 , n2166 , n1638 );
not ( n2168 , n2167 );
or ( n2169 , n2163 , n2168 );
not ( n2170 , n1491 );
nand ( n2171 , n2170 , n31 );
and ( n2172 , n2171 , n1662 );
nand ( n2173 , n2169 , n2172 );
nand ( n2174 , n32 , n2173 );
nand ( n2175 , n2161 , n2174 );
not ( n2176 , n2175 );
or ( n2177 , n2154 , n2176 );
not ( n2178 , n33 );
not ( n2179 , n32 );
not ( n2180 , n31 );
nor ( n2181 , n2180 , n2101 );
nand ( n2182 , n2179 , n2181 );
not ( n2183 , n1618 );
nand ( n2184 , n2182 , n2183 , n2018 );
nand ( n2185 , n2178 , n2184 );
nand ( n2186 , n2177 , n2185 );
not ( n2187 , n33 );
and ( n2188 , n32 , n2187 );
not ( n2189 , n2188 );
or ( n2190 , n31 , n2091 );
not ( n2191 , n2032 );
nand ( n2192 , n31 , n2191 );
nand ( n2193 , n2190 , n2192 , n2133 );
not ( n2194 , n2193 );
or ( n2195 , n2189 , n2194 );
not ( n2196 , n1493 );
not ( n2197 , n31 );
nand ( n2198 , n2196 , n2197 );
not ( n2199 , n2198 );
not ( n2200 , n2042 );
nand ( n2201 , n31 , n2200 );
not ( n2202 , n2201 );
or ( n2203 , n2199 , n2202 );
not ( n2204 , n32 );
nand ( n2205 , n2203 , n2204 );
nand ( n2206 , n2195 , n2205 );
nor ( n2207 , n2186 , n2206 );
nand ( n2208 , n2153 , n2207 );
buf ( n2209 , n2208 );
not ( n2210 , n2209 );
not ( n2211 , n2210 );
not ( n2212 , n992 );
nand ( n2213 , n3 , n1235 );
buf ( n2214 , n1317 );
nand ( n2215 , n1229 , n2214 );
and ( n2216 , n2213 , n1221 , n2215 );
not ( n2217 , n1115 );
not ( n2218 , n2217 );
nand ( n2219 , n3 , n2218 );
not ( n2220 , n1142 );
nand ( n2221 , n2220 , n3 );
nand ( n2222 , n2219 , n1124 , n2221 );
nand ( n2223 , n7 , n2222 );
not ( n2224 , n7 );
nand ( n2225 , n1339 , n1066 , n1375 );
nand ( n2226 , n2224 , n2225 );
nand ( n2227 , n2216 , n2223 , n2226 );
not ( n2228 , n2227 );
or ( n2229 , n2212 , n2228 );
not ( n2230 , n1355 );
or ( n2231 , n3 , n2230 );
nand ( n2232 , n2231 , n1293 );
nand ( n2233 , n1425 , n2232 );
nand ( n2234 , n2229 , n2233 );
not ( n2235 , n7 );
or ( n2236 , n1097 , n2214 );
nand ( n2237 , n2236 , n1277 );
or ( n2238 , n2235 , n2237 );
nand ( n2239 , n2238 , n1223 );
nor ( n2240 , n2234 , n2239 );
and ( n2241 , n7 , n1111 );
not ( n2242 , n7 );
and ( n2243 , n2242 , n996 );
nor ( n2244 , n2241 , n2243 );
nand ( n2245 , n1136 , n1063 );
not ( n2246 , n2245 );
nand ( n2247 , n7 , n2246 );
nand ( n2248 , n2244 , n1018 , n2247 );
not ( n2249 , n2248 );
not ( n2250 , n1306 );
nor ( n2251 , n2250 , n1248 );
nor ( n2252 , n7 , n1293 );
nor ( n2253 , n1318 , n3 );
nor ( n2254 , n2252 , n2253 );
nand ( n2255 , n2249 , n2251 , n2254 );
nand ( n2256 , n992 , n2255 );
not ( n2257 , n8 );
not ( n2258 , n7 );
not ( n2259 , n5 );
not ( n2260 , n1391 );
or ( n2261 , n2259 , n2260 );
nand ( n2262 , n2261 , n1233 );
nand ( n2263 , n2258 , n2262 );
not ( n2264 , n995 );
nor ( n2265 , n2264 , n4 );
nand ( n2266 , n7 , n2265 );
not ( n2267 , n7 );
not ( n2268 , n6 );
nor ( n2269 , n2268 , n1049 );
nand ( n2270 , n2267 , n1429 , n2269 );
nand ( n2271 , n2263 , n2266 , n2270 );
not ( n2272 , n2271 );
or ( n2273 , n2257 , n2272 );
nand ( n2274 , n1159 , n1017 );
nand ( n2275 , n2273 , n2274 );
not ( n2276 , n1058 );
not ( n2277 , n2276 );
nand ( n2278 , n2277 , n1277 );
nand ( n2279 , n1277 , n2214 );
nand ( n2280 , n2278 , n2279 );
nor ( n2281 , n2275 , n2280 );
not ( n2282 , n1252 );
not ( n2283 , n2282 );
nand ( n2284 , n1365 , n1077 , n2283 );
nand ( n2285 , n1170 , n2284 );
nand ( n2286 , n2256 , n2281 , n2285 );
nand ( n2287 , n9 , n2286 );
not ( n2288 , n2287 );
not ( n2289 , n3 );
nor ( n2290 , n2289 , n1138 );
and ( n2291 , n1425 , n2290 );
not ( n2292 , n8 );
not ( n2293 , n7 );
not ( n2294 , n1075 );
and ( n2295 , n3 , n2294 );
not ( n2296 , n2295 );
nand ( n2297 , n3 , n1396 );
nand ( n2298 , n2296 , n2297 , n1173 );
nand ( n2299 , n2293 , n2298 );
not ( n2300 , n1433 );
nand ( n2301 , n3 , n1230 );
not ( n2302 , n2301 );
or ( n2303 , n2300 , n2302 );
nand ( n2304 , n2303 , n7 );
nand ( n2305 , n2299 , n1409 , n2304 );
not ( n2306 , n2305 );
or ( n2307 , n2292 , n2306 );
not ( n2308 , n1452 );
not ( n2309 , n1164 );
or ( n2310 , n2308 , n2309 );
nand ( n2311 , n2310 , n1122 );
nand ( n2312 , n992 , n2311 );
nand ( n2313 , n2307 , n2312 );
nand ( n2314 , n1170 , n1294 );
not ( n2315 , n7 );
not ( n2316 , n3 );
nor ( n2317 , n2316 , n1339 );
nand ( n2318 , n2315 , n2317 );
nand ( n2319 , n2314 , n1126 , n2318 );
nor ( n2320 , n2313 , n2319 );
or ( n2321 , n2320 , n9 );
not ( n2322 , n7 );
not ( n2323 , n2322 );
not ( n2324 , n1392 );
nand ( n2325 , n2324 , n1063 );
not ( n2326 , n1196 );
nand ( n2327 , n2325 , n1270 , n2326 );
not ( n2328 , n2327 );
or ( n2329 , n2323 , n2328 );
not ( n2330 , n1025 );
not ( n2331 , n2330 );
nand ( n2332 , n2329 , n2331 );
nand ( n2333 , n8 , n2332 );
nand ( n2334 , n2321 , n2333 );
nor ( n2335 , n2288 , n2291 , n2334 );
nand ( n2336 , n2240 , n2335 );
not ( n2337 , n2336 );
not ( n2338 , n2337 );
and ( n2339 , n2211 , n2338 );
not ( n2340 , n2209 );
not ( n2341 , n2336 );
and ( n2342 , n2340 , n2341 );
nor ( n2343 , n2339 , n2342 );
and ( n2344 , n2011 , n2343 );
not ( n2345 , n2011 );
not ( n2346 , n2343 );
and ( n2347 , n2345 , n2346 );
nor ( n2348 , n2344 , n2347 );
nor ( n2349 , n1482 , n2348 );
not ( n2350 , n2349 );
nand ( n2351 , n1482 , n2348 );
not ( n2352 , n1 );
nand ( n2353 , n2350 , n2351 , n2352 );
nand ( n2354 , n742 , n2353 );
not ( n2355 , n1 );
and ( n2356 , n267 , n104 );
not ( n2357 , n267 );
not ( n2358 , n104 );
and ( n2359 , n2357 , n2358 );
nor ( n2360 , n2356 , n2359 );
not ( n2361 , n2360 );
or ( n2362 , n2355 , n2361 );
not ( n2363 , n2358 );
not ( n2364 , n195 );
not ( n2365 , n194 );
not ( n2366 , n2365 );
not ( n2367 , n188 );
nand ( n2368 , n2367 , n190 );
not ( n2369 , n2368 );
not ( n2370 , n2369 );
not ( n2371 , n191 );
nor ( n2372 , n2370 , n2371 );
nand ( n2373 , n192 , n2372 );
not ( n2374 , n2373 );
not ( n2375 , n192 );
not ( n2376 , n190 );
nand ( n2377 , n188 , n2376 );
nor ( n2378 , n2377 , n189 );
nand ( n2379 , n2375 , n2378 );
not ( n2380 , n2379 );
nor ( n2381 , n2374 , n2380 );
nand ( n2382 , n191 , n192 );
not ( n2383 , n2382 );
not ( n2384 , n190 );
nand ( n2385 , n2384 , n189 );
not ( n2386 , n2385 );
nand ( n2387 , n2383 , n2386 );
not ( n2388 , n193 );
nand ( n2389 , n2388 , n2372 );
not ( n2390 , n191 );
nand ( n2391 , n2369 , n189 );
not ( n2392 , n2391 );
not ( n2393 , n192 );
and ( n2394 , n2392 , n2393 );
nand ( n2395 , n2390 , n2394 );
nand ( n2396 , n2381 , n2387 , n2389 , n2395 );
not ( n2397 , n2396 );
or ( n2398 , n2366 , n2397 );
not ( n2399 , n191 );
nand ( n2400 , n188 , n190 );
nor ( n2401 , n189 , n2400 );
nand ( n2402 , n192 , n2401 );
not ( n2403 , n2402 );
nand ( n2404 , n2399 , n2403 );
nand ( n2405 , n2398 , n2404 );
not ( n2406 , n2405 );
not ( n2407 , n192 );
not ( n2408 , n189 );
nand ( n2409 , n2408 , n188 );
nor ( n2410 , n2407 , n2409 );
not ( n2411 , n2410 );
buf ( n2412 , n2400 );
not ( n2413 , n2412 );
nand ( n2414 , n191 , n2413 );
not ( n2415 , n192 );
not ( n2416 , n190 );
nor ( n2417 , n2416 , n189 );
nand ( n2418 , n2415 , n2417 );
nand ( n2419 , n2411 , n2414 , n2418 );
nand ( n2420 , n193 , n2419 );
nor ( n2421 , n189 , n2400 );
not ( n2422 , n2421 );
nor ( n2423 , n192 , n2422 );
not ( n2424 , n2423 );
nand ( n2425 , n188 , n190 );
not ( n2426 , n2425 );
nand ( n2427 , n2426 , n189 );
not ( n2428 , n2427 );
nand ( n2429 , n2428 , n192 );
not ( n2430 , n2429 );
nand ( n2431 , n191 , n2430 );
nand ( n2432 , n2420 , n2424 , n2431 );
nand ( n2433 , n194 , n2432 );
not ( n2434 , n193 );
not ( n2435 , n191 );
nand ( n2436 , n2435 , n2421 );
or ( n2437 , n2434 , n2436 );
not ( n2438 , n193 );
not ( n2439 , n2438 );
not ( n2440 , n191 );
nand ( n2441 , n188 , n189 );
not ( n2442 , n2441 );
nand ( n2443 , n2376 , n2442 );
not ( n2444 , n2443 );
nand ( n2445 , n2440 , n2444 );
nor ( n2446 , n188 , n190 );
not ( n2447 , n2446 );
not ( n2448 , n2447 );
nand ( n2449 , n2448 , n189 );
not ( n2450 , n2449 );
nand ( n2451 , n2450 , n192 );
not ( n2452 , n2391 );
nand ( n2453 , n191 , n2452 );
nand ( n2454 , n2445 , n2451 , n2453 , n2379 );
not ( n2455 , n2454 );
or ( n2456 , n2439 , n2455 );
not ( n2457 , n191 );
not ( n2458 , n2451 );
nand ( n2459 , n2457 , n2458 );
nand ( n2460 , n2456 , n2459 );
not ( n2461 , n2460 );
nand ( n2462 , n2406 , n2433 , n2437 , n2461 );
not ( n2463 , n2462 );
or ( n2464 , n2364 , n2463 );
not ( n2465 , n193 );
not ( n2466 , n189 );
nand ( n2467 , n2466 , n2369 );
not ( n2468 , n2467 );
nand ( n2469 , n2383 , n2468 );
nor ( n2470 , n2465 , n2469 );
not ( n2471 , n189 );
and ( n2472 , n191 , n193 );
not ( n2473 , n192 );
not ( n2474 , n2447 );
nand ( n2475 , n2473 , n2474 );
not ( n2476 , n2475 );
and ( n2477 , n2471 , n2472 , n2476 );
nor ( n2478 , n2470 , n2477 );
not ( n2479 , n193 );
not ( n2480 , n2479 );
not ( n2481 , n2449 );
not ( n2482 , n2481 );
nor ( n2483 , n191 , n2482 );
not ( n2484 , n2483 );
not ( n2485 , n192 );
nand ( n2486 , n2485 , n2444 );
not ( n2487 , n191 );
not ( n2488 , n188 );
nand ( n2489 , n2488 , n189 );
nor ( n2490 , n192 , n2489 );
nand ( n2491 , n2487 , n2490 );
and ( n2492 , n2486 , n2491 );
nand ( n2493 , n2471 , n2474 );
not ( n2494 , n2493 );
not ( n2495 , n2494 );
not ( n2496 , n2495 );
not ( n2497 , n192 );
nand ( n2498 , n2496 , n2497 );
nand ( n2499 , n2484 , n2492 , n2498 );
not ( n2500 , n2499 );
or ( n2501 , n2480 , n2500 );
not ( n2502 , n193 );
nand ( n2503 , n191 , n2502 );
not ( n2504 , n2503 );
nand ( n2505 , n2504 , n2494 );
nand ( n2506 , n2501 , n2505 );
and ( n2507 , n194 , n2506 );
not ( n2508 , n192 );
not ( n2509 , n2442 );
nor ( n2510 , n2508 , n2509 );
not ( n2511 , n2510 );
not ( n2512 , n2511 );
or ( n2513 , n2512 , n2423 );
nand ( n2514 , n2513 , n191 );
and ( n2515 , n2404 , n2514 );
and ( n2516 , n193 , n194 );
not ( n2517 , n2516 );
nor ( n2518 , n2515 , n2517 );
nor ( n2519 , n2507 , n2518 );
nand ( n2520 , n2464 , n2478 , n2519 );
not ( n2521 , n194 );
not ( n2522 , n2521 );
not ( n2523 , n193 );
not ( n2524 , n2523 );
nand ( n2525 , n189 , n190 );
nor ( n2526 , n192 , n2525 );
nand ( n2527 , n191 , n2526 );
buf ( n2528 , n2378 );
nand ( n2529 , n191 , n2528 );
not ( n2530 , n2493 );
nand ( n2531 , n2530 , n192 );
not ( n2532 , n2531 );
not ( n2533 , n191 );
nand ( n2534 , n2532 , n2533 );
nand ( n2535 , n2527 , n2529 , n2534 );
not ( n2536 , n2535 );
or ( n2537 , n2524 , n2536 );
not ( n2538 , n191 );
nor ( n2539 , n2451 , n2538 );
not ( n2540 , n2539 );
and ( n2541 , n2469 , n2540 );
nand ( n2542 , n2537 , n2541 );
not ( n2543 , n2542 );
or ( n2544 , n2522 , n2543 );
not ( n2545 , n194 );
and ( n2546 , n193 , n2545 );
not ( n2547 , n2467 );
not ( n2548 , n2547 );
or ( n2549 , n191 , n2548 );
nor ( n2550 , n191 , n2475 );
not ( n2551 , n2550 );
not ( n2552 , n191 );
not ( n2553 , n2429 );
nand ( n2554 , n2552 , n2553 );
nand ( n2555 , n2549 , n2551 , n2554 );
nand ( n2556 , n2546 , n2555 );
nand ( n2557 , n2544 , n2556 );
not ( n2558 , n194 );
not ( n2559 , n191 );
nand ( n2560 , n193 , n2559 );
not ( n2561 , n2560 );
nand ( n2562 , n2561 , n2444 );
nand ( n2563 , n192 , n2378 );
not ( n2564 , n2563 );
nand ( n2565 , n191 , n2564 );
and ( n2566 , n2562 , n2565 );
and ( n2567 , n191 , n2401 );
nand ( n2568 , n193 , n2567 );
not ( n2569 , n2427 );
not ( n2570 , n192 );
nand ( n2571 , n2569 , n2570 );
not ( n2572 , n2571 );
nand ( n2573 , n191 , n2572 );
not ( n2574 , n2563 );
nor ( n2575 , n191 , n192 );
nand ( n2576 , n2575 , n2401 );
not ( n2577 , n2576 );
or ( n2578 , n2574 , n2577 );
not ( n2579 , n193 );
nand ( n2580 , n2578 , n2579 );
nand ( n2581 , n2568 , n2573 , n2580 );
not ( n2582 , n2581 );
nand ( n2583 , n2566 , n2582 );
and ( n2584 , n2558 , n2583 );
nor ( n2585 , n191 , n193 );
not ( n2586 , n2585 );
not ( n2587 , n2391 );
nand ( n2588 , n2587 , n192 );
buf ( n2589 , n2588 );
nor ( n2590 , n2586 , n2589 );
not ( n2591 , n2590 );
not ( n2592 , n193 );
nor ( n2593 , n2592 , n2540 );
not ( n2594 , n2593 );
nand ( n2595 , n2591 , n2594 );
nor ( n2596 , n2584 , n2595 );
not ( n2597 , n193 );
not ( n2598 , n2376 );
nor ( n2599 , n191 , n192 );
not ( n2600 , n2599 );
or ( n2601 , n2598 , n2600 );
not ( n2602 , n2495 );
not ( n2603 , n191 );
nand ( n2604 , n2602 , n2603 );
nand ( n2605 , n2601 , n2604 );
not ( n2606 , n2605 );
or ( n2607 , n2597 , n2606 );
nand ( n2608 , n2607 , n2551 );
not ( n2609 , n194 );
not ( n2610 , n192 );
nor ( n2611 , n2610 , n2525 );
not ( n2612 , n2611 );
not ( n2613 , n191 );
not ( n2614 , n2427 );
nand ( n2615 , n2613 , n2614 );
nand ( n2616 , n2612 , n2615 );
and ( n2617 , n193 , n2616 );
not ( n2618 , n193 );
and ( n2619 , n191 , n2410 );
not ( n2620 , n191 );
not ( n2621 , n2370 );
and ( n2622 , n2620 , n2621 );
nor ( n2623 , n2619 , n2622 );
not ( n2624 , n192 );
nor ( n2625 , n188 , n189 );
nand ( n2626 , n2624 , n2625 );
nand ( n2627 , n2623 , n2626 );
and ( n2628 , n2618 , n2627 );
nor ( n2629 , n2617 , n2628 );
not ( n2630 , n2493 );
nand ( n2631 , n2630 , n191 );
not ( n2632 , n2443 );
nand ( n2633 , n2632 , n191 );
nor ( n2634 , n192 , n2377 );
nand ( n2635 , n191 , n2634 );
nand ( n2636 , n2633 , n2635 );
not ( n2637 , n2636 );
nand ( n2638 , n2629 , n2631 , n2637 );
not ( n2639 , n2638 );
or ( n2640 , n2609 , n2639 );
not ( n2641 , n193 );
not ( n2642 , n2573 );
nand ( n2643 , n2641 , n2642 );
nand ( n2644 , n2640 , n2643 );
nor ( n2645 , n2608 , n2644 );
and ( n2646 , n2596 , n2645 );
nor ( n2647 , n2646 , n195 );
nor ( n2648 , n2557 , n2647 );
not ( n2649 , n2648 );
nor ( n2650 , n2520 , n2649 );
not ( n2651 , n2650 );
and ( n2652 , n2363 , n2651 );
nand ( n2653 , n195 , n2462 );
and ( n2654 , n2648 , n2478 , n2519 , n2653 );
and ( n2655 , n2358 , n2654 );
nor ( n2656 , n2652 , n2655 );
not ( n2657 , n194 );
not ( n2658 , n191 );
not ( n2659 , n2658 );
not ( n2660 , n2379 );
nor ( n2661 , n2660 , n2572 );
not ( n2662 , n2661 );
not ( n2663 , n2662 );
or ( n2664 , n2659 , n2663 );
nand ( n2665 , n2383 , n2474 );
nor ( n2666 , n193 , n2665 );
not ( n2667 , n2666 );
nand ( n2668 , n2664 , n2667 );
nand ( n2669 , n2657 , n2668 );
not ( n2670 , n2417 );
or ( n2671 , n2670 , n2586 );
not ( n2672 , n193 );
or ( n2673 , n2672 , n2633 );
nand ( n2674 , n2671 , n2673 , n2475 );
not ( n2675 , n191 );
nand ( n2676 , n2675 , n2474 );
not ( n2677 , n2676 );
nor ( n2678 , n2412 , n2382 );
or ( n2679 , n2674 , n2677 , n2678 );
nand ( n2680 , n2679 , n194 );
not ( n2681 , n2546 );
or ( n2682 , n191 , n2525 );
not ( n2683 , n2452 );
nand ( n2684 , n2682 , n2683 );
not ( n2685 , n2684 );
or ( n2686 , n2681 , n2685 );
nand ( n2687 , n191 , n2614 );
not ( n2688 , n2687 );
nand ( n2689 , n2625 , n2599 );
not ( n2690 , n2689 );
or ( n2691 , n2688 , n2690 );
not ( n2692 , n193 );
nand ( n2693 , n2691 , n2692 );
nand ( n2694 , n2686 , n2693 );
not ( n2695 , n2409 );
not ( n2696 , n2695 );
and ( n2697 , n2696 , n2482 );
not ( n2698 , n191 );
not ( n2699 , n192 );
nand ( n2700 , n2699 , n193 );
nor ( n2701 , n2697 , n2698 , n2700 );
nor ( n2702 , n2694 , n2590 , n2701 );
and ( n2703 , n2669 , n2680 , n2702 );
nor ( n2704 , n2703 , n195 );
not ( n2705 , n2704 );
not ( n2706 , n193 );
and ( n2707 , n2706 , n2678 );
not ( n2708 , n2495 );
nand ( n2709 , n2708 , n2599 );
not ( n2710 , n191 );
nor ( n2711 , n2710 , n2467 );
nand ( n2712 , n193 , n2711 );
not ( n2713 , n192 );
nand ( n2714 , n2713 , n2481 );
not ( n2715 , n2714 );
nand ( n2716 , n191 , n2715 );
and ( n2717 , n2712 , n2716 );
not ( n2718 , n193 );
not ( n2719 , n191 );
nand ( n2720 , n2719 , n2611 );
not ( n2721 , n2720 );
and ( n2722 , n2718 , n2721 );
not ( n2723 , n2718 );
not ( n2724 , n191 );
not ( n2725 , n2563 );
nand ( n2726 , n2724 , n2725 );
not ( n2727 , n2726 );
and ( n2728 , n2723 , n2727 );
nor ( n2729 , n2722 , n2728 );
nand ( n2730 , n194 , n2709 , n2717 , n2729 );
not ( n2731 , n2730 );
not ( n2732 , n194 );
not ( n2733 , n193 );
not ( n2734 , n191 );
nor ( n2735 , n2734 , n2486 );
nand ( n2736 , n2733 , n2735 );
not ( n2737 , n2736 );
nor ( n2738 , n2593 , n2737 );
not ( n2739 , n2509 );
nand ( n2740 , n2739 , n2575 );
not ( n2741 , n2740 );
nand ( n2742 , n2599 , n2547 );
not ( n2743 , n2742 );
or ( n2744 , n2741 , n2743 );
nand ( n2745 , n2744 , n193 );
not ( n2746 , n193 );
not ( n2747 , n191 );
nand ( n2748 , n2747 , n2528 );
not ( n2749 , n2377 );
nand ( n2750 , n2749 , n192 );
not ( n2751 , n2750 );
not ( n2752 , n191 );
nand ( n2753 , n2751 , n2752 );
not ( n2754 , n2714 );
not ( n2755 , n191 );
nand ( n2756 , n2754 , n2755 );
nand ( n2757 , n2748 , n2753 , n2756 );
nand ( n2758 , n2746 , n2757 );
nand ( n2759 , n2732 , n2738 , n2745 , n2758 );
not ( n2760 , n2759 );
or ( n2761 , n2731 , n2760 );
not ( n2762 , n2740 );
nand ( n2763 , n2762 , n193 , n2376 );
nand ( n2764 , n2761 , n2763 );
nor ( n2765 , n2707 , n2764 );
nor ( n2766 , n192 , n2467 );
nand ( n2767 , n191 , n2766 );
not ( n2768 , n2430 );
not ( n2769 , n2768 );
not ( n2770 , n191 );
nand ( n2771 , n2770 , n192 );
or ( n2772 , n2385 , n2771 );
not ( n2773 , n2772 );
or ( n2774 , n2769 , n2773 );
not ( n2775 , n193 );
nand ( n2776 , n2774 , n2775 );
and ( n2777 , n2767 , n2445 , n2776 );
not ( n2778 , n193 );
not ( n2779 , n191 );
nor ( n2780 , n2779 , n192 );
not ( n2781 , n2780 );
or ( n2782 , n190 , n2781 );
nand ( n2783 , n191 , n2695 );
nand ( n2784 , n2782 , n2783 );
and ( n2785 , n2778 , n2784 );
not ( n2786 , n2778 );
not ( n2787 , n2766 );
nor ( n2788 , n191 , n2588 );
not ( n2789 , n2788 );
not ( n2790 , n2527 );
nor ( n2791 , n2790 , n2539 );
nand ( n2792 , n2787 , n2789 , n2791 );
and ( n2793 , n2786 , n2792 );
nor ( n2794 , n2785 , n2793 );
not ( n2795 , n2739 );
or ( n2796 , n193 , n2795 );
not ( n2797 , n2564 );
not ( n2798 , n2494 );
nor ( n2799 , n2798 , n193 );
not ( n2800 , n2799 );
nand ( n2801 , n2796 , n2797 , n2800 );
nand ( n2802 , n194 , n2801 );
not ( n2803 , n2621 );
nor ( n2804 , n192 , n2803 );
nand ( n2805 , n191 , n2804 );
not ( n2806 , n191 );
nor ( n2807 , n192 , n2385 );
nand ( n2808 , n2806 , n2807 );
nand ( n2809 , n2805 , n2808 );
nand ( n2810 , n2471 , n2780 );
nand ( n2811 , n192 , n2468 );
not ( n2812 , n2811 );
nand ( n2813 , n2585 , n2812 );
nand ( n2814 , n2444 , n192 );
not ( n2815 , n2814 );
not ( n2816 , n2815 );
not ( n2817 , n2403 );
nand ( n2818 , n2816 , n2817 , n2604 );
nand ( n2819 , n193 , n2818 );
nand ( n2820 , n2810 , n2813 , n2819 );
or ( n2821 , n2809 , n2820 );
not ( n2822 , n194 );
nand ( n2823 , n2821 , n2822 );
nand ( n2824 , n2777 , n2794 , n2802 , n2823 );
nand ( n2825 , n195 , n2824 );
nand ( n2826 , n2705 , n2765 , n2825 );
not ( n2827 , n2826 );
nand ( n2828 , n191 , n2481 );
not ( n2829 , n2828 );
not ( n2830 , n192 );
nor ( n2831 , n2830 , n2489 );
not ( n2832 , n2831 );
not ( n2833 , n2832 );
not ( n2834 , n2661 );
or ( n2835 , n2833 , n2834 );
nand ( n2836 , n2835 , n191 );
not ( n2837 , n2836 );
or ( n2838 , n2829 , n2837 );
not ( n2839 , n194 );
nor ( n2840 , n2839 , n193 );
nand ( n2841 , n2838 , n2840 );
not ( n2842 , n2546 );
not ( n2843 , n191 );
nand ( n2844 , n2843 , n2512 );
nand ( n2845 , n2403 , n191 );
nand ( n2846 , n2844 , n2631 , n2845 );
not ( n2847 , n2846 );
or ( n2848 , n2842 , n2847 );
nand ( n2849 , n2599 , n2444 );
not ( n2850 , n2849 );
nand ( n2851 , n2383 , n2494 );
not ( n2852 , n2851 );
or ( n2853 , n2850 , n2852 );
not ( n2854 , n193 );
nand ( n2855 , n2853 , n2854 );
nand ( n2856 , n2848 , n2855 );
not ( n2857 , n2856 );
not ( n2858 , n194 );
not ( n2859 , n193 );
not ( n2860 , n191 );
nor ( n2861 , n2860 , n2418 );
nand ( n2862 , n2859 , n2861 );
not ( n2863 , n2808 );
not ( n2864 , n2615 );
or ( n2865 , n2863 , n2864 );
not ( n2866 , n193 );
nand ( n2867 , n2865 , n2866 );
nand ( n2868 , n2862 , n2720 , n2867 );
nand ( n2869 , n2858 , n2868 );
not ( n2870 , n191 );
not ( n2871 , n2870 );
nor ( n2872 , n2412 , n192 );
not ( n2873 , n2872 );
nand ( n2874 , n2873 , n2811 , n2714 );
not ( n2875 , n2874 );
or ( n2876 , n2871 , n2875 );
and ( n2877 , n2633 , n2424 );
nand ( n2878 , n2876 , n2877 );
nand ( n2879 , n2516 , n2878 );
nand ( n2880 , n2841 , n2857 , n2869 , n2879 );
not ( n2881 , n2880 );
or ( n2882 , n2430 , n2458 );
nand ( n2883 , n2882 , n2472 );
and ( n2884 , n2867 , n2883 );
not ( n2885 , n2531 );
not ( n2886 , n2814 );
nand ( n2887 , n2886 , n191 );
not ( n2888 , n2887 );
or ( n2889 , n2885 , n2888 );
not ( n2890 , n193 );
nand ( n2891 , n2889 , n2890 );
not ( n2892 , n193 );
not ( n2893 , n2892 );
not ( n2894 , n188 );
not ( n2895 , n2894 );
not ( n2896 , n2383 );
or ( n2897 , n2895 , n2896 );
nand ( n2898 , n2897 , n2529 );
not ( n2899 , n2898 );
or ( n2900 , n2893 , n2899 );
not ( n2901 , n2411 );
nand ( n2902 , n2561 , n2901 );
nand ( n2903 , n2900 , n2902 );
nand ( n2904 , n2453 , n2404 );
or ( n2905 , n2903 , n2904 );
nand ( n2906 , n2905 , n194 );
nand ( n2907 , n2884 , n2891 , n2906 );
not ( n2908 , n194 );
not ( n2909 , n2908 );
not ( n2910 , n2472 );
nand ( n2911 , n192 , n2417 );
not ( n2912 , n2911 );
not ( n2913 , n2912 );
or ( n2914 , n2910 , n2913 );
nand ( n2915 , n193 , n2494 );
nand ( n2916 , n2914 , n2915 );
not ( n2917 , n2916 );
or ( n2918 , n2909 , n2917 );
not ( n2919 , n194 );
or ( n2920 , n193 , n2376 , n192 );
nand ( n2921 , n2920 , n2527 );
and ( n2922 , n2919 , n2921 );
nor ( n2923 , n2922 , n2477 );
nand ( n2924 , n2918 , n2923 );
or ( n2925 , n2907 , n2924 );
nand ( n2926 , n2925 , n2364 );
not ( n2927 , n193 );
not ( n2928 , n191 );
nand ( n2929 , n2928 , n2872 );
not ( n2930 , n2815 );
not ( n2931 , n191 );
nand ( n2932 , n2931 , n2831 );
nand ( n2933 , n2929 , n2930 , n2932 );
not ( n2934 , n2933 );
or ( n2935 , n2927 , n2934 );
nand ( n2936 , n2935 , n2772 );
not ( n2937 , n2936 );
not ( n2938 , n2585 );
not ( n2939 , n2547 );
or ( n2940 , n2938 , n2939 );
nand ( n2941 , n2940 , n2845 );
nand ( n2942 , n194 , n2941 );
not ( n2943 , n194 );
nand ( n2944 , n191 , n2490 );
and ( n2945 , n2753 , n2944 );
not ( n2946 , n193 );
nand ( n2947 , n2946 , n2444 );
not ( n2948 , n2947 );
not ( n2949 , n191 );
nand ( n2950 , n2949 , n2749 );
nor ( n2951 , n193 , n2950 );
nor ( n2952 , n2948 , n2951 );
not ( n2953 , n2418 );
nand ( n2954 , n2953 , n2561 );
not ( n2955 , n2750 );
nand ( n2956 , n192 , n2625 );
nand ( n2957 , n2511 , n2956 );
or ( n2958 , n2955 , n2957 );
not ( n2959 , n193 );
nand ( n2960 , n2958 , n2959 );
nand ( n2961 , n2945 , n2952 , n2954 , n2960 );
nand ( n2962 , n2943 , n2961 );
nand ( n2963 , n2937 , n2942 , n2962 );
not ( n2964 , n2516 );
not ( n2965 , n2894 );
not ( n2966 , n192 );
and ( n2967 , n2965 , n2966 );
and ( n2968 , n191 , n2749 );
nor ( n2969 , n2967 , n2968 );
nand ( n2970 , n2969 , n2956 , n2676 );
not ( n2971 , n2970 );
or ( n2972 , n2964 , n2971 );
not ( n2973 , n193 );
not ( n2974 , n2753 );
and ( n2975 , n2973 , n2974 );
not ( n2976 , n192 );
nand ( n2977 , n2976 , n2695 );
not ( n2978 , n2977 );
and ( n2979 , n2472 , n2978 );
nor ( n2980 , n2975 , n2979 );
nand ( n2981 , n2972 , n2980 );
or ( n2982 , n2963 , n2981 );
nand ( n2983 , n2982 , n195 );
nand ( n2984 , n2881 , n2926 , n2983 );
buf ( n2985 , n2984 );
not ( n2986 , n2985 );
not ( n2987 , n2986 );
and ( n2988 , n2827 , n2987 );
not ( n2989 , n2827 );
not ( n2990 , n2984 );
not ( n2991 , n2990 );
not ( n2992 , n2991 );
and ( n2993 , n2989 , n2992 );
nor ( n2994 , n2988 , n2993 );
and ( n2995 , n2656 , n2994 );
not ( n2996 , n2656 );
not ( n2997 , n2994 );
and ( n2998 , n2996 , n2997 );
nor ( n2999 , n2995 , n2998 );
not ( n3000 , n2999 );
not ( n3001 , n180 );
nand ( n3002 , n3001 , n182 );
not ( n3003 , n180 );
not ( n3004 , n3003 );
nor ( n3005 , n181 , n182 );
nand ( n3006 , n3004 , n3005 );
buf ( n3007 , n3006 );
not ( n3008 , n3007 );
not ( n3009 , n3008 );
and ( n3010 , n3002 , n3009 );
nand ( n3011 , n184 , n185 );
nor ( n3012 , n3010 , n183 , n3011 );
not ( n3013 , n186 );
not ( n3014 , n3013 );
not ( n3015 , n184 );
not ( n3016 , n3015 );
not ( n3017 , n180 );
nand ( n3018 , n181 , n182 );
nor ( n3019 , n3017 , n3018 );
not ( n3020 , n3019 );
not ( n3021 , n3020 );
not ( n3022 , n183 );
nand ( n3023 , n3021 , n3022 );
not ( n3024 , n183 );
not ( n3025 , n181 );
nand ( n3026 , n3025 , n182 );
not ( n3027 , n3026 );
not ( n3028 , n180 );
nand ( n3029 , n3027 , n3028 );
not ( n3030 , n3029 );
nand ( n3031 , n3024 , n3030 );
nand ( n3032 , n3023 , n3031 );
not ( n3033 , n3032 );
or ( n3034 , n3016 , n3033 );
nand ( n3035 , n183 , n184 );
nor ( n3036 , n181 , n182 );
not ( n3037 , n3036 );
or ( n3038 , n3035 , n3037 );
not ( n3039 , n3038 );
not ( n3040 , n185 );
nand ( n3041 , n3039 , n3040 );
nand ( n3042 , n3034 , n3041 );
not ( n3043 , n3042 );
or ( n3044 , n3014 , n3043 );
nand ( n3045 , n185 , n3013 );
not ( n3046 , n3045 );
nand ( n3047 , n180 , n181 );
or ( n3048 , n184 , n3047 );
not ( n3049 , n181 );
nor ( n3050 , n3049 , n182 );
nand ( n3051 , n180 , n3050 );
not ( n3052 , n3051 );
not ( n3053 , n3052 );
not ( n3054 , n3053 );
not ( n3055 , n3054 );
nand ( n3056 , n3048 , n3055 );
nand ( n3057 , n3046 , n3056 );
nand ( n3058 , n3044 , n3057 );
nor ( n3059 , n3012 , n3058 );
not ( n3060 , n185 );
not ( n3061 , n184 );
not ( n3062 , n183 );
nor ( n3063 , n180 , n182 );
nand ( n3064 , n3062 , n3063 );
not ( n3065 , n3064 );
nand ( n3066 , n3061 , n3065 );
not ( n3067 , n184 );
not ( n3068 , n3020 );
not ( n3069 , n3068 );
or ( n3070 , n3067 , n3069 );
nand ( n3071 , n183 , n3052 );
not ( n3072 , n3071 );
not ( n3073 , n184 );
nand ( n3074 , n3072 , n3073 );
nand ( n3075 , n3070 , n3074 );
not ( n3076 , n3075 );
nand ( n3077 , n3066 , n3076 );
and ( n3078 , n3060 , n3077 );
nor ( n3079 , n3078 , n187 );
not ( n3080 , n183 );
not ( n3081 , n3037 );
nand ( n3082 , n3080 , n3081 );
not ( n3083 , n184 );
nand ( n3084 , n3083 , n3081 );
nand ( n3085 , n3082 , n3084 );
not ( n3086 , n181 );
nor ( n3087 , n3086 , n180 );
not ( n3088 , n3087 );
not ( n3089 , n3088 );
nor ( n3090 , n184 , n185 );
not ( n3091 , n3090 );
not ( n3092 , n3091 );
nand ( n3093 , n3089 , n3092 );
not ( n3094 , n183 );
nand ( n3095 , n181 , n182 );
not ( n3096 , n3095 );
nand ( n3097 , n184 , n3096 );
nor ( n3098 , n3094 , n3097 );
not ( n3099 , n3098 );
not ( n3100 , n3026 );
nand ( n3101 , n3100 , n180 );
not ( n3102 , n3101 );
not ( n3103 , n3102 );
not ( n3104 , n184 );
nor ( n3105 , n3103 , n3104 );
nand ( n3106 , n185 , n3105 );
nand ( n3107 , n3093 , n3099 , n3106 );
or ( n3108 , n3085 , n3107 );
nand ( n3109 , n3108 , n186 );
nand ( n3110 , n3059 , n3079 , n3109 );
not ( n3111 , n3110 );
nand ( n3112 , n180 , n182 );
or ( n3113 , n185 , n3112 );
and ( n3114 , n183 , n3030 );
not ( n3115 , n3114 );
nand ( n3116 , n3028 , n3005 );
or ( n3117 , n185 , n3116 );
nand ( n3118 , n3113 , n3115 , n3117 );
and ( n3119 , n186 , n3118 );
not ( n3120 , n3102 );
not ( n3121 , n3120 );
not ( n3122 , n184 );
nand ( n3123 , n3121 , n3122 );
not ( n3124 , n3123 );
nor ( n3125 , n3119 , n3124 );
not ( n3126 , n3003 );
not ( n3127 , n3126 );
not ( n3128 , n183 );
nand ( n3129 , n3128 , n184 );
not ( n3130 , n3129 );
nand ( n3131 , n3127 , n3130 );
not ( n3132 , n3050 );
nor ( n3133 , n183 , n3132 );
nand ( n3134 , n184 , n3133 );
not ( n3135 , n184 );
not ( n3136 , n181 );
nand ( n3137 , n3136 , n180 );
nor ( n3138 , n183 , n3137 );
nand ( n3139 , n3135 , n3138 );
and ( n3140 , n3131 , n3134 , n3139 );
nand ( n3141 , n3050 , n3003 );
not ( n3142 , n3141 );
nand ( n3143 , n183 , n3142 );
not ( n3144 , n3143 );
nand ( n3145 , n3092 , n3144 );
nor ( n3146 , n181 , n184 );
nand ( n3147 , n3063 , n3146 );
nor ( n3148 , n180 , n3018 );
nand ( n3149 , n183 , n3148 );
nand ( n3150 , n183 , n3102 );
nand ( n3151 , n3147 , n3149 , n3150 );
nand ( n3152 , n185 , n3151 );
nand ( n3153 , n3140 , n3145 , n3152 );
nand ( n3154 , n3013 , n3153 );
not ( n3155 , n185 );
not ( n3156 , n3155 );
or ( n3157 , n181 , n3129 );
not ( n3158 , n3002 );
nand ( n3159 , n184 , n3158 );
nand ( n3160 , n3157 , n3159 );
not ( n3161 , n3160 );
or ( n3162 , n3156 , n3161 );
nand ( n3163 , n183 , n3019 );
not ( n3164 , n3163 );
not ( n3165 , n3137 );
not ( n3166 , n183 );
nor ( n3167 , n3166 , n184 );
nand ( n3168 , n3165 , n3167 );
not ( n3169 , n3168 );
or ( n3170 , n3164 , n3169 );
not ( n3171 , n185 );
nand ( n3172 , n3170 , n3171 );
nand ( n3173 , n3162 , n3172 );
not ( n3174 , n183 );
not ( n3175 , n3141 );
nand ( n3176 , n3174 , n3175 );
not ( n3177 , n3176 );
nand ( n3178 , n184 , n3177 );
not ( n3179 , n3177 );
nor ( n3180 , n183 , n3047 );
nand ( n3181 , n184 , n3180 );
not ( n3182 , n183 );
nor ( n3183 , n3182 , n3006 );
nand ( n3184 , n184 , n3183 );
nand ( n3185 , n3179 , n3074 , n3181 , n3184 );
nand ( n3186 , n185 , n3185 );
nand ( n3187 , n3178 , n3186 );
nor ( n3188 , n3173 , n3187 );
nand ( n3189 , n187 , n3125 , n3154 , n3188 );
not ( n3190 , n3189 );
or ( n3191 , n3111 , n3190 );
not ( n3192 , n184 );
not ( n3193 , n183 );
and ( n3194 , n3102 , n3193 );
nand ( n3195 , n3192 , n3194 );
not ( n3196 , n3195 );
and ( n3197 , n185 , n3196 );
not ( n3198 , n185 );
and ( n3199 , n3198 , n3098 );
nor ( n3200 , n3197 , n3199 );
not ( n3201 , n185 );
not ( n3202 , n3030 );
not ( n3203 , n3202 );
nand ( n3204 , n3167 , n3203 );
not ( n3205 , n3204 );
or ( n3206 , n3201 , n3205 );
not ( n3207 , n185 );
nand ( n3208 , n180 , n181 );
not ( n3209 , n3208 );
nand ( n3210 , n3209 , n183 );
not ( n3211 , n3210 );
not ( n3212 , n184 );
nand ( n3213 , n3211 , n3212 );
nand ( n3214 , n3207 , n3213 );
nand ( n3215 , n3206 , n3214 );
nand ( n3216 , n3130 , n3008 );
not ( n3217 , n3116 );
nor ( n3218 , n183 , n184 );
not ( n3219 , n3218 );
not ( n3220 , n3219 );
nand ( n3221 , n3217 , n3220 );
nand ( n3222 , n3142 , n184 );
not ( n3223 , n185 );
nor ( n3224 , n3222 , n3223 );
not ( n3225 , n3224 );
nand ( n3226 , n3215 , n3216 , n3221 , n3225 );
nand ( n3227 , n186 , n3226 );
not ( n3228 , n185 );
not ( n3229 , n3228 );
not ( n3230 , n184 );
nand ( n3231 , n3230 , n3203 );
not ( n3232 , n3026 );
not ( n3233 , n3232 );
not ( n3234 , n3233 );
nand ( n3235 , n3234 , n183 );
not ( n3236 , n3235 );
not ( n3237 , n184 );
nand ( n3238 , n3236 , n3237 );
not ( n3239 , n3238 );
not ( n3240 , n3239 );
not ( n3241 , n183 );
not ( n3242 , n3006 );
nand ( n3243 , n3241 , n3242 );
not ( n3244 , n3243 );
not ( n3245 , n184 );
nand ( n3246 , n3244 , n3245 );
nand ( n3247 , n3231 , n3240 , n3246 );
not ( n3248 , n3247 );
or ( n3249 , n3229 , n3248 );
not ( n3250 , n3112 );
nand ( n3251 , n3250 , n3218 );
not ( n3252 , n3251 );
nand ( n3253 , n3220 , n3175 );
not ( n3254 , n3253 );
or ( n3255 , n3252 , n3254 );
nand ( n3256 , n3255 , n185 );
nand ( n3257 , n3249 , n3256 );
not ( n3258 , n3011 );
not ( n3259 , n3183 );
not ( n3260 , n3259 );
nand ( n3261 , n3258 , n3260 );
not ( n3262 , n185 );
not ( n3263 , n3194 );
not ( n3264 , n184 );
nor ( n3265 , n3263 , n3264 );
nand ( n3266 , n3262 , n3265 );
nand ( n3267 , n3261 , n3266 );
or ( n3268 , n3257 , n3267 );
nand ( n3269 , n3268 , n3013 );
nand ( n3270 , n3200 , n3227 , n3269 );
not ( n3271 , n3270 );
nand ( n3272 , n3191 , n3271 );
not ( n3273 , n3272 );
not ( n3274 , n3273 );
not ( n3275 , n187 );
nand ( n3276 , n183 , n3063 );
not ( n3277 , n3112 );
and ( n3278 , n183 , n3277 );
not ( n3279 , n3278 );
and ( n3280 , n3276 , n3279 , n3235 );
nor ( n3281 , n3280 , n185 );
not ( n3282 , n185 );
nor ( n3283 , n3282 , n184 );
not ( n3284 , n3283 );
not ( n3285 , n3087 );
nor ( n3286 , n3285 , n183 );
not ( n3287 , n3286 );
or ( n3288 , n3284 , n3287 );
not ( n3289 , n180 );
nor ( n3290 , n3289 , n182 );
not ( n3291 , n3290 );
nor ( n3292 , n183 , n3291 );
nand ( n3293 , n184 , n3292 );
nand ( n3294 , n3288 , n3293 );
not ( n3295 , n3294 );
not ( n3296 , n3102 );
not ( n3297 , n3296 );
not ( n3298 , n185 );
nand ( n3299 , n3297 , n3298 );
not ( n3300 , n3233 );
nand ( n3301 , n3300 , n3090 );
nand ( n3302 , n3238 , n3295 , n3299 , n3301 );
or ( n3303 , n3281 , n3302 );
nand ( n3304 , n3303 , n3013 );
not ( n3305 , n184 );
nor ( n3306 , n183 , n3095 );
nand ( n3307 , n3305 , n3306 );
nand ( n3308 , n183 , n3290 );
not ( n3309 , n3308 );
not ( n3310 , n184 );
nand ( n3311 , n3309 , n3310 );
nand ( n3312 , n3307 , n3150 , n3311 );
nand ( n3313 , n185 , n3312 );
not ( n3314 , n3091 );
not ( n3315 , n3314 );
not ( n3316 , n3175 );
or ( n3317 , n3315 , n3316 );
not ( n3318 , n3149 );
nand ( n3319 , n3318 , n184 );
nand ( n3320 , n3317 , n3319 );
and ( n3321 , n186 , n3320 );
not ( n3322 , n185 );
and ( n3323 , n3239 , n3322 );
nor ( n3324 , n3321 , n3323 );
nand ( n3325 , n3304 , n3313 , n3324 );
or ( n3326 , n183 , n3002 );
not ( n3327 , n3326 );
nand ( n3328 , n3327 , n3258 );
and ( n3329 , n185 , n186 );
and ( n3330 , n184 , n3300 );
not ( n3331 , n182 );
nor ( n3332 , n3331 , n183 );
nor ( n3333 , n3330 , n3332 );
nand ( n3334 , n3333 , n3276 , n3084 );
nand ( n3335 , n3329 , n3334 );
nand ( n3336 , n3328 , n3168 , n3335 );
nor ( n3337 , n3325 , n3336 );
or ( n3338 , n3275 , n3337 );
nand ( n3339 , n184 , n3054 );
nor ( n3340 , n3126 , n3095 );
nand ( n3341 , n3167 , n3340 );
and ( n3342 , n3339 , n3341 );
not ( n3343 , n183 );
nor ( n3344 , n3343 , n3002 );
not ( n3345 , n3344 );
not ( n3346 , n3345 );
buf ( n3347 , n3283 );
nand ( n3348 , n3346 , n3347 );
not ( n3349 , n184 );
nor ( n3350 , n3349 , n182 );
nand ( n3351 , n183 , n3350 );
not ( n3352 , n3351 );
nand ( n3353 , n184 , n3030 );
not ( n3354 , n3353 );
or ( n3355 , n3352 , n3354 );
not ( n3356 , n185 );
nand ( n3357 , n3355 , n3356 );
nand ( n3358 , n3342 , n3348 , n3357 );
nand ( n3359 , n3358 , n186 , n3275 );
not ( n3360 , n3045 );
not ( n3361 , n184 );
nand ( n3362 , n3361 , n3278 );
not ( n3363 , n3116 );
nand ( n3364 , n184 , n3363 );
nand ( n3365 , n3362 , n3364 , n3319 );
nand ( n3366 , n3360 , n3365 );
not ( n3367 , n3013 );
not ( n3368 , n184 );
not ( n3369 , n3020 );
nand ( n3370 , n3368 , n3369 );
not ( n3371 , n3370 );
not ( n3372 , n3139 );
or ( n3373 , n3371 , n3372 );
not ( n3374 , n185 );
nand ( n3375 , n3373 , n3374 );
not ( n3376 , n3286 );
not ( n3377 , n3376 );
not ( n3378 , n185 );
nand ( n3379 , n3377 , n184 , n3378 );
nand ( n3380 , n3375 , n3213 , n3379 );
not ( n3381 , n3380 );
or ( n3382 , n3367 , n3381 );
not ( n3383 , n3195 );
nand ( n3384 , n183 , n3363 );
not ( n3385 , n3384 );
nand ( n3386 , n184 , n3385 );
not ( n3387 , n3386 );
or ( n3388 , n3383 , n3387 );
not ( n3389 , n185 );
nand ( n3390 , n3388 , n3389 );
nand ( n3391 , n3382 , n3390 );
not ( n3392 , n3391 );
and ( n3393 , n3359 , n3366 , n3392 );
nand ( n3394 , n3338 , n3393 );
not ( n3395 , n3394 );
not ( n3396 , n184 );
nor ( n3397 , n3396 , n3007 );
not ( n3398 , n3397 );
not ( n3399 , n3398 );
not ( n3400 , n3308 );
not ( n3401 , n3032 );
not ( n3402 , n3401 );
or ( n3403 , n3400 , n3402 );
nand ( n3404 , n3403 , n184 );
not ( n3405 , n3404 );
or ( n3406 , n3399 , n3405 );
not ( n3407 , n185 );
nand ( n3408 , n3406 , n3407 );
not ( n3409 , n184 );
not ( n3410 , n3409 );
not ( n3411 , n3306 );
nand ( n3412 , n3411 , n3143 , n3243 );
not ( n3413 , n3412 );
or ( n3414 , n3410 , n3413 );
not ( n3415 , n3105 );
not ( n3416 , n183 );
nand ( n3417 , n3416 , n3340 );
and ( n3418 , n3415 , n3417 );
nand ( n3419 , n3414 , n3418 );
nand ( n3420 , n185 , n3419 );
nand ( n3421 , n3408 , n3420 );
and ( n3422 , n186 , n3421 );
not ( n3423 , n3163 );
or ( n3424 , n3423 , n3183 );
nand ( n3425 , n3424 , n3258 );
not ( n3426 , n3384 );
not ( n3427 , n3426 );
not ( n3428 , n3427 );
not ( n3429 , n3102 );
not ( n3430 , n183 );
nor ( n3431 , n3429 , n3430 );
nand ( n3432 , n184 , n3431 );
not ( n3433 , n3432 );
or ( n3434 , n3428 , n3433 );
not ( n3435 , n185 );
nand ( n3436 , n3434 , n3435 );
not ( n3437 , n3013 );
nand ( n3438 , n185 , n3363 );
nand ( n3439 , n183 , n3087 );
not ( n3440 , n3439 );
nand ( n3441 , n3258 , n3440 );
nand ( n3442 , n3438 , n3441 );
not ( n3443 , n3442 );
or ( n3444 , n3437 , n3443 );
not ( n3445 , n185 );
not ( n3446 , n183 );
nand ( n3447 , n3445 , n181 , n3446 );
not ( n3448 , n3447 );
not ( n3449 , n3181 );
or ( n3450 , n3448 , n3449 );
nand ( n3451 , n3450 , n3013 );
nand ( n3452 , n3444 , n3451 );
not ( n3453 , n183 );
nand ( n3454 , n3453 , n3363 );
not ( n3455 , n3454 );
and ( n3456 , n3258 , n3455 );
not ( n3457 , n3375 );
nor ( n3458 , n3452 , n3456 , n3457 );
and ( n3459 , n3425 , n3436 , n3458 );
nor ( n3460 , n3459 , n187 );
nor ( n3461 , n3422 , n3460 );
nand ( n3462 , n3395 , n3461 );
not ( n3463 , n3462 );
not ( n3464 , n3463 );
and ( n3465 , n3274 , n3464 );
not ( n3466 , n3462 );
and ( n3467 , n3273 , n3466 );
nor ( n3468 , n3465 , n3467 );
not ( n3469 , n212 );
not ( n3470 , n209 );
not ( n3471 , n205 );
nor ( n3472 , n3471 , n206 );
nand ( n3473 , n207 , n3472 );
buf ( n3474 , n3473 );
nor ( n3475 , n210 , n3474 );
not ( n3476 , n3475 );
nor ( n3477 , n205 , n206 );
nand ( n3478 , n207 , n3477 );
not ( n3479 , n3478 );
nand ( n3480 , n3479 , n208 );
nand ( n3481 , n206 , n207 );
nor ( n3482 , n3481 , n205 );
nand ( n3483 , n210 , n3482 );
not ( n3484 , n207 );
not ( n3485 , n205 );
nor ( n3486 , n3485 , n206 );
nand ( n3487 , n3484 , n3486 );
not ( n3488 , n3487 );
not ( n3489 , n208 );
nand ( n3490 , n3488 , n3489 );
nand ( n3491 , n3476 , n3480 , n3483 , n3490 );
nand ( n3492 , n3470 , n3491 );
not ( n3493 , n207 );
nand ( n3494 , n3493 , n205 );
not ( n3495 , n3494 );
nand ( n3496 , n208 , n3495 );
nand ( n3497 , n205 , n206 );
not ( n3498 , n3497 );
not ( n3499 , n3498 );
not ( n3500 , n3499 );
nand ( n3501 , n210 , n3500 );
not ( n3502 , n208 );
not ( n3503 , n206 );
nor ( n3504 , n3503 , n207 );
nand ( n3505 , n3502 , n3504 );
nand ( n3506 , n3496 , n3501 , n3505 );
nand ( n3507 , n209 , n3506 );
not ( n3508 , n207 );
nand ( n3509 , n3508 , n3498 );
not ( n3510 , n3509 );
not ( n3511 , n3510 );
nor ( n3512 , n3511 , n208 );
not ( n3513 , n3512 );
not ( n3514 , n3513 );
not ( n3515 , n3514 );
not ( n3516 , n210 );
not ( n3517 , n3497 );
nand ( n3518 , n3517 , n207 );
not ( n3519 , n3518 );
nand ( n3520 , n208 , n3519 );
nor ( n3521 , n3516 , n3520 );
not ( n3522 , n3521 );
nand ( n3523 , n3507 , n3515 , n3522 );
nand ( n3524 , n211 , n3523 );
nand ( n3525 , n3492 , n3524 );
not ( n3526 , n210 );
not ( n3527 , n3480 );
and ( n3528 , n3526 , n3527 );
or ( n3529 , n210 , n3509 );
not ( n3530 , n3529 );
and ( n3531 , n209 , n3530 );
nor ( n3532 , n3528 , n3531 );
not ( n3533 , n3509 );
nand ( n3534 , n3533 , n208 );
not ( n3535 , n3534 );
not ( n3536 , n210 );
nand ( n3537 , n3535 , n3536 );
buf ( n3538 , n3537 );
buf ( n3539 , n3538 );
not ( n3540 , n211 );
not ( n3541 , n210 );
not ( n3542 , n206 );
nor ( n3543 , n3542 , n205 );
not ( n3544 , n3543 );
nor ( n3545 , n3541 , n3544 );
nand ( n3546 , n208 , n3545 );
nand ( n3547 , n3546 , n3490 );
not ( n3548 , n3547 );
not ( n3549 , n3545 );
not ( n3550 , n3549 );
not ( n3551 , n209 );
nand ( n3552 , n3550 , n3551 );
not ( n3553 , n210 );
not ( n3554 , n208 );
and ( n3555 , n3554 , n3482 );
nand ( n3556 , n3553 , n3555 );
nand ( n3557 , n208 , n210 );
not ( n3558 , n3557 );
not ( n3559 , n206 );
nand ( n3560 , n3559 , n207 );
not ( n3561 , n3560 );
nand ( n3562 , n3558 , n3561 );
nand ( n3563 , n3548 , n3552 , n3556 , n3562 );
nand ( n3564 , n3540 , n3563 );
nand ( n3565 , n3532 , n3539 , n3564 );
nor ( n3566 , n3525 , n3565 );
nor ( n3567 , n3469 , n3566 );
not ( n3568 , n3567 );
not ( n3569 , n210 );
nor ( n3570 , n206 , n208 );
nand ( n3571 , n3569 , n3570 );
not ( n3572 , n210 );
nand ( n3573 , n3508 , n3477 );
not ( n3574 , n3573 );
nand ( n3575 , n3572 , n3574 );
and ( n3576 , n3571 , n3575 );
not ( n3577 , n209 );
nor ( n3578 , n3576 , n3577 );
nand ( n3579 , n209 , n210 );
or ( n3580 , n3579 , n3480 );
not ( n3581 , n208 );
nor ( n3582 , n205 , n206 );
nand ( n3583 , n3581 , n3582 );
nor ( n3584 , n210 , n3583 );
not ( n3585 , n3584 );
not ( n3586 , n208 );
nand ( n3587 , n3586 , n3519 );
not ( n3588 , n3587 );
nand ( n3589 , n210 , n3588 );
not ( n3590 , n3589 );
nand ( n3591 , n208 , n3482 );
not ( n3592 , n3591 );
not ( n3593 , n210 );
nand ( n3594 , n3592 , n3593 );
not ( n3595 , n3594 );
or ( n3596 , n3590 , n3595 );
not ( n3597 , n209 );
nand ( n3598 , n3596 , n3597 );
and ( n3599 , n3585 , n3598 );
not ( n3600 , n211 );
not ( n3601 , n3510 );
not ( n3602 , n210 );
nor ( n3603 , n3601 , n3602 );
nand ( n3604 , n209 , n3603 );
not ( n3605 , n3487 );
nand ( n3606 , n3558 , n3605 );
nand ( n3607 , n209 , n3475 );
and ( n3608 , n3604 , n3606 , n3607 );
not ( n3609 , n3487 );
nand ( n3610 , n3609 , n208 );
not ( n3611 , n3610 );
not ( n3612 , n210 );
nand ( n3613 , n3612 , n3512 );
not ( n3614 , n3613 );
or ( n3615 , n3611 , n3614 );
not ( n3616 , n209 );
nand ( n3617 , n3615 , n3616 );
nand ( n3618 , n3608 , n3589 , n3617 );
and ( n3619 , n3600 , n3618 );
not ( n3620 , n3600 );
not ( n3621 , n208 );
nor ( n3622 , n205 , n207 );
nand ( n3623 , n3621 , n3622 );
not ( n3624 , n3623 );
not ( n3625 , n210 );
not ( n3626 , n3496 );
or ( n3627 , n3625 , n3626 );
not ( n3628 , n210 );
not ( n3629 , n3543 );
nand ( n3630 , n3628 , n3629 );
nand ( n3631 , n3627 , n3630 );
not ( n3632 , n3631 );
or ( n3633 , n3624 , n3632 );
not ( n3634 , n209 );
nand ( n3635 , n3633 , n3634 );
not ( n3636 , n210 );
nor ( n3637 , n3636 , n3474 );
not ( n3638 , n3637 );
not ( n3639 , n208 );
buf ( n3640 , n3486 );
nand ( n3641 , n3639 , n3640 );
not ( n3642 , n3641 );
nand ( n3643 , n3642 , n210 );
nand ( n3644 , n3638 , n3643 );
not ( n3645 , n3644 );
not ( n3646 , n208 );
nor ( n3647 , n3646 , n3481 );
not ( n3648 , n3647 );
not ( n3649 , n3648 );
not ( n3650 , n210 );
nand ( n3651 , n3650 , n3519 );
not ( n3652 , n3651 );
or ( n3653 , n3649 , n3652 );
nand ( n3654 , n3653 , n209 );
buf ( n3655 , n3573 );
not ( n3656 , n3655 );
nand ( n3657 , n210 , n3656 );
nand ( n3658 , n3635 , n3645 , n3654 , n3657 );
and ( n3659 , n3620 , n3658 );
nor ( n3660 , n3619 , n3659 );
nand ( n3661 , n3580 , n3599 , n3660 );
or ( n3662 , n3578 , n3661 );
nand ( n3663 , n3662 , n3469 );
not ( n3664 , n211 );
not ( n3665 , n3664 );
not ( n3666 , n209 );
not ( n3667 , n3666 );
nand ( n3668 , n206 , n207 );
nor ( n3669 , n208 , n3668 );
nand ( n3670 , n210 , n3669 );
not ( n3671 , n3670 );
not ( n3672 , n3671 );
not ( n3673 , n3487 );
nand ( n3674 , n3673 , n210 );
not ( n3675 , n3573 );
nand ( n3676 , n208 , n3675 );
not ( n3677 , n3676 );
not ( n3678 , n210 );
nand ( n3679 , n3677 , n3678 );
nand ( n3680 , n3672 , n3674 , n3679 );
not ( n3681 , n3680 );
or ( n3682 , n3667 , n3681 );
nor ( n3683 , n3542 , n205 );
and ( n3684 , n3508 , n3683 );
nand ( n3685 , n208 , n3684 );
not ( n3686 , n3685 );
nand ( n3687 , n3686 , n210 );
not ( n3688 , n210 );
nor ( n3689 , n3688 , n3480 );
not ( n3690 , n3689 );
and ( n3691 , n3687 , n3690 );
nand ( n3692 , n3682 , n3691 );
not ( n3693 , n3692 );
or ( n3694 , n3665 , n3693 );
not ( n3695 , n211 );
and ( n3696 , n209 , n3695 );
nand ( n3697 , n3508 , n3683 );
not ( n3698 , n3697 );
not ( n3699 , n3698 );
or ( n3700 , n210 , n3699 );
not ( n3701 , n210 );
not ( n3702 , n3520 );
nand ( n3703 , n3701 , n3702 );
nand ( n3704 , n3700 , n3585 , n3703 );
nand ( n3705 , n3696 , n3704 );
nand ( n3706 , n3694 , n3705 );
not ( n3707 , n3538 );
nand ( n3708 , n205 , n207 );
not ( n3709 , n3708 );
nand ( n3710 , n208 , n3709 );
not ( n3711 , n3710 );
not ( n3712 , n3513 );
or ( n3713 , n3711 , n3712 );
nand ( n3714 , n3713 , n210 );
not ( n3715 , n3714 );
or ( n3716 , n3707 , n3715 );
and ( n3717 , n209 , n211 );
nand ( n3718 , n3716 , n3717 );
not ( n3719 , n209 );
not ( n3720 , n210 );
not ( n3721 , n207 );
nor ( n3722 , n3721 , n208 , n205 );
nand ( n3723 , n3720 , n3722 );
not ( n3724 , n210 );
not ( n3725 , n3478 );
nand ( n3726 , n3724 , n3725 );
not ( n3727 , n208 );
not ( n3728 , n3474 );
nand ( n3729 , n3727 , n3728 );
nor ( n3730 , n205 , n207 );
nand ( n3731 , n3730 , n3570 );
nand ( n3732 , n3723 , n3726 , n3729 , n3731 );
and ( n3733 , n211 , n3719 , n3732 );
nor ( n3734 , n3579 , n3731 );
not ( n3735 , n3734 );
not ( n3736 , n3735 );
nor ( n3737 , n3733 , n3736 );
not ( n3738 , n209 );
nand ( n3739 , n3738 , n3656 );
not ( n3740 , n3739 );
and ( n3741 , n210 , n211 );
nand ( n3742 , n3740 , n3741 );
not ( n3743 , n209 );
or ( n3744 , n3743 , n3687 );
nand ( n3745 , n3718 , n3737 , n3742 , n3744 );
nor ( n3746 , n3706 , n3745 );
nand ( n3747 , n3568 , n3663 , n3746 );
not ( n3748 , n3747 );
not ( n3749 , n3748 );
not ( n3750 , n201 );
not ( n3751 , n197 );
nand ( n3752 , n3751 , n200 );
not ( n3753 , n3752 );
not ( n3754 , n3753 );
nor ( n3755 , n3750 , n3754 );
nand ( n3756 , n199 , n3755 );
not ( n3757 , n3756 );
not ( n3758 , n199 );
not ( n3759 , n198 );
not ( n3760 , n197 );
nor ( n3761 , n3760 , n200 );
nand ( n3762 , n3759 , n3761 );
not ( n3763 , n3762 );
nand ( n3764 , n3758 , n3763 );
not ( n3765 , n3764 );
nor ( n3766 , n3757 , n3765 );
not ( n3767 , n201 );
nand ( n3768 , n198 , n3753 );
not ( n3769 , n3768 );
nand ( n3770 , n3758 , n3769 );
not ( n3771 , n3770 );
nand ( n3772 , n3767 , n3771 );
not ( n3773 , n202 );
and ( n3774 , n3773 , n3755 );
nand ( n3775 , n199 , n201 );
not ( n3776 , n3775 );
not ( n3777 , n198 );
nor ( n3778 , n3777 , n200 );
and ( n3779 , n3776 , n3778 );
nor ( n3780 , n3774 , n3779 );
and ( n3781 , n3766 , n3772 , n3780 );
nor ( n3782 , n3781 , n203 );
not ( n3783 , n3782 );
not ( n3784 , n202 );
not ( n3785 , n3769 );
not ( n3786 , n3785 );
nand ( n3787 , n201 , n3786 );
not ( n3788 , n201 );
nand ( n3789 , n198 , n3761 );
not ( n3790 , n3789 );
nand ( n3791 , n3788 , n3790 );
nor ( n3792 , n197 , n200 );
nand ( n3793 , n198 , n3792 );
nor ( n3794 , n3758 , n3793 );
not ( n3795 , n3794 );
nand ( n3796 , n3787 , n3791 , n3795 , n3764 );
nand ( n3797 , n3784 , n3796 );
not ( n3798 , n201 );
nand ( n3799 , n197 , n200 );
nor ( n3800 , n198 , n3799 );
nand ( n3801 , n3798 , n3800 );
not ( n3802 , n3801 );
nand ( n3803 , n202 , n3802 );
not ( n3804 , n201 );
nand ( n3805 , n199 , n3800 );
not ( n3806 , n3805 );
nand ( n3807 , n3804 , n3806 );
not ( n3808 , n201 );
nand ( n3809 , n3808 , n3794 );
and ( n3810 , n3803 , n3807 , n3809 );
nand ( n3811 , n197 , n200 );
nor ( n3812 , n198 , n3811 );
and ( n3813 , n3758 , n3812 );
not ( n3814 , n3813 );
not ( n3815 , n3814 );
not ( n3816 , n198 );
nor ( n3817 , n3816 , n3799 );
nand ( n3818 , n199 , n3817 );
not ( n3819 , n3818 );
nand ( n3820 , n3819 , n201 );
not ( n3821 , n3820 );
or ( n3822 , n3815 , n3821 );
nand ( n3823 , n3822 , n203 );
nand ( n3824 , n202 , n203 );
not ( n3825 , n3824 );
not ( n3826 , n200 );
nor ( n3827 , n3826 , n198 );
nand ( n3828 , n3758 , n3827 );
not ( n3829 , n201 );
nor ( n3830 , n3829 , n3811 );
not ( n3831 , n3830 );
not ( n3832 , n198 );
nand ( n3833 , n3832 , n197 );
not ( n3834 , n3833 );
nand ( n3835 , n3834 , n199 );
nand ( n3836 , n3828 , n3831 , n3835 );
nand ( n3837 , n3825 , n3836 );
and ( n3838 , n3810 , n3823 , n3837 );
nand ( n3839 , n3783 , n3797 , n3838 );
nand ( n3840 , n204 , n3839 );
not ( n3841 , n3824 );
nand ( n3842 , n197 , n198 );
not ( n3843 , n3842 );
and ( n3844 , n199 , n3843 );
and ( n3845 , n201 , n3844 );
not ( n3846 , n3807 );
not ( n3847 , n201 );
nor ( n3848 , n3847 , n3814 );
nor ( n3849 , n3845 , n3846 , n3848 );
not ( n3850 , n3849 );
and ( n3851 , n3841 , n3850 );
not ( n3852 , n203 );
nand ( n3853 , n202 , n3852 );
not ( n3854 , n3853 );
nand ( n3855 , n3753 , n3759 );
buf ( n3856 , n3855 );
not ( n3857 , n3856 );
not ( n3858 , n3857 );
or ( n3859 , n201 , n3858 );
nor ( n3860 , n199 , n201 );
not ( n3861 , n3860 );
buf ( n3862 , n3792 );
not ( n3863 , n3862 );
nor ( n3864 , n3861 , n3863 );
not ( n3865 , n3864 );
not ( n3866 , n3818 );
not ( n3867 , n201 );
nand ( n3868 , n3866 , n3867 );
nand ( n3869 , n3859 , n3865 , n3868 );
and ( n3870 , n3854 , n3869 );
nor ( n3871 , n3851 , n3870 );
not ( n3872 , n3776 );
nor ( n3873 , n3872 , n3856 );
nand ( n3874 , n201 , n3794 );
not ( n3875 , n3874 );
or ( n3876 , n3873 , n3875 );
not ( n3877 , n203 );
nand ( n3878 , n3876 , n3877 );
not ( n3879 , n203 );
nor ( n3880 , n3879 , n202 );
nand ( n3881 , n3758 , n3790 );
nor ( n3882 , n201 , n3793 );
not ( n3883 , n3882 );
not ( n3884 , n201 );
not ( n3885 , n197 );
nand ( n3886 , n3885 , n198 );
nor ( n3887 , n199 , n3886 );
nand ( n3888 , n3884 , n3887 );
not ( n3889 , n197 );
nor ( n3890 , n198 , n200 );
nand ( n3891 , n3889 , n3890 );
not ( n3892 , n3891 );
and ( n3893 , n3758 , n3892 );
not ( n3894 , n3893 );
nand ( n3895 , n3881 , n3883 , n3888 , n3894 );
nand ( n3896 , n3880 , n3895 );
and ( n3897 , n201 , n202 );
not ( n3898 , n3897 );
nand ( n3899 , n199 , n3857 );
or ( n3900 , n3898 , n3899 );
nand ( n3901 , n3897 , n3893 );
and ( n3902 , n3900 , n3901 );
not ( n3903 , n201 );
nor ( n3904 , n3903 , n202 );
and ( n3905 , n203 , n3904 , n3892 );
nor ( n3906 , n202 , n203 );
not ( n3907 , n201 );
nand ( n3908 , n3907 , n199 );
not ( n3909 , n3908 );
nand ( n3910 , n3909 , n3892 );
nand ( n3911 , n198 , n200 );
nor ( n3912 , n199 , n3911 );
nand ( n3913 , n201 , n3912 );
not ( n3914 , n3762 );
nand ( n3915 , n201 , n3914 );
not ( n3916 , n3915 );
not ( n3917 , n3916 );
nand ( n3918 , n3910 , n3913 , n3917 );
and ( n3919 , n3906 , n3918 );
nor ( n3920 , n3905 , n3919 );
and ( n3921 , n3878 , n3896 , n3902 , n3920 );
not ( n3922 , n3817 );
not ( n3923 , n3922 );
nand ( n3924 , n3923 , n3758 );
not ( n3925 , n3924 );
nand ( n3926 , n201 , n3925 );
not ( n3927 , n3926 );
not ( n3928 , n3768 );
nand ( n3929 , n3928 , n199 );
not ( n3930 , n3929 );
not ( n3931 , n201 );
nand ( n3932 , n3930 , n3931 );
not ( n3933 , n3932 );
or ( n3934 , n3927 , n3933 );
not ( n3935 , n202 );
nand ( n3936 , n3934 , n3935 );
not ( n3937 , n203 );
not ( n3938 , n3762 );
nand ( n3939 , n199 , n3938 );
not ( n3940 , n3939 );
not ( n3941 , n3860 );
not ( n3942 , n3941 );
nand ( n3943 , n3942 , n3812 );
not ( n3944 , n3943 );
or ( n3945 , n3940 , n3944 );
not ( n3946 , n202 );
nand ( n3947 , n3945 , n3946 );
nand ( n3948 , n3776 , n3763 );
nand ( n3949 , n3947 , n3926 , n3948 );
nand ( n3950 , n3937 , n3949 );
nand ( n3951 , n3936 , n3950 );
not ( n3952 , n199 );
nor ( n3953 , n197 , n198 );
nand ( n3954 , n3952 , n3953 );
not ( n3955 , n3954 );
and ( n3956 , n201 , n3835 );
not ( n3957 , n201 );
not ( n3958 , n3753 );
and ( n3959 , n3957 , n3958 );
or ( n3960 , n3956 , n3959 );
not ( n3961 , n3960 );
or ( n3962 , n3955 , n3961 );
not ( n3963 , n202 );
nand ( n3964 , n3962 , n3963 );
nand ( n3965 , n201 , n3892 );
not ( n3966 , n3789 );
nand ( n3967 , n201 , n3966 );
not ( n3968 , n200 );
and ( n3969 , n197 , n3968 );
not ( n3970 , n3969 );
nor ( n3971 , n199 , n3970 );
nand ( n3972 , n201 , n3971 );
and ( n3973 , n3967 , n3972 );
nand ( n3974 , n3964 , n3965 , n3973 );
nand ( n3975 , n203 , n3974 );
nor ( n3976 , n3758 , n3911 );
not ( n3977 , n3976 );
not ( n3978 , n201 );
not ( n3979 , n3922 );
nand ( n3980 , n3978 , n3979 );
nand ( n3981 , n3977 , n3980 );
and ( n3982 , n3825 , n3981 );
not ( n3983 , n201 );
not ( n3984 , n3983 );
nor ( n3985 , n199 , n200 );
not ( n3986 , n3985 );
or ( n3987 , n3984 , n3986 );
not ( n3988 , n201 );
nand ( n3989 , n3988 , n3892 );
nand ( n3990 , n3987 , n3989 );
and ( n3991 , n202 , n3990 );
nor ( n3992 , n3982 , n3991 );
not ( n3993 , n203 );
not ( n3994 , n202 );
nand ( n3995 , n201 , n3812 );
or ( n3996 , n3994 , n3995 );
not ( n3997 , n201 );
nand ( n3998 , n3997 , n202 );
not ( n3999 , n3998 );
nand ( n4000 , n3999 , n3790 );
nand ( n4001 , n3996 , n4000 );
nand ( n4002 , n3993 , n4001 );
not ( n4003 , n3874 );
nand ( n4004 , n4003 , n202 );
and ( n4005 , n4002 , n3865 , n4004 );
nand ( n4006 , n3975 , n3992 , n4005 );
or ( n4007 , n3951 , n4006 );
not ( n4008 , n204 );
nand ( n4009 , n4007 , n4008 );
nand ( n4010 , n3840 , n3871 , n3921 , n4009 );
not ( n4011 , n4010 );
not ( n4012 , n4011 );
or ( n4013 , n3749 , n4012 );
nand ( n4014 , n3747 , n4010 );
nand ( n4015 , n4013 , n4014 );
and ( n4016 , n3468 , n4015 );
not ( n4017 , n3468 );
not ( n4018 , n4015 );
and ( n4019 , n4017 , n4018 );
nor ( n4020 , n4016 , n4019 );
not ( n4021 , n4020 );
or ( n4022 , n3000 , n4021 );
nor ( n4023 , n2999 , n4020 );
nor ( n4024 , n4023 , n1 );
nand ( n4025 , n4022 , n4024 );
nand ( n4026 , n2362 , n4025 );
xnor ( n4027 , n386 , n387 );
or ( n4028 , n2352 , n4027 );
not ( n4029 , n161 );
not ( n4030 , n157 );
nand ( n4031 , n4030 , n155 );
not ( n4032 , n4031 );
not ( n4033 , n154 );
nand ( n4034 , n4032 , n4033 );
not ( n4035 , n4034 );
nand ( n4036 , n158 , n4035 );
nand ( n4037 , n155 , n157 );
nor ( n4038 , n4037 , n156 );
not ( n4039 , n4038 );
not ( n4040 , n4039 );
nand ( n4041 , n4040 , n158 );
nor ( n4042 , n154 , n158 );
not ( n4043 , n4042 );
not ( n4044 , n4043 );
not ( n4045 , n156 );
nor ( n4046 , n155 , n157 );
and ( n4047 , n4045 , n4046 );
not ( n4048 , n4047 );
not ( n4049 , n4048 );
nand ( n4050 , n4044 , n4049 );
and ( n4051 , n4036 , n4041 , n4050 );
nor ( n4052 , n4051 , n159 );
not ( n4053 , n4052 );
not ( n4054 , n160 );
not ( n4055 , n159 );
not ( n4056 , n154 );
nand ( n4057 , n156 , n157 );
not ( n4058 , n4057 );
nand ( n4059 , n4056 , n4058 );
not ( n4060 , n4059 );
and ( n4061 , n4055 , n4060 );
and ( n4062 , n158 , n4058 );
nand ( n4063 , n154 , n158 );
not ( n4064 , n4063 );
nor ( n4065 , n155 , n157 );
buf ( n4066 , n4065 );
nand ( n4067 , n4064 , n4066 );
nor ( n4068 , n159 , n4067 );
nor ( n4069 , n4061 , n4062 , n4068 );
not ( n4070 , n4037 );
not ( n4071 , n4070 );
nor ( n4072 , n154 , n4071 );
nand ( n4073 , n158 , n4072 );
not ( n4074 , n155 );
nand ( n4075 , n157 , n4074 );
not ( n4076 , n4075 );
nand ( n4077 , n4076 , n156 );
not ( n4078 , n4077 );
nand ( n4079 , n4078 , n154 );
not ( n4080 , n4079 );
nand ( n4081 , n159 , n4080 );
nand ( n4082 , n4069 , n4073 , n4081 );
and ( n4083 , n4054 , n4082 );
not ( n4084 , n4054 );
nand ( n4085 , n154 , n4047 );
nor ( n4086 , n158 , n4085 );
not ( n4087 , n4086 );
nand ( n4088 , n157 , n4074 );
not ( n4089 , n4088 );
not ( n4090 , n4089 );
nor ( n4091 , n154 , n4090 );
nand ( n4092 , n159 , n4091 );
not ( n4093 , n4035 );
not ( n4094 , n4093 );
not ( n4095 , n154 );
not ( n4096 , n4088 );
not ( n4097 , n156 );
nand ( n4098 , n4096 , n4097 );
nor ( n4099 , n4095 , n4098 );
not ( n4100 , n4099 );
not ( n4101 , n4100 );
or ( n4102 , n4094 , n4101 );
not ( n4103 , n159 );
nand ( n4104 , n4102 , n4103 );
not ( n4105 , n154 );
nand ( n4106 , n156 , n4065 );
not ( n4107 , n4106 );
nand ( n4108 , n4105 , n4107 );
not ( n4109 , n4108 );
nand ( n4110 , n158 , n4109 );
nand ( n4111 , n4087 , n4092 , n4104 , n4110 );
and ( n4112 , n4084 , n4111 );
nor ( n4113 , n4083 , n4112 );
not ( n4114 , n154 );
nor ( n4115 , n4114 , n158 );
not ( n4116 , n4115 );
or ( n4117 , n157 , n4116 );
not ( n4118 , n4037 );
nand ( n4119 , n4118 , n156 );
not ( n4120 , n4119 );
not ( n4121 , n154 );
nand ( n4122 , n4120 , n4121 );
not ( n4123 , n4122 );
not ( n4124 , n4123 );
nand ( n4125 , n4117 , n4124 );
nand ( n4126 , n159 , n4125 );
not ( n4127 , n154 );
nand ( n4128 , n4127 , n158 );
not ( n4129 , n4128 );
buf ( n4130 , n4129 );
not ( n4131 , n4130 );
or ( n4132 , n155 , n4131 );
not ( n4133 , n158 );
not ( n4134 , n4075 );
not ( n4135 , n156 );
nand ( n4136 , n4134 , n4135 );
nor ( n4137 , n4133 , n4136 );
not ( n4138 , n4137 );
nand ( n4139 , n4132 , n4138 );
nand ( n4140 , n159 , n4139 );
nand ( n4141 , n4053 , n4113 , n4126 , n4140 );
not ( n4142 , n4141 );
or ( n4143 , n4029 , n4142 );
not ( n4144 , n161 );
not ( n4145 , n158 );
not ( n4146 , n159 );
nand ( n4147 , n4145 , n4146 );
not ( n4148 , n4147 );
and ( n4149 , n154 , n4038 );
nand ( n4150 , n4148 , n4149 );
not ( n4151 , n4107 );
or ( n4152 , n4043 , n4151 );
nand ( n4153 , n155 , n156 );
nor ( n4154 , n157 , n4153 );
and ( n4155 , n4148 , n4154 );
not ( n4156 , n154 );
nand ( n4157 , n155 , n156 );
nor ( n4158 , n4156 , n4157 );
and ( n4159 , n159 , n4158 );
nor ( n4160 , n4155 , n4159 );
not ( n4161 , n158 );
not ( n4162 , n154 );
nand ( n4163 , n4162 , n4066 );
nor ( n4164 , n4161 , n4163 );
not ( n4165 , n4164 );
nand ( n4166 , n159 , n4049 );
nand ( n4167 , n4160 , n4165 , n4166 );
nand ( n4168 , n4054 , n4167 );
and ( n4169 , n4150 , n4152 , n4168 );
not ( n4170 , n154 );
not ( n4171 , n156 );
nand ( n4172 , n4171 , n155 );
not ( n4173 , n4172 );
nand ( n4174 , n4170 , n4173 );
or ( n4175 , n158 , n4174 );
nand ( n4176 , n4064 , n4049 );
nand ( n4177 , n4175 , n4176 );
nand ( n4178 , n159 , n4177 );
not ( n4179 , n159 );
not ( n4180 , n4179 );
not ( n4181 , n158 );
not ( n4182 , n4078 );
not ( n4183 , n4182 );
nand ( n4184 , n4181 , n4183 );
nor ( n4185 , n154 , n4098 );
not ( n4186 , n4185 );
nand ( n4187 , n4184 , n4079 , n4186 );
not ( n4188 , n4187 );
or ( n4189 , n4180 , n4188 );
not ( n4190 , n156 );
nand ( n4191 , n4190 , n157 );
not ( n4192 , n4191 );
nand ( n4193 , n154 , n4192 );
not ( n4194 , n4193 );
not ( n4195 , n159 );
nor ( n4196 , n4195 , n158 );
not ( n4197 , n4196 );
not ( n4198 , n4197 );
nand ( n4199 , n4194 , n4198 );
nand ( n4200 , n4189 , n4199 );
nand ( n4201 , n159 , n4154 );
not ( n4202 , n4031 );
not ( n4203 , n4202 );
not ( n4204 , n154 );
nor ( n4205 , n4203 , n4204 );
not ( n4206 , n4205 );
not ( n4207 , n4206 );
nand ( n4208 , n158 , n4207 );
nand ( n4209 , n4201 , n4208 );
or ( n4210 , n4200 , n4209 );
nand ( n4211 , n4210 , n160 );
nand ( n4212 , n4169 , n4178 , n4211 );
and ( n4213 , n4144 , n4212 );
not ( n4214 , n159 );
not ( n4215 , n4031 );
not ( n4216 , n156 );
nand ( n4217 , n4215 , n4216 );
not ( n4218 , n4217 );
not ( n4219 , n154 );
nand ( n4220 , n4218 , n4219 );
not ( n4221 , n4220 );
nand ( n4222 , n158 , n4221 );
not ( n4223 , n4222 );
and ( n4224 , n4214 , n4223 );
nand ( n4225 , n158 , n159 );
not ( n4226 , n4225 );
not ( n4227 , n4158 );
not ( n4228 , n4227 );
and ( n4229 , n4226 , n4228 );
nor ( n4230 , n4224 , n4229 );
not ( n4231 , n4205 );
nor ( n4232 , n4231 , n158 );
nand ( n4233 , n159 , n4232 );
not ( n4234 , n158 );
not ( n4235 , n4107 );
nor ( n4236 , n4234 , n4235 );
nand ( n4237 , n159 , n4236 );
nand ( n4238 , n158 , n4185 );
and ( n4239 , n4233 , n4237 , n4238 );
not ( n4240 , n158 );
not ( n4241 , n4149 );
nor ( n4242 , n4240 , n4241 );
not ( n4243 , n4242 );
not ( n4244 , n159 );
nor ( n4245 , n4173 , n4192 );
not ( n4246 , n4245 );
nand ( n4247 , n4246 , n158 );
not ( n4248 , n158 );
nand ( n4249 , n4248 , n4123 );
nand ( n4250 , n4247 , n4249 , n4050 );
nand ( n4251 , n4244 , n4250 );
nand ( n4252 , n4239 , n4243 , n4251 );
and ( n4253 , n160 , n4252 );
not ( n4254 , n160 );
nor ( n4255 , n157 , n4153 );
nand ( n4256 , n154 , n4255 );
buf ( n4257 , n4256 );
not ( n4258 , n4257 );
nand ( n4259 , n4258 , n158 );
nand ( n4260 , n4259 , n4152 );
not ( n4261 , n4260 );
not ( n4262 , n159 );
not ( n4263 , n158 );
nor ( n4264 , n4263 , n4122 );
not ( n4265 , n4264 );
not ( n4266 , n158 );
not ( n4267 , n154 );
nor ( n4268 , n4267 , n4172 );
nand ( n4269 , n4266 , n4268 );
not ( n4270 , n4039 );
not ( n4271 , n158 );
nand ( n4272 , n4270 , n4271 );
nand ( n4273 , n4265 , n4269 , n4272 );
nand ( n4274 , n4262 , n4273 );
nor ( n4275 , n158 , n4151 );
not ( n4276 , n4275 );
not ( n4277 , n4063 );
not ( n4278 , n4042 );
not ( n4279 , n4278 );
or ( n4280 , n4277 , n4279 );
not ( n4281 , n4098 );
nand ( n4282 , n4280 , n4281 );
nand ( n4283 , n158 , n4154 );
not ( n4284 , n156 );
nor ( n4285 , n4284 , n155 );
not ( n4286 , n4285 );
nor ( n4287 , n154 , n4286 );
nand ( n4288 , n158 , n4287 );
nand ( n4289 , n4276 , n4282 , n4283 , n4288 );
nand ( n4290 , n4289 , n159 );
nand ( n4291 , n4261 , n4274 , n4290 );
and ( n4292 , n4254 , n4291 );
nor ( n4293 , n4253 , n4292 );
nand ( n4294 , n4230 , n4293 );
nor ( n4295 , n4213 , n4294 );
nand ( n4296 , n4143 , n4295 );
not ( n4297 , n4296 );
not ( n4298 , n4297 );
and ( n4299 , n386 , n4298 );
not ( n4300 , n386 );
not ( n4301 , n4296 );
and ( n4302 , n4300 , n4301 );
nor ( n4303 , n4299 , n4302 );
not ( n4304 , n4303 );
nand ( n4305 , n147 , n151 );
not ( n4306 , n4305 );
nand ( n4307 , n150 , n4306 );
not ( n4308 , n4307 );
not ( n4309 , n149 );
nand ( n4310 , n150 , n4309 );
nor ( n4311 , n146 , n151 );
nand ( n4312 , n148 , n4311 );
nor ( n4313 , n4310 , n4312 );
nor ( n4314 , n4308 , n4313 );
not ( n4315 , n149 );
not ( n4316 , n148 );
nand ( n4317 , n4316 , n4306 );
not ( n4318 , n4317 );
nand ( n4319 , n4315 , n4318 );
nand ( n4320 , n146 , n151 );
nor ( n4321 , n148 , n4320 );
nand ( n4322 , n150 , n4321 );
not ( n4323 , n146 );
nand ( n4324 , n4323 , n151 );
not ( n4325 , n4324 );
nand ( n4326 , n4325 , n147 );
not ( n4327 , n4326 );
nand ( n4328 , n4327 , n148 );
not ( n4329 , n4328 );
nand ( n4330 , n149 , n4329 );
and ( n4331 , n4314 , n4319 , n4322 , n4330 );
or ( n4332 , n152 , n4331 );
not ( n4333 , n151 );
not ( n4334 , n148 );
nor ( n4335 , n4334 , n150 );
buf ( n4336 , n4335 );
and ( n4337 , n4333 , n4336 );
not ( n4338 , n148 );
not ( n4339 , n150 );
nor ( n4340 , n4339 , n146 );
and ( n4341 , n4338 , n4340 );
nor ( n4342 , n4337 , n4341 );
not ( n4343 , n4320 );
nand ( n4344 , n4343 , n147 );
not ( n4345 , n4344 );
not ( n4346 , n148 );
nand ( n4347 , n4345 , n4346 );
not ( n4348 , n4347 );
not ( n4349 , n4348 );
not ( n4350 , n147 );
nand ( n4351 , n4350 , n4325 );
not ( n4352 , n4351 );
and ( n4353 , n150 , n4352 );
not ( n4354 , n4353 );
nand ( n4355 , n4342 , n4349 , n4354 );
nand ( n4356 , n149 , n4355 );
nand ( n4357 , n4332 , n4356 );
not ( n4358 , n152 );
not ( n4359 , n149 );
not ( n4360 , n151 );
nand ( n4361 , n146 , n4360 );
nor ( n4362 , n148 , n4361 );
not ( n4363 , n4362 );
not ( n4364 , n4351 );
nand ( n4365 , n4364 , n148 );
nand ( n4366 , n4363 , n4365 );
and ( n4367 , n4359 , n4366 );
not ( n4368 , n4325 );
nor ( n4369 , n148 , n4368 );
nand ( n4370 , n149 , n4369 );
not ( n4371 , n4370 );
nor ( n4372 , n4367 , n4371 );
nor ( n4373 , n146 , n151 );
and ( n4374 , n147 , n4373 );
not ( n4375 , n4374 );
not ( n4376 , n4375 );
not ( n4377 , n148 );
nand ( n4378 , n4376 , n4377 );
not ( n4379 , n4378 );
nand ( n4380 , n150 , n4379 );
not ( n4381 , n147 );
nand ( n4382 , n4381 , n4373 );
not ( n4383 , n4382 );
nand ( n4384 , n148 , n4383 );
nor ( n4385 , n150 , n4384 );
not ( n4386 , n4385 );
nand ( n4387 , n4372 , n4380 , n4386 );
not ( n4388 , n4387 );
or ( n4389 , n4358 , n4388 );
not ( n4390 , n149 );
buf ( n4391 , n4382 );
not ( n4392 , n4391 );
nor ( n4393 , n148 , n150 );
nand ( n4394 , n4392 , n4393 );
nand ( n4395 , n146 , n151 );
not ( n4396 , n4395 );
nand ( n4397 , n4396 , n4350 );
not ( n4398 , n4397 );
nand ( n4399 , n150 , n4398 );
nand ( n4400 , n150 , n4362 );
nand ( n4401 , n4394 , n4399 , n4400 );
nand ( n4402 , n4390 , n4401 );
nand ( n4403 , n4389 , n4402 );
nor ( n4404 , n4357 , n4403 );
not ( n4405 , n153 );
nor ( n4406 , n4404 , n4405 );
not ( n4407 , n4406 );
not ( n4408 , n4361 );
nand ( n4409 , n148 , n4408 );
not ( n4410 , n4409 );
not ( n4411 , n150 );
nand ( n4412 , n4410 , n4411 );
not ( n4413 , n4412 );
nand ( n4414 , n4413 , n149 );
not ( n4415 , n4374 );
not ( n4416 , n4415 );
and ( n4417 , n150 , n4416 );
nand ( n4418 , n149 , n4417 );
buf ( n4419 , n4351 );
not ( n4420 , n4419 );
not ( n4421 , n148 );
nand ( n4422 , n4420 , n4421 );
not ( n4423 , n4422 );
nand ( n4424 , n150 , n4423 );
and ( n4425 , n4414 , n4418 , n4424 );
not ( n4426 , n149 );
not ( n4427 , n4426 );
not ( n4428 , n150 );
not ( n4429 , n147 );
nand ( n4430 , n4429 , n146 );
not ( n4431 , n151 );
nor ( n4432 , n4431 , n147 );
not ( n4433 , n4432 );
nand ( n4434 , n4430 , n4433 );
not ( n4435 , n4434 );
or ( n4436 , n4428 , n4435 );
not ( n4437 , n150 );
nand ( n4438 , n4437 , n4348 );
nand ( n4439 , n4436 , n4438 , n4394 );
not ( n4440 , n4439 );
or ( n4441 , n4427 , n4440 );
nand ( n4442 , n148 , n4398 );
not ( n4443 , n4442 );
nand ( n4444 , n4443 , n150 );
nand ( n4445 , n4441 , n4444 );
not ( n4446 , n4445 );
nand ( n4447 , n4425 , n4446 );
and ( n4448 , n152 , n4447 );
not ( n4449 , n148 );
not ( n4450 , n151 );
nand ( n4451 , n4450 , n146 );
not ( n4452 , n4451 );
nand ( n4453 , n4350 , n4452 );
not ( n4454 , n4453 );
nand ( n4455 , n4449 , n4454 );
not ( n4456 , n4455 );
nand ( n4457 , n150 , n4456 );
or ( n4458 , n149 , n4457 );
nand ( n4459 , n149 , n150 );
not ( n4460 , n4459 );
not ( n4461 , n4460 );
not ( n4462 , n4461 );
not ( n4463 , n4462 );
nand ( n4464 , n146 , n147 );
not ( n4465 , n4464 );
nand ( n4466 , n4465 , n148 );
not ( n4467 , n4466 );
not ( n4468 , n4467 );
or ( n4469 , n4463 , n4468 );
nand ( n4470 , n4458 , n4469 );
nor ( n4471 , n4448 , n4470 );
not ( n4472 , n149 );
nand ( n4473 , n147 , n4452 );
or ( n4474 , n4472 , n4473 );
not ( n4475 , n4474 );
not ( n4476 , n150 );
nor ( n4477 , n4476 , n4409 );
nor ( n4478 , n4475 , n4477 );
not ( n4479 , n149 );
nor ( n4480 , n4479 , n150 );
nand ( n4481 , n148 , n4432 );
not ( n4482 , n4481 );
nand ( n4483 , n4480 , n4482 );
not ( n4484 , n149 );
not ( n4485 , n150 );
not ( n4486 , n4326 );
nand ( n4487 , n4485 , n4486 );
not ( n4488 , n4329 );
nand ( n4489 , n4487 , n4488 , n4422 );
nand ( n4490 , n4484 , n4489 );
nand ( n4491 , n4478 , n4483 , n4490 );
nand ( n4492 , n152 , n4491 );
not ( n4493 , n4492 );
not ( n4494 , n149 );
not ( n4495 , n150 );
not ( n4496 , n4495 );
not ( n4497 , n148 );
not ( n4498 , n4430 );
nand ( n4499 , n4497 , n4498 );
not ( n4500 , n4499 );
not ( n4501 , n4500 );
or ( n4502 , n4496 , n4501 );
not ( n4503 , n4384 );
nand ( n4504 , n4503 , n150 );
nand ( n4505 , n4502 , n4504 );
not ( n4506 , n4505 );
or ( n4507 , n4494 , n4506 );
not ( n4508 , n4375 );
nand ( n4509 , n4508 , n4393 );
nand ( n4510 , n4507 , n4509 );
not ( n4511 , n4391 );
nand ( n4512 , n149 , n4511 );
not ( n4513 , n148 );
and ( n4514 , n4513 , n4311 );
nand ( n4515 , n150 , n4514 );
nand ( n4516 , n4512 , n4515 );
and ( n4517 , n149 , n4468 );
not ( n4518 , n149 );
nor ( n4519 , n150 , n4473 );
not ( n4520 , n4519 );
and ( n4521 , n4518 , n4520 );
nor ( n4522 , n4517 , n4521 );
nor ( n4523 , n4516 , n4522 );
or ( n4524 , n4523 , n152 );
nand ( n4525 , n4336 , n4398 );
or ( n4526 , n149 , n4525 );
nand ( n4527 , n4524 , n4526 );
nor ( n4528 , n4510 , n4527 );
not ( n4529 , n4528 );
or ( n4530 , n4493 , n4529 );
nand ( n4531 , n4530 , n4405 );
not ( n4532 , n152 );
nand ( n4533 , n147 , n4452 );
not ( n4534 , n148 );
nor ( n4535 , n4533 , n4534 );
nand ( n4536 , n150 , n4535 );
and ( n4537 , n4536 , n4509 );
not ( n4538 , n149 );
not ( n4539 , n148 );
nor ( n4540 , n4539 , n4430 );
not ( n4541 , n4540 );
or ( n4542 , n150 , n4541 );
not ( n4543 , n150 );
nand ( n4544 , n4543 , n4398 );
not ( n4545 , n4544 );
not ( n4546 , n4545 );
not ( n4547 , n4347 );
nand ( n4548 , n150 , n4547 );
nand ( n4549 , n4542 , n4546 , n4548 );
nand ( n4550 , n4538 , n4549 );
not ( n4551 , n148 );
not ( n4552 , n147 );
nor ( n4553 , n4552 , n146 );
nand ( n4554 , n4551 , n4553 );
not ( n4555 , n4554 );
nand ( n4556 , n150 , n4555 );
not ( n4557 , n4375 );
not ( n4558 , n150 );
nand ( n4559 , n4557 , n4558 );
nand ( n4560 , n4556 , n4559 );
not ( n4561 , n4533 );
nand ( n4562 , n150 , n4561 );
not ( n4563 , n4365 );
nand ( n4564 , n150 , n4563 );
not ( n4565 , n4419 );
nand ( n4566 , n4565 , n4393 );
nand ( n4567 , n4562 , n4564 , n4566 );
or ( n4568 , n4560 , n4567 );
nand ( n4569 , n4568 , n149 );
nand ( n4570 , n4537 , n4550 , n4569 );
nand ( n4571 , n4532 , n4570 );
nand ( n4572 , n4407 , n4471 , n4531 , n4571 );
not ( n4573 , n177 );
not ( n4574 , n174 );
nor ( n4575 , n4574 , n171 );
and ( n4576 , n4575 , n175 );
nand ( n4577 , n4576 , n173 );
not ( n4578 , n4577 );
nand ( n4579 , n172 , n4578 );
not ( n4580 , n4579 );
or ( n4581 , n172 , n173 );
not ( n4582 , n4581 );
nor ( n4583 , n171 , n174 );
not ( n4584 , n4583 );
not ( n4585 , n4584 );
nand ( n4586 , n4585 , n175 );
not ( n4587 , n4586 );
nand ( n4588 , n4582 , n4587 );
not ( n4589 , n4588 );
nor ( n4590 , n4580 , n4589 );
not ( n4591 , n176 );
not ( n4592 , n175 );
nand ( n4593 , n4592 , n174 );
not ( n4594 , n4593 );
nand ( n4595 , n4594 , n173 );
or ( n4596 , n172 , n4595 );
not ( n4597 , n172 );
nand ( n4598 , n171 , n174 );
nor ( n4599 , n175 , n4598 );
buf ( n4600 , n4599 );
nand ( n4601 , n4597 , n4600 );
not ( n4602 , n173 );
not ( n4603 , n175 );
nand ( n4604 , n171 , n174 );
nor ( n4605 , n4603 , n4604 );
nand ( n4606 , n4602 , n4605 );
not ( n4607 , n4606 );
nand ( n4608 , n172 , n4607 );
nand ( n4609 , n4596 , n4601 , n4608 );
and ( n4610 , n4591 , n4609 );
not ( n4611 , n4591 );
not ( n4612 , n4576 );
not ( n4613 , n4612 );
nand ( n4614 , n172 , n4613 );
not ( n4615 , n4614 );
not ( n4616 , n4586 );
not ( n4617 , n172 );
nand ( n4618 , n4616 , n4617 );
not ( n4619 , n4618 );
nor ( n4620 , n4615 , n4619 );
not ( n4621 , n4581 );
not ( n4622 , n175 );
not ( n4623 , n174 );
nand ( n4624 , n4623 , n171 );
not ( n4625 , n4624 );
nand ( n4626 , n4622 , n4625 );
not ( n4627 , n4626 );
buf ( n4628 , n4627 );
nand ( n4629 , n4621 , n4628 );
not ( n4630 , n174 );
nand ( n4631 , n4630 , n175 );
nor ( n4632 , n173 , n4631 );
nand ( n4633 , n172 , n4632 );
not ( n4634 , n4626 );
nand ( n4635 , n4634 , n173 );
not ( n4636 , n4635 );
nand ( n4637 , n4636 , n172 );
nand ( n4638 , n4620 , n4629 , n4633 , n4637 );
and ( n4639 , n4611 , n4638 );
nor ( n4640 , n4610 , n4639 );
nand ( n4641 , n4590 , n4640 );
and ( n4642 , n4573 , n4641 );
not ( n4643 , n176 );
not ( n4644 , n4643 );
not ( n4645 , n175 );
nand ( n4646 , n4645 , n171 );
nand ( n4647 , n4646 , n4593 );
nand ( n4648 , n172 , n4647 );
not ( n4649 , n172 );
not ( n4650 , n4606 );
nand ( n4651 , n4649 , n4650 );
not ( n4652 , n172 );
not ( n4653 , n171 );
nor ( n4654 , n174 , n175 );
nand ( n4655 , n4653 , n4654 );
not ( n4656 , n4655 );
not ( n4657 , n173 );
nand ( n4658 , n4656 , n4657 );
not ( n4659 , n4658 );
nand ( n4660 , n4652 , n4659 );
nand ( n4661 , n4648 , n4651 , n4660 );
not ( n4662 , n4661 );
or ( n4663 , n4644 , n4662 );
nand ( n4664 , n173 , n4599 );
not ( n4665 , n4664 );
nand ( n4666 , n172 , n4665 );
not ( n4667 , n173 );
nand ( n4668 , n4628 , n4667 );
not ( n4669 , n172 );
nor ( n4670 , n4668 , n4669 );
not ( n4671 , n4670 );
and ( n4672 , n4666 , n4671 );
nand ( n4673 , n4663 , n4672 );
nand ( n4674 , n177 , n4673 );
not ( n4675 , n4674 );
nor ( n4676 , n4642 , n4675 );
not ( n4677 , n177 );
not ( n4678 , n176 );
nand ( n4679 , n172 , n173 );
not ( n4680 , n4679 );
not ( n4681 , n4584 );
not ( n4682 , n4681 );
not ( n4683 , n4682 );
nand ( n4684 , n4680 , n4683 );
not ( n4685 , n4684 );
nand ( n4686 , n4678 , n4685 );
not ( n4687 , n4686 );
nand ( n4688 , n171 , n175 );
nor ( n4689 , n173 , n4688 );
not ( n4690 , n4689 );
nor ( n4691 , n176 , n4690 );
nand ( n4692 , n171 , n175 );
not ( n4693 , n4692 );
nand ( n4694 , n4693 , n172 );
not ( n4695 , n4694 );
nor ( n4696 , n4687 , n4691 , n4695 );
not ( n4697 , n172 );
not ( n4698 , n173 );
buf ( n4699 , n4604 );
not ( n4700 , n4699 );
nand ( n4701 , n4698 , n4700 );
nor ( n4702 , n4697 , n4701 );
not ( n4703 , n4702 );
nor ( n4704 , n4622 , n4624 );
and ( n4705 , n173 , n4704 );
not ( n4706 , n4705 );
not ( n4707 , n4706 );
nand ( n4708 , n176 , n4707 );
nand ( n4709 , n4696 , n4703 , n4708 );
and ( n4710 , n4677 , n4709 );
not ( n4711 , n4677 );
not ( n4712 , n4625 );
nor ( n4713 , n173 , n4712 );
nand ( n4714 , n176 , n4713 );
not ( n4715 , n4714 );
not ( n4716 , n4715 );
not ( n4717 , n4655 );
nand ( n4718 , n173 , n4717 );
nor ( n4719 , n172 , n4718 );
not ( n4720 , n4719 );
not ( n4721 , n173 );
not ( n4722 , n174 );
nor ( n4723 , n4722 , n171 );
nand ( n4724 , n4721 , n4723 );
not ( n4725 , n4724 );
not ( n4726 , n4635 );
or ( n4727 , n4725 , n4726 );
not ( n4728 , n176 );
nand ( n4729 , n4727 , n4728 );
not ( n4730 , n173 );
not ( n4731 , n4586 );
nand ( n4732 , n4730 , n4731 );
not ( n4733 , n4732 );
nand ( n4734 , n172 , n4733 );
nand ( n4735 , n4716 , n4720 , n4729 , n4734 );
and ( n4736 , n4711 , n4735 );
nor ( n4737 , n4710 , n4736 );
not ( n4738 , n172 );
nand ( n4739 , n4738 , n173 );
or ( n4740 , n171 , n4739 );
not ( n4741 , n4607 );
nand ( n4742 , n4740 , n4741 );
and ( n4743 , n176 , n4742 );
not ( n4744 , n176 );
not ( n4745 , n4600 );
not ( n4746 , n172 );
nor ( n4747 , n4745 , n4746 );
not ( n4748 , n4747 );
not ( n4749 , n4724 );
nand ( n4750 , n172 , n4749 );
nand ( n4751 , n4748 , n4750 , n4660 );
and ( n4752 , n4744 , n4751 );
nor ( n4753 , n4743 , n4752 );
not ( n4754 , n173 );
nand ( n4755 , n4754 , n172 );
or ( n4756 , n174 , n4755 );
not ( n4757 , n4627 );
not ( n4758 , n172 );
nor ( n4759 , n4757 , n4758 );
not ( n4760 , n4759 );
nand ( n4761 , n4756 , n4760 );
nand ( n4762 , n176 , n4761 );
nand ( n4763 , n4737 , n4753 , n4762 );
nand ( n4764 , n178 , n4763 );
not ( n4765 , n178 );
not ( n4766 , n4723 );
not ( n4767 , n4766 );
nand ( n4768 , n173 , n4767 );
not ( n4769 , n4768 );
nand ( n4770 , n172 , n4769 );
not ( n4771 , n176 );
nor ( n4772 , n4771 , n4612 );
not ( n4773 , n4772 );
and ( n4774 , n4770 , n4773 );
not ( n4775 , n176 );
nor ( n4776 , n4775 , n172 );
not ( n4777 , n173 );
nor ( n4778 , n4777 , n4646 );
nand ( n4779 , n4776 , n4778 );
not ( n4780 , n176 );
not ( n4781 , n172 );
not ( n4782 , n4704 );
not ( n4783 , n4782 );
nand ( n4784 , n4781 , n4783 );
nand ( n4785 , n4784 , n4706 , n4668 );
nand ( n4786 , n4780 , n4785 );
nand ( n4787 , n4774 , n4779 , n4786 );
nand ( n4788 , n177 , n4787 );
not ( n4789 , n176 );
nor ( n4790 , n172 , n4664 );
and ( n4791 , n4789 , n4790 );
nor ( n4792 , n4791 , n4589 );
not ( n4793 , n172 );
not ( n4794 , n4793 );
or ( n4795 , n173 , n4593 );
not ( n4796 , n4795 );
not ( n4797 , n4796 );
or ( n4798 , n4794 , n4797 );
not ( n4799 , n4718 );
nand ( n4800 , n172 , n4799 );
nand ( n4801 , n4798 , n4800 );
and ( n4802 , n176 , n4801 );
nand ( n4803 , n174 , n175 );
not ( n4804 , n4803 );
nand ( n4805 , n4804 , n173 );
not ( n4806 , n4805 );
and ( n4807 , n176 , n4806 );
not ( n4808 , n176 );
nor ( n4809 , n172 , n4612 );
and ( n4810 , n4808 , n4809 );
nor ( n4811 , n4807 , n4810 );
not ( n4812 , n173 );
nand ( n4813 , n4812 , n4681 );
not ( n4814 , n4813 );
nand ( n4815 , n172 , n4814 );
not ( n4816 , n4655 );
nand ( n4817 , n4816 , n176 );
and ( n4818 , n4811 , n4815 , n4817 );
nor ( n4819 , n4818 , n177 );
nor ( n4820 , n4802 , n4819 );
nand ( n4821 , n4788 , n4792 , n4820 );
nand ( n4822 , n4765 , n4821 );
not ( n4823 , n176 );
not ( n4824 , n172 );
nand ( n4825 , n4824 , n4769 );
or ( n4826 , n4823 , n4825 );
nand ( n4827 , n172 , n176 );
not ( n4828 , n4827 );
nand ( n4829 , n4828 , n4587 );
nand ( n4830 , n4826 , n4829 );
and ( n4831 , n177 , n4830 );
not ( n4832 , n176 );
nand ( n4833 , n174 , n175 );
or ( n4834 , n4832 , n4679 , n4833 );
not ( n4835 , n172 );
nor ( n4836 , n4835 , n176 );
not ( n4837 , n4836 );
not ( n4838 , n173 );
nand ( n4839 , n4622 , n4723 );
not ( n4840 , n4839 );
nand ( n4841 , n4838 , n4840 );
not ( n4842 , n4841 );
not ( n4843 , n4842 );
or ( n4844 , n4837 , n4843 );
nand ( n4845 , n4834 , n4844 );
nor ( n4846 , n4831 , n4845 );
nand ( n4847 , n4676 , n4764 , n4822 , n4846 );
not ( n4848 , n4847 );
and ( n4849 , n4572 , n4848 );
not ( n4850 , n4572 );
and ( n4851 , n4850 , n4847 );
or ( n4852 , n4849 , n4851 );
not ( n4853 , n4852 );
or ( n4854 , n4304 , n4853 );
or ( n4855 , n4303 , n4852 );
nand ( n4856 , n4854 , n4855 );
or ( n4857 , n176 , n4612 );
nand ( n4858 , n4825 , n4857 );
nor ( n4859 , n173 , n4646 );
nand ( n4860 , n4776 , n4859 );
not ( n4861 , n176 );
not ( n4862 , n172 );
not ( n4863 , n4766 );
nand ( n4864 , n4862 , n4863 );
not ( n4865 , n4864 );
nand ( n4866 , n4861 , n4865 );
and ( n4867 , n4633 , n4866 );
buf ( n4868 , n4654 );
nand ( n4869 , n173 , n4868 );
nand ( n4870 , n4805 , n4869 );
or ( n4871 , n4769 , n4870 );
not ( n4872 , n176 );
nand ( n4873 , n4871 , n4872 );
nand ( n4874 , n4860 , n4867 , n4873 );
or ( n4875 , n4858 , n4874 );
not ( n4876 , n177 );
nand ( n4877 , n4875 , n4876 );
nand ( n4878 , n176 , n177 );
not ( n4879 , n4878 );
not ( n4880 , n4879 );
not ( n4881 , n174 );
not ( n4882 , n4881 );
not ( n4883 , n173 );
and ( n4884 , n4882 , n4883 );
and ( n4885 , n172 , n4767 );
nor ( n4886 , n4884 , n4885 );
not ( n4887 , n172 );
not ( n4888 , n4682 );
nand ( n4889 , n4887 , n4888 );
nand ( n4890 , n4886 , n4869 , n4889 );
not ( n4891 , n4890 );
or ( n4892 , n4880 , n4891 );
nand ( n4893 , n4892 , n178 );
or ( n4894 , n176 , n4825 );
nand ( n4895 , n4828 , n4796 );
not ( n4896 , n171 );
nand ( n4897 , n4896 , n175 );
not ( n4898 , n4897 );
not ( n4899 , n4739 );
nand ( n4900 , n4898 , n4899 );
nand ( n4901 , n4894 , n4895 , n4900 );
nor ( n4902 , n4893 , n4901 );
not ( n4903 , n4666 );
nor ( n4904 , n172 , n176 );
not ( n4905 , n4904 );
not ( n4906 , n4905 );
nand ( n4907 , n4906 , n4628 );
not ( n4908 , n4907 );
or ( n4909 , n4903 , n4908 );
nand ( n4910 , n4909 , n177 );
or ( n4911 , n172 , n4701 );
not ( n4912 , n172 );
not ( n4913 , n173 );
nor ( n4914 , n4913 , n4631 );
nand ( n4915 , n4912 , n4914 );
nand ( n4916 , n4911 , n4577 , n4915 );
nand ( n4917 , n176 , n4916 );
nand ( n4918 , n4910 , n4917 );
not ( n4919 , n4918 );
nand ( n4920 , n4877 , n4902 , n4919 );
nand ( n4921 , n4828 , n4659 );
not ( n4922 , n172 );
not ( n4923 , n175 );
nor ( n4924 , n4923 , n4699 );
nand ( n4925 , n4922 , n4924 );
not ( n4926 , n4925 );
not ( n4927 , n172 );
nor ( n4928 , n173 , n4897 );
nand ( n4929 , n4927 , n4928 );
not ( n4930 , n4929 );
or ( n4931 , n4926 , n4930 );
not ( n4932 , n176 );
nand ( n4933 , n4931 , n4932 );
nand ( n4934 , n4765 , n4921 , n4933 );
not ( n4935 , n177 );
not ( n4936 , n4935 );
not ( n4937 , n4828 );
not ( n4938 , n4778 );
or ( n4939 , n4937 , n4938 );
nand ( n4940 , n4939 , n4817 );
not ( n4941 , n4940 );
or ( n4942 , n4936 , n4941 );
not ( n4943 , n173 );
nand ( n4944 , n4943 , n171 );
not ( n4945 , n4944 );
not ( n4946 , n176 );
nand ( n4947 , n4945 , n4946 );
not ( n4948 , n4947 );
nand ( n4949 , n172 , n4689 );
not ( n4950 , n4949 );
or ( n4951 , n4948 , n4950 );
not ( n4952 , n177 );
nand ( n4953 , n4951 , n4952 );
nand ( n4954 , n4942 , n4953 );
nor ( n4955 , n4934 , n4954 );
not ( n4956 , n4782 );
nand ( n4957 , n4956 , n172 );
not ( n4958 , n172 );
nand ( n4959 , n4958 , n4665 );
nand ( n4960 , n4957 , n4959 );
not ( n4961 , n176 );
not ( n4962 , n4961 );
not ( n4963 , n174 );
not ( n4964 , n4963 );
not ( n4965 , n4680 );
or ( n4966 , n4964 , n4965 );
nand ( n4967 , n172 , n4840 );
nand ( n4968 , n4966 , n4967 );
not ( n4969 , n4968 );
or ( n4970 , n4962 , n4969 );
not ( n4971 , n4595 );
nand ( n4972 , n4971 , n4776 );
nand ( n4973 , n4970 , n4972 );
or ( n4974 , n4960 , n4973 );
nand ( n4975 , n4974 , n177 );
nand ( n4976 , n173 , n4605 );
not ( n4977 , n4976 );
not ( n4978 , n4586 );
nand ( n4979 , n4978 , n173 );
not ( n4980 , n4979 );
or ( n4981 , n4977 , n4980 );
buf ( n4982 , n4828 );
nand ( n4983 , n4981 , n4982 );
not ( n4984 , n4718 );
not ( n4985 , n4579 );
or ( n4986 , n4984 , n4985 );
not ( n4987 , n176 );
nand ( n4988 , n4986 , n4987 );
nand ( n4989 , n4955 , n4975 , n4983 , n4988 );
nand ( n4990 , n4920 , n4989 );
not ( n4991 , n172 );
not ( n4992 , n4576 );
nor ( n4993 , n173 , n4992 );
nand ( n4994 , n4991 , n4993 );
not ( n4995 , n4994 );
not ( n4996 , n4995 );
nand ( n4997 , n4996 , n4800 );
not ( n4998 , n176 );
and ( n4999 , n4997 , n4998 );
not ( n5000 , n172 );
nand ( n5001 , n5000 , n4806 );
not ( n5002 , n4655 );
nand ( n5003 , n5002 , n172 );
and ( n5004 , n5001 , n5003 , n4666 );
not ( n5005 , n177 );
and ( n5006 , n176 , n5005 );
not ( n5007 , n5006 );
nor ( n5008 , n5004 , n5007 );
nor ( n5009 , n4999 , n5008 );
not ( n5010 , n177 );
nand ( n5011 , n172 , n4859 );
or ( n5012 , n176 , n5011 );
not ( n5013 , n4692 );
nand ( n5014 , n5013 , n173 );
not ( n5015 , n5014 );
not ( n5016 , n172 );
nand ( n5017 , n5015 , n5016 );
nand ( n5018 , n5012 , n5017 , n4933 );
nand ( n5019 , n5010 , n5018 );
not ( n5020 , n176 );
not ( n5021 , n172 );
not ( n5022 , n5021 );
nand ( n5023 , n4701 , n4635 , n4732 );
not ( n5024 , n5023 );
or ( n5025 , n5022 , n5024 );
not ( n5026 , n173 );
nand ( n5027 , n5026 , n4600 );
not ( n5028 , n5027 );
not ( n5029 , n5028 );
and ( n5030 , n4614 , n5029 );
nand ( n5031 , n5025 , n5030 );
not ( n5032 , n5031 );
or ( n5033 , n5020 , n5032 );
not ( n5034 , n4587 );
not ( n5035 , n4914 );
nand ( n5036 , n5034 , n5035 , n4741 , n4843 );
nand ( n5037 , n4836 , n5036 );
nand ( n5038 , n5033 , n5037 );
nand ( n5039 , n177 , n5038 );
nand ( n5040 , n4990 , n5009 , n5019 , n5039 );
buf ( n5041 , n5040 );
not ( n5042 , n5041 );
not ( n5043 , n5042 );
not ( n5044 , n177 );
not ( n5045 , n176 );
not ( n5046 , n172 );
not ( n5047 , n4631 );
nand ( n5048 , n5046 , n5047 );
not ( n5049 , n4778 );
nand ( n5050 , n5048 , n4782 , n5049 );
not ( n5051 , n5050 );
or ( n5052 , n5045 , n5051 );
nand ( n5053 , n5052 , n4748 );
not ( n5054 , n5053 );
not ( n5055 , n176 );
nand ( n5056 , n5055 , n4717 );
and ( n5057 , n5017 , n4706 , n4866 , n5056 );
nand ( n5058 , n5054 , n5057 );
not ( n5059 , n5058 );
or ( n5060 , n5044 , n5059 );
nor ( n5061 , n173 , n4612 );
nand ( n5062 , n172 , n5061 );
not ( n5063 , n5062 );
not ( n5064 , n5063 );
nand ( n5065 , n5060 , n5064 );
not ( n5066 , n4712 );
nand ( n5067 , n172 , n5066 );
not ( n5068 , n173 );
nor ( n5069 , n5067 , n5068 );
not ( n5070 , n5069 );
buf ( n5071 , n4839 );
not ( n5072 , n5071 );
not ( n5073 , n5072 );
not ( n5074 , n4628 );
nand ( n5075 , n5073 , n5074 );
nand ( n5076 , n173 , n5075 );
and ( n5077 , n5070 , n5076 );
not ( n5078 , n176 );
nor ( n5079 , n5077 , n5078 );
not ( n5080 , n5079 );
not ( n5081 , n176 );
not ( n5082 , n172 );
nand ( n5083 , n5082 , n4859 );
buf ( n5084 , n4924 );
nand ( n5085 , n172 , n5084 );
not ( n5086 , n172 );
and ( n5087 , n5086 , n4705 );
not ( n5088 , n5087 );
nand ( n5089 , n5083 , n5085 , n5088 );
nand ( n5090 , n5081 , n5089 );
nand ( n5091 , n176 , n4759 );
not ( n5092 , n176 );
not ( n5093 , n4928 );
or ( n5094 , n5092 , n5093 );
or ( n5095 , n4833 , n4581 );
nand ( n5096 , n5091 , n5094 , n5095 );
not ( n5097 , n172 );
nand ( n5098 , n5097 , n4814 );
not ( n5099 , n4601 );
not ( n5100 , n4967 );
or ( n5101 , n5099 , n5100 );
not ( n5102 , n176 );
nand ( n5103 , n5101 , n5102 );
nand ( n5104 , n4773 , n4637 , n5098 , n5103 );
or ( n5105 , n5096 , n5104 );
not ( n5106 , n177 );
nand ( n5107 , n5105 , n5106 );
nand ( n5108 , n5080 , n5090 , n5107 );
nor ( n5109 , n5065 , n5108 );
nor ( n5110 , n5109 , n4765 );
not ( n5111 , n5110 );
not ( n5112 , n5071 );
nand ( n5113 , n4680 , n5112 );
not ( n5114 , n4637 );
nand ( n5115 , n176 , n5114 );
nand ( n5116 , n5113 , n5115 );
not ( n5117 , n5116 );
not ( n5118 , n176 );
not ( n5119 , n5118 );
not ( n5120 , n4976 );
not ( n5121 , n172 );
nand ( n5122 , n5120 , n5121 );
nand ( n5123 , n4770 , n5122 );
not ( n5124 , n5123 );
or ( n5125 , n5119 , n5124 );
not ( n5126 , n173 );
nor ( n5127 , n171 , n175 );
nand ( n5128 , n5126 , n5127 );
not ( n5129 , n5128 );
nand ( n5130 , n4982 , n5129 );
nand ( n5131 , n5125 , n5130 );
not ( n5132 , n5131 );
nand ( n5133 , n176 , n4607 );
not ( n5134 , n172 );
nand ( n5135 , n5134 , n4842 );
and ( n5136 , n5133 , n5135 );
not ( n5137 , n177 );
not ( n5138 , n4706 );
nand ( n5139 , n5138 , n4836 );
and ( n5140 , n176 , n173 , n4888 );
nand ( n5141 , n4699 , n4688 );
and ( n5142 , n4776 , n5141 );
nor ( n5143 , n5140 , n5142 );
and ( n5144 , n4718 , n5143 );
nand ( n5145 , n5139 , n5083 , n5144 );
nand ( n5146 , n5137 , n5145 );
not ( n5147 , n4704 );
not ( n5148 , n5147 );
not ( n5149 , n173 );
nand ( n5150 , n5148 , n5149 );
or ( n5151 , n176 , n5150 );
not ( n5152 , n4976 );
nand ( n5153 , n5152 , n172 );
nand ( n5154 , n5151 , n4760 , n5153 );
not ( n5155 , n5128 );
not ( n5156 , n172 );
nand ( n5157 , n5156 , n4578 );
not ( n5158 , n5157 );
or ( n5159 , n5155 , n5158 );
nand ( n5160 , n5159 , n176 );
nand ( n5161 , n5160 , n4651 );
or ( n5162 , n5154 , n5161 );
nand ( n5163 , n5162 , n177 );
nand ( n5164 , n5132 , n5136 , n5146 , n5163 );
nand ( n5165 , n5164 , n4765 );
nor ( n5166 , n176 , n177 );
and ( n5167 , n5166 , n4702 );
not ( n5168 , n5028 );
not ( n5169 , n5168 );
and ( n5170 , n4982 , n5169 );
nor ( n5171 , n5167 , n5170 );
nand ( n5172 , n5117 , n5165 , n5171 );
not ( n5173 , n5172 );
not ( n5174 , n4833 );
not ( n5175 , n4755 );
nand ( n5176 , n5174 , n5175 );
and ( n5177 , n5176 , n4748 );
nor ( n5178 , n5177 , n4878 );
not ( n5179 , n4905 );
nand ( n5180 , n4869 , n4724 , n5150 );
nand ( n5181 , n5179 , n5180 );
not ( n5182 , n176 );
nand ( n5183 , n5182 , n4670 );
nand ( n5184 , n5181 , n4708 , n5183 );
nand ( n5185 , n177 , n5184 );
not ( n5186 , n5185 );
nor ( n5187 , n5178 , n5186 );
not ( n5188 , n177 );
not ( n5189 , n176 );
not ( n5190 , n4719 );
or ( n5191 , n5189 , n5190 );
not ( n5192 , n4841 );
nand ( n5193 , n4776 , n5192 );
nand ( n5194 , n5191 , n5193 );
nand ( n5195 , n5188 , n5194 );
nand ( n5196 , n5111 , n5173 , n5187 , n5195 );
not ( n5197 , n5196 );
not ( n5198 , n5197 );
and ( n5199 , n5043 , n5198 );
not ( n5200 , n5041 );
not ( n5201 , n5172 );
not ( n5202 , n5195 );
nor ( n5203 , n5202 , n5110 );
nand ( n5204 , n5201 , n5187 , n5203 );
not ( n5205 , n5204 );
and ( n5206 , n5200 , n5205 );
nor ( n5207 , n5199 , n5206 );
not ( n5208 , n5207 );
not ( n5209 , n166 );
nor ( n5210 , n5209 , n165 );
not ( n5211 , n5210 );
not ( n5212 , n168 );
nor ( n5213 , n5212 , n163 );
nand ( n5214 , n164 , n5213 );
not ( n5215 , n5214 );
not ( n5216 , n5215 );
nor ( n5217 , n5211 , n5216 );
not ( n5218 , n167 );
not ( n5219 , n5218 );
not ( n5220 , n165 );
not ( n5221 , n163 );
nor ( n5222 , n5221 , n164 );
nand ( n5223 , n5220 , n5222 );
nor ( n5224 , n166 , n5223 );
not ( n5225 , n5224 );
nand ( n5226 , n163 , n168 );
not ( n5227 , n5226 );
nand ( n5228 , n5227 , n164 );
not ( n5229 , n5228 );
nand ( n5230 , n166 , n5229 );
not ( n5231 , n166 );
not ( n5232 , n163 );
nor ( n5233 , n5232 , n168 );
and ( n5234 , n164 , n5233 );
nand ( n5235 , n165 , n5234 );
not ( n5236 , n5235 );
nand ( n5237 , n5231 , n5236 );
nand ( n5238 , n5225 , n5230 , n5237 );
not ( n5239 , n5238 );
or ( n5240 , n5219 , n5239 );
not ( n5241 , n165 );
not ( n5242 , n164 );
nand ( n5243 , n5242 , n5213 );
not ( n5244 , n5243 );
not ( n5245 , n5244 );
not ( n5246 , n5233 );
not ( n5247 , n5246 );
not ( n5248 , n164 );
nand ( n5249 , n5247 , n5248 );
buf ( n5250 , n5249 );
nand ( n5251 , n5245 , n5250 );
not ( n5252 , n5251 );
or ( n5253 , n5241 , n5252 );
not ( n5254 , n5246 );
not ( n5255 , n5254 );
not ( n5256 , n5255 );
nand ( n5257 , n5256 , n166 );
not ( n5258 , n5257 );
nand ( n5259 , n165 , n5258 );
nand ( n5260 , n5253 , n5259 );
nand ( n5261 , n167 , n5260 );
nand ( n5262 , n5240 , n5261 );
nor ( n5263 , n5217 , n5262 );
not ( n5264 , n5263 );
not ( n5265 , n167 );
not ( n5266 , n168 );
nand ( n5267 , n5266 , n164 );
not ( n5268 , n5267 );
not ( n5269 , n166 );
nand ( n5270 , n5268 , n5269 );
not ( n5271 , n164 );
nand ( n5272 , n5271 , n163 );
nor ( n5273 , n5220 , n5272 );
not ( n5274 , n5273 );
not ( n5275 , n5234 );
not ( n5276 , n5275 );
not ( n5277 , n5276 );
nand ( n5278 , n5270 , n5274 , n5277 );
not ( n5279 , n5278 );
or ( n5280 , n5265 , n5279 );
not ( n5281 , n5226 );
nand ( n5282 , n5248 , n5281 );
not ( n5283 , n5282 );
nand ( n5284 , n166 , n5283 );
nand ( n5285 , n5280 , n5284 );
not ( n5286 , n5285 );
not ( n5287 , n166 );
not ( n5288 , n165 );
nand ( n5289 , n163 , n164 );
nor ( n5290 , n5288 , n5289 );
nand ( n5291 , n5287 , n5290 );
not ( n5292 , n166 );
not ( n5293 , n163 );
and ( n5294 , n168 , n5293 );
nand ( n5295 , n5292 , n5294 );
nor ( n5296 , n167 , n5295 );
not ( n5297 , n5296 );
not ( n5298 , n167 );
not ( n5299 , n164 );
nor ( n5300 , n163 , n168 );
buf ( n5301 , n5300 );
nand ( n5302 , n5299 , n5301 );
not ( n5303 , n5302 );
nand ( n5304 , n5298 , n5303 );
and ( n5305 , n5291 , n5235 , n5297 , n5304 );
nand ( n5306 , n5286 , n5305 );
and ( n5307 , n169 , n5306 );
not ( n5308 , n169 );
not ( n5309 , n5215 );
not ( n5310 , n5309 );
nand ( n5311 , n167 , n5310 );
nand ( n5312 , n164 , n168 );
nor ( n5313 , n165 , n166 );
not ( n5314 , n5313 );
nor ( n5315 , n5312 , n5314 );
not ( n5316 , n5315 );
not ( n5317 , n165 );
nand ( n5318 , n5317 , n5301 );
nor ( n5319 , n166 , n5318 );
not ( n5320 , n5319 );
and ( n5321 , n5311 , n5316 , n5320 );
not ( n5322 , n167 );
not ( n5323 , n163 );
nand ( n5324 , n5323 , n164 );
nor ( n5325 , n165 , n5324 );
not ( n5326 , n5325 );
or ( n5327 , n5322 , n5326 );
not ( n5328 , n166 );
nand ( n5329 , n5328 , n5283 );
not ( n5330 , n5329 );
not ( n5331 , n5243 );
nand ( n5332 , n166 , n5331 );
not ( n5333 , n5332 );
or ( n5334 , n5330 , n5333 );
not ( n5335 , n167 );
nand ( n5336 , n5334 , n5335 );
nand ( n5337 , n165 , n166 );
not ( n5338 , n5337 );
not ( n5339 , n5250 );
nand ( n5340 , n5338 , n5339 );
not ( n5341 , n166 );
nor ( n5342 , n5341 , n5249 );
nand ( n5343 , n167 , n5342 );
and ( n5344 , n5340 , n5343 );
nand ( n5345 , n5321 , n5327 , n5336 , n5344 );
and ( n5346 , n5308 , n5345 );
nor ( n5347 , n5307 , n5346 );
not ( n5348 , n5347 );
or ( n5349 , n5264 , n5348 );
nand ( n5350 , n5349 , n170 );
not ( n5351 , n5281 );
nor ( n5352 , n165 , n5351 );
nand ( n5353 , n166 , n5352 );
not ( n5354 , n5353 );
nor ( n5355 , n167 , n169 );
nand ( n5356 , n5354 , n5355 );
nand ( n5357 , n5338 , n5244 );
nand ( n5358 , n166 , n167 );
not ( n5359 , n5249 );
nand ( n5360 , n165 , n5359 );
or ( n5361 , n5358 , n5360 );
and ( n5362 , n5356 , n5357 , n5361 );
not ( n5363 , n169 );
not ( n5364 , n167 );
not ( n5365 , n166 );
nand ( n5366 , n5365 , n165 );
not ( n5367 , n5366 );
not ( n5368 , n5302 );
nand ( n5369 , n5367 , n5368 );
or ( n5370 , n5364 , n5369 );
not ( n5371 , n167 );
nor ( n5372 , n5371 , n166 );
not ( n5373 , n5372 );
nand ( n5374 , n5220 , n5331 );
nor ( n5375 , n5373 , n5374 );
not ( n5376 , n5375 );
nand ( n5377 , n5370 , n5376 );
and ( n5378 , n5363 , n5377 );
and ( n5379 , n167 , n169 );
or ( n5380 , n5312 , n5211 );
nand ( n5381 , n5380 , n5284 );
and ( n5382 , n5379 , n5381 );
nor ( n5383 , n5378 , n5382 );
and ( n5384 , n5362 , n5383 );
nand ( n5385 , n5350 , n5384 );
not ( n5386 , n167 );
not ( n5387 , n5228 );
nand ( n5388 , n5387 , n5220 );
or ( n5389 , n5386 , n5388 );
not ( n5390 , n5389 );
not ( n5391 , n166 );
nand ( n5392 , n165 , n5294 );
nor ( n5393 , n5391 , n5392 );
not ( n5394 , n5228 );
nand ( n5395 , n5394 , n165 );
nor ( n5396 , n166 , n5395 );
nor ( n5397 , n5393 , n5396 );
or ( n5398 , n167 , n5397 );
not ( n5399 , n166 );
not ( n5400 , n5374 );
nand ( n5401 , n5399 , n5400 );
nand ( n5402 , n5398 , n5401 );
nor ( n5403 , n5390 , n5402 );
not ( n5404 , n165 );
nor ( n5405 , n163 , n164 );
nand ( n5406 , n5404 , n5405 );
or ( n5407 , n5358 , n5406 );
not ( n5408 , n169 );
not ( n5409 , n5408 );
not ( n5410 , n167 );
nand ( n5411 , n166 , n5410 );
not ( n5412 , n5411 );
not ( n5413 , n5235 );
nand ( n5414 , n5412 , n5413 );
not ( n5415 , n167 );
not ( n5416 , n5415 );
nand ( n5417 , n165 , n5301 );
not ( n5418 , n5417 );
and ( n5419 , n5416 , n5418 );
nor ( n5420 , n5419 , n5224 );
not ( n5421 , n5372 );
buf ( n5422 , n5289 );
nand ( n5423 , n5422 , n5351 );
not ( n5424 , n5423 );
or ( n5425 , n5421 , n5424 );
not ( n5426 , n5302 );
nand ( n5427 , n5426 , n165 );
nand ( n5428 , n5425 , n5427 );
not ( n5429 , n5428 );
and ( n5430 , n5414 , n5420 , n5429 );
not ( n5431 , n5430 );
or ( n5432 , n5409 , n5431 );
not ( n5433 , n167 );
nor ( n5434 , n165 , n5275 );
nand ( n5435 , n5433 , n5434 );
not ( n5436 , n5342 );
not ( n5437 , n166 );
or ( n5438 , n5437 , n5395 );
and ( n5439 , n5435 , n5436 , n5438 );
or ( n5440 , n166 , n5388 );
nand ( n5441 , n165 , n5215 );
or ( n5442 , n5441 , n166 );
nand ( n5443 , n5442 , n5406 );
nand ( n5444 , n167 , n5443 );
and ( n5445 , n5440 , n5444 );
nand ( n5446 , n169 , n5439 , n5445 );
nand ( n5447 , n5432 , n5446 );
nand ( n5448 , n5403 , n5407 , n5447 );
not ( n5449 , n170 );
nand ( n5450 , n5448 , n5449 );
nor ( n5451 , n166 , n167 );
nor ( n5452 , n164 , n168 );
not ( n5453 , n5452 );
not ( n5454 , n5453 );
nand ( n5455 , n5454 , n165 );
not ( n5456 , n5294 );
nor ( n5457 , n165 , n5456 );
not ( n5458 , n5457 );
not ( n5459 , n5434 );
nand ( n5460 , n5455 , n5458 , n5459 );
nand ( n5461 , n5451 , n5460 );
nand ( n5462 , n167 , n5413 );
not ( n5463 , n167 );
not ( n5464 , n166 );
nand ( n5465 , n5220 , n5359 );
nor ( n5466 , n5464 , n5465 );
nand ( n5467 , n5463 , n5466 );
nand ( n5468 , n5461 , n5462 , n5467 );
nand ( n5469 , n169 , n5468 );
not ( n5470 , n167 );
not ( n5471 , n5282 );
and ( n5472 , n5220 , n5471 );
nand ( n5473 , n166 , n5472 );
or ( n5474 , n5470 , n5473 );
nand ( n5475 , n5450 , n5469 , n5474 );
nor ( n5476 , n5385 , n5475 );
not ( n5477 , n169 );
and ( n5478 , n167 , n5477 );
not ( n5479 , n5478 );
not ( n5480 , n166 );
not ( n5481 , n165 );
nor ( n5482 , n5481 , n5312 );
nand ( n5483 , n5480 , n5482 );
not ( n5484 , n5302 );
nand ( n5485 , n166 , n5484 );
not ( n5486 , n5282 );
nand ( n5487 , n5486 , n165 );
not ( n5488 , n5487 );
nand ( n5489 , n5488 , n166 );
nand ( n5490 , n5483 , n5485 , n5489 );
not ( n5491 , n5490 );
or ( n5492 , n5479 , n5491 );
nor ( n5493 , n5314 , n5216 );
not ( n5494 , n5427 );
nand ( n5495 , n5494 , n166 );
not ( n5496 , n5495 );
or ( n5497 , n5493 , n5496 );
not ( n5498 , n167 );
nand ( n5499 , n5497 , n5498 );
nand ( n5500 , n5492 , n5499 );
not ( n5501 , n5500 );
not ( n5502 , n5358 );
not ( n5503 , n5302 );
nand ( n5504 , n5503 , n5220 );
not ( n5505 , n5504 );
nand ( n5506 , n5502 , n5505 );
not ( n5507 , n169 );
not ( n5508 , n5507 );
not ( n5509 , n5502 );
not ( n5510 , n5273 );
or ( n5511 , n5509 , n5510 );
nand ( n5512 , n5484 , n167 );
nand ( n5513 , n5511 , n5512 );
not ( n5514 , n5513 );
or ( n5515 , n5508 , n5514 );
not ( n5516 , n167 );
not ( n5517 , n163 );
nor ( n5518 , n5517 , n165 );
nand ( n5519 , n5516 , n5518 );
not ( n5520 , n5519 );
nor ( n5521 , n165 , n5422 );
nand ( n5522 , n166 , n5521 );
not ( n5523 , n5522 );
or ( n5524 , n5520 , n5523 );
not ( n5525 , n169 );
nand ( n5526 , n5524 , n5525 );
nand ( n5527 , n5515 , n5526 );
not ( n5528 , n5527 );
not ( n5529 , n166 );
nand ( n5530 , n5529 , n5325 );
not ( n5531 , n5530 );
not ( n5532 , n166 );
nand ( n5533 , n5532 , n5229 );
not ( n5534 , n5533 );
or ( n5535 , n5531 , n5534 );
not ( n5536 , n167 );
nand ( n5537 , n5535 , n5536 );
not ( n5538 , n5395 );
nand ( n5539 , n164 , n5300 );
not ( n5540 , n5539 );
nand ( n5541 , n5540 , n165 );
not ( n5542 , n5541 );
or ( n5543 , n5538 , n5542 );
nand ( n5544 , n5543 , n5502 );
and ( n5545 , n5449 , n5537 , n5544 );
and ( n5546 , n5506 , n5528 , n5545 );
not ( n5547 , n5427 );
not ( n5548 , n5441 );
nand ( n5549 , n166 , n5548 );
not ( n5550 , n5549 );
or ( n5551 , n5547 , n5550 );
not ( n5552 , n167 );
nand ( n5553 , n5551 , n5552 );
not ( n5554 , n5372 );
not ( n5555 , n164 );
nand ( n5556 , n5555 , n168 );
nor ( n5557 , n5220 , n5556 );
not ( n5558 , n5557 );
or ( n5559 , n5554 , n5558 );
not ( n5560 , n166 );
nor ( n5561 , n5560 , n168 );
nand ( n5562 , n165 , n5561 );
not ( n5563 , n5562 );
not ( n5564 , n5332 );
or ( n5565 , n5563 , n5564 );
not ( n5566 , n167 );
nand ( n5567 , n5565 , n5566 );
nand ( n5568 , n5559 , n5567 );
not ( n5569 , n5568 );
nand ( n5570 , n166 , n5276 );
not ( n5571 , n5487 );
not ( n5572 , n166 );
nand ( n5573 , n5571 , n5572 );
nand ( n5574 , n5569 , n5570 , n5573 );
nand ( n5575 , n169 , n5574 );
nand ( n5576 , n5546 , n5553 , n5575 );
not ( n5577 , n169 );
not ( n5578 , n5451 );
not ( n5579 , n5339 );
or ( n5580 , n5578 , n5579 );
nand ( n5581 , n5580 , n5489 );
not ( n5582 , n5581 );
or ( n5583 , n5577 , n5582 );
and ( n5584 , n166 , n5294 );
not ( n5585 , n168 );
nor ( n5586 , n5585 , n165 );
nor ( n5587 , n5584 , n5586 );
not ( n5588 , n166 );
nand ( n5589 , n5588 , n5301 );
nand ( n5590 , n5587 , n5455 , n5589 );
nand ( n5591 , n5379 , n5590 );
nand ( n5592 , n5583 , n5591 );
not ( n5593 , n5592 );
nor ( n5594 , n165 , n5556 );
nand ( n5595 , n5502 , n5594 );
not ( n5596 , n5324 );
nand ( n5597 , n5596 , n5367 );
not ( n5598 , n167 );
nor ( n5599 , n166 , n5392 );
nand ( n5600 , n5598 , n5599 );
and ( n5601 , n5597 , n170 , n5600 );
not ( n5602 , n169 );
not ( n5603 , n5602 );
not ( n5604 , n167 );
not ( n5605 , n5482 );
nand ( n5606 , n5455 , n5605 , n5392 );
nand ( n5607 , n5604 , n5606 );
nand ( n5608 , n167 , n5224 );
not ( n5609 , n165 );
not ( n5610 , n5267 );
nand ( n5611 , n5609 , n5610 );
not ( n5612 , n166 );
nor ( n5613 , n5611 , n5612 );
nor ( n5614 , n5599 , n5613 );
nor ( n5615 , n167 , n5309 );
nor ( n5616 , n5615 , n5296 );
nand ( n5617 , n5607 , n5608 , n5614 , n5616 );
not ( n5618 , n5617 );
or ( n5619 , n5603 , n5618 );
not ( n5620 , n166 );
nand ( n5621 , n5620 , n5352 );
not ( n5622 , n166 );
nor ( n5623 , n5220 , n5267 );
nand ( n5624 , n5622 , n5623 );
nand ( n5625 , n5621 , n5441 , n5624 );
nand ( n5626 , n167 , n5625 );
nand ( n5627 , n5619 , n5626 );
not ( n5628 , n5627 );
nand ( n5629 , n5593 , n5595 , n5601 , n5628 );
nand ( n5630 , n5576 , n5629 );
not ( n5631 , n5539 );
nand ( n5632 , n166 , n5631 );
not ( n5633 , n5632 );
nand ( n5634 , n5388 , n5374 );
or ( n5635 , n5623 , n5634 );
nand ( n5636 , n5635 , n166 );
not ( n5637 , n5636 );
or ( n5638 , n5633 , n5637 );
not ( n5639 , n167 );
nand ( n5640 , n5638 , n5639 );
not ( n5641 , n166 );
not ( n5642 , n5641 );
not ( n5643 , n5352 );
nor ( n5644 , n165 , n5539 );
not ( n5645 , n5644 );
nand ( n5646 , n5360 , n5643 , n5645 );
not ( n5647 , n5646 );
or ( n5648 , n5642 , n5647 );
nand ( n5649 , n166 , n5215 );
not ( n5650 , n5472 );
and ( n5651 , n5649 , n5650 );
nand ( n5652 , n5648 , n5651 );
nand ( n5653 , n167 , n5652 );
nand ( n5654 , n5640 , n5653 );
and ( n5655 , n169 , n5654 );
not ( n5656 , n169 );
not ( n5657 , n166 );
nor ( n5658 , n5657 , n5223 );
not ( n5659 , n5658 );
or ( n5660 , n5659 , n167 );
nand ( n5661 , n5660 , n5291 , n5537 );
and ( n5662 , n5656 , n5661 );
nor ( n5663 , n5655 , n5662 );
nand ( n5664 , n5501 , n5630 , n5663 );
buf ( n5665 , n5664 );
and ( n5666 , n5476 , n5665 );
not ( n5667 , n5476 );
not ( n5668 , n5500 );
and ( n5669 , n5630 , n5668 , n5663 );
not ( n5670 , n5669 );
not ( n5671 , n5670 );
and ( n5672 , n5667 , n5671 );
nor ( n5673 , n5666 , n5672 );
nand ( n5674 , n5208 , n5673 );
not ( n5675 , n5673 );
nand ( n5676 , n5675 , n5207 );
nand ( n5677 , n5674 , n5676 );
or ( n5678 , n4856 , n5677 );
nand ( n5679 , n4856 , n5677 );
nand ( n5680 , n5678 , n5679 , n2352 );
nand ( n5681 , n4028 , n5680 );
not ( n5682 , n946 );
not ( n5683 , n5682 );
not ( n5684 , n782 );
or ( n5685 , n5683 , n5684 );
nand ( n5686 , n5685 , n970 );
and ( n5687 , n793 , n5686 );
nor ( n5688 , n5687 , n10 );
not ( n5689 , n5688 );
not ( n5690 , n17 );
not ( n5691 , n16 );
not ( n5692 , n15 );
nand ( n5693 , n5692 , n14 );
not ( n5694 , n5693 );
nand ( n5695 , n13 , n5694 );
not ( n5696 , n769 );
nand ( n5697 , n13 , n5696 );
nand ( n5698 , n5695 , n5697 , n856 );
nand ( n5699 , n5691 , n5698 );
not ( n5700 , n13 );
nor ( n5701 , n5700 , n960 );
not ( n5702 , n5701 );
not ( n5703 , n13 );
nand ( n5704 , n5703 , n866 );
not ( n5705 , n5704 );
nand ( n5706 , n13 , n753 );
not ( n5707 , n5706 );
or ( n5708 , n5705 , n5707 );
nand ( n5709 , n5708 , n16 );
nand ( n5710 , n5699 , n5702 , n5709 );
not ( n5711 , n5710 );
or ( n5712 , n5690 , n5711 );
not ( n5713 , n12 );
nand ( n5714 , n15 , n865 );
not ( n5715 , n5714 );
nand ( n5716 , n5713 , n5715 );
not ( n5717 , n5716 );
nand ( n5718 , n5717 , n13 );
nor ( n5719 , n16 , n5718 );
nand ( n5720 , n12 , n770 );
or ( n5721 , n809 , n5720 );
buf ( n5722 , n923 );
nand ( n5723 , n5721 , n5722 );
nor ( n5724 , n5719 , n5723 );
nand ( n5725 , n5712 , n5724 );
not ( n5726 , n5725 );
not ( n5727 , n5726 );
or ( n5728 , n5689 , n5727 );
not ( n5729 , n17 );
not ( n5730 , n16 );
not ( n5731 , n14 );
or ( n5732 , n5731 , n858 );
nand ( n5733 , n5732 , n748 );
nand ( n5734 , n5730 , n5733 );
nand ( n5735 , n16 , n940 );
not ( n5736 , n861 );
not ( n5737 , n16 );
nand ( n5738 , n5736 , n5737 );
not ( n5739 , n5738 );
nand ( n5740 , n929 , n5739 );
nand ( n5741 , n5734 , n5735 , n5740 );
not ( n5742 , n5741 );
or ( n5743 , n5729 , n5742 );
not ( n5744 , n846 );
nor ( n5745 , n5744 , n935 );
not ( n5746 , n5745 );
not ( n5747 , n13 );
not ( n5748 , n5716 );
nand ( n5749 , n5747 , n5748 );
and ( n5750 , n5746 , n5749 );
nand ( n5751 , n5743 , n5750 );
not ( n5752 , n5751 );
not ( n5753 , n12 );
nor ( n5754 , n5753 , n5714 );
not ( n5755 , n5754 );
not ( n5756 , n849 );
nand ( n5757 , n12 , n800 );
nand ( n5758 , n5755 , n5756 , n5757 );
nand ( n5759 , n810 , n5758 );
not ( n5760 , n743 );
not ( n5761 , n940 );
or ( n5762 , n5760 , n5761 );
nand ( n5763 , n5762 , n931 );
not ( n5764 , n5763 );
not ( n5765 , n12 );
nand ( n5766 , n5765 , n914 );
not ( n5767 , n5766 );
nand ( n5768 , n5767 , n16 );
not ( n5769 , n13 );
nand ( n5770 , n5769 , n947 );
and ( n5771 , n5768 , n820 , n5770 );
not ( n5772 , n974 );
nand ( n5773 , n16 , n5772 );
not ( n5774 , n5714 );
not ( n5775 , n5774 );
nor ( n5776 , n13 , n5775 );
nor ( n5777 , n16 , n5720 );
nor ( n5778 , n5776 , n5777 );
nand ( n5779 , n5764 , n5771 , n5773 , n5778 );
nand ( n5780 , n793 , n5779 );
not ( n5781 , n13 );
nand ( n5782 , n5781 , n862 );
not ( n5783 , n5782 );
nand ( n5784 , n16 , n5783 );
not ( n5785 , n5784 );
nor ( n5786 , n841 , n5785 );
nand ( n5787 , n5752 , n5759 , n5780 , n5786 );
nand ( n5788 , n5728 , n5787 );
nand ( n5789 , n743 , n5774 );
and ( n5790 , n789 , n5789 );
not ( n5791 , n746 );
nand ( n5792 , n13 , n5791 );
not ( n5793 , n902 );
nand ( n5794 , n13 , n5793 );
nand ( n5795 , n5792 , n970 , n5794 );
nand ( n5796 , n16 , n5795 );
not ( n5797 , n748 );
nand ( n5798 , n13 , n5797 );
not ( n5799 , n16 );
not ( n5800 , n862 );
not ( n5801 , n12 );
nor ( n5802 , n5800 , n5801 );
nand ( n5803 , n5802 , n13 );
nand ( n5804 , n5716 , n917 , n5803 );
nand ( n5805 , n5799 , n5804 );
nand ( n5806 , n5790 , n5796 , n5798 , n5805 );
and ( n5807 , n793 , n5806 );
not ( n5808 , n793 );
not ( n5809 , n13 );
not ( n5810 , n835 );
nor ( n5811 , n5809 , n5810 );
and ( n5812 , n16 , n5811 );
not ( n5813 , n13 );
nand ( n5814 , n5813 , n813 );
not ( n5815 , n5814 );
nor ( n5816 , n5812 , n5815 );
not ( n5817 , n12 );
nand ( n5818 , n5817 , n11 );
or ( n5819 , n13 , n5818 );
nand ( n5820 , n5819 , n5720 );
nand ( n5821 , n16 , n5820 );
not ( n5822 , n16 );
not ( n5823 , n859 );
not ( n5824 , n914 );
or ( n5825 , n5823 , n5824 );
nand ( n5826 , n5825 , n816 , n854 );
nand ( n5827 , n5822 , n5826 );
nand ( n5828 , n5816 , n5821 , n5827 );
and ( n5829 , n5808 , n5828 );
nor ( n5830 , n5807 , n5829 );
not ( n5831 , n5774 );
nand ( n5832 , n876 , n5831 );
nand ( n5833 , n5832 , n16 , n846 );
and ( n5834 , n791 , n5833 );
nand ( n5835 , n5788 , n5830 , n5834 );
not ( n5836 , n1134 );
nand ( n5837 , n1243 , n1249 , n1274 , n5836 );
xor ( n5838 , n5835 , n5837 );
and ( n5839 , n16 , n17 );
not ( n5840 , n13 );
not ( n5841 , n5840 );
not ( n5842 , n819 );
not ( n5843 , n786 );
nand ( n5844 , n5843 , n12 );
nand ( n5845 , n5842 , n5844 , n5716 );
not ( n5846 , n5845 );
or ( n5847 , n5841 , n5846 );
nand ( n5848 , n13 , n862 );
and ( n5849 , n5848 , n816 );
nand ( n5850 , n5847 , n5849 );
nand ( n5851 , n5839 , n5850 );
not ( n5852 , n13 );
not ( n5853 , n16 );
nand ( n5854 , n17 , n5853 );
nor ( n5855 , n5852 , n5854 );
not ( n5856 , n12 );
nor ( n5857 , n957 , n5856 );
not ( n5858 , n5857 );
nand ( n5859 , n5831 , n5858 , n902 , n884 );
and ( n5860 , n5855 , n5859 );
nand ( n5861 , n796 , n977 );
and ( n5862 , n862 , n846 );
not ( n5863 , n862 );
and ( n5864 , n5863 , n5744 );
nor ( n5865 , n5862 , n5864 );
nand ( n5866 , n5861 , n5865 );
not ( n5867 , n16 );
and ( n5868 , n5866 , n5867 );
nor ( n5869 , n5860 , n5868 );
not ( n5870 , n16 );
nand ( n5871 , n5870 , n13 , n879 );
not ( n5872 , n13 );
nand ( n5873 , n5872 , n849 );
not ( n5874 , n5873 );
not ( n5875 , n5770 );
or ( n5876 , n5874 , n5875 );
not ( n5877 , n16 );
nand ( n5878 , n5876 , n5877 );
nand ( n5879 , n5871 , n970 , n5878 );
nand ( n5880 , n793 , n5879 );
and ( n5881 , n16 , n793 );
not ( n5882 , n13 );
not ( n5883 , n763 );
nand ( n5884 , n5883 , n12 );
not ( n5885 , n5884 );
nand ( n5886 , n5882 , n5885 );
nand ( n5887 , n13 , n977 );
nand ( n5888 , n12 , n770 );
not ( n5889 , n5888 );
nand ( n5890 , n5889 , n13 );
nand ( n5891 , n5886 , n5887 , n5890 );
nand ( n5892 , n5881 , n5891 );
nand ( n5893 , n5851 , n5869 , n5880 , n5892 );
not ( n5894 , n5893 );
or ( n5895 , n16 , n5818 );
nor ( n5896 , n12 , n868 );
nand ( n5897 , n13 , n5896 );
nand ( n5898 , n5895 , n5897 );
and ( n5899 , n793 , n5898 );
not ( n5900 , n793 );
nor ( n5901 , n13 , n5888 );
nor ( n5902 , n5701 , n5901 );
nand ( n5903 , n12 , n5694 );
not ( n5904 , n5903 );
nand ( n5905 , n5904 , n833 );
not ( n5906 , n13 );
nor ( n5907 , n5906 , n14 );
nand ( n5908 , n12 , n5907 );
not ( n5909 , n5908 );
not ( n5910 , n799 );
nand ( n5911 , n13 , n5910 );
not ( n5912 , n5911 );
or ( n5913 , n5909 , n5912 );
not ( n5914 , n16 );
nand ( n5915 , n5913 , n5914 );
nand ( n5916 , n5902 , n5905 , n5915 );
and ( n5917 , n5900 , n5916 );
nor ( n5918 , n5899 , n5917 );
not ( n5919 , n864 );
not ( n5920 , n5803 );
or ( n5921 , n5919 , n5920 );
not ( n5922 , n16 );
nand ( n5923 , n5921 , n5922 );
nand ( n5924 , n5918 , n5878 , n5923 );
not ( n5925 , n961 );
and ( n5926 , n810 , n5925 );
not ( n5927 , n16 );
not ( n5928 , n827 );
nor ( n5929 , n5927 , n5928 );
nor ( n5930 , n5926 , n5929 );
or ( n5931 , n17 , n5930 );
nand ( n5932 , n810 , n866 , n834 );
not ( n5933 , n852 );
not ( n5934 , n5755 );
or ( n5935 , n5933 , n5934 );
nand ( n5936 , n5935 , n810 );
nand ( n5937 , n5931 , n5932 , n5936 );
or ( n5938 , n5924 , n5937 );
nand ( n5939 , n5938 , n841 );
not ( n5940 , n12 );
nand ( n5941 , n5940 , n14 );
nand ( n5942 , n13 , n752 );
nand ( n5943 , n5941 , n5942 , n748 , n5704 );
and ( n5944 , n5839 , n5943 );
and ( n5945 , n5682 , n859 );
nor ( n5946 , n5944 , n5945 );
not ( n5947 , n12 );
nand ( n5948 , n5947 , n5694 );
not ( n5949 , n5948 );
nand ( n5950 , n5949 , n810 );
not ( n5951 , n13 );
nand ( n5952 , n5951 , n819 );
not ( n5953 , n861 );
nand ( n5954 , n5953 , n12 );
not ( n5955 , n13 );
nand ( n5956 , n5955 , n5857 );
nand ( n5957 , n5952 , n5954 , n5956 );
nand ( n5958 , n16 , n5957 );
nand ( n5959 , n5946 , n5950 , n5958 );
not ( n5960 , n5959 );
not ( n5961 , n890 );
nor ( n5962 , n5961 , n13 );
not ( n5963 , n5962 );
or ( n5964 , n16 , n5963 );
not ( n5965 , n16 );
not ( n5966 , n890 );
nand ( n5967 , n5966 , n5884 , n748 );
nand ( n5968 , n5965 , n5967 );
nor ( n5969 , n5962 , n975 );
and ( n5970 , n879 , n833 );
not ( n5971 , n13 );
not ( n5972 , n12 );
nand ( n5973 , n5972 , n958 );
nor ( n5974 , n5971 , n5973 );
nor ( n5975 , n5970 , n5974 );
nand ( n5976 , n5968 , n5738 , n5969 , n5975 );
and ( n5977 , n793 , n5976 );
not ( n5978 , n793 );
not ( n5979 , n744 );
not ( n5980 , n935 );
not ( n5981 , n5980 );
or ( n5982 , n5979 , n5981 );
nand ( n5983 , n5982 , n5890 );
and ( n5984 , n5978 , n5983 );
nor ( n5985 , n5977 , n5984 );
nand ( n5986 , n5960 , n5964 , n5985 );
nand ( n5987 , n10 , n5986 );
nand ( n5988 , n5894 , n5939 , n5987 );
buf ( n5989 , n5988 );
not ( n5990 , n5989 );
not ( n5991 , n65 );
and ( n5992 , n5990 , n5991 );
not ( n5993 , n5990 );
and ( n5994 , n5993 , n65 );
nor ( n5995 , n5992 , n5994 );
xor ( n5996 , n5838 , n5995 );
not ( n5997 , n32 );
nand ( n5998 , n5997 , n2033 );
nand ( n5999 , n2096 , n5998 );
not ( n6000 , n5999 );
nand ( n6001 , n31 , n1659 );
not ( n6002 , n1685 );
and ( n6003 , n6001 , n6002 );
not ( n6004 , n31 );
not ( n6005 , n2107 );
nand ( n6006 , n6004 , n6005 );
nand ( n6007 , n6006 , n1710 , n2026 );
nand ( n6008 , n32 , n6007 );
nand ( n6009 , n6000 , n6003 , n2183 , n6008 );
and ( n6010 , n33 , n6009 );
not ( n6011 , n27 );
not ( n6012 , n1545 );
nand ( n6013 , n1532 , n6012 );
not ( n6014 , n6013 );
or ( n6015 , n6011 , n6014 );
nand ( n6016 , n6015 , n1635 );
nand ( n6017 , n32 , n6016 );
not ( n6018 , n6017 );
nor ( n6019 , n6010 , n6018 );
not ( n6020 , n32 );
not ( n6021 , n31 );
nand ( n6022 , n6021 , n1685 );
nand ( n6023 , n31 , n1526 );
not ( n6024 , n2102 );
and ( n6025 , n6023 , n6024 );
nand ( n6026 , n6022 , n6025 );
and ( n6027 , n6020 , n6026 );
nor ( n6028 , n6027 , n1494 );
not ( n6029 , n33 );
not ( n6030 , n1668 );
not ( n6031 , n2069 );
or ( n6032 , n6030 , n6031 );
not ( n6033 , n32 );
nand ( n6034 , n6032 , n6033 );
not ( n6035 , n2166 );
nand ( n6036 , n6035 , n31 );
not ( n6037 , n32 );
nand ( n6038 , n31 , n1545 );
nor ( n6039 , n6037 , n6038 );
nor ( n6040 , n1593 , n6039 );
nand ( n6041 , n32 , n1573 );
not ( n6042 , n2089 );
nand ( n6043 , n6042 , n1539 );
and ( n6044 , n6041 , n6043 , n1562 );
nand ( n6045 , n6034 , n6036 , n6040 , n6044 );
nand ( n6046 , n6029 , n6045 );
nand ( n6047 , n6019 , n6028 , n6046 );
nand ( n6048 , n34 , n6047 );
not ( n6049 , n33 );
not ( n6050 , n32 );
not ( n6051 , n31 );
nand ( n6052 , n6051 , n2200 );
or ( n6053 , n6050 , n6052 );
not ( n6054 , n1749 );
nand ( n6055 , n2074 , n6054 );
nand ( n6056 , n6053 , n6055 );
nand ( n6057 , n6049 , n6056 );
not ( n6058 , n33 );
not ( n6059 , n1716 );
not ( n6060 , n1604 );
not ( n6061 , n1709 );
not ( n6062 , n6061 );
not ( n6063 , n27 );
nand ( n6064 , n6062 , n6063 );
nand ( n6065 , n6059 , n6060 , n6064 );
nand ( n6066 , n1608 , n6065 );
nand ( n6067 , n32 , n1686 );
nand ( n6068 , n6066 , n6067 , n1729 );
not ( n6069 , n6068 );
or ( n6070 , n6058 , n6069 );
not ( n6071 , n31 );
nor ( n6072 , n6071 , n27 );
not ( n6073 , n6072 );
or ( n6074 , n2089 , n6073 );
not ( n6075 , n6001 );
not ( n6076 , n6075 );
nand ( n6077 , n6074 , n6076 );
nand ( n6078 , n1739 , n6077 );
nand ( n6079 , n6070 , n6078 );
not ( n6080 , n6079 );
nand ( n6081 , n6048 , n6057 , n6080 );
not ( n6082 , n6081 );
nand ( n6083 , n1629 , n2068 );
not ( n6084 , n6036 );
nand ( n6085 , n6084 , n32 );
and ( n6086 , n6083 , n6085 );
not ( n6087 , n1662 );
not ( n6088 , n6087 );
not ( n6089 , n6088 );
and ( n6090 , n1515 , n6089 );
nor ( n6091 , n32 , n33 );
not ( n6092 , n6091 );
nor ( n6093 , n6092 , n1569 );
nor ( n6094 , n6090 , n6093 );
not ( n6095 , n32 );
not ( n6096 , n6095 );
nand ( n6097 , n31 , n2114 );
not ( n6098 , n31 );
nand ( n6099 , n6098 , n1651 );
not ( n6100 , n6099 );
not ( n6101 , n6100 );
nand ( n6102 , n6097 , n6101 );
not ( n6103 , n6102 );
or ( n6104 , n6096 , n6103 );
nand ( n6105 , n1515 , n1705 );
nand ( n6106 , n6104 , n6105 );
not ( n6107 , n6106 );
not ( n6108 , n2158 );
nand ( n6109 , n32 , n6108 );
not ( n6110 , n31 );
nand ( n6111 , n6110 , n6054 );
and ( n6112 , n6109 , n6111 );
not ( n6113 , n33 );
and ( n6114 , n32 , n27 , n1497 );
nand ( n6115 , n1567 , n1615 );
and ( n6116 , n2074 , n6115 );
nor ( n6117 , n6114 , n6116 );
and ( n6118 , n2042 , n6117 );
nand ( n6119 , n2155 , n1686 );
nand ( n6120 , n6118 , n6024 , n6119 );
and ( n6121 , n6113 , n6120 );
not ( n6122 , n6113 );
not ( n6123 , n6038 );
not ( n6124 , n6123 );
not ( n6125 , n6124 );
not ( n6126 , n31 );
nand ( n6127 , n6126 , n1623 );
not ( n6128 , n6127 );
nor ( n6129 , n6125 , n6128 );
not ( n6130 , n32 );
not ( n6131 , n6064 );
nand ( n6132 , n6130 , n6131 );
not ( n6133 , n1706 );
not ( n6134 , n2142 );
not ( n6135 , n31 );
nand ( n6136 , n6134 , n6135 );
not ( n6137 , n6136 );
or ( n6138 , n6133 , n6137 );
nand ( n6139 , n6138 , n32 );
nand ( n6140 , n6129 , n6132 , n1654 , n6139 );
and ( n6141 , n6122 , n6140 );
nor ( n6142 , n6121 , n6141 );
nand ( n6143 , n6107 , n6112 , n6142 );
nand ( n6144 , n1673 , n6143 );
nand ( n6145 , n6082 , n6086 , n6094 , n6144 );
not ( n6146 , n6145 );
not ( n6147 , n2006 );
or ( n6148 , n6146 , n6147 );
nand ( n6149 , n6082 , n6086 , n6094 , n6144 );
not ( n6150 , n6149 );
nor ( n6151 , n2004 , n1879 );
nand ( n6152 , n6150 , n6151 );
nand ( n6153 , n6148 , n6152 );
not ( n6154 , n26 );
not ( n6155 , n6154 );
not ( n6156 , n23 );
not ( n6157 , n6156 );
not ( n6158 , n1860 );
and ( n6159 , n6157 , n6158 );
not ( n6160 , n1867 );
not ( n6161 , n25 );
not ( n6162 , n23 );
and ( n6163 , n24 , n1771 );
and ( n6164 , n6162 , n6163 );
nand ( n6165 , n6161 , n6164 );
nand ( n6166 , n6160 , n6165 );
nor ( n6167 , n6159 , n6166 );
nand ( n6168 , n23 , n1859 );
not ( n6169 , n1901 );
nand ( n6170 , n23 , n1837 );
nand ( n6171 , n6168 , n6169 , n6170 );
nand ( n6172 , n25 , n6171 );
nand ( n6173 , n1812 , n6163 );
not ( n6174 , n6173 );
not ( n6175 , n1969 );
not ( n6176 , n1820 );
nand ( n6177 , n23 , n6176 );
not ( n6178 , n6177 );
or ( n6179 , n6174 , n6175 , n6178 );
not ( n6180 , n25 );
nand ( n6181 , n6179 , n6180 );
nand ( n6182 , n6167 , n6172 , n6181 );
not ( n6183 , n6182 );
or ( n6184 , n6155 , n6183 );
nand ( n6185 , n22 , n1874 );
not ( n6186 , n6185 );
not ( n6187 , n6186 );
not ( n6188 , n6187 );
nand ( n6189 , n1800 , n6188 );
not ( n6190 , n25 );
nand ( n6191 , n23 , n6174 );
not ( n6192 , n6191 );
nand ( n6193 , n6190 , n6192 );
nand ( n6194 , n6189 , n1766 , n6193 );
not ( n6195 , n26 );
not ( n6196 , n6195 );
not ( n6197 , n1925 );
not ( n6198 , n6197 );
not ( n6199 , n1768 );
or ( n6200 , n6198 , n6199 );
nand ( n6201 , n6200 , n6169 );
not ( n6202 , n6201 );
or ( n6203 , n6196 , n6202 );
not ( n6204 , n25 );
not ( n6205 , n24 );
nand ( n6206 , n6205 , n20 );
not ( n6207 , n6206 );
nand ( n6208 , n23 , n6207 );
not ( n6209 , n23 );
nor ( n6210 , n6209 , n1787 );
not ( n6211 , n6210 );
nand ( n6212 , n6208 , n6211 , n1803 );
nand ( n6213 , n6204 , n6212 );
not ( n6214 , n1887 );
nand ( n6215 , n6214 , n23 );
not ( n6216 , n1920 );
nor ( n6217 , n6216 , n23 );
not ( n6218 , n6217 );
nand ( n6219 , n23 , n1857 );
not ( n6220 , n6219 );
or ( n6221 , n6218 , n6220 );
nand ( n6222 , n6221 , n25 );
nand ( n6223 , n6213 , n6215 , n6222 );
nand ( n6224 , n26 , n6223 );
nand ( n6225 , n6203 , n6224 );
or ( n6226 , n6194 , n6225 );
nand ( n6227 , n6226 , n1853 );
nand ( n6228 , n6184 , n6227 );
not ( n6229 , n6228 );
not ( n6230 , n22 );
nand ( n6231 , n6230 , n21 );
or ( n6232 , n23 , n6231 );
nand ( n6233 , n6232 , n6187 );
and ( n6234 , n1987 , n6233 );
not ( n6235 , n6163 );
and ( n6236 , n1779 , n6235 );
not ( n6237 , n25 );
nor ( n6238 , n6236 , n6237 , n1918 );
nor ( n6239 , n6234 , n6238 );
not ( n6240 , n26 );
nor ( n6241 , n6240 , n1799 , n1813 );
nor ( n6242 , n1869 , n6241 );
or ( n6243 , n25 , n1827 );
not ( n6244 , n25 );
not ( n6245 , n1967 );
not ( n6246 , n6245 );
not ( n6247 , n1996 );
not ( n6248 , n6247 );
or ( n6249 , n6246 , n6248 );
nand ( n6250 , n6249 , n1875 );
nand ( n6251 , n6244 , n6250 );
not ( n6252 , n1931 );
not ( n6253 , n6252 );
nand ( n6254 , n6243 , n6251 , n6253 );
nand ( n6255 , n26 , n6254 );
and ( n6256 , n6239 , n6242 , n6255 );
not ( n6257 , n26 );
not ( n6258 , n6257 );
not ( n6259 , n25 );
and ( n6260 , n6259 , n1922 );
not ( n6261 , n1904 );
and ( n6262 , n25 , n6261 );
nor ( n6263 , n6260 , n6262 );
not ( n6264 , n25 );
nand ( n6265 , n6264 , n6188 );
nor ( n6266 , n1915 , n6164 );
nor ( n6267 , n22 , n1967 );
nand ( n6268 , n25 , n6267 );
not ( n6269 , n23 );
nand ( n6270 , n6269 , n1926 );
and ( n6271 , n1979 , n6268 , n6270 );
nand ( n6272 , n6263 , n6265 , n6266 , n6271 );
not ( n6273 , n6272 );
or ( n6274 , n6258 , n6273 );
not ( n6275 , n1918 );
nand ( n6276 , n6275 , n6163 );
nand ( n6277 , n22 , n1933 );
not ( n6278 , n6277 );
nand ( n6279 , n22 , n6163 );
not ( n6280 , n6279 );
nor ( n6281 , n1952 , n6280 );
not ( n6282 , n6281 );
or ( n6283 , n6278 , n6282 );
nand ( n6284 , n6283 , n1800 );
nand ( n6285 , n6276 , n6284 );
not ( n6286 , n26 );
not ( n6287 , n25 );
not ( n6288 , n20 );
or ( n6289 , n6288 , n1996 );
nand ( n6290 , n6289 , n1860 );
nand ( n6291 , n6287 , n6290 );
not ( n6292 , n1921 );
nand ( n6293 , n25 , n6292 );
not ( n6294 , n1913 );
nor ( n6295 , n25 , n6294 );
nand ( n6296 , n1960 , n6295 );
nand ( n6297 , n6291 , n6293 , n6296 );
not ( n6298 , n6297 );
or ( n6299 , n6286 , n6298 );
nand ( n6300 , n1794 , n1913 );
not ( n6301 , n6300 );
nor ( n6302 , n1918 , n1963 );
nor ( n6303 , n6301 , n6302 );
nand ( n6304 , n6299 , n6303 );
nor ( n6305 , n6285 , n6304 );
nand ( n6306 , n6274 , n6305 );
nand ( n6307 , n19 , n6306 );
nand ( n6308 , n6229 , n6256 , n6307 );
not ( n6309 , n6308 );
not ( n6310 , n19 );
nand ( n6311 , n1812 , n6207 );
not ( n6312 , n6311 );
nand ( n6313 , n6312 , n1800 );
nand ( n6314 , n6197 , n1997 );
not ( n6315 , n23 );
nand ( n6316 , n6315 , n1977 );
buf ( n6317 , n1820 );
not ( n6318 , n23 );
nor ( n6319 , n1812 , n1884 );
nand ( n6320 , n6318 , n6319 );
nand ( n6321 , n6316 , n6317 , n6320 );
nand ( n6322 , n25 , n6321 );
nand ( n6323 , n6313 , n6314 , n6322 );
not ( n6324 , n1987 );
nor ( n6325 , n6288 , n22 );
nand ( n6326 , n23 , n1809 );
nand ( n6327 , n1860 , n6217 );
nand ( n6328 , n6325 , n6326 , n6327 );
not ( n6329 , n6328 );
or ( n6330 , n6324 , n6329 );
nand ( n6331 , n23 , n6186 );
not ( n6332 , n6331 );
not ( n6333 , n1963 );
nand ( n6334 , n1855 , n6333 );
not ( n6335 , n6334 );
or ( n6336 , n6332 , n6335 );
nand ( n6337 , n6336 , n26 );
nand ( n6338 , n6330 , n6337 );
nor ( n6339 , n6323 , n6338 );
not ( n6340 , n1843 );
not ( n6341 , n23 );
nand ( n6342 , n6340 , n6341 );
not ( n6343 , n6342 );
not ( n6344 , n25 );
nand ( n6345 , n6343 , n6344 );
not ( n6346 , n26 );
not ( n6347 , n25 );
not ( n6348 , n1916 );
and ( n6349 , n22 , n6348 );
not ( n6350 , n6349 );
nand ( n6351 , n1843 , n6350 , n1860 );
nand ( n6352 , n6347 , n6351 );
nand ( n6353 , n25 , n1950 );
nor ( n6354 , n22 , n1884 );
nand ( n6355 , n23 , n6354 );
and ( n6356 , n6342 , n6355 );
nor ( n6357 , n6295 , n1905 );
nand ( n6358 , n6352 , n6353 , n6356 , n6357 );
nand ( n6359 , n6346 , n6358 );
nand ( n6360 , n6339 , n6345 , n6359 );
not ( n6361 , n6360 );
or ( n6362 , n6310 , n6361 );
and ( n6363 , n1812 , n1785 );
nand ( n6364 , n1800 , n6363 );
not ( n6365 , n6231 );
not ( n6366 , n25 );
nand ( n6367 , n6365 , n6366 );
not ( n6368 , n6367 );
nor ( n6369 , n22 , n1789 );
nand ( n6370 , n23 , n6369 );
not ( n6371 , n6370 );
or ( n6372 , n6368 , n6371 );
not ( n6373 , n26 );
nand ( n6374 , n6372 , n6373 );
nand ( n6375 , n6364 , n6374 );
not ( n6376 , n25 );
not ( n6377 , n6376 );
nand ( n6378 , n1786 , n6177 );
not ( n6379 , n6378 );
or ( n6380 , n6377 , n6379 );
nand ( n6381 , n25 , n1785 );
not ( n6382 , n6381 );
not ( n6383 , n1889 );
nand ( n6384 , n1800 , n6383 );
not ( n6385 , n6384 );
or ( n6386 , n6382 , n6385 );
not ( n6387 , n26 );
nand ( n6388 , n6386 , n6387 );
nand ( n6389 , n6380 , n6388 );
nor ( n6390 , n6375 , n6389 );
not ( n6391 , n23 );
nand ( n6392 , n6391 , n1952 );
not ( n6393 , n6392 );
not ( n6394 , n6270 );
or ( n6395 , n6393 , n6394 );
not ( n6396 , n25 );
nand ( n6397 , n6395 , n6396 );
not ( n6398 , n6397 );
not ( n6399 , n1825 );
not ( n6400 , n6279 );
or ( n6401 , n6399 , n6400 );
nand ( n6402 , n6401 , n1800 );
not ( n6403 , n6402 );
nor ( n6404 , n6398 , n6403 );
not ( n6405 , n23 );
nand ( n6406 , n6405 , n6186 );
nand ( n6407 , n6215 , n6406 );
not ( n6408 , n1794 );
not ( n6409 , n22 );
nor ( n6410 , n6409 , n6206 );
not ( n6411 , n6410 );
or ( n6412 , n6408 , n6411 );
not ( n6413 , n23 );
nor ( n6414 , n6413 , n20 );
nand ( n6415 , n22 , n6414 );
not ( n6416 , n6415 );
not ( n6417 , n1934 );
or ( n6418 , n6416 , n6417 );
not ( n6419 , n25 );
nand ( n6420 , n6418 , n6419 );
nand ( n6421 , n6412 , n6420 );
or ( n6422 , n6407 , n6421 );
nand ( n6423 , n6422 , n26 );
and ( n6424 , n6390 , n6404 , n6423 );
nor ( n6425 , n6424 , n19 );
not ( n6426 , n25 );
nand ( n6427 , n23 , n1780 );
not ( n6428 , n6427 );
nand ( n6429 , n6426 , n6428 );
and ( n6430 , n6429 , n6169 , n6397 );
nor ( n6431 , n6430 , n26 );
not ( n6432 , n6431 );
not ( n6433 , n1768 );
not ( n6434 , n6319 );
nand ( n6435 , n6434 , n6235 , n1836 , n1813 );
not ( n6436 , n6435 );
or ( n6437 , n6433 , n6436 );
not ( n6438 , n23 );
not ( n6439 , n6438 );
nand ( n6440 , n1978 , n1984 , n6173 );
not ( n6441 , n6440 );
or ( n6442 , n6439 , n6441 );
nand ( n6443 , n23 , n1913 );
not ( n6444 , n6443 );
nor ( n6445 , n6444 , n1876 );
nand ( n6446 , n6442 , n6445 );
nand ( n6447 , n25 , n6446 );
nand ( n6448 , n6437 , n6447 );
nand ( n6449 , n26 , n6448 );
not ( n6450 , n23 );
not ( n6451 , n1913 );
nor ( n6452 , n22 , n6451 );
nand ( n6453 , n6450 , n6452 );
not ( n6454 , n6453 );
not ( n6455 , n1786 );
nand ( n6456 , n6455 , n23 );
not ( n6457 , n6456 );
or ( n6458 , n6454 , n6457 );
not ( n6459 , n25 );
nand ( n6460 , n6458 , n6459 );
not ( n6461 , n26 );
and ( n6462 , n25 , n6461 );
not ( n6463 , n23 );
nand ( n6464 , n6463 , n6349 );
nand ( n6465 , n23 , n1785 );
nand ( n6466 , n6464 , n6465 , n6331 );
nand ( n6467 , n6462 , n6466 );
nand ( n6468 , n6460 , n6467 );
not ( n6469 , n6468 );
nand ( n6470 , n6432 , n6449 , n6469 );
nor ( n6471 , n6425 , n6470 );
nand ( n6472 , n6362 , n6471 );
buf ( n6473 , n6472 );
not ( n6474 , n6473 );
or ( n6475 , n6309 , n6474 );
not ( n6476 , n19 );
not ( n6477 , n6306 );
or ( n6478 , n6476 , n6477 );
nand ( n6479 , n6478 , n6256 );
nor ( n6480 , n6479 , n6228 );
not ( n6481 , n6472 );
nand ( n6482 , n6480 , n6481 );
nand ( n6483 , n6475 , n6482 );
xor ( n6484 , n6153 , n6483 );
nor ( n6485 , n5996 , n6484 );
not ( n6486 , n5996 );
not ( n6487 , n6484 );
or ( n6488 , n6486 , n6487 );
nand ( n6489 , n6488 , n2352 );
or ( n6490 , n6485 , n6489 );
and ( n6491 , n66 , n5991 );
not ( n6492 , n66 );
and ( n6493 , n6492 , n65 );
nor ( n6494 , n6491 , n6493 );
or ( n6495 , n2352 , n6494 );
nand ( n6496 , n6490 , n6495 );
not ( n6497 , n67 );
and ( n6498 , n68 , n6497 );
not ( n6499 , n68 );
and ( n6500 , n6499 , n67 );
nor ( n6501 , n6498 , n6500 );
or ( n6502 , n2352 , n6501 );
not ( n6503 , n5837 );
not ( n6504 , n6149 );
or ( n6505 , n6503 , n6504 );
nand ( n6506 , n1276 , n6150 );
nand ( n6507 , n6505 , n6506 );
and ( n6508 , n987 , n6497 );
not ( n6509 , n987 );
and ( n6510 , n6509 , n67 );
nor ( n6511 , n6508 , n6510 );
not ( n6512 , n6511 );
and ( n6513 , n6507 , n6512 );
not ( n6514 , n6507 );
and ( n6515 , n6514 , n6511 );
nor ( n6516 , n6513 , n6515 );
not ( n6517 , n6516 );
and ( n6518 , n1758 , n2209 );
not ( n6519 , n1758 );
and ( n6520 , n6519 , n2210 );
nor ( n6521 , n6518 , n6520 );
not ( n6522 , n6521 );
not ( n6523 , n6483 );
and ( n6524 , n6522 , n6523 );
and ( n6525 , n6521 , n6483 );
nor ( n6526 , n6524 , n6525 );
not ( n6527 , n6526 );
nand ( n6528 , n6517 , n6527 );
nand ( n6529 , n6516 , n6526 );
nand ( n6530 , n6528 , n2352 , n6529 );
nand ( n6531 , n6502 , n6530 );
not ( n6532 , n228 );
and ( n6533 , n229 , n6532 );
not ( n6534 , n229 );
and ( n6535 , n6534 , n228 );
nor ( n6536 , n6533 , n6535 );
or ( n6537 , n2352 , n6536 );
not ( n6538 , n144 );
nand ( n6539 , n138 , n143 );
not ( n6540 , n6539 );
nand ( n6541 , n142 , n6540 );
not ( n6542 , n141 );
nand ( n6543 , n6542 , n142 );
not ( n6544 , n6543 );
nor ( n6545 , n139 , n143 );
not ( n6546 , n6545 );
not ( n6547 , n6546 );
nand ( n6548 , n140 , n6547 );
not ( n6549 , n6548 );
nand ( n6550 , n6544 , n6549 );
and ( n6551 , n6541 , n6550 );
not ( n6552 , n141 );
nor ( n6553 , n140 , n6539 );
nand ( n6554 , n6552 , n6553 );
not ( n6555 , n142 );
nand ( n6556 , n139 , n143 );
nor ( n6557 , n140 , n6556 );
not ( n6558 , n6557 );
or ( n6559 , n6555 , n6558 );
not ( n6560 , n139 );
nand ( n6561 , n6560 , n143 );
not ( n6562 , n6561 );
nand ( n6563 , n138 , n6562 );
not ( n6564 , n6563 );
nand ( n6565 , n140 , n6564 );
not ( n6566 , n6565 );
not ( n6567 , n6566 );
not ( n6568 , n6567 );
nand ( n6569 , n141 , n6568 );
nand ( n6570 , n6551 , n6554 , n6559 , n6569 );
and ( n6571 , n6538 , n6570 );
not ( n6572 , n143 );
not ( n6573 , n142 );
nand ( n6574 , n6573 , n140 );
not ( n6575 , n6574 );
and ( n6576 , n6572 , n6575 );
not ( n6577 , n140 );
not ( n6578 , n142 );
nor ( n6579 , n6578 , n139 );
and ( n6580 , n6577 , n6579 );
nor ( n6581 , n6576 , n6580 );
nand ( n6582 , n139 , n143 );
not ( n6583 , n6582 );
nand ( n6584 , n6583 , n138 );
not ( n6585 , n6584 );
not ( n6586 , n140 );
nand ( n6587 , n6585 , n6586 );
not ( n6588 , n138 );
nand ( n6589 , n6562 , n6588 );
not ( n6590 , n6589 );
and ( n6591 , n142 , n6590 );
not ( n6592 , n6591 );
and ( n6593 , n6581 , n6587 , n6592 );
not ( n6594 , n141 );
nor ( n6595 , n6593 , n6594 );
nor ( n6596 , n6571 , n6595 );
not ( n6597 , n144 );
not ( n6598 , n140 );
and ( n6599 , n138 , n6545 );
not ( n6600 , n6599 );
not ( n6601 , n6600 );
nand ( n6602 , n6598 , n6601 );
not ( n6603 , n6602 );
nand ( n6604 , n6603 , n142 );
and ( n6605 , n6588 , n6545 );
not ( n6606 , n6605 );
not ( n6607 , n140 );
nor ( n6608 , n6606 , n6607 );
not ( n6609 , n6608 );
nor ( n6610 , n6609 , n142 );
not ( n6611 , n6610 );
not ( n6612 , n140 );
and ( n6613 , n6612 , n6562 );
not ( n6614 , n6613 );
not ( n6615 , n141 );
nor ( n6616 , n6614 , n6615 );
not ( n6617 , n6616 );
not ( n6618 , n140 );
not ( n6619 , n139 );
nor ( n6620 , n6619 , n143 );
not ( n6621 , n6620 );
not ( n6622 , n6621 );
nand ( n6623 , n6618 , n6622 );
not ( n6624 , n6623 );
not ( n6625 , n6589 );
nand ( n6626 , n6625 , n140 );
not ( n6627 , n6626 );
or ( n6628 , n6624 , n6627 );
not ( n6629 , n141 );
nand ( n6630 , n6628 , n6629 );
nand ( n6631 , n6604 , n6611 , n6617 , n6630 );
not ( n6632 , n6631 );
or ( n6633 , n6597 , n6632 );
not ( n6634 , n141 );
buf ( n6635 , n6605 );
not ( n6636 , n6635 );
not ( n6637 , n6636 );
not ( n6638 , n142 );
not ( n6639 , n140 );
nand ( n6640 , n6638 , n6639 );
not ( n6641 , n6640 );
nand ( n6642 , n6637 , n6641 );
nor ( n6643 , n138 , n6582 );
and ( n6644 , n142 , n6643 );
not ( n6645 , n6644 );
not ( n6646 , n6623 );
nand ( n6647 , n6646 , n142 );
nand ( n6648 , n6642 , n6645 , n6647 );
nand ( n6649 , n6634 , n6648 );
nand ( n6650 , n6633 , n6649 );
not ( n6651 , n6650 );
nand ( n6652 , n6596 , n6651 );
and ( n6653 , n137 , n6652 );
not ( n6654 , n140 );
nand ( n6655 , n6588 , n6620 );
not ( n6656 , n6655 );
nand ( n6657 , n6654 , n6656 );
not ( n6658 , n6657 );
nand ( n6659 , n142 , n6658 );
or ( n6660 , n141 , n6659 );
nand ( n6661 , n141 , n142 );
nand ( n6662 , n138 , n139 );
not ( n6663 , n6662 );
nand ( n6664 , n6663 , n140 );
or ( n6665 , n6661 , n6664 );
nand ( n6666 , n6660 , n6665 );
nor ( n6667 , n6653 , n6666 );
not ( n6668 , n144 );
not ( n6669 , n139 );
nor ( n6670 , n6669 , n143 );
and ( n6671 , n138 , n6670 );
nand ( n6672 , n140 , n6671 );
not ( n6673 , n6672 );
nand ( n6674 , n6673 , n142 );
not ( n6675 , n6674 );
not ( n6676 , n6600 );
nand ( n6677 , n6641 , n6676 );
not ( n6678 , n6677 );
nor ( n6679 , n6675 , n6678 );
not ( n6680 , n141 );
not ( n6681 , n140 );
not ( n6682 , n138 );
nand ( n6683 , n6682 , n139 );
nor ( n6684 , n6681 , n6683 );
not ( n6685 , n6684 );
or ( n6686 , n142 , n6685 );
not ( n6687 , n142 );
nand ( n6688 , n6687 , n6643 );
not ( n6689 , n6587 );
nand ( n6690 , n6689 , n142 );
nand ( n6691 , n6686 , n6688 , n6690 );
nand ( n6692 , n6680 , n6691 );
not ( n6693 , n6600 );
not ( n6694 , n142 );
nand ( n6695 , n6693 , n6694 );
not ( n6696 , n6590 );
not ( n6697 , n6696 );
nand ( n6698 , n6697 , n6641 );
nand ( n6699 , n6695 , n6698 );
not ( n6700 , n6671 );
not ( n6701 , n6700 );
nand ( n6702 , n142 , n6701 );
not ( n6703 , n139 );
nand ( n6704 , n6703 , n138 );
nor ( n6705 , n140 , n6704 );
nand ( n6706 , n142 , n6705 );
not ( n6707 , n6626 );
nand ( n6708 , n142 , n6707 );
nand ( n6709 , n6702 , n6706 , n6708 );
or ( n6710 , n6699 , n6709 );
nand ( n6711 , n6710 , n141 );
nand ( n6712 , n6679 , n6692 , n6711 );
nand ( n6713 , n6668 , n6712 );
not ( n6714 , n142 );
not ( n6715 , n6621 );
nand ( n6716 , n140 , n6715 );
not ( n6717 , n6716 );
nand ( n6718 , n6714 , n6717 );
not ( n6719 , n6718 );
not ( n6720 , n6719 );
not ( n6721 , n6720 );
nand ( n6722 , n141 , n6721 );
nand ( n6723 , n142 , n6676 );
not ( n6724 , n6723 );
nand ( n6725 , n6724 , n141 );
not ( n6726 , n140 );
and ( n6727 , n6590 , n6726 );
nand ( n6728 , n142 , n6727 );
and ( n6729 , n6722 , n6725 , n6728 );
not ( n6730 , n142 );
nand ( n6731 , n140 , n6643 );
nor ( n6732 , n6730 , n6731 );
not ( n6733 , n6732 );
not ( n6734 , n141 );
not ( n6735 , n143 );
nor ( n6736 , n6735 , n138 );
not ( n6737 , n6736 );
nand ( n6738 , n6683 , n6737 );
nand ( n6739 , n142 , n6738 );
not ( n6740 , n6587 );
not ( n6741 , n142 );
nand ( n6742 , n6740 , n6741 );
nand ( n6743 , n6739 , n6742 , n6642 );
nand ( n6744 , n6734 , n6743 );
nand ( n6745 , n6729 , n6733 , n6744 );
nand ( n6746 , n144 , n6745 );
not ( n6747 , n141 );
nor ( n6748 , n138 , n6556 );
not ( n6749 , n6748 );
not ( n6750 , n6749 );
nand ( n6751 , n6575 , n6750 );
not ( n6752 , n6751 );
and ( n6753 , n6747 , n6752 );
not ( n6754 , n144 );
not ( n6755 , n141 );
nor ( n6756 , n142 , n6700 );
not ( n6757 , n6756 );
and ( n6758 , n6755 , n6757 );
not ( n6759 , n6755 );
and ( n6760 , n6759 , n6664 );
or ( n6761 , n6758 , n6760 );
nand ( n6762 , n141 , n6635 );
not ( n6763 , n140 );
nand ( n6764 , n6763 , n6547 );
not ( n6765 , n6764 );
nand ( n6766 , n142 , n6765 );
nand ( n6767 , n6761 , n6762 , n6766 );
and ( n6768 , n6754 , n6767 );
nor ( n6769 , n6753 , n6768 );
not ( n6770 , n140 );
not ( n6771 , n6683 );
nand ( n6772 , n6770 , n6771 );
not ( n6773 , n6772 );
not ( n6774 , n142 );
nand ( n6775 , n6773 , n6774 );
not ( n6776 , n6775 );
not ( n6777 , n6608 );
not ( n6778 , n6777 );
nand ( n6779 , n142 , n6778 );
not ( n6780 , n6779 );
or ( n6781 , n6776 , n6780 );
nand ( n6782 , n6781 , n141 );
not ( n6783 , n141 );
not ( n6784 , n6783 );
not ( n6785 , n6727 );
not ( n6786 , n142 );
not ( n6787 , n6563 );
not ( n6788 , n6787 );
not ( n6789 , n6788 );
nand ( n6790 , n6786 , n6789 );
nand ( n6791 , n6785 , n6567 , n6790 );
not ( n6792 , n6791 );
or ( n6793 , n6784 , n6792 );
not ( n6794 , n141 );
nor ( n6795 , n6794 , n142 );
not ( n6796 , n6737 );
nand ( n6797 , n140 , n6796 );
not ( n6798 , n6797 );
nand ( n6799 , n6795 , n6798 );
nand ( n6800 , n6793 , n6799 );
nand ( n6801 , n141 , n6701 );
nand ( n6802 , n142 , n6717 );
nand ( n6803 , n6801 , n6802 );
or ( n6804 , n6800 , n6803 );
nand ( n6805 , n6804 , n144 );
nand ( n6806 , n6769 , n6782 , n6805 );
or ( n6807 , n6806 , n6678 );
not ( n6808 , n137 );
nand ( n6809 , n6807 , n6808 );
nand ( n6810 , n6667 , n6713 , n6746 , n6809 );
not ( n6811 , n6810 );
not ( n6812 , n6811 );
not ( n6813 , n134 );
not ( n6814 , n6813 );
not ( n6815 , n133 );
not ( n6816 , n132 );
not ( n6817 , n129 );
nor ( n6818 , n128 , n130 );
nand ( n6819 , n6817 , n6818 );
not ( n6820 , n6819 );
not ( n6821 , n6820 );
not ( n6822 , n131 );
nor ( n6823 , n6821 , n6822 );
nand ( n6824 , n6816 , n6823 );
or ( n6825 , n6815 , n6824 );
not ( n6826 , n133 );
nor ( n6827 , n6826 , n132 );
not ( n6828 , n128 );
nor ( n6829 , n6828 , n130 );
nand ( n6830 , n6829 , n6817 );
not ( n6831 , n6830 );
nand ( n6832 , n6831 , n6822 );
not ( n6833 , n6832 );
nand ( n6834 , n6827 , n6833 );
nand ( n6835 , n6825 , n6834 );
not ( n6836 , n6835 );
or ( n6837 , n6814 , n6836 );
not ( n6838 , n133 );
nand ( n6839 , n131 , n132 );
not ( n6840 , n6839 );
not ( n6841 , n128 );
nand ( n6842 , n130 , n6841 );
not ( n6843 , n6842 );
nand ( n6844 , n6817 , n6843 );
not ( n6845 , n6844 );
nand ( n6846 , n6840 , n6845 );
or ( n6847 , n6838 , n6846 );
nand ( n6848 , n6837 , n6847 );
not ( n6849 , n134 );
nor ( n6850 , n128 , n129 );
nand ( n6851 , n131 , n6850 );
not ( n6852 , n6851 );
not ( n6853 , n6852 );
not ( n6854 , n6829 );
nor ( n6855 , n6854 , n131 );
not ( n6856 , n6855 );
nand ( n6857 , n129 , n130 );
nor ( n6858 , n128 , n6857 );
nand ( n6859 , n6822 , n6858 );
and ( n6860 , n6853 , n6856 , n6859 );
not ( n6861 , n6860 );
nor ( n6862 , n132 , n133 );
not ( n6863 , n6862 );
not ( n6864 , n6863 );
not ( n6865 , n6864 );
not ( n6866 , n6865 );
and ( n6867 , n6861 , n6866 );
nand ( n6868 , n128 , n129 );
not ( n6869 , n6868 );
not ( n6870 , n6869 );
not ( n6871 , n131 );
nand ( n6872 , n6871 , n132 );
not ( n6873 , n6872 );
not ( n6874 , n6873 );
or ( n6875 , n6870 , n6874 );
nand ( n6876 , n128 , n130 );
not ( n6877 , n6876 );
nand ( n6878 , n6877 , n6817 );
not ( n6879 , n6878 );
not ( n6880 , n6879 );
not ( n6881 , n6880 );
nand ( n6882 , n6881 , n132 );
nand ( n6883 , n6875 , n6882 );
and ( n6884 , n133 , n6883 );
nor ( n6885 , n6867 , n6884 );
nand ( n6886 , n131 , n6858 );
not ( n6887 , n6886 );
nand ( n6888 , n133 , n6887 );
nand ( n6889 , n6817 , n6843 );
nor ( n6890 , n131 , n6889 );
nand ( n6891 , n132 , n6890 );
or ( n6892 , n133 , n6891 );
nand ( n6893 , n6885 , n6888 , n6892 );
not ( n6894 , n6893 );
or ( n6895 , n6849 , n6894 );
not ( n6896 , n134 );
not ( n6897 , n133 );
not ( n6898 , n132 );
nor ( n6899 , n131 , n6876 );
not ( n6900 , n6899 );
nor ( n6901 , n6898 , n6900 );
nand ( n6902 , n6896 , n6897 , n6901 );
nand ( n6903 , n6895 , n6902 );
nor ( n6904 , n6848 , n6903 );
nand ( n6905 , n132 , n133 );
not ( n6906 , n6905 );
not ( n6907 , n6880 );
nand ( n6908 , n6907 , n6822 );
not ( n6909 , n6908 );
nand ( n6910 , n6906 , n6909 );
not ( n6911 , n132 );
not ( n6912 , n6830 );
nand ( n6913 , n6912 , n131 );
or ( n6914 , n6911 , n6913 );
not ( n6915 , n131 );
not ( n6916 , n6889 );
not ( n6917 , n6916 );
nand ( n6918 , n6917 , n6830 );
not ( n6919 , n6918 );
or ( n6920 , n6915 , n6919 );
not ( n6921 , n132 );
not ( n6922 , n6843 );
nor ( n6923 , n6921 , n6922 );
nand ( n6924 , n131 , n6923 );
nand ( n6925 , n6920 , n6924 );
and ( n6926 , n133 , n6925 );
not ( n6927 , n133 );
not ( n6928 , n132 );
nand ( n6929 , n6928 , n6887 );
nand ( n6930 , n128 , n130 );
not ( n6931 , n6930 );
nand ( n6932 , n6931 , n129 );
not ( n6933 , n6932 );
nand ( n6934 , n132 , n6933 );
not ( n6935 , n132 );
not ( n6936 , n129 );
nand ( n6937 , n6936 , n130 );
nor ( n6938 , n6937 , n131 );
nand ( n6939 , n6935 , n6938 );
and ( n6940 , n6934 , n6939 );
nand ( n6941 , n6929 , n6940 );
and ( n6942 , n6927 , n6941 );
nor ( n6943 , n6926 , n6942 );
not ( n6944 , n6887 );
not ( n6945 , n133 );
nor ( n6946 , n132 , n6854 );
nand ( n6947 , n6945 , n6946 );
and ( n6948 , n6944 , n6947 );
not ( n6949 , n132 );
not ( n6950 , n131 );
buf ( n6951 , n6857 );
nor ( n6952 , n6950 , n6951 );
nand ( n6953 , n6949 , n6952 );
buf ( n6954 , n6953 );
not ( n6955 , n6820 );
not ( n6956 , n6955 );
not ( n6957 , n133 );
nand ( n6958 , n6956 , n6957 );
nand ( n6959 , n6948 , n6954 , n6958 );
not ( n6960 , n133 );
not ( n6961 , n129 );
nor ( n6962 , n6961 , n128 );
not ( n6963 , n6962 );
or ( n6964 , n132 , n6963 );
not ( n6965 , n6858 );
not ( n6966 , n6965 );
not ( n6967 , n6966 );
buf ( n6968 , n6937 );
nor ( n6969 , n6822 , n6968 );
not ( n6970 , n6969 );
nand ( n6971 , n6964 , n6967 , n6970 );
not ( n6972 , n6971 );
or ( n6973 , n6960 , n6972 );
nand ( n6974 , n6973 , n6882 );
or ( n6975 , n6959 , n6974 );
nand ( n6976 , n6975 , n134 );
not ( n6977 , n132 );
nand ( n6978 , n128 , n129 );
nor ( n6979 , n6978 , n130 );
not ( n6980 , n6979 );
not ( n6981 , n6980 );
nand ( n6982 , n6822 , n6981 );
nor ( n6983 , n6977 , n6982 );
not ( n6984 , n6983 );
not ( n6985 , n134 );
not ( n6986 , n132 );
nor ( n6987 , n128 , n130 );
not ( n6988 , n6987 );
nor ( n6989 , n6988 , n131 );
nand ( n6990 , n6986 , n6989 );
not ( n6991 , n6990 );
not ( n6992 , n133 );
not ( n6993 , n132 );
nor ( n6994 , n6993 , n6844 );
not ( n6995 , n6994 );
nor ( n6996 , n6992 , n6995 );
nor ( n6997 , n6991 , n6996 );
not ( n6998 , n6980 );
nand ( n6999 , n133 , n6998 );
not ( n7000 , n133 );
nand ( n7001 , n132 , n7000 );
not ( n7002 , n7001 );
not ( n7003 , n7002 );
not ( n7004 , n6830 );
not ( n7005 , n7004 );
or ( n7006 , n7003 , n7005 );
nand ( n7007 , n6862 , n6879 );
nand ( n7008 , n7006 , n7007 );
not ( n7009 , n130 );
nand ( n7010 , n7009 , n129 );
nor ( n7011 , n131 , n7010 );
nand ( n7012 , n133 , n7011 );
nor ( n7013 , n131 , n132 );
nand ( n7014 , n6869 , n7013 );
nand ( n7015 , n7012 , n7014 , n6846 );
nor ( n7016 , n7008 , n7015 );
nand ( n7017 , n6997 , n6999 , n7016 );
nand ( n7018 , n6985 , n7017 );
nand ( n7019 , n6943 , n6976 , n6984 , n7018 );
and ( n7020 , n135 , n7019 );
not ( n7021 , n135 );
not ( n7022 , n132 );
not ( n7023 , n7022 );
not ( n7024 , n6833 );
or ( n7025 , n7023 , n7024 );
not ( n7026 , n131 );
nor ( n7027 , n129 , n130 );
nand ( n7028 , n7026 , n7027 );
not ( n7029 , n7028 );
nand ( n7030 , n6906 , n7029 );
nand ( n7031 , n7025 , n7030 );
not ( n7032 , n133 );
not ( n7033 , n7032 );
nand ( n7034 , n131 , n6829 );
not ( n7035 , n7034 );
nand ( n7036 , n132 , n7035 );
not ( n7037 , n6932 );
nand ( n7038 , n7037 , n131 );
not ( n7039 , n7038 );
not ( n7040 , n132 );
nand ( n7041 , n7039 , n7040 );
nand ( n7042 , n7036 , n7041 );
not ( n7043 , n7042 );
or ( n7044 , n7033 , n7043 );
not ( n7045 , n6932 );
nand ( n7046 , n7045 , n6822 );
not ( n7047 , n7046 );
nand ( n7048 , n133 , n7047 );
nand ( n7049 , n7044 , n7048 );
nor ( n7050 , n7031 , n7049 );
not ( n7051 , n134 );
not ( n7052 , n6823 );
nand ( n7053 , n7002 , n6887 );
nand ( n7054 , n133 , n131 , n6987 );
not ( n7055 , n6876 );
not ( n7056 , n6951 );
or ( n7057 , n7055 , n7056 );
nand ( n7058 , n7057 , n6827 );
and ( n7059 , n7054 , n7058 );
nand ( n7060 , n6939 , n7052 , n7053 , n7059 );
and ( n7061 , n7051 , n7060 );
not ( n7062 , n7051 );
not ( n7063 , n133 );
not ( n7064 , n6859 );
nand ( n7065 , n7063 , n7064 );
not ( n7066 , n6994 );
not ( n7067 , n7038 );
nand ( n7068 , n7067 , n132 );
nand ( n7069 , n7065 , n7066 , n7068 );
not ( n7070 , n7069 );
not ( n7071 , n132 );
nand ( n7072 , n7071 , n7047 );
not ( n7073 , n7028 );
not ( n7074 , n132 );
nand ( n7075 , n131 , n6979 );
not ( n7076 , n7075 );
nand ( n7077 , n7074 , n7076 );
not ( n7078 , n7077 );
or ( n7079 , n7073 , n7078 );
nand ( n7080 , n7079 , n133 );
nand ( n7081 , n7072 , n7080 );
not ( n7082 , n7081 );
nand ( n7083 , n7070 , n7082 );
and ( n7084 , n7062 , n7083 );
nor ( n7085 , n7061 , n7084 );
nand ( n7086 , n7050 , n7085 );
and ( n7087 , n7021 , n7086 );
nor ( n7088 , n7020 , n7087 );
and ( n7089 , n6904 , n6910 , n6914 , n7088 );
not ( n7090 , n7089 );
or ( n7091 , n6812 , n7090 );
nand ( n7092 , n6667 , n6713 , n6746 , n6809 );
not ( n7093 , n7092 );
not ( n7094 , n6904 );
nor ( n7095 , n7031 , n7049 );
not ( n7096 , n7095 );
not ( n7097 , n7085 );
or ( n7098 , n7096 , n7097 );
not ( n7099 , n135 );
nand ( n7100 , n7098 , n7099 );
not ( n7101 , n6943 );
nand ( n7102 , n6976 , n6984 , n7018 );
or ( n7103 , n7101 , n7102 );
nand ( n7104 , n7103 , n135 );
nand ( n7105 , n6910 , n6914 , n7100 , n7104 );
nor ( n7106 , n7094 , n7105 );
buf ( n7107 , n7106 );
or ( n7108 , n7093 , n7107 );
nand ( n7109 , n7091 , n7108 );
nand ( n7110 , n133 , n6820 );
not ( n7111 , n7110 );
nand ( n7112 , n6906 , n6969 );
not ( n7113 , n7112 );
or ( n7114 , n7111 , n7113 );
not ( n7115 , n134 );
nand ( n7116 , n7114 , n7115 );
not ( n7117 , n132 );
nand ( n7118 , n7117 , n6933 );
not ( n7119 , n7118 );
not ( n7120 , n132 );
nand ( n7121 , n7120 , n7011 );
not ( n7122 , n7121 );
or ( n7123 , n7119 , n7122 );
not ( n7124 , n133 );
nand ( n7125 , n7123 , n7124 );
not ( n7126 , n7038 );
nand ( n7127 , n129 , n6818 );
not ( n7128 , n7127 );
nand ( n7129 , n7128 , n131 );
not ( n7130 , n7129 );
or ( n7131 , n7126 , n7130 );
nand ( n7132 , n7131 , n6906 );
and ( n7133 , n7116 , n7125 , n7132 );
nand ( n7134 , n6822 , n6820 );
nor ( n7135 , n6905 , n7134 );
not ( n7136 , n133 );
nand ( n7137 , n7136 , n130 , n6822 );
nor ( n7138 , n131 , n6951 );
nand ( n7139 , n132 , n7138 );
and ( n7140 , n7137 , n7139 );
nor ( n7141 , n7140 , n134 );
nor ( n7142 , n7135 , n7141 );
not ( n7143 , n7052 );
not ( n7144 , n7075 );
nand ( n7145 , n132 , n7144 );
not ( n7146 , n7145 );
or ( n7147 , n7143 , n7146 );
not ( n7148 , n133 );
nand ( n7149 , n7147 , n7148 );
not ( n7150 , n6965 );
nand ( n7151 , n7150 , n132 );
not ( n7152 , n6878 );
nand ( n7153 , n7152 , n131 );
not ( n7154 , n7153 );
not ( n7155 , n132 );
nand ( n7156 , n7154 , n7155 );
nand ( n7157 , n7151 , n7156 );
not ( n7158 , n133 );
not ( n7159 , n7158 );
not ( n7160 , n6841 );
not ( n7161 , n6840 );
or ( n7162 , n7160 , n7161 );
nand ( n7163 , n132 , n7004 );
nand ( n7164 , n7162 , n7163 );
not ( n7165 , n7164 );
or ( n7166 , n7159 , n7165 );
not ( n7167 , n131 );
not ( n7168 , n129 );
nand ( n7169 , n7168 , n128 );
nor ( n7170 , n7167 , n7169 );
nand ( n7171 , n6827 , n7170 );
nand ( n7172 , n7166 , n7171 );
or ( n7173 , n7157 , n7172 );
nand ( n7174 , n7173 , n134 );
and ( n7175 , n7133 , n7142 , n7149 , n7174 );
or ( n7176 , n7175 , n135 );
not ( n7177 , n134 );
and ( n7178 , n133 , n7177 );
not ( n7179 , n132 );
not ( n7180 , n131 );
nor ( n7181 , n7180 , n6868 );
nand ( n7182 , n7179 , n7181 );
not ( n7183 , n6820 );
not ( n7184 , n7183 );
nand ( n7185 , n7184 , n132 );
buf ( n7186 , n7185 );
not ( n7187 , n7153 );
nand ( n7188 , n7187 , n132 );
not ( n7189 , n7188 );
not ( n7190 , n7189 );
nand ( n7191 , n7182 , n7186 , n7190 );
nand ( n7192 , n7178 , n7191 );
nand ( n7193 , n7176 , n7192 );
not ( n7194 , n135 );
and ( n7195 , n133 , n134 );
not ( n7196 , n6841 );
not ( n7197 , n131 );
and ( n7198 , n7196 , n7197 );
not ( n7199 , n6854 );
and ( n7200 , n7199 , n132 );
nor ( n7201 , n7198 , n7200 );
not ( n7202 , n132 );
nand ( n7203 , n7202 , n6987 );
nand ( n7204 , n7201 , n6853 , n7203 );
nand ( n7205 , n7195 , n7204 );
not ( n7206 , n7010 );
not ( n7207 , n131 );
nor ( n7208 , n7207 , n132 );
nand ( n7209 , n7206 , n7208 );
not ( n7210 , n7188 );
nand ( n7211 , n6862 , n6916 );
not ( n7212 , n7211 );
or ( n7213 , n7210 , n7212 );
nand ( n7214 , n7213 , n134 );
nand ( n7215 , n7205 , n7209 , n7214 );
not ( n7216 , n7215 );
not ( n7217 , n133 );
not ( n7218 , n132 );
nand ( n7219 , n7218 , n6899 );
not ( n7220 , n7144 );
not ( n7221 , n132 );
nor ( n7222 , n6822 , n6963 );
nand ( n7223 , n7221 , n7222 );
nand ( n7224 , n7219 , n7220 , n7223 );
not ( n7225 , n7224 );
or ( n7226 , n7217 , n7225 );
not ( n7227 , n131 );
not ( n7228 , n128 );
nor ( n7229 , n7228 , n129 );
nand ( n7230 , n7227 , n7229 );
not ( n7231 , n7230 );
nand ( n7232 , n6906 , n7231 );
nand ( n7233 , n7226 , n7232 );
not ( n7234 , n7233 );
not ( n7235 , n134 );
not ( n7236 , n132 );
nand ( n7237 , n7236 , n7035 );
nand ( n7238 , n7237 , n6947 );
nand ( n7239 , n6827 , n6938 );
nor ( n7240 , n133 , n6980 );
not ( n7241 , n132 );
not ( n7242 , n131 );
nand ( n7243 , n7242 , n6962 );
nor ( n7244 , n7241 , n7243 );
nor ( n7245 , n7240 , n7244 );
not ( n7246 , n7034 );
not ( n7247 , n6851 );
nor ( n7248 , n7247 , n7181 );
not ( n7249 , n7248 );
or ( n7250 , n7246 , n7249 );
not ( n7251 , n133 );
nand ( n7252 , n7250 , n7251 );
nand ( n7253 , n7239 , n7245 , n7252 );
nor ( n7254 , n7238 , n7253 );
not ( n7255 , n7254 );
and ( n7256 , n7235 , n7255 );
not ( n7257 , n133 );
not ( n7258 , n7237 );
not ( n7259 , n7258 );
not ( n7260 , n7259 );
and ( n7261 , n7257 , n7260 );
nor ( n7262 , n7256 , n7261 );
nand ( n7263 , n7216 , n7234 , n7262 );
not ( n7264 , n7263 );
or ( n7265 , n7194 , n7264 );
not ( n7266 , n134 );
not ( n7267 , n7266 );
not ( n7268 , n133 );
nand ( n7269 , n7268 , n132 , n6938 );
nand ( n7270 , n7269 , n6954 , n7125 );
not ( n7271 , n7270 );
or ( n7272 , n7267 , n7271 );
nand ( n7273 , n7013 , n6998 );
not ( n7274 , n7273 );
not ( n7275 , n6955 );
nand ( n7276 , n6840 , n7275 );
not ( n7277 , n7276 );
or ( n7278 , n7274 , n7277 );
not ( n7279 , n133 );
nand ( n7280 , n7278 , n7279 );
nand ( n7281 , n7272 , n7280 );
not ( n7282 , n7281 );
not ( n7283 , n132 );
buf ( n7284 , n7127 );
nor ( n7285 , n7283 , n7284 );
not ( n7286 , n7285 );
not ( n7287 , n7286 );
not ( n7288 , n7222 );
not ( n7289 , n7288 );
nand ( n7290 , n7046 , n6832 );
not ( n7291 , n7290 );
not ( n7292 , n7291 );
or ( n7293 , n7289 , n7292 );
nand ( n7294 , n7293 , n132 );
not ( n7295 , n7294 );
or ( n7296 , n7287 , n7295 );
not ( n7297 , n134 );
nor ( n7298 , n7297 , n133 );
nand ( n7299 , n7296 , n7298 );
not ( n7300 , n132 );
not ( n7301 , n7300 );
nor ( n7302 , n6822 , n6889 );
not ( n7303 , n7302 );
not ( n7304 , n7127 );
nand ( n7305 , n7304 , n6822 );
nand ( n7306 , n6900 , n7303 , n7305 );
not ( n7307 , n7306 );
or ( n7308 , n7301 , n7307 );
nand ( n7309 , n132 , n6998 );
and ( n7310 , n7309 , n6908 );
nand ( n7311 , n7308 , n7310 );
nand ( n7312 , n7195 , n7311 );
nand ( n7313 , n7282 , n7299 , n7312 );
not ( n7314 , n7313 );
nand ( n7315 , n7265 , n7314 );
nor ( n7316 , n7193 , n7315 );
buf ( n7317 , n7316 );
xor ( n7318 , n6532 , n7317 );
not ( n7319 , n7318 );
and ( n7320 , n7109 , n7319 );
not ( n7321 , n7109 );
and ( n7322 , n7321 , n7318 );
nor ( n7323 , n7320 , n7322 );
not ( n7324 , n7323 );
not ( n7325 , n119 );
not ( n7326 , n7325 );
not ( n7327 , n117 );
not ( n7328 , n7327 );
not ( n7329 , n112 );
not ( n7330 , n113 );
nand ( n7331 , n7330 , n114 );
not ( n7332 , n7331 );
nand ( n7333 , n7329 , n7332 );
not ( n7334 , n7333 );
nand ( n7335 , n7334 , n115 );
nor ( n7336 , n116 , n7335 );
not ( n7337 , n7336 );
not ( n7338 , n7337 );
not ( n7339 , n7338 );
or ( n7340 , n7328 , n7339 );
not ( n7341 , n114 );
nand ( n7342 , n7341 , n113 );
not ( n7343 , n7342 );
nand ( n7344 , n112 , n7343 );
not ( n7345 , n7344 );
not ( n7346 , n7345 );
not ( n7347 , n7346 );
nor ( n7348 , n115 , n116 );
buf ( n7349 , n7348 );
nand ( n7350 , n7347 , n7349 );
nand ( n7351 , n7340 , n7350 );
not ( n7352 , n7351 );
nand ( n7353 , n113 , n114 );
not ( n7354 , n7353 );
nand ( n7355 , n7354 , n112 );
not ( n7356 , n7355 );
not ( n7357 , n7356 );
not ( n7358 , n7357 );
nand ( n7359 , n7358 , n117 );
buf ( n7360 , n7353 );
not ( n7361 , n7360 );
nand ( n7362 , n7361 , n115 );
not ( n7363 , n7362 );
nand ( n7364 , n116 , n7363 );
nand ( n7365 , n7359 , n7364 );
not ( n7366 , n117 );
not ( n7367 , n7366 );
not ( n7368 , n116 );
nor ( n7369 , n113 , n114 );
nand ( n7370 , n112 , n7369 );
not ( n7371 , n7370 );
nand ( n7372 , n7368 , n7371 );
not ( n7373 , n7370 );
nand ( n7374 , n7373 , n115 );
buf ( n7375 , n7374 );
nor ( n7376 , n113 , n114 );
nand ( n7377 , n7329 , n7376 );
not ( n7378 , n7377 );
not ( n7379 , n115 );
nand ( n7380 , n7378 , n7379 );
not ( n7381 , n7380 );
not ( n7382 , n7381 );
nand ( n7383 , n7372 , n7375 , n7382 );
not ( n7384 , n7383 );
or ( n7385 , n7367 , n7384 );
not ( n7386 , n116 );
nand ( n7387 , n7386 , n117 );
not ( n7388 , n7387 );
nor ( n7389 , n112 , n113 );
nand ( n7390 , n115 , n7389 );
not ( n7391 , n7390 );
nand ( n7392 , n7388 , n7391 );
nand ( n7393 , n7385 , n7392 );
or ( n7394 , n7365 , n7393 );
nand ( n7395 , n7394 , n118 );
not ( n7396 , n116 );
not ( n7397 , n7396 );
not ( n7398 , n115 );
not ( n7399 , n114 );
nor ( n7400 , n7399 , n112 );
nand ( n7401 , n7398 , n7400 );
not ( n7402 , n7401 );
not ( n7403 , n7402 );
or ( n7404 , n7397 , n7403 );
not ( n7405 , n7342 );
nand ( n7406 , n7405 , n7329 );
not ( n7407 , n7406 );
nand ( n7408 , n115 , n7407 );
not ( n7409 , n7408 );
nand ( n7410 , n116 , n7409 );
nand ( n7411 , n7404 , n7410 );
and ( n7412 , n117 , n7411 );
not ( n7413 , n7407 );
not ( n7414 , n117 );
nor ( n7415 , n7413 , n7414 );
not ( n7416 , n116 );
not ( n7417 , n115 );
and ( n7418 , n7417 , n7343 );
not ( n7419 , n7418 );
nor ( n7420 , n7416 , n7419 );
nor ( n7421 , n7415 , n7420 );
not ( n7422 , n117 );
not ( n7423 , n7355 );
not ( n7424 , n116 );
nand ( n7425 , n7423 , n7424 );
not ( n7426 , n7425 );
not ( n7427 , n7426 );
and ( n7428 , n7422 , n7427 );
not ( n7429 , n7422 );
nand ( n7430 , n112 , n114 );
not ( n7431 , n7430 );
nand ( n7432 , n115 , n7431 );
and ( n7433 , n7429 , n7432 );
or ( n7434 , n7428 , n7433 );
and ( n7435 , n7421 , n7434 );
nor ( n7436 , n7435 , n118 );
nor ( n7437 , n7412 , n7436 );
nand ( n7438 , n7352 , n7395 , n7437 );
not ( n7439 , n7438 );
or ( n7440 , n7326 , n7439 );
not ( n7441 , n7335 );
nand ( n7442 , n116 , n7441 );
not ( n7443 , n7442 );
not ( n7444 , n7381 );
not ( n7445 , n116 );
nor ( n7446 , n7444 , n7445 );
nor ( n7447 , n7443 , n7446 );
not ( n7448 , n7447 );
not ( n7449 , n117 );
not ( n7450 , n7400 );
not ( n7451 , n7389 );
nand ( n7452 , n7450 , n7451 );
nand ( n7453 , n116 , n7452 );
not ( n7454 , n115 );
not ( n7455 , n112 );
nor ( n7456 , n7455 , n7331 );
nand ( n7457 , n7454 , n7456 );
nor ( n7458 , n116 , n7457 );
not ( n7459 , n7458 );
not ( n7460 , n7406 );
nand ( n7461 , n7460 , n7349 );
nand ( n7462 , n7453 , n7459 , n7461 );
nand ( n7463 , n7449 , n7462 );
not ( n7464 , n7463 );
or ( n7465 , n7448 , n7464 );
nand ( n7466 , n7465 , n118 );
nand ( n7467 , n115 , n116 );
not ( n7468 , n7467 );
nand ( n7469 , n117 , n7431 , n7468 );
not ( n7470 , n117 );
not ( n7471 , n116 );
nand ( n7472 , n7471 , n7363 );
not ( n7473 , n7472 );
not ( n7474 , n7473 );
or ( n7475 , n7470 , n7474 );
not ( n7476 , n7346 );
not ( n7477 , n7476 );
nand ( n7478 , n116 , n117 );
nor ( n7479 , n7477 , n7478 );
not ( n7480 , n7479 );
nand ( n7481 , n7475 , n7480 );
and ( n7482 , n118 , n7481 );
not ( n7483 , n117 );
nand ( n7484 , n116 , n7483 );
not ( n7485 , n7484 );
not ( n7486 , n7353 );
nand ( n7487 , n7486 , n7329 );
not ( n7488 , n7487 );
not ( n7489 , n115 );
and ( n7490 , n7488 , n7489 );
and ( n7491 , n7485 , n7490 );
nor ( n7492 , n7482 , n7491 );
nand ( n7493 , n7466 , n7469 , n7492 );
not ( n7494 , n7493 );
nand ( n7495 , n7440 , n7494 );
not ( n7496 , n119 );
not ( n7497 , n116 );
nor ( n7498 , n7497 , n115 );
not ( n7499 , n7498 );
or ( n7500 , n114 , n7499 );
not ( n7501 , n7377 );
nand ( n7502 , n116 , n7501 );
not ( n7503 , n7502 );
not ( n7504 , n7503 );
nand ( n7505 , n7500 , n7504 );
nand ( n7506 , n117 , n7505 );
not ( n7507 , n113 );
not ( n7508 , n116 );
nand ( n7509 , n7508 , n115 );
not ( n7510 , n7509 );
not ( n7511 , n7510 );
not ( n7512 , n7511 );
not ( n7513 , n7512 );
or ( n7514 , n7507 , n7513 );
nand ( n7515 , n7514 , n7457 );
and ( n7516 , n117 , n7515 );
not ( n7517 , n117 );
nor ( n7518 , n115 , n7360 );
nand ( n7519 , n116 , n7518 );
not ( n7520 , n7333 );
nand ( n7521 , n7520 , n116 );
not ( n7522 , n7521 );
not ( n7523 , n7522 );
nand ( n7524 , n7461 , n7519 , n7523 );
and ( n7525 , n7517 , n7524 );
nor ( n7526 , n7516 , n7525 );
not ( n7527 , n118 );
not ( n7528 , n117 );
not ( n7529 , n115 );
not ( n7530 , n112 );
nor ( n7531 , n7530 , n113 );
nand ( n7532 , n7529 , n7531 );
not ( n7533 , n7532 );
nand ( n7534 , n7528 , n7533 );
nand ( n7535 , n116 , n7531 );
not ( n7536 , n117 );
not ( n7537 , n7467 );
nand ( n7538 , n7537 , n7343 );
not ( n7539 , n7538 );
nand ( n7540 , n7536 , n7539 );
and ( n7541 , n7534 , n7535 , n7540 );
not ( n7542 , n7332 );
nor ( n7543 , n115 , n7542 );
nand ( n7544 , n116 , n7543 );
not ( n7545 , n7375 );
nand ( n7546 , n117 , n7545 );
nand ( n7547 , n7541 , n7544 , n7546 );
and ( n7548 , n7527 , n7547 );
not ( n7549 , n7527 );
not ( n7550 , n115 );
and ( n7551 , n7550 , n7376 );
nand ( n7552 , n117 , n7551 );
not ( n7553 , n7552 );
not ( n7554 , n116 );
not ( n7555 , n115 );
nand ( n7556 , n7555 , n7345 );
nor ( n7557 , n7554 , n7556 );
nor ( n7558 , n7553 , n7557 );
not ( n7559 , n7408 );
not ( n7560 , n116 );
nand ( n7561 , n7559 , n7560 );
not ( n7562 , n7518 );
not ( n7563 , n7562 );
not ( n7564 , n7377 );
nand ( n7565 , n115 , n7564 );
not ( n7566 , n7565 );
not ( n7567 , n7566 );
not ( n7568 , n7567 );
or ( n7569 , n7563 , n7568 );
not ( n7570 , n117 );
nand ( n7571 , n7569 , n7570 );
nand ( n7572 , n7558 , n7561 , n7571 );
and ( n7573 , n7549 , n7572 );
nor ( n7574 , n7548 , n7573 );
nand ( n7575 , n7506 , n7526 , n7574 );
not ( n7576 , n7575 );
or ( n7577 , n7496 , n7576 );
not ( n7578 , n7355 );
nand ( n7579 , n7578 , n115 );
not ( n7580 , n7579 );
nand ( n7581 , n7580 , n116 );
and ( n7582 , n7581 , n7350 );
not ( n7583 , n7582 );
not ( n7584 , n117 );
nand ( n7585 , n115 , n7400 );
or ( n7586 , n116 , n7585 );
not ( n7587 , n7457 );
nand ( n7588 , n116 , n7587 );
buf ( n7589 , n7588 );
not ( n7590 , n116 );
nand ( n7591 , n7590 , n7520 );
not ( n7592 , n7591 );
not ( n7593 , n7592 );
nand ( n7594 , n7586 , n7589 , n7593 );
and ( n7595 , n7584 , n7594 );
not ( n7596 , n7584 );
not ( n7597 , n116 );
nand ( n7598 , n7597 , n7345 );
not ( n7599 , n7598 );
not ( n7600 , n116 );
not ( n7601 , n112 );
nor ( n7602 , n7601 , n115 , n114 );
not ( n7603 , n7602 );
nor ( n7604 , n7600 , n7603 );
nor ( n7605 , n7599 , n7604 );
not ( n7606 , n7356 );
not ( n7607 , n116 );
nor ( n7608 , n7606 , n7607 );
not ( n7609 , n7608 );
nand ( n7610 , n116 , n7566 );
not ( n7611 , n7382 );
not ( n7612 , n116 );
nand ( n7613 , n7611 , n7612 );
nand ( n7614 , n7605 , n7609 , n7610 , n7613 );
and ( n7615 , n7596 , n7614 );
nor ( n7616 , n7595 , n7615 );
not ( n7617 , n7616 );
or ( n7618 , n7583 , n7617 );
not ( n7619 , n118 );
nand ( n7620 , n7618 , n7619 );
nand ( n7621 , n7577 , n7620 );
nor ( n7622 , n7495 , n7621 );
not ( n7623 , n127 );
nand ( n7624 , n123 , n124 );
nor ( n7625 , n7624 , n122 );
not ( n7626 , n7625 );
not ( n7627 , n7626 );
nand ( n7628 , n7627 , n121 );
not ( n7629 , n7628 );
not ( n7630 , n7629 );
not ( n7631 , n124 );
not ( n7632 , n121 );
nand ( n7633 , n7632 , n125 );
buf ( n7634 , n7633 );
not ( n7635 , n7634 );
and ( n7636 , n7631 , n7635 );
not ( n7637 , n125 );
not ( n7638 , n123 );
nand ( n7639 , n7637 , n121 , n7638 );
not ( n7640 , n7639 );
nor ( n7641 , n7636 , n7640 );
not ( n7642 , n125 );
not ( n7643 , n123 );
nand ( n7644 , n7643 , n122 , n124 );
nor ( n7645 , n7642 , n7644 );
not ( n7646 , n7645 );
buf ( n7647 , n7646 );
nand ( n7648 , n7630 , n7641 , n7647 );
and ( n7649 , n120 , n7648 );
not ( n7650 , n120 );
nor ( n7651 , n123 , n124 );
buf ( n7652 , n7651 );
nand ( n7653 , n7652 , n125 );
not ( n7654 , n121 );
nor ( n7655 , n7653 , n7654 );
not ( n7656 , n7655 );
not ( n7657 , n121 );
not ( n7658 , n123 );
not ( n7659 , n122 );
nand ( n7660 , n7658 , n7659 , n124 );
not ( n7661 , n7660 );
not ( n7662 , n7661 );
nor ( n7663 , n7657 , n7662 );
not ( n7664 , n7663 );
not ( n7665 , n123 );
nor ( n7666 , n7665 , n124 );
not ( n7667 , n7666 );
nand ( n7668 , n7667 , n7659 );
not ( n7669 , n7668 );
not ( n7670 , n7633 );
nand ( n7671 , n7669 , n7670 );
nand ( n7672 , n7656 , n7664 , n7671 );
and ( n7673 , n7650 , n7672 );
nor ( n7674 , n7649 , n7673 );
not ( n7675 , n121 );
not ( n7676 , n124 );
nor ( n7677 , n7676 , n123 );
nand ( n7678 , n7642 , n7677 );
nor ( n7679 , n7675 , n7678 );
not ( n7680 , n124 );
nand ( n7681 , n7680 , n123 );
not ( n7682 , n7681 );
nor ( n7683 , n7682 , n125 );
nand ( n7684 , n121 , n7683 );
nor ( n7685 , n120 , n7684 );
nor ( n7686 , n7679 , n7685 );
not ( n7687 , n120 );
not ( n7688 , n125 );
nand ( n7689 , n122 , n124 );
not ( n7690 , n7689 );
nand ( n7691 , n7688 , n7690 );
not ( n7692 , n7691 );
nand ( n7693 , n7687 , n7692 );
not ( n7694 , n121 );
not ( n7695 , n7690 );
nor ( n7696 , n7694 , n7695 );
not ( n7697 , n120 );
not ( n7698 , n122 );
nand ( n7699 , n123 , n124 );
nor ( n7700 , n7698 , n7699 );
nand ( n7701 , n125 , n7700 );
not ( n7702 , n7701 );
not ( n7703 , n7702 );
nor ( n7704 , n7697 , n7703 );
nor ( n7705 , n7696 , n7704 );
nand ( n7706 , n7686 , n7693 , n7705 );
and ( n7707 , n126 , n7706 );
not ( n7708 , n126 );
not ( n7709 , n7653 );
nand ( n7710 , n125 , n7625 );
not ( n7711 , n7710 );
or ( n7712 , n7709 , n7711 );
not ( n7713 , n120 );
nand ( n7714 , n7712 , n7713 );
and ( n7715 , n7671 , n7714 );
not ( n7716 , n125 );
nor ( n7717 , n7716 , n7624 );
nand ( n7718 , n120 , n7717 );
not ( n7719 , n7666 );
nand ( n7720 , n7719 , n122 );
nor ( n7721 , n125 , n7720 );
and ( n7722 , n121 , n7721 );
not ( n7723 , n7722 );
nand ( n7724 , n7715 , n7718 , n7723 );
and ( n7725 , n7708 , n7724 );
nor ( n7726 , n7707 , n7725 );
nand ( n7727 , n7674 , n7726 );
not ( n7728 , n7727 );
or ( n7729 , n7623 , n7728 );
not ( n7730 , n122 );
nand ( n7731 , n7730 , n7652 );
not ( n7732 , n7731 );
not ( n7733 , n7732 );
not ( n7734 , n7733 );
nand ( n7735 , n7734 , n7642 );
not ( n7736 , n7735 );
not ( n7737 , n7736 );
or ( n7738 , n120 , n7737 );
nand ( n7739 , n122 , n123 );
not ( n7740 , n7739 );
nand ( n7741 , n7740 , n125 );
not ( n7742 , n7741 );
nand ( n7743 , n120 , n7742 );
nand ( n7744 , n7738 , n7743 );
nand ( n7745 , n121 , n7744 );
nand ( n7746 , n7729 , n7745 );
not ( n7747 , n7746 );
not ( n7748 , n127 );
not ( n7749 , n126 );
not ( n7750 , n120 );
nor ( n7751 , n7750 , n121 );
not ( n7752 , n7751 );
not ( n7753 , n125 );
not ( n7754 , n124 );
nor ( n7755 , n7754 , n122 );
nor ( n7756 , n7753 , n7755 );
not ( n7757 , n7756 );
or ( n7758 , n7752 , n7757 );
nand ( n7759 , n122 , n7651 );
not ( n7760 , n7759 );
nand ( n7761 , n7760 , n120 );
nand ( n7762 , n7758 , n7761 );
and ( n7763 , n7749 , n7762 );
not ( n7764 , n7720 );
not ( n7765 , n7764 );
nor ( n7766 , n7765 , n7634 );
nor ( n7767 , n7763 , n7766 );
not ( n7768 , n126 );
not ( n7769 , n125 );
nand ( n7770 , n7769 , n7652 );
not ( n7771 , n7770 );
nand ( n7772 , n7771 , n121 );
not ( n7773 , n7772 );
nand ( n7774 , n7768 , n7773 );
not ( n7775 , n7743 );
not ( n7776 , n7668 );
not ( n7777 , n7776 );
not ( n7778 , n7777 );
nand ( n7779 , n120 , n7778 );
not ( n7780 , n7779 );
or ( n7781 , n7775 , n7780 );
nand ( n7782 , n7781 , n126 );
nand ( n7783 , n7767 , n7774 , n7782 );
not ( n7784 , n7783 );
not ( n7785 , n120 );
not ( n7786 , n121 );
not ( n7787 , n7661 );
nor ( n7788 , n7642 , n7787 );
nand ( n7789 , n7786 , n7788 );
not ( n7790 , n7789 );
and ( n7791 , n7785 , n7790 );
not ( n7792 , n7785 );
not ( n7793 , n121 );
not ( n7794 , n7793 );
not ( n7795 , n125 );
not ( n7796 , n122 );
nand ( n7797 , n7796 , n123 );
nor ( n7798 , n7795 , n7797 );
not ( n7799 , n7798 );
or ( n7800 , n7794 , n7799 );
not ( n7801 , n7668 );
nand ( n7802 , n7801 , n7642 );
not ( n7803 , n7802 );
nand ( n7804 , n121 , n7803 );
nand ( n7805 , n7800 , n7804 );
and ( n7806 , n7792 , n7805 );
nor ( n7807 , n7791 , n7806 );
not ( n7808 , n126 );
not ( n7809 , n7808 );
not ( n7810 , n121 );
nand ( n7811 , n125 , n7681 );
nor ( n7812 , n7810 , n7811 );
nor ( n7813 , n120 , n121 );
not ( n7814 , n7759 );
and ( n7815 , n7813 , n7814 );
nor ( n7816 , n7812 , n7815 );
not ( n7817 , n7816 );
and ( n7818 , n7809 , n7817 );
or ( n7819 , n120 , n126 );
not ( n7820 , n7819 );
not ( n7821 , n121 );
buf ( n7822 , n7700 );
nand ( n7823 , n7821 , n7822 );
not ( n7824 , n7710 );
not ( n7825 , n7824 );
nand ( n7826 , n7823 , n7703 , n7825 );
and ( n7827 , n7820 , n7826 );
nor ( n7828 , n7818 , n7827 );
nand ( n7829 , n7784 , n7807 , n7828 );
nand ( n7830 , n7748 , n7829 );
not ( n7831 , n120 );
not ( n7832 , n7770 );
not ( n7833 , n121 );
nand ( n7834 , n7832 , n7833 );
or ( n7835 , n7831 , n7834 );
nand ( n7836 , n120 , n121 );
not ( n7837 , n7836 );
nand ( n7838 , n7837 , n7764 );
not ( n7839 , n121 );
nor ( n7840 , n7839 , n7710 );
not ( n7841 , n7840 );
nand ( n7842 , n7835 , n7838 , n7841 );
not ( n7843 , n120 );
not ( n7844 , n7843 );
nand ( n7845 , n7797 , n7755 );
nand ( n7846 , n121 , n7845 );
not ( n7847 , n121 );
not ( n7848 , n7646 );
nand ( n7849 , n7847 , n7848 );
not ( n7850 , n7849 );
not ( n7851 , n7850 );
nand ( n7852 , n7846 , n7671 , n7851 );
not ( n7853 , n7852 );
or ( n7854 , n7844 , n7853 );
nand ( n7855 , n121 , n7788 );
nand ( n7856 , n7854 , n7855 );
or ( n7857 , n7842 , n7856 );
not ( n7858 , n126 );
nand ( n7859 , n7857 , n7858 );
nor ( n7860 , n125 , n7759 );
nand ( n7861 , n121 , n7860 );
not ( n7862 , n7861 );
not ( n7863 , n7766 );
not ( n7864 , n7863 );
nor ( n7865 , n7862 , n7864 );
not ( n7866 , n7865 );
not ( n7867 , n7759 );
nand ( n7868 , n7867 , n121 );
nand ( n7869 , n121 , n125 );
not ( n7870 , n7869 );
not ( n7871 , n7633 );
or ( n7872 , n7870 , n7871 );
not ( n7873 , n7625 );
not ( n7874 , n7873 );
nand ( n7875 , n7872 , n7874 );
nand ( n7876 , n7868 , n7875 );
not ( n7877 , n7876 );
not ( n7878 , n7720 );
not ( n7879 , n7878 );
nor ( n7880 , n7879 , n121 );
not ( n7881 , n7880 );
not ( n7882 , n125 );
not ( n7883 , n123 );
nand ( n7884 , n7883 , n122 );
nor ( n7885 , n7882 , n7884 );
nand ( n7886 , n121 , n7885 );
nand ( n7887 , n7877 , n7881 , n7886 );
and ( n7888 , n120 , n7887 );
not ( n7889 , n120 );
not ( n7890 , n121 );
nor ( n7891 , n125 , n7797 );
nand ( n7892 , n7890 , n7891 );
not ( n7893 , n121 );
nand ( n7894 , n7893 , n7661 );
not ( n7895 , n7894 );
not ( n7896 , n7895 );
and ( n7897 , n121 , n7645 );
not ( n7898 , n7897 );
nand ( n7899 , n7892 , n7896 , n7898 );
and ( n7900 , n7889 , n7899 );
nor ( n7901 , n7888 , n7900 );
not ( n7902 , n7901 );
or ( n7903 , n7866 , n7902 );
nand ( n7904 , n7903 , n126 );
nand ( n7905 , n7830 , n7859 , n7904 );
not ( n7906 , n7905 );
nand ( n7907 , n7747 , n7906 );
and ( n7908 , n7622 , n7907 );
not ( n7909 , n7622 );
nor ( n7910 , n7746 , n7905 );
and ( n7911 , n7909 , n7910 );
nor ( n7912 , n7908 , n7911 );
not ( n7913 , n7912 );
not ( n7914 , n126 );
not ( n7915 , n120 );
not ( n7916 , n7756 );
not ( n7917 , n7916 );
nand ( n7918 , n7915 , n121 , n7917 );
not ( n7919 , n7691 );
not ( n7920 , n121 );
nand ( n7921 , n7919 , n7920 );
not ( n7922 , n121 );
not ( n7923 , n7644 );
nand ( n7924 , n7922 , n7923 );
not ( n7925 , n7924 );
not ( n7926 , n121 );
not ( n7927 , n124 );
nand ( n7928 , n7927 , n122 );
nor ( n7929 , n125 , n7928 );
nand ( n7930 , n7926 , n7929 );
not ( n7931 , n7930 );
or ( n7932 , n7925 , n7931 );
not ( n7933 , n120 );
nand ( n7934 , n7932 , n7933 );
nand ( n7935 , n7918 , n7921 , n7934 );
not ( n7936 , n7935 );
or ( n7937 , n7914 , n7936 );
not ( n7938 , n7804 );
not ( n7939 , n121 );
nor ( n7940 , n125 , n7759 );
nand ( n7941 , n7939 , n7940 );
not ( n7942 , n7941 );
or ( n7943 , n7938 , n7942 );
not ( n7944 , n120 );
nand ( n7945 , n7943 , n7944 );
nand ( n7946 , n7937 , n7945 );
not ( n7947 , n7946 );
nand ( n7948 , n120 , n126 );
not ( n7949 , n7948 );
not ( n7950 , n7742 );
or ( n7951 , n121 , n7950 );
not ( n7952 , n121 );
nor ( n7953 , n7952 , n7777 );
not ( n7954 , n7953 );
nand ( n7955 , n7951 , n7954 , n7855 );
nand ( n7956 , n7949 , n7955 );
not ( n7957 , n126 );
not ( n7958 , n120 );
not ( n7959 , n121 );
not ( n7960 , n7959 );
not ( n7961 , n7721 );
nand ( n7962 , n7678 , n7961 , n7710 );
not ( n7963 , n7962 );
or ( n7964 , n7960 , n7963 );
nand ( n7965 , n7642 , n7661 );
and ( n7966 , n7868 , n7965 );
nand ( n7967 , n7964 , n7966 );
not ( n7968 , n7967 );
or ( n7969 , n7958 , n7968 );
not ( n7970 , n120 );
nand ( n7971 , n121 , n7970 );
not ( n7972 , n7971 );
nor ( n7973 , n125 , n7884 );
not ( n7974 , n7973 );
not ( n7975 , n7764 );
nand ( n7976 , n7974 , n7975 , n7647 , n7735 );
nand ( n7977 , n7972 , n7976 );
nand ( n7978 , n7969 , n7977 );
nand ( n7979 , n7957 , n7978 );
nand ( n7980 , n7947 , n7956 , n7979 );
not ( n7981 , n7748 );
not ( n7982 , n126 );
not ( n7983 , n7836 );
not ( n7984 , n7983 );
not ( n7985 , n7756 );
or ( n7986 , n7984 , n7985 );
not ( n7987 , n120 );
or ( n7988 , n7987 , n7777 );
nand ( n7989 , n7986 , n7988 );
not ( n7990 , n7989 );
or ( n7991 , n7982 , n7990 );
not ( n7992 , n7836 );
not ( n7993 , n7776 );
nor ( n7994 , n7993 , n7642 );
nand ( n7995 , n7992 , n7994 );
nand ( n7996 , n7991 , n7995 );
not ( n7997 , n120 );
not ( n7998 , n7997 );
nand ( n7999 , n7802 , n7861 );
not ( n8000 , n7999 );
or ( n8001 , n7998 , n8000 );
nand ( n8002 , n8001 , n7934 );
nor ( n8003 , n7996 , n8002 );
not ( n8004 , n7992 );
not ( n8005 , n7764 );
nor ( n8006 , n8005 , n7642 );
not ( n8007 , n7647 );
nor ( n8008 , n8006 , n8007 );
or ( n8009 , n8004 , n8008 );
not ( n8010 , n125 );
nand ( n8011 , n8010 , n124 );
not ( n8012 , n8011 );
not ( n8013 , n120 );
nand ( n8014 , n8012 , n8013 );
not ( n8015 , n8014 );
not ( n8016 , n7691 );
nand ( n8017 , n8016 , n121 );
not ( n8018 , n8017 );
or ( n8019 , n8015 , n8018 );
nand ( n8020 , n8019 , n126 );
nand ( n8021 , n8009 , n8020 );
not ( n8022 , n8021 );
not ( n8023 , n126 );
not ( n8024 , n7751 );
not ( n8025 , n7891 );
or ( n8026 , n8024 , n8025 );
not ( n8027 , n7639 );
not ( n8028 , n7731 );
nand ( n8029 , n8028 , n121 );
not ( n8030 , n8029 );
or ( n8031 , n8027 , n8030 );
not ( n8032 , n120 );
nand ( n8033 , n8031 , n8032 );
nand ( n8034 , n8026 , n8033 );
not ( n8035 , n8034 );
nand ( n8036 , n121 , n7822 );
nand ( n8037 , n8035 , n8036 , n7789 );
nand ( n8038 , n8023 , n8037 );
nand ( n8039 , n8003 , n8022 , n8038 );
not ( n8040 , n8039 );
or ( n8041 , n7981 , n8040 );
or ( n8042 , n120 , n7834 );
not ( n8043 , n7855 );
nand ( n8044 , n7813 , n7874 );
not ( n8045 , n8044 );
or ( n8046 , n8043 , n8045 );
not ( n8047 , n126 );
nand ( n8048 , n8046 , n8047 );
not ( n8049 , n126 );
and ( n8050 , n120 , n8049 );
not ( n8051 , n7638 );
not ( n8052 , n125 );
and ( n8053 , n8051 , n8052 );
and ( n8054 , n121 , n7652 );
nor ( n8055 , n8053 , n8054 );
not ( n8056 , n7681 );
nor ( n8057 , n8056 , n121 );
not ( n8058 , n8057 );
nor ( n8059 , n122 , n123 );
nand ( n8060 , n125 , n8059 );
nand ( n8061 , n8055 , n8058 , n8060 );
nand ( n8062 , n8050 , n8061 );
nand ( n8063 , n8042 , n8048 , n8062 );
not ( n8064 , n126 );
and ( n8065 , n7886 , n7834 );
nor ( n8066 , n7759 , n120 );
not ( n8067 , n121 );
nand ( n8068 , n8067 , n7652 );
nor ( n8069 , n120 , n8068 );
nor ( n8070 , n8066 , n8069 );
not ( n8071 , n120 );
nand ( n8072 , n8060 , n7741 , n7770 );
and ( n8073 , n8071 , n8072 );
not ( n8074 , n8071 );
not ( n8075 , n7756 );
nor ( n8076 , n8075 , n121 );
and ( n8077 , n8074 , n8076 );
nor ( n8078 , n8073 , n8077 );
nand ( n8079 , n8065 , n8070 , n8078 );
not ( n8080 , n8079 );
or ( n8081 , n8064 , n8080 );
not ( n8082 , n120 );
nor ( n8083 , n121 , n7678 );
not ( n8084 , n121 );
nand ( n8085 , n8084 , n7973 );
not ( n8086 , n7940 );
nand ( n8087 , n8085 , n8086 );
nor ( n8088 , n8083 , n8087 );
or ( n8089 , n8082 , n8088 );
nand ( n8090 , n7837 , n7798 );
not ( n8091 , n7928 );
nand ( n8092 , n8091 , n7635 );
nand ( n8093 , n8089 , n8090 , n8092 );
not ( n8094 , n8093 );
nand ( n8095 , n8081 , n8094 );
or ( n8096 , n8063 , n8095 );
nand ( n8097 , n8096 , n127 );
nand ( n8098 , n8041 , n8097 );
nor ( n8099 , n7980 , n8098 );
not ( n8100 , n8099 );
not ( n8101 , n7965 );
nand ( n8102 , n121 , n8101 );
not ( n8103 , n8102 );
nand ( n8104 , n8103 , n120 );
not ( n8105 , n126 );
not ( n8106 , n7702 );
nand ( n8107 , n8060 , n7653 , n8106 );
nand ( n8108 , n7813 , n8107 );
not ( n8109 , n7704 );
not ( n8110 , n120 );
nand ( n8111 , n8110 , n7840 );
nand ( n8112 , n8108 , n8109 , n8111 );
nand ( n8113 , n8105 , n8112 );
not ( n8114 , n121 );
nand ( n8115 , n8114 , n7736 );
not ( n8116 , n7647 );
nand ( n8117 , n120 , n8116 );
not ( n8118 , n120 );
nand ( n8119 , n7772 , n7849 );
nand ( n8120 , n8118 , n8119 );
nand ( n8121 , n8115 , n8117 , n8120 );
not ( n8122 , n7695 );
not ( n8123 , n7677 );
not ( n8124 , n8123 );
or ( n8125 , n8122 , n8124 );
nand ( n8126 , n8125 , n7751 );
and ( n8127 , n7802 , n8126 );
not ( n8128 , n7701 );
nand ( n8129 , n7972 , n8128 );
not ( n8130 , n8076 );
nand ( n8131 , n120 , n7683 );
and ( n8132 , n8130 , n8131 );
nand ( n8133 , n8127 , n8129 , n8132 , n126 );
not ( n8134 , n8133 );
nor ( n8135 , n122 , n124 );
nand ( n8136 , n125 , n8135 );
not ( n8137 , n8136 );
not ( n8138 , n8137 );
nand ( n8139 , n8138 , n7941 );
and ( n8140 , n120 , n8139 );
nor ( n8141 , n8140 , n126 );
nor ( n8142 , n7850 , n7629 );
nor ( n8143 , n120 , n7701 );
nor ( n8144 , n8143 , n7897 );
nand ( n8145 , n8141 , n8142 , n8144 );
not ( n8146 , n8145 );
or ( n8147 , n8134 , n8146 );
not ( n8148 , n8004 );
not ( n8149 , n8138 );
nand ( n8150 , n8148 , n8149 );
nand ( n8151 , n8147 , n8150 );
or ( n8152 , n8121 , n8151 );
nand ( n8153 , n8152 , n7748 );
and ( n8154 , n8104 , n8113 , n8153 );
not ( n8155 , n127 );
not ( n8156 , n120 );
not ( n8157 , n8156 );
nand ( n8158 , n121 , n7923 );
not ( n8159 , n121 );
nand ( n8160 , n8159 , n7702 );
nand ( n8161 , n8130 , n8158 , n8160 );
not ( n8162 , n8161 );
or ( n8163 , n8157 , n8162 );
not ( n8164 , n125 );
not ( n8165 , n7732 );
nand ( n8166 , n7873 , n8165 );
not ( n8167 , n8166 );
or ( n8168 , n8164 , n8167 );
not ( n8169 , n7624 );
nand ( n8170 , n8169 , n121 );
or ( n8171 , n7642 , n8170 );
nand ( n8172 , n8168 , n8171 );
nand ( n8173 , n8172 , n120 );
nand ( n8174 , n8163 , n8173 );
not ( n8175 , n7869 );
and ( n8176 , n8175 , n7814 );
nor ( n8177 , n8174 , n8176 );
not ( n8178 , n8069 );
and ( n8179 , n7703 , n8178 );
not ( n8180 , n120 );
not ( n8181 , n7777 );
nand ( n8182 , n8180 , n8181 );
nand ( n8183 , n8179 , n7921 , n8182 );
not ( n8184 , n120 );
or ( n8185 , n121 , n7884 );
not ( n8186 , n7822 );
nand ( n8187 , n8185 , n8186 , n7916 );
not ( n8188 , n8187 );
or ( n8189 , n8184 , n8188 );
nand ( n8190 , n8189 , n7664 );
or ( n8191 , n8183 , n8190 );
not ( n8192 , n126 );
nand ( n8193 , n8191 , n8192 );
not ( n8194 , n120 );
not ( n8195 , n8194 );
nand ( n8196 , n7894 , n8029 );
not ( n8197 , n8196 );
or ( n8198 , n8195 , n8197 );
nor ( n8199 , n121 , n7811 );
not ( n8200 , n8199 );
nand ( n8201 , n8198 , n8200 );
not ( n8202 , n8201 );
not ( n8203 , n7739 );
nand ( n8204 , n8203 , n7670 );
not ( n8205 , n8204 );
not ( n8206 , n7761 );
nor ( n8207 , n8205 , n8206 );
not ( n8208 , n120 );
not ( n8209 , n7929 );
or ( n8210 , n8208 , n8209 );
not ( n8211 , n7873 );
nand ( n8212 , n8175 , n8211 );
not ( n8213 , n8212 );
not ( n8214 , n120 );
nor ( n8215 , n8214 , n7628 );
nor ( n8216 , n8213 , n8215 );
nand ( n8217 , n8202 , n8207 , n8210 , n8216 );
nand ( n8218 , n126 , n8217 );
nand ( n8219 , n8177 , n8193 , n8218 );
not ( n8220 , n8219 );
or ( n8221 , n8155 , n8220 );
not ( n8222 , n126 );
nor ( n8223 , n8222 , n120 );
and ( n8224 , n8223 , n7679 );
not ( n8225 , n8165 );
and ( n8226 , n8175 , n8225 );
not ( n8227 , n7992 );
buf ( n8228 , n7710 );
nor ( n8229 , n8227 , n8228 );
nor ( n8230 , n8224 , n8226 , n8229 );
or ( n8231 , n7739 , n7869 );
nand ( n8232 , n8231 , n7664 );
nand ( n8233 , n8050 , n8232 );
not ( n8234 , n120 );
not ( n8235 , n7671 );
not ( n8236 , n8235 );
or ( n8237 , n8234 , n8236 );
not ( n8238 , n7751 );
nor ( n8239 , n8238 , n7735 );
not ( n8240 , n8239 );
nand ( n8241 , n8237 , n8240 );
nand ( n8242 , n126 , n8241 );
and ( n8243 , n8230 , n8233 , n8242 );
nand ( n8244 , n8221 , n8243 );
not ( n8245 , n8244 );
nand ( n8246 , n8154 , n8245 );
not ( n8247 , n8246 );
and ( n8248 , n8100 , n8247 );
not ( n8249 , n8100 );
and ( n8250 , n8249 , n8246 );
or ( n8251 , n8248 , n8250 );
not ( n8252 , n8251 );
or ( n8253 , n7913 , n8252 );
or ( n8254 , n8251 , n7912 );
nand ( n8255 , n8253 , n8254 );
not ( n8256 , n8255 );
nand ( n8257 , n7324 , n8256 );
nand ( n8258 , n8255 , n7323 );
nand ( n8259 , n8257 , n2352 , n8258 );
nand ( n8260 , n6537 , n8259 );
not ( n8261 , n270 );
and ( n8262 , n271 , n8261 );
not ( n8263 , n271 );
and ( n8264 , n8263 , n270 );
nor ( n8265 , n8262 , n8264 );
or ( n8266 , n2352 , n8265 );
and ( n8267 , n3968 , n3909 );
nand ( n8268 , n201 , n3889 );
not ( n8269 , n8268 );
and ( n8270 , n3758 , n8269 );
nor ( n8271 , n8267 , n8270 );
not ( n8272 , n201 );
nor ( n8273 , n8272 , n3856 );
not ( n8274 , n8273 );
and ( n8275 , n8271 , n3924 , n8274 );
not ( n8276 , n202 );
nor ( n8277 , n8275 , n8276 );
not ( n8278 , n8277 );
not ( n8279 , n3971 );
not ( n8280 , n8279 );
not ( n8281 , n3899 );
or ( n8282 , n8280 , n8281 );
not ( n8283 , n202 );
nand ( n8284 , n8282 , n8283 );
nor ( n8285 , n199 , n3958 );
nand ( n8286 , n202 , n8285 );
nor ( n8287 , n199 , n3793 );
and ( n8288 , n201 , n8287 );
not ( n8289 , n8288 );
and ( n8290 , n8286 , n8289 );
nand ( n8291 , n8284 , n3910 , n8290 );
and ( n8292 , n203 , n8291 );
not ( n8293 , n3941 );
nand ( n8294 , n8293 , n3892 );
and ( n8295 , n8294 , n3995 , n3972 );
nor ( n8296 , n8295 , n202 );
nor ( n8297 , n8292 , n8296 );
nor ( n8298 , n199 , n3811 );
nand ( n8299 , n201 , n8298 );
not ( n8300 , n8299 );
not ( n8301 , n8300 );
not ( n8302 , n202 );
not ( n8303 , n201 );
nand ( n8304 , n199 , n3862 );
nor ( n8305 , n8303 , n8304 );
nand ( n8306 , n8302 , n8305 );
nand ( n8307 , n8301 , n8306 );
not ( n8308 , n202 );
nand ( n8309 , n8308 , n3912 );
not ( n8310 , n3911 );
nand ( n8311 , n201 , n8310 );
buf ( n8312 , n3929 );
not ( n8313 , n8312 );
nand ( n8314 , n202 , n8313 );
nand ( n8315 , n8309 , n8311 , n8314 );
or ( n8316 , n8307 , n8315 );
not ( n8317 , n203 );
nand ( n8318 , n8316 , n8317 );
nand ( n8319 , n8278 , n8297 , n8318 );
nand ( n8320 , n204 , n8319 );
not ( n8321 , n4008 );
not ( n8322 , n3880 );
not ( n8323 , n201 );
not ( n8324 , n3785 );
nand ( n8325 , n8323 , n8324 );
nor ( n8326 , n3856 , n199 );
not ( n8327 , n8326 );
nand ( n8328 , n8325 , n8312 , n8327 );
not ( n8329 , n8328 );
or ( n8330 , n8322 , n8329 );
not ( n8331 , n201 );
nor ( n8332 , n199 , n3833 );
nand ( n8333 , n8331 , n8332 );
not ( n8334 , n8333 );
nand ( n8335 , n199 , n3892 );
not ( n8336 , n8335 );
nand ( n8337 , n201 , n8336 );
not ( n8338 , n8337 );
or ( n8339 , n8334 , n8338 );
nand ( n8340 , n8339 , n202 );
nand ( n8341 , n8330 , n8340 );
not ( n8342 , n8341 );
not ( n8343 , n3941 );
not ( n8344 , n3793 );
nand ( n8345 , n8343 , n8344 );
nand ( n8346 , n199 , n3969 );
not ( n8347 , n8346 );
nand ( n8348 , n201 , n8347 );
not ( n8349 , n8348 );
nand ( n8350 , n8349 , n203 );
nand ( n8351 , n202 , n3844 );
not ( n8352 , n8351 );
nand ( n8353 , n202 , n3892 );
not ( n8354 , n8353 );
or ( n8355 , n8352 , n8354 );
not ( n8356 , n203 );
nand ( n8357 , n8355 , n8356 );
and ( n8358 , n8345 , n8350 , n8357 );
not ( n8359 , n202 );
nand ( n8360 , n8359 , n3846 );
not ( n8361 , n198 );
nand ( n8362 , n8361 , n200 );
not ( n8363 , n8362 );
nand ( n8364 , n8363 , n199 );
or ( n8365 , n3998 , n8364 );
not ( n8366 , n202 );
not ( n8367 , n3789 );
not ( n8368 , n8367 );
nor ( n8369 , n8366 , n8368 );
not ( n8370 , n8369 );
nand ( n8371 , n8365 , n8370 );
and ( n8372 , n203 , n8371 );
not ( n8373 , n203 );
nor ( n8374 , n201 , n202 );
not ( n8375 , n8374 );
not ( n8376 , n8367 );
or ( n8377 , n8375 , n8376 );
not ( n8378 , n199 );
nand ( n8379 , n8378 , n3862 );
not ( n8380 , n8379 );
nand ( n8381 , n201 , n8380 );
nand ( n8382 , n8377 , n8381 );
and ( n8383 , n8373 , n8382 );
nor ( n8384 , n8372 , n8383 );
nand ( n8385 , n8342 , n8358 , n8360 , n8384 );
not ( n8386 , n8385 );
or ( n8387 , n8321 , n8386 );
not ( n8388 , n201 );
nand ( n8389 , n8388 , n8347 );
not ( n8390 , n8389 );
nand ( n8391 , n202 , n8390 );
not ( n8392 , n201 );
nor ( n8393 , n8392 , n3793 );
and ( n8394 , n202 , n8393 );
not ( n8395 , n8394 );
nand ( n8396 , n201 , n8326 );
and ( n8397 , n8391 , n8395 , n8396 );
nand ( n8398 , n201 , n3806 );
not ( n8399 , n202 );
nand ( n8400 , n3833 , n8362 );
nand ( n8401 , n201 , n8400 );
not ( n8402 , n201 );
nand ( n8403 , n8402 , n3925 );
nand ( n8404 , n8401 , n8403 , n8294 );
nand ( n8405 , n8399 , n8404 );
nand ( n8406 , n8397 , n8398 , n8405 );
nand ( n8407 , n203 , n8406 );
nand ( n8408 , n8387 , n8407 );
not ( n8409 , n203 );
not ( n8410 , n8409 );
nor ( n8411 , n3789 , n3758 );
nand ( n8412 , n201 , n8411 );
and ( n8413 , n8412 , n8345 );
not ( n8414 , n202 );
not ( n8415 , n3835 );
not ( n8416 , n201 );
nand ( n8417 , n8415 , n8416 );
not ( n8418 , n3802 );
nand ( n8419 , n8417 , n8418 , n3926 );
nand ( n8420 , n8414 , n8419 );
not ( n8421 , n3883 );
nor ( n8422 , n8421 , n3873 );
nand ( n8423 , n201 , n3887 );
not ( n8424 , n3856 );
nand ( n8425 , n8293 , n8424 );
nand ( n8426 , n8422 , n3967 , n8423 , n8425 );
nand ( n8427 , n202 , n8426 );
nand ( n8428 , n8413 , n8420 , n8427 );
not ( n8429 , n8428 );
or ( n8430 , n8410 , n8429 );
or ( n8431 , n202 , n3764 );
nand ( n8432 , n8431 , n8351 );
nand ( n8433 , n201 , n8432 );
nand ( n8434 , n8430 , n8433 );
nor ( n8435 , n8408 , n8434 );
nand ( n8436 , n8320 , n8435 );
not ( n8437 , n8436 );
not ( n8438 , n212 );
not ( n8439 , n208 );
nand ( n8440 , n8439 , n210 );
or ( n8441 , n205 , n8440 );
not ( n8442 , n210 );
nor ( n8443 , n8442 , n3699 );
not ( n8444 , n8443 );
nand ( n8445 , n8441 , n8444 );
nand ( n8446 , n209 , n8445 );
not ( n8447 , n210 );
nand ( n8448 , n208 , n8447 );
or ( n8449 , n206 , n8448 );
nand ( n8450 , n8449 , n3587 );
and ( n8451 , n209 , n8450 );
not ( n8452 , n209 );
nor ( n8453 , n208 , n210 );
not ( n8454 , n8453 );
or ( n8455 , n8454 , n3655 );
not ( n8456 , n3603 );
buf ( n8457 , n8456 );
nand ( n8458 , n8455 , n8457 , n3643 );
and ( n8459 , n8452 , n8458 );
nor ( n8460 , n8451 , n8459 );
not ( n8461 , n211 );
nor ( n8462 , n208 , n3499 );
nand ( n8463 , n210 , n8462 );
not ( n8464 , n8463 );
not ( n8465 , n3557 );
nand ( n8466 , n8465 , n3582 );
nor ( n8467 , n8466 , n209 );
nor ( n8468 , n8464 , n8467 );
not ( n8469 , n209 );
nand ( n8470 , n8469 , n3669 );
not ( n8471 , n3668 );
nand ( n8472 , n210 , n8471 );
not ( n8473 , n3591 );
nand ( n8474 , n209 , n8473 );
nand ( n8475 , n8468 , n8470 , n8472 , n8474 );
and ( n8476 , n8461 , n8475 );
not ( n8477 , n8461 );
not ( n8478 , n3641 );
not ( n8479 , n3685 );
or ( n8480 , n8478 , n8479 );
not ( n8481 , n209 );
nand ( n8482 , n8480 , n8481 );
not ( n8483 , n208 );
nand ( n8484 , n8483 , n3543 );
not ( n8485 , n8484 );
nand ( n8486 , n209 , n8485 );
not ( n8487 , n3478 );
not ( n8488 , n208 );
nand ( n8489 , n8487 , n8488 );
not ( n8490 , n8489 );
nand ( n8491 , n210 , n8490 );
nand ( n8492 , n8482 , n3679 , n8486 , n8491 );
and ( n8493 , n8477 , n8492 );
nor ( n8494 , n8476 , n8493 );
nand ( n8495 , n8446 , n8460 , n8494 );
not ( n8496 , n8495 );
or ( n8497 , n8438 , n8496 );
not ( n8498 , n209 );
not ( n8499 , n3504 );
nand ( n8500 , n3494 , n8499 );
nand ( n8501 , n210 , n8500 );
not ( n8502 , n210 );
nand ( n8503 , n8502 , n3588 );
nand ( n8504 , n8501 , n8503 , n8455 );
nand ( n8505 , n8498 , n8504 );
not ( n8506 , n3534 );
nand ( n8507 , n8506 , n210 );
not ( n8508 , n208 );
nand ( n8509 , n3684 , n8508 );
not ( n8510 , n8509 );
nand ( n8511 , n8510 , n210 );
nand ( n8512 , n8505 , n8507 , n8511 );
nand ( n8513 , n211 , n8512 );
nand ( n8514 , n8497 , n8513 );
not ( n8515 , n8514 );
not ( n8516 , n211 );
nand ( n8517 , n3640 , n208 );
nor ( n8518 , n210 , n8517 );
and ( n8519 , n209 , n8518 );
nand ( n8520 , n210 , n3725 );
not ( n8521 , n8520 );
nand ( n8522 , n209 , n8521 );
not ( n8523 , n8522 );
nor ( n8524 , n8519 , n8523 );
not ( n8525 , n8524 );
or ( n8526 , n8516 , n8525 );
not ( n8527 , n211 );
not ( n8528 , n208 );
nor ( n8529 , n8528 , n3473 );
nand ( n8530 , n210 , n8529 );
nand ( n8531 , n8453 , n3725 );
and ( n8532 , n8527 , n8530 , n8531 );
not ( n8533 , n209 );
or ( n8534 , n210 , n3496 );
nand ( n8535 , n8534 , n3529 , n3589 );
nand ( n8536 , n8533 , n8535 );
nand ( n8537 , n3638 , n3726 );
nor ( n8538 , n8454 , n3699 );
not ( n8539 , n8538 );
not ( n8540 , n210 );
not ( n8541 , n3722 );
nor ( n8542 , n8540 , n8541 );
not ( n8543 , n8542 );
nand ( n8544 , n8539 , n8543 , n3687 );
or ( n8545 , n8537 , n8544 );
nand ( n8546 , n8545 , n209 );
nand ( n8547 , n8532 , n8536 , n8546 );
nand ( n8548 , n8526 , n8547 );
not ( n8549 , n209 );
not ( n8550 , n3537 );
and ( n8551 , n8549 , n8550 );
not ( n8552 , n8531 );
nor ( n8553 , n8551 , n8552 );
nand ( n8554 , n209 , n3728 );
not ( n8555 , n8517 );
nand ( n8556 , n8555 , n210 );
and ( n8557 , n8554 , n8556 );
nand ( n8558 , n208 , n3504 );
not ( n8559 , n8558 );
not ( n8560 , n209 );
nor ( n8561 , n8560 , n210 );
nand ( n8562 , n8559 , n8561 );
not ( n8563 , n209 );
not ( n8564 , n210 );
not ( n8565 , n3482 );
not ( n8566 , n8565 );
nand ( n8567 , n8564 , n8566 );
not ( n8568 , n3591 );
not ( n8569 , n8568 );
nand ( n8570 , n8567 , n8569 , n8509 );
nand ( n8571 , n8563 , n8570 );
nand ( n8572 , n8557 , n8562 , n8571 );
nand ( n8573 , n211 , n8572 );
not ( n8574 , n210 );
not ( n8575 , n8574 );
not ( n8576 , n208 );
nand ( n8577 , n8576 , n3495 );
not ( n8578 , n8577 );
not ( n8579 , n8578 );
or ( n8580 , n8575 , n8579 );
nand ( n8581 , n208 , n3675 );
not ( n8582 , n8581 );
nand ( n8583 , n210 , n8582 );
nand ( n8584 , n8580 , n8583 );
and ( n8585 , n209 , n8584 );
not ( n8586 , n3710 );
and ( n8587 , n209 , n8586 );
not ( n8588 , n209 );
and ( n8589 , n8588 , n3475 );
nor ( n8590 , n8587 , n8589 );
not ( n8591 , n209 );
nor ( n8592 , n8591 , n3655 );
not ( n8593 , n8592 );
not ( n8594 , n210 );
nor ( n8595 , n8594 , n3583 );
not ( n8596 , n8595 );
and ( n8597 , n8590 , n8593 , n8596 );
nor ( n8598 , n8597 , n211 );
nor ( n8599 , n8585 , n8598 );
nand ( n8600 , n8553 , n8573 , n8599 );
nand ( n8601 , n3469 , n8600 );
and ( n8602 , n209 , n3709 , n3558 );
not ( n8603 , n210 );
nor ( n8604 , n8603 , n209 );
not ( n8605 , n3490 );
and ( n8606 , n8604 , n8605 );
nor ( n8607 , n8602 , n8606 );
nand ( n8608 , n8515 , n8548 , n8601 , n8607 );
not ( n8609 , n8608 );
not ( n8610 , n8609 );
or ( n8611 , n8437 , n8610 );
not ( n8612 , n8436 );
nand ( n8613 , n8608 , n8612 );
nand ( n8614 , n8611 , n8613 );
not ( n8615 , n8614 );
not ( n8616 , n8615 );
or ( n8617 , n209 , n211 );
not ( n8618 , n8617 );
not ( n8619 , n210 );
and ( n8620 , n8619 , n3669 );
not ( n8621 , n3534 );
not ( n8622 , n8530 );
nor ( n8623 , n8620 , n8621 , n8622 );
not ( n8624 , n8623 );
and ( n8625 , n8618 , n8624 );
not ( n8626 , n211 );
not ( n8627 , n209 );
not ( n8628 , n8448 );
not ( n8629 , n3698 );
and ( n8630 , n8629 , n3487 );
not ( n8631 , n8630 );
and ( n8632 , n8628 , n8631 );
not ( n8633 , n3703 );
nor ( n8634 , n8632 , n8633 );
or ( n8635 , n8627 , n8634 );
not ( n8636 , n3579 );
not ( n8637 , n205 );
nand ( n8638 , n8637 , n208 , n207 );
not ( n8639 , n8638 );
and ( n8640 , n8636 , n8639 );
nor ( n8641 , n8640 , n3584 );
nand ( n8642 , n8635 , n8641 );
and ( n8643 , n8626 , n8642 );
nor ( n8644 , n8625 , n8643 );
not ( n8645 , n210 );
or ( n8646 , n8645 , n3731 );
not ( n8647 , n8473 );
or ( n8648 , n209 , n8647 );
nand ( n8649 , n8646 , n8648 );
and ( n8650 , n211 , n8649 );
not ( n8651 , n210 );
nand ( n8652 , n8651 , n8529 );
not ( n8653 , n8652 );
and ( n8654 , n3717 , n8653 );
nor ( n8655 , n8650 , n8654 );
not ( n8656 , n209 );
nand ( n8657 , n8656 , n3530 );
not ( n8658 , n209 );
not ( n8659 , n8491 );
nand ( n8660 , n8658 , n8659 );
nand ( n8661 , n8655 , n8657 , n3580 , n8660 );
not ( n8662 , n8661 );
not ( n8663 , n210 );
not ( n8664 , n8663 );
not ( n8665 , n208 );
nor ( n8666 , n206 , n207 );
nand ( n8667 , n8665 , n8666 );
not ( n8668 , n8667 );
and ( n8669 , n8664 , n8668 );
not ( n8670 , n3583 );
nor ( n8671 , n8669 , n8670 );
nand ( n8672 , n210 , n3647 );
not ( n8673 , n8448 );
nand ( n8674 , n8673 , n3605 );
nand ( n8675 , n8671 , n8672 , n8674 );
nand ( n8676 , n209 , n8675 );
nor ( n8677 , n209 , n8569 );
nand ( n8678 , n8604 , n208 , n8666 );
not ( n8679 , n8678 );
nor ( n8680 , n8677 , n8679 );
not ( n8681 , n209 );
nand ( n8682 , n8681 , n3514 );
and ( n8683 , n8676 , n8680 , n3731 , n8682 );
not ( n8684 , n211 );
not ( n8685 , n3623 );
nand ( n8686 , n8685 , n8636 );
not ( n8687 , n210 );
not ( n8688 , n3685 );
nand ( n8689 , n8687 , n8688 );
nand ( n8690 , n8561 , n3656 );
nand ( n8691 , n8686 , n8689 , n8503 , n8690 );
nand ( n8692 , n8684 , n8691 );
not ( n8693 , n209 );
not ( n8694 , n8693 );
not ( n8695 , n210 );
nand ( n8696 , n8695 , n3642 );
not ( n8697 , n8638 );
not ( n8698 , n210 );
nand ( n8699 , n8697 , n8698 );
nand ( n8700 , n8696 , n3549 , n8699 );
not ( n8701 , n8700 );
or ( n8702 , n8694 , n8701 );
not ( n8703 , n3555 );
not ( n8704 , n8472 );
not ( n8705 , n8529 );
not ( n8706 , n8705 );
or ( n8707 , n8704 , n8706 );
nand ( n8708 , n8707 , n209 );
nand ( n8709 , n8703 , n8708 );
not ( n8710 , n8709 );
nand ( n8711 , n8702 , n8710 );
not ( n8712 , n208 );
not ( n8713 , n3640 );
nor ( n8714 , n8713 , n210 );
nand ( n8715 , n8712 , n207 , n8714 );
nand ( n8716 , n8672 , n3657 , n3529 , n8715 );
or ( n8717 , n8711 , n8716 );
nand ( n8718 , n8717 , n211 );
nand ( n8719 , n8683 , n8692 , n8718 );
and ( n8720 , n3469 , n8719 );
not ( n8721 , n3469 );
not ( n8722 , n211 );
not ( n8723 , n8722 );
nor ( n8724 , n209 , n3474 );
not ( n8725 , n8724 );
nand ( n8726 , n8577 , n8466 );
and ( n8727 , n209 , n8726 );
not ( n8728 , n209 );
not ( n8729 , n210 );
nor ( n8730 , n8729 , n3697 );
and ( n8731 , n8728 , n8730 );
nor ( n8732 , n8727 , n8731 );
nand ( n8733 , n8725 , n3703 , n3638 , n8732 );
not ( n8734 , n8733 );
or ( n8735 , n8723 , n8734 );
nor ( n8736 , n208 , n3560 );
or ( n8737 , n8736 , n3644 );
not ( n8738 , n209 );
nand ( n8739 , n8737 , n8738 );
nand ( n8740 , n8735 , n8739 );
not ( n8741 , n8740 );
not ( n8742 , n210 );
nor ( n8743 , n8742 , n8484 );
not ( n8744 , n3594 );
nor ( n8745 , n8743 , n8744 );
nand ( n8746 , n8745 , n3690 , n3679 );
nand ( n8747 , n211 , n8746 );
not ( n8748 , n209 );
nand ( n8749 , n8748 , n8621 );
or ( n8750 , n3508 , n8440 );
nand ( n8751 , n208 , n8666 );
nand ( n8752 , n8750 , n8751 , n3623 );
not ( n8753 , n209 );
nand ( n8754 , n8752 , n211 , n8753 );
nand ( n8755 , n8749 , n8754 );
nand ( n8756 , n209 , n8633 );
not ( n8757 , n210 );
nor ( n8758 , n8757 , n3729 );
not ( n8759 , n8758 );
nand ( n8760 , n8561 , n8605 );
nand ( n8761 , n8756 , n8759 , n8760 );
nor ( n8762 , n8755 , n8761 );
nand ( n8763 , n8741 , n8747 , n8762 );
and ( n8764 , n8721 , n8763 );
nor ( n8765 , n8720 , n8764 );
and ( n8766 , n8644 , n8662 , n8765 );
not ( n8767 , n8766 );
or ( n8768 , n185 , n186 );
not ( n8769 , n8768 );
not ( n8770 , n8769 );
not ( n8771 , n3180 );
or ( n8772 , n184 , n8771 );
nand ( n8773 , n8772 , n3149 , n3432 );
not ( n8774 , n8773 );
or ( n8775 , n8770 , n8774 );
nor ( n8776 , n184 , n3082 );
not ( n8777 , n8776 );
not ( n8778 , n3308 );
nand ( n8779 , n8778 , n3258 );
not ( n8780 , n184 );
nand ( n8781 , n8780 , n3423 );
not ( n8782 , n8781 );
not ( n8783 , n3175 );
nand ( n8784 , n3202 , n8783 );
and ( n8785 , n3167 , n8784 );
or ( n8786 , n8782 , n8785 );
nand ( n8787 , n8786 , n185 );
nand ( n8788 , n8777 , n8779 , n8787 );
nand ( n8789 , n3013 , n8788 );
nand ( n8790 , n8775 , n8789 );
not ( n8791 , n185 );
not ( n8792 , n3071 );
nand ( n8793 , n8791 , n8792 );
not ( n8794 , n184 );
nor ( n8795 , n8794 , n185 );
nor ( n8796 , n180 , n181 );
nand ( n8797 , n183 , n8796 );
not ( n8798 , n8797 );
nand ( n8799 , n8795 , n8798 );
nand ( n8800 , n8793 , n8799 );
not ( n8801 , n183 );
nand ( n8802 , n8801 , n8796 );
not ( n8803 , n8802 );
and ( n8804 , n184 , n8803 );
not ( n8805 , n3082 );
nor ( n8806 , n8804 , n8805 );
not ( n8807 , n3210 );
nand ( n8808 , n184 , n8807 );
and ( n8809 , n8806 , n8808 , n3204 );
not ( n8810 , n185 );
nor ( n8811 , n8809 , n8810 );
not ( n8812 , n8811 );
not ( n8813 , n185 );
nand ( n8814 , n8813 , n3127 , n3306 );
and ( n8815 , n3454 , n8814 );
not ( n8816 , n3013 );
or ( n8817 , n184 , n3143 );
or ( n8818 , n3011 , n3064 );
nand ( n8819 , n8817 , n8818 );
not ( n8820 , n3219 );
nand ( n8821 , n3068 , n8820 );
nand ( n8822 , n3347 , n3363 );
nand ( n8823 , n8821 , n8822 );
nor ( n8824 , n8819 , n8823 );
not ( n8825 , n8824 );
or ( n8826 , n8816 , n8825 );
not ( n8827 , n184 );
nand ( n8828 , n8827 , n3148 );
nand ( n8829 , n8828 , n3364 );
not ( n8830 , n8829 );
nand ( n8831 , n8830 , n8808 , n3195 );
not ( n8832 , n8831 );
not ( n8833 , n184 );
or ( n8834 , n8833 , n3047 );
and ( n8835 , n8834 , n3150 );
not ( n8836 , n185 );
nor ( n8837 , n8835 , n8836 );
not ( n8838 , n185 );
not ( n8839 , n8838 );
not ( n8840 , n184 );
not ( n8841 , n3232 );
nor ( n8842 , n8841 , n183 );
nand ( n8843 , n8840 , n8842 );
not ( n8844 , n3132 );
nand ( n8845 , n184 , n8844 );
nand ( n8846 , n8843 , n8845 , n3311 );
not ( n8847 , n8846 );
or ( n8848 , n8839 , n8847 );
not ( n8849 , n183 );
nand ( n8850 , n3052 , n8849 );
nand ( n8851 , n8848 , n8850 );
nor ( n8852 , n8837 , n8851 );
nand ( n8853 , n8832 , n186 , n8852 );
nand ( n8854 , n8826 , n8853 );
nand ( n8855 , n8812 , n8815 , n8854 );
nor ( n8856 , n8800 , n8855 );
or ( n8857 , n187 , n8856 );
not ( n8858 , n3138 );
not ( n8859 , n8858 );
not ( n8860 , n3105 );
not ( n8861 , n8842 );
not ( n8862 , n184 );
or ( n8863 , n8861 , n8862 );
and ( n8864 , n8860 , n8863 );
not ( n8865 , n8864 );
or ( n8866 , n8859 , n8865 );
not ( n8867 , n185 );
nand ( n8868 , n8866 , n8867 );
not ( n8869 , n3299 );
or ( n8870 , n185 , n3222 );
not ( n8871 , n3326 );
not ( n8872 , n3038 );
or ( n8873 , n8871 , n8872 );
nand ( n8874 , n8873 , n185 );
nand ( n8875 , n8870 , n8874 );
nor ( n8876 , n8869 , n8875 );
nand ( n8877 , n8876 , n3415 , n8781 );
nand ( n8878 , n3013 , n8877 );
and ( n8879 , n8868 , n8878 );
nand ( n8880 , n3134 , n3074 );
not ( n8881 , n184 );
nand ( n8882 , n8881 , n3426 );
nand ( n8883 , n3184 , n8882 );
or ( n8884 , n8880 , n8883 );
nand ( n8885 , n8884 , n186 );
nor ( n8886 , n185 , n3149 );
not ( n8887 , n8886 );
or ( n8888 , n3127 , n3129 );
nand ( n8889 , n8888 , n8797 , n3064 );
not ( n8890 , n185 );
nand ( n8891 , n8889 , n186 , n8890 );
and ( n8892 , n8887 , n8891 );
nand ( n8893 , n185 , n8782 );
not ( n8894 , n3265 );
not ( n8895 , n3031 );
nand ( n8896 , n3347 , n8895 );
and ( n8897 , n8892 , n8893 , n8894 , n8896 );
nand ( n8898 , n8879 , n8885 , n8897 );
nand ( n8899 , n187 , n8898 );
not ( n8900 , n185 );
not ( n8901 , n8828 );
nand ( n8902 , n8900 , n8901 );
nor ( n8903 , n185 , n3216 );
not ( n8904 , n8903 );
and ( n8905 , n8902 , n3261 , n8904 );
not ( n8906 , n3329 );
not ( n8907 , n184 );
nand ( n8908 , n8907 , n3431 );
not ( n8909 , n8908 );
not ( n8910 , n8909 );
or ( n8911 , n8906 , n8910 );
not ( n8912 , n184 );
not ( n8913 , n3455 );
or ( n8914 , n8912 , n8913 );
nand ( n8915 , n8914 , n8793 );
nand ( n8916 , n186 , n8915 );
nand ( n8917 , n8911 , n8916 );
not ( n8918 , n8917 );
and ( n8919 , n8905 , n8918 );
nand ( n8920 , n8857 , n8899 , n8919 );
nor ( n8921 , n8790 , n8920 );
not ( n8922 , n8921 );
or ( n8923 , n8767 , n8922 );
not ( n8924 , n8661 );
nand ( n8925 , n8924 , n8765 , n8644 );
not ( n8926 , n8790 );
or ( n8927 , n8800 , n8855 );
nand ( n8928 , n8927 , n3275 );
nand ( n8929 , n8926 , n8899 , n8919 , n8928 );
nand ( n8930 , n8925 , n8929 );
nand ( n8931 , n8923 , n8930 );
not ( n8932 , n194 );
not ( n8933 , n8932 );
not ( n8934 , n2472 );
not ( n8935 , n8934 );
not ( n8936 , n2832 );
and ( n8937 , n8935 , n8936 );
not ( n8938 , n2551 );
nor ( n8939 , n8937 , n8938 );
nor ( n8940 , n2547 , n2528 );
or ( n8941 , n2771 , n8940 );
nand ( n8942 , n8941 , n2554 );
nand ( n8943 , n193 , n8942 );
not ( n8944 , n193 );
not ( n8945 , n191 );
nand ( n8946 , n8945 , n2526 );
nand ( n8947 , n8946 , n2817 , n2887 );
nand ( n8948 , n8944 , n8947 );
nand ( n8949 , n8939 , n8943 , n8948 );
not ( n8950 , n8949 );
or ( n8951 , n8933 , n8950 );
not ( n8952 , n194 );
not ( n8953 , n191 );
or ( n8954 , n8953 , n2498 );
not ( n8955 , n193 );
not ( n8956 , n2588 );
nand ( n8957 , n8955 , n8956 );
nand ( n8958 , n8954 , n8957 );
not ( n8959 , n8958 );
or ( n8960 , n8952 , n8959 );
not ( n8961 , n2716 );
not ( n8962 , n193 );
nand ( n8963 , n8961 , n8962 );
nand ( n8964 , n8960 , n8963 );
not ( n8965 , n191 );
nand ( n8966 , n8965 , n2815 );
not ( n8967 , n8966 );
nand ( n8968 , n2516 , n8967 );
nand ( n8969 , n2585 , n2421 );
nand ( n8970 , n8968 , n8969 , n2594 );
nor ( n8971 , n8964 , n8970 );
nand ( n8972 , n8951 , n8971 );
not ( n8973 , n8972 );
nor ( n8974 , n193 , n2817 );
not ( n8975 , n194 );
nor ( n8976 , n2788 , n2539 );
nand ( n8977 , n8976 , n2805 , n2534 );
not ( n8978 , n8977 );
or ( n8979 , n8975 , n8978 );
nand ( n8980 , n2561 , n2380 );
nand ( n8981 , n8979 , n8980 );
nor ( n8982 , n8974 , n8981 );
not ( n8983 , n193 );
nor ( n8984 , n8983 , n2554 );
not ( n8985 , n2840 );
nand ( n8986 , n189 , n2780 );
nor ( n8987 , n189 , n190 );
nand ( n8988 , n192 , n8987 );
nand ( n8989 , n8986 , n8988 , n2626 );
not ( n8990 , n8989 );
or ( n8991 , n8985 , n8990 );
or ( n8992 , n2807 , n2636 );
not ( n8993 , n193 );
nand ( n8994 , n8992 , n8993 );
nand ( n8995 , n8991 , n8994 );
not ( n8996 , n8995 );
not ( n8997 , n2735 );
nand ( n8998 , n2977 , n2665 );
and ( n8999 , n193 , n8998 );
not ( n9000 , n193 );
nand ( n9001 , n9000 , n2711 );
and ( n9002 , n2633 , n2947 );
nand ( n9003 , n9001 , n2554 , n9002 );
or ( n9004 , n8999 , n9003 );
not ( n9005 , n194 );
nand ( n9006 , n9004 , n9005 );
nand ( n9007 , n8996 , n8997 , n9006 );
nor ( n9008 , n8984 , n9007 );
nand ( n9009 , n8982 , n9008 );
and ( n9010 , n195 , n9009 );
not ( n9011 , n195 );
not ( n9012 , n193 );
not ( n9013 , n192 );
nand ( n9014 , n9013 , n8987 );
not ( n9015 , n9014 );
and ( n9016 , n191 , n9015 );
nor ( n9017 , n9016 , n2476 );
nand ( n9018 , n191 , n2611 );
nand ( n9019 , n9017 , n9018 , n2726 );
not ( n9020 , n9019 );
or ( n9021 , n9012 , n9020 );
nand ( n9022 , n9021 , n8957 );
not ( n9023 , n9022 );
not ( n9024 , n2498 );
nor ( n9025 , n2503 , n8988 );
nor ( n9026 , n9024 , n9025 );
not ( n9027 , n193 );
nand ( n9028 , n9027 , n2471 , n2872 );
not ( n9029 , n2525 );
nand ( n9030 , n191 , n9029 );
and ( n9031 , n9030 , n2816 );
not ( n9032 , n193 );
nor ( n9033 , n9031 , n9032 );
not ( n9034 , n193 );
not ( n9035 , n9034 );
not ( n9036 , n191 );
nand ( n9037 , n9036 , n2634 );
not ( n9038 , n2372 );
nand ( n9039 , n9037 , n9038 , n2932 );
not ( n9040 , n9039 );
or ( n9041 , n9035 , n9040 );
nand ( n9042 , n9041 , n2436 );
not ( n9043 , n9042 );
not ( n9044 , n2394 );
and ( n9045 , n9018 , n2631 , n9044 , n2849 );
nand ( n9046 , n9043 , n194 , n9045 );
or ( n9047 , n9033 , n9046 );
not ( n9048 , n194 );
not ( n9049 , n8934 );
not ( n9050 , n2626 );
and ( n9051 , n9049 , n9050 );
not ( n9052 , n191 );
and ( n9053 , n9052 , n2812 );
nor ( n9054 , n9051 , n9053 );
not ( n9055 , n191 );
nand ( n9056 , n9055 , n2572 );
nand ( n9057 , n2561 , n2494 );
nand ( n9058 , n9048 , n9054 , n9056 , n9057 );
nand ( n9059 , n9047 , n9058 );
nand ( n9060 , n9023 , n9026 , n9028 , n9059 );
and ( n9061 , n9011 , n9060 );
nor ( n9062 , n9010 , n9061 );
nand ( n9063 , n8973 , n9062 );
not ( n9064 , n9063 );
and ( n9065 , n9064 , n270 );
not ( n9066 , n9064 );
and ( n9067 , n9066 , n8261 );
nor ( n9068 , n9065 , n9067 );
not ( n9069 , n9068 );
and ( n9070 , n8931 , n9069 );
not ( n9071 , n8931 );
and ( n9072 , n9071 , n9068 );
nor ( n9073 , n9070 , n9072 );
not ( n9074 , n9073 );
nand ( n9075 , n8616 , n9074 );
nand ( n9076 , n8615 , n9073 );
nand ( n9077 , n9075 , n2352 , n9076 );
nand ( n9078 , n8266 , n9077 );
not ( n9079 , n95 );
and ( n9080 , n987 , n9079 );
not ( n9081 , n987 );
and ( n9082 , n9081 , n95 );
nor ( n9083 , n9080 , n9082 );
not ( n9084 , n5835 );
not ( n9085 , n9084 );
not ( n9086 , n5989 );
not ( n9087 , n9086 );
and ( n9088 , n9085 , n9087 );
not ( n9089 , n5989 );
and ( n9090 , n9084 , n9089 );
nor ( n9091 , n9088 , n9090 );
xor ( n9092 , n9083 , n9091 );
not ( n9093 , n9092 );
not ( n9094 , n2337 );
not ( n9095 , n1313 );
and ( n9096 , n1133 , n1413 );
not ( n9097 , n1133 );
and ( n9098 , n9097 , n1469 );
nor ( n9099 , n9096 , n9098 );
nand ( n9100 , n9095 , n1349 , n9099 );
buf ( n9101 , n9100 );
not ( n9102 , n9101 );
and ( n9103 , n9094 , n9102 );
not ( n9104 , n9101 );
not ( n9105 , n9104 );
and ( n9106 , n2341 , n9105 );
nor ( n9107 , n9103 , n9106 );
xor ( n9108 , n9107 , n6153 );
not ( n9109 , n9108 );
or ( n9110 , n9093 , n9109 );
nand ( n9111 , n9110 , n2352 );
nor ( n9112 , n9092 , n9108 );
or ( n9113 , n9111 , n9112 );
and ( n9114 , n96 , n9079 );
not ( n9115 , n96 );
and ( n9116 , n9115 , n95 );
nor ( n9117 , n9114 , n9116 );
or ( n9118 , n2352 , n9117 );
nand ( n9119 , n9113 , n9118 );
xnor ( n9120 , n322 , n323 );
or ( n9121 , n2352 , n9120 );
not ( n9122 , n2654 );
not ( n9123 , n9122 );
not ( n9124 , n322 );
and ( n9125 , n9123 , n9124 );
not ( n9126 , n2654 );
and ( n9127 , n322 , n9126 );
nor ( n9128 , n9125 , n9127 );
not ( n9129 , n3023 );
nand ( n9130 , n184 , n9129 );
and ( n9131 , n9130 , n3074 );
nor ( n9132 , n9131 , n185 );
not ( n9133 , n9132 );
nand ( n9134 , n185 , n3124 );
nand ( n9135 , n184 , n3340 );
not ( n9136 , n9135 );
nand ( n9137 , n185 , n9136 );
nand ( n9138 , n184 , n3114 );
nand ( n9139 , n9134 , n9137 , n9138 );
not ( n9140 , n9139 );
not ( n9141 , n185 );
nand ( n9142 , n3218 , n3148 );
nand ( n9143 , n3115 , n9142 );
and ( n9144 , n9141 , n9143 );
not ( n9145 , n9130 );
nor ( n9146 , n9144 , n9145 );
nand ( n9147 , n9140 , n3013 , n9146 );
nand ( n9148 , n3210 , n3370 );
and ( n9149 , n185 , n9148 );
not ( n9150 , n185 );
nand ( n9151 , n184 , n3344 );
nor ( n9152 , n3132 , n184 );
nor ( n9153 , n9152 , n3065 );
nand ( n9154 , n9151 , n9153 );
and ( n9155 , n9150 , n9154 );
nor ( n9156 , n9149 , n9155 );
nand ( n9157 , n186 , n9156 , n3364 , n8864 );
nand ( n9158 , n9147 , n9157 );
not ( n9159 , n3146 );
or ( n9160 , n183 , n9159 );
nand ( n9161 , n9160 , n3147 );
nand ( n9162 , n185 , n9161 );
and ( n9163 , n8777 , n3261 , n9162 );
nand ( n9164 , n9133 , n9158 , n9163 );
and ( n9165 , n3275 , n9164 );
not ( n9166 , n3275 );
not ( n9167 , n185 );
not ( n9168 , n9167 );
not ( n9169 , n3339 );
not ( n9170 , n9169 );
nand ( n9171 , n9170 , n3123 , n3259 , n3031 );
not ( n9172 , n9171 );
or ( n9173 , n9168 , n9172 );
nand ( n9174 , n9173 , n3341 );
not ( n9175 , n9174 );
nand ( n9176 , n185 , n8901 );
or ( n9177 , n184 , n8850 );
or ( n9178 , n185 , n8845 );
or ( n9179 , n3035 , n3137 );
nand ( n9180 , n9177 , n9178 , n9179 );
not ( n9181 , n183 );
or ( n9182 , n9181 , n8845 );
not ( n9183 , n9182 );
or ( n9184 , n9180 , n9183 , n8895 );
nand ( n9185 , n9184 , n3013 );
not ( n9186 , n186 );
nand ( n9187 , n3345 , n3097 , n3376 );
nand ( n9188 , n185 , n9187 );
nand ( n9189 , n184 , n3423 );
nand ( n9190 , n9188 , n3417 , n9189 );
not ( n9191 , n9190 );
or ( n9192 , n9186 , n9191 );
not ( n9193 , n184 );
not ( n9194 , n3259 );
nand ( n9195 , n9193 , n9194 );
nand ( n9196 , n9192 , n9195 );
not ( n9197 , n9196 );
nand ( n9198 , n9175 , n9176 , n9185 , n9197 );
and ( n9199 , n9166 , n9198 );
nor ( n9200 , n9165 , n9199 );
not ( n9201 , n184 );
not ( n9202 , n8783 );
nand ( n9203 , n9201 , n9202 );
and ( n9204 , n9203 , n8777 , n8781 );
or ( n9205 , n3045 , n9204 );
not ( n9206 , n185 );
nand ( n9207 , n184 , n3144 );
or ( n9208 , n9206 , n9207 );
not ( n9209 , n3456 );
nand ( n9210 , n9205 , n9208 , n9209 );
not ( n9211 , n186 );
not ( n9212 , n184 );
nand ( n9213 , n9212 , n3292 );
not ( n9214 , n184 );
nand ( n9215 , n9214 , n3008 );
and ( n9216 , n3263 , n9213 , n9215 , n3454 );
or ( n9217 , n185 , n9216 );
not ( n9218 , n8795 );
or ( n9219 , n9218 , n3116 );
nand ( n9220 , n9217 , n9219 );
not ( n9221 , n9220 );
or ( n9222 , n9211 , n9221 );
not ( n9223 , n3341 );
not ( n9224 , n3279 );
not ( n9225 , n3417 );
or ( n9226 , n9224 , n9225 );
nand ( n9227 , n9226 , n184 );
not ( n9228 , n9227 );
or ( n9229 , n9223 , n9228 );
nand ( n9230 , n9229 , n3329 );
nand ( n9231 , n9222 , n9230 );
nor ( n9232 , n9210 , n9231 );
and ( n9233 , n3181 , n3353 , n8882 );
or ( n9234 , n185 , n9233 );
and ( n9235 , n9207 , n3184 );
nand ( n9236 , n9234 , n9235 );
nand ( n9237 , n3013 , n9236 );
nand ( n9238 , n9200 , n9232 , n9237 );
not ( n9239 , n9238 );
not ( n9240 , n3747 );
and ( n9241 , n9239 , n9240 );
not ( n9242 , n9239 );
not ( n9243 , n9240 );
and ( n9244 , n9242 , n9243 );
nor ( n9245 , n9241 , n9244 );
not ( n9246 , n9245 );
and ( n9247 , n9128 , n9246 );
not ( n9248 , n9128 );
and ( n9249 , n9248 , n9245 );
nor ( n9250 , n9247 , n9249 );
not ( n9251 , n9250 );
not ( n9252 , n209 );
nand ( n9253 , n210 , n3519 );
not ( n9254 , n3623 );
not ( n9255 , n210 );
nand ( n9256 , n9254 , n9255 );
nand ( n9257 , n3594 , n9253 , n9256 );
nand ( n9258 , n9252 , n9257 );
not ( n9259 , n211 );
not ( n9260 , n9259 );
not ( n9261 , n210 );
not ( n9262 , n9261 );
nand ( n9263 , n3587 , n3490 );
not ( n9264 , n9263 );
or ( n9265 , n9262 , n9264 );
not ( n9266 , n8467 );
nand ( n9267 , n9265 , n9266 );
not ( n9268 , n9267 );
or ( n9269 , n9260 , n9268 );
or ( n9270 , n3495 , n3725 );
not ( n9271 , n8440 );
nand ( n9272 , n9270 , n209 , n9271 );
nand ( n9273 , n9269 , n9272 );
not ( n9274 , n211 );
nor ( n9275 , n3499 , n3557 );
not ( n9276 , n9275 );
not ( n9277 , n210 );
nand ( n9278 , n9277 , n3582 );
nand ( n9279 , n9276 , n9278 );
not ( n9280 , n210 );
not ( n9281 , n209 );
nand ( n9282 , n9280 , n9281 );
nor ( n9283 , n8499 , n9282 );
not ( n9284 , n209 );
not ( n9285 , n3637 );
or ( n9286 , n9284 , n9285 );
not ( n9287 , n8670 );
nand ( n9288 , n9286 , n9287 );
nor ( n9289 , n9279 , n9283 , n9288 );
or ( n9290 , n9274 , n9289 );
not ( n9291 , n8471 );
or ( n9292 , n210 , n9291 );
nand ( n9293 , n9292 , n8565 );
nand ( n9294 , n3696 , n9293 );
nand ( n9295 , n9290 , n9294 );
nor ( n9296 , n9273 , n9295 );
and ( n9297 , n9258 , n9296 );
nor ( n9298 , n9297 , n212 );
not ( n9299 , n9298 );
not ( n9300 , n211 );
not ( n9301 , n8674 );
and ( n9302 , n209 , n9301 );
not ( n9303 , n9282 );
and ( n9304 , n9303 , n3647 );
nor ( n9305 , n9302 , n9304 );
nand ( n9306 , n209 , n8730 );
and ( n9307 , n9305 , n9306 , n8491 , n8455 );
or ( n9308 , n9300 , n9307 );
not ( n9309 , n209 );
not ( n9310 , n8715 );
or ( n9311 , n9309 , n9310 );
or ( n9312 , n209 , n9275 );
nand ( n9313 , n9311 , n9312 );
nand ( n9314 , n9308 , n9313 );
not ( n9315 , n211 );
not ( n9316 , n9315 );
not ( n9317 , n209 );
nand ( n9318 , n9317 , n8758 );
not ( n9319 , n209 );
not ( n9320 , n210 );
nand ( n9321 , n9320 , n3605 );
not ( n9322 , n8518 );
nand ( n9323 , n9321 , n9322 , n8531 );
nand ( n9324 , n9319 , n9323 );
nand ( n9325 , n3580 , n9318 , n9324 );
not ( n9326 , n9325 );
or ( n9327 , n9316 , n9326 );
nand ( n9328 , n3709 , n8453 );
not ( n9329 , n9328 );
or ( n9330 , n9329 , n8538 );
nand ( n9331 , n9330 , n3696 );
nand ( n9332 , n9327 , n9331 );
nor ( n9333 , n9314 , n9332 );
and ( n9334 , n3476 , n8511 );
not ( n9335 , n3520 );
nand ( n9336 , n3561 , n8673 );
not ( n9337 , n9336 );
or ( n9338 , n9335 , n9337 );
not ( n9339 , n209 );
nand ( n9340 , n9338 , n9339 );
nor ( n9341 , n3671 , n3689 );
nand ( n9342 , n3594 , n8509 , n9341 );
nand ( n9343 , n209 , n9342 );
nand ( n9344 , n9334 , n9340 , n9343 );
not ( n9345 , n8743 );
not ( n9346 , n210 );
nor ( n9347 , n208 , n3560 );
nand ( n9348 , n9346 , n9347 );
nand ( n9349 , n9345 , n9348 );
nand ( n9350 , n3508 , n9271 );
nand ( n9351 , n9303 , n8688 );
nand ( n9352 , n8705 , n3534 , n3575 );
nand ( n9353 , n209 , n9352 );
nand ( n9354 , n9350 , n9351 , n9353 );
nor ( n9355 , n9349 , n9354 );
or ( n9356 , n211 , n9355 );
and ( n9357 , n210 , n3570 );
nand ( n9358 , n210 , n3495 );
not ( n9359 , n9358 );
nor ( n9360 , n9357 , n9359 );
or ( n9361 , n209 , n9360 );
or ( n9362 , n209 , n3708 );
nand ( n9363 , n9362 , n3610 , n3739 );
nand ( n9364 , n211 , n9363 );
nand ( n9365 , n9356 , n9361 , n9364 );
or ( n9366 , n9344 , n9365 );
nand ( n9367 , n9366 , n212 );
nand ( n9368 , n9299 , n9333 , n9367 );
not ( n9369 , n9368 );
not ( n9370 , n9369 );
not ( n9371 , n211 );
nand ( n9372 , n3483 , n3537 );
not ( n9373 , n8561 );
not ( n9374 , n3496 );
not ( n9375 , n9374 );
or ( n9376 , n9373 , n9375 );
not ( n9377 , n205 );
nand ( n9378 , n9377 , n3558 );
not ( n9379 , n9378 );
not ( n9380 , n3674 );
or ( n9381 , n9379 , n9380 );
not ( n9382 , n209 );
nand ( n9383 , n9381 , n9382 );
nand ( n9384 , n9376 , n9383 );
nor ( n9385 , n9372 , n9384 );
or ( n9386 , n9371 , n9385 );
not ( n9387 , n3520 );
not ( n9388 , n3480 );
or ( n9389 , n9387 , n9388 );
nand ( n9390 , n9389 , n8636 );
not ( n9391 , n8581 );
not ( n9392 , n8530 );
or ( n9393 , n9391 , n9392 );
not ( n9394 , n209 );
nand ( n9395 , n9393 , n9394 );
nand ( n9396 , n9390 , n9395 );
not ( n9397 , n9396 );
nor ( n9398 , n3579 , n8558 );
nor ( n9399 , n8592 , n9398 );
or ( n9400 , n211 , n9399 );
nand ( n9401 , n9400 , n3735 );
not ( n9402 , n211 );
not ( n9403 , n9402 );
not ( n9404 , n209 );
not ( n9405 , n9404 );
not ( n9406 , n208 );
nand ( n9407 , n9406 , n206 );
not ( n9408 , n9407 );
not ( n9409 , n9408 );
or ( n9410 , n9405 , n9409 );
nand ( n9411 , n9410 , n3670 );
not ( n9412 , n9411 );
or ( n9413 , n9403 , n9412 );
not ( n9414 , n3651 );
not ( n9415 , n9348 );
or ( n9416 , n9414 , n9415 );
not ( n9417 , n209 );
nand ( n9418 , n9416 , n9417 );
nand ( n9419 , n9413 , n9418 );
nor ( n9420 , n9401 , n9419 );
nand ( n9421 , n9386 , n9397 , n9420 );
nand ( n9422 , n9421 , n3469 );
not ( n9423 , n211 );
not ( n9424 , n3505 );
nand ( n9425 , n210 , n9424 );
or ( n9426 , n209 , n9425 );
not ( n9427 , n210 );
nand ( n9428 , n9427 , n3647 );
nand ( n9429 , n9426 , n9428 , n9418 );
nand ( n9430 , n9423 , n9429 );
not ( n9431 , n3696 );
not ( n9432 , n210 );
nand ( n9433 , n9432 , n8586 );
nand ( n9434 , n9433 , n3657 , n8507 );
not ( n9435 , n9434 );
or ( n9436 , n9431 , n9435 );
not ( n9437 , n8715 );
not ( n9438 , n8583 );
or ( n9439 , n9437 , n9438 );
not ( n9440 , n209 );
nand ( n9441 , n9439 , n9440 );
nand ( n9442 , n9436 , n9441 );
not ( n9443 , n9442 );
nand ( n9444 , n9422 , n9430 , n9443 );
not ( n9445 , n211 );
not ( n9446 , n9445 );
not ( n9447 , n209 );
nand ( n9448 , n208 , n3730 );
nand ( n9449 , n9448 , n3710 , n8517 );
nand ( n9450 , n9447 , n9449 );
nor ( n9451 , n210 , n3505 );
nand ( n9452 , n209 , n9451 );
nor ( n9453 , n8518 , n8542 );
not ( n9454 , n209 );
nand ( n9455 , n9454 , n8714 );
not ( n9456 , n9455 );
nor ( n9457 , n8724 , n9456 );
nand ( n9458 , n9450 , n9452 , n9453 , n9457 );
not ( n9459 , n9458 );
or ( n9460 , n9446 , n9459 );
not ( n9461 , n209 );
nand ( n9462 , n9461 , n8518 );
nand ( n9463 , n9460 , n9462 );
and ( n9464 , n8636 , n8578 );
not ( n9465 , n209 );
not ( n9466 , n210 );
nand ( n9467 , n9466 , n8462 );
nand ( n9468 , n9467 , n8705 , n8699 );
not ( n9469 , n9468 );
or ( n9470 , n9465 , n9469 );
nand ( n9471 , n9470 , n9336 );
nor ( n9472 , n9464 , n9471 );
not ( n9473 , n8507 );
nand ( n9474 , n9303 , n3684 );
not ( n9475 , n9474 );
or ( n9476 , n9473 , n9475 );
nand ( n9477 , n9476 , n211 );
and ( n9478 , n210 , n3640 );
not ( n9479 , n205 );
nor ( n9480 , n9479 , n208 );
nor ( n9481 , n9478 , n9480 );
nand ( n9482 , n9481 , n9448 , n9278 );
nand ( n9483 , n3717 , n9482 );
nand ( n9484 , n9472 , n9477 , n9483 );
nor ( n9485 , n9463 , n9484 );
or ( n9486 , n3469 , n9485 );
not ( n9487 , n209 );
not ( n9488 , n210 );
nor ( n9489 , n8639 , n9263 );
or ( n9490 , n9488 , n9489 );
nand ( n9491 , n9490 , n8520 );
nand ( n9492 , n9487 , n9491 );
not ( n9493 , n9492 );
not ( n9494 , n210 );
not ( n9495 , n9494 );
not ( n9496 , n8462 );
nand ( n9497 , n9496 , n3685 , n8489 );
not ( n9498 , n9497 );
or ( n9499 , n9495 , n9498 );
and ( n9500 , n3638 , n3513 );
nand ( n9501 , n9499 , n9500 );
nand ( n9502 , n209 , n9501 );
not ( n9503 , n9502 );
or ( n9504 , n9493 , n9503 );
nand ( n9505 , n9504 , n211 );
nand ( n9506 , n9486 , n9505 );
nor ( n9507 , n9444 , n9506 );
not ( n9508 , n9507 );
not ( n9509 , n9508 );
not ( n9510 , n9509 );
or ( n9511 , n9370 , n9510 );
buf ( n9512 , n9507 );
not ( n9513 , n9512 );
not ( n9514 , n9513 );
or ( n9515 , n9369 , n9514 );
nand ( n9516 , n9511 , n9515 );
not ( n9517 , n202 );
nand ( n9518 , n8335 , n8412 );
and ( n9519 , n9517 , n9518 );
and ( n9520 , n3818 , n3795 );
nor ( n9521 , n9520 , n3898 );
nor ( n9522 , n9519 , n9521 );
not ( n9523 , n3758 );
not ( n9524 , n8268 );
and ( n9525 , n9523 , n9524 );
nor ( n9526 , n9525 , n3916 );
or ( n9527 , n202 , n9526 );
or ( n9528 , n3998 , n3835 );
nand ( n9529 , n9527 , n9528 );
nand ( n9530 , n3787 , n3807 );
or ( n9531 , n9529 , n9530 );
nand ( n9532 , n9531 , n203 );
not ( n9533 , n3980 );
not ( n9534 , n201 );
not ( n9535 , n199 );
nand ( n9536 , n9535 , n3778 );
not ( n9537 , n9536 );
nand ( n9538 , n9534 , n9537 );
not ( n9539 , n9538 );
or ( n9540 , n9533 , n9539 );
not ( n9541 , n202 );
nand ( n9542 , n9540 , n9541 );
nand ( n9543 , n4008 , n3901 , n9542 );
not ( n9544 , n203 );
not ( n9545 , n9544 );
not ( n9546 , n202 );
not ( n9547 , n9546 );
not ( n9548 , n200 );
nor ( n9549 , n9548 , n199 );
not ( n9550 , n9549 );
or ( n9551 , n9547 , n9550 );
nand ( n9552 , n9551 , n3913 );
not ( n9553 , n9552 );
or ( n9554 , n9545 , n9553 );
not ( n9555 , n203 );
not ( n9556 , n3897 );
not ( n9557 , n8364 );
not ( n9558 , n9557 );
or ( n9559 , n9556 , n9558 );
nand ( n9560 , n9559 , n8353 );
nand ( n9561 , n9555 , n9560 );
nand ( n9562 , n9554 , n9561 );
nor ( n9563 , n9543 , n9562 );
nand ( n9564 , n9522 , n9532 , n9563 );
not ( n9565 , n9564 );
not ( n9566 , n202 );
not ( n9567 , n8298 );
or ( n9568 , n201 , n9567 );
not ( n9569 , n8411 );
not ( n9570 , n201 );
nor ( n9571 , n3758 , n3886 );
nand ( n9572 , n9570 , n9571 );
nand ( n9573 , n9568 , n9569 , n9572 );
not ( n9574 , n9573 );
or ( n9575 , n9566 , n9574 );
nor ( n9576 , n8376 , n202 );
not ( n9577 , n9576 );
nand ( n9578 , n3969 , n8374 );
and ( n9579 , n8423 , n9578 );
nor ( n9580 , n3828 , n201 );
nand ( n9581 , n202 , n9580 );
nand ( n9582 , n9577 , n9579 , n8389 , n9581 );
nand ( n9583 , n199 , n3953 );
not ( n9584 , n3844 );
and ( n9585 , n9583 , n9584 , n8346 );
nor ( n9586 , n9585 , n202 );
or ( n9587 , n9582 , n9586 );
not ( n9588 , n203 );
nand ( n9589 , n9587 , n9588 );
nand ( n9590 , n9575 , n9589 );
not ( n9591 , n9590 );
not ( n9592 , n202 );
and ( n9593 , n9592 , n8390 );
and ( n9594 , n3778 , n3909 );
nor ( n9595 , n9593 , n9594 , n4008 );
nand ( n9596 , n3897 , n8332 );
not ( n9597 , n3857 );
or ( n9598 , n8375 , n9597 );
nand ( n9599 , n9598 , n8398 );
and ( n9600 , n203 , n9599 );
and ( n9601 , n201 , n3969 );
and ( n9602 , n197 , n3758 );
nor ( n9603 , n9601 , n9602 );
not ( n9604 , n201 );
nand ( n9605 , n9604 , n3862 );
and ( n9606 , n9603 , n9583 , n9605 );
nor ( n9607 , n9606 , n3824 );
nor ( n9608 , n9600 , n9607 );
nand ( n9609 , n9591 , n9595 , n9596 , n9608 );
not ( n9610 , n9609 );
or ( n9611 , n9565 , n9610 );
not ( n9612 , n3854 );
or ( n9613 , n201 , n9584 );
nand ( n9614 , n9613 , n3965 , n8398 );
not ( n9615 , n9614 );
or ( n9616 , n9612 , n9615 );
nand ( n9617 , n8343 , n3790 );
not ( n9618 , n9617 );
not ( n9619 , n8337 );
or ( n9620 , n9618 , n9619 );
not ( n9621 , n202 );
nand ( n9622 , n9620 , n9621 );
nand ( n9623 , n9616 , n9622 );
not ( n9624 , n203 );
not ( n9625 , n202 );
not ( n9626 , n201 );
nor ( n9627 , n9626 , n3828 );
nand ( n9628 , n9625 , n9627 );
not ( n9629 , n201 );
nand ( n9630 , n9629 , n3976 );
and ( n9631 , n9628 , n9630 , n9542 );
and ( n9632 , n9624 , n9631 );
not ( n9633 , n9624 );
not ( n9634 , n202 );
not ( n9635 , n201 );
not ( n9636 , n9571 );
nand ( n9637 , n9636 , n3924 , n3764 );
not ( n9638 , n9637 );
or ( n9639 , n9635 , n9638 );
not ( n9640 , n8393 );
nand ( n9641 , n9639 , n9640 );
and ( n9642 , n9634 , n9641 );
not ( n9643 , n9634 );
not ( n9644 , n201 );
not ( n9645 , n9644 );
not ( n9646 , n8287 );
nand ( n9647 , n3899 , n9567 , n9646 );
not ( n9648 , n9647 );
or ( n9649 , n9645 , n9648 );
and ( n9650 , n3967 , n3814 );
nand ( n9651 , n9649 , n9650 );
and ( n9652 , n9643 , n9651 );
nor ( n9653 , n9642 , n9652 );
and ( n9654 , n9633 , n9653 );
nor ( n9655 , n9632 , n9654 );
nor ( n9656 , n9623 , n9655 );
nand ( n9657 , n9611 , n9656 );
buf ( n9658 , n9657 );
not ( n9659 , n9658 );
not ( n9660 , n203 );
not ( n9661 , n3842 );
nand ( n9662 , n9661 , n3860 );
nand ( n9663 , n9662 , n8425 );
and ( n9664 , n202 , n9663 );
not ( n9665 , n202 );
not ( n9666 , n201 );
nand ( n9667 , n9666 , n3938 );
nand ( n9668 , n9667 , n8389 , n8345 );
and ( n9669 , n9665 , n9668 );
nor ( n9670 , n9664 , n9669 );
not ( n9671 , n201 );
nor ( n9672 , n9671 , n199 );
nand ( n9673 , n9672 , n9576 );
nand ( n9674 , n9670 , n4004 , n9673 );
nand ( n9675 , n9660 , n9674 );
not ( n9676 , n202 );
nor ( n9677 , n8274 , n9676 );
not ( n9678 , n9677 );
nand ( n9679 , n3909 , n3938 );
not ( n9680 , n9679 );
and ( n9681 , n202 , n9680 );
not ( n9682 , n202 );
not ( n9683 , n9630 );
and ( n9684 , n9682 , n9683 );
nor ( n9685 , n9681 , n9684 );
nand ( n9686 , n9678 , n8289 , n8294 , n9685 );
nand ( n9687 , n203 , n9686 );
not ( n9688 , n202 );
nand ( n9689 , n199 , n3830 );
and ( n9690 , n9688 , n9689 );
not ( n9691 , n9688 );
and ( n9692 , n9691 , n9617 );
or ( n9693 , n9690 , n9692 );
nand ( n9694 , n9675 , n9687 , n9693 );
not ( n9695 , n9694 );
not ( n9696 , n3967 );
nand ( n9697 , n202 , n9696 );
nand ( n9698 , n3827 , n8374 );
and ( n9699 , n9698 , n9605 , n9689 );
nand ( n9700 , n9697 , n8379 , n9699 );
nand ( n9701 , n203 , n9700 );
or ( n9702 , n201 , n3911 );
not ( n9703 , n3786 );
nand ( n9704 , n9702 , n9703 );
nand ( n9705 , n3854 , n9704 );
not ( n9706 , n203 );
not ( n9707 , n201 );
not ( n9708 , n9707 );
nand ( n9709 , n3924 , n3764 );
not ( n9710 , n9709 );
or ( n9711 , n9708 , n9710 );
nand ( n9712 , n9711 , n8306 );
nand ( n9713 , n9706 , n9712 );
nand ( n9714 , n9701 , n9705 , n9713 );
not ( n9715 , n9714 );
not ( n9716 , n202 );
not ( n9717 , n9716 );
not ( n9718 , n3954 );
not ( n9719 , n201 );
nand ( n9720 , n9718 , n9719 );
nand ( n9721 , n201 , n3979 );
nand ( n9722 , n9720 , n9721 , n3932 );
not ( n9723 , n9722 );
or ( n9724 , n9717 , n9723 );
not ( n9725 , n8344 );
nand ( n9726 , n3833 , n9725 );
nand ( n9727 , n9726 , n202 , n9672 );
nand ( n9728 , n9724 , n9727 );
not ( n9729 , n9728 );
and ( n9730 , n9715 , n9729 );
nor ( n9731 , n9730 , n204 );
not ( n9732 , n9731 );
and ( n9733 , n3791 , n8396 );
not ( n9734 , n3818 );
or ( n9735 , n9734 , n9594 );
not ( n9736 , n202 );
nand ( n9737 , n9735 , n9736 );
not ( n9738 , n8326 );
nand ( n9739 , n3913 , n3874 );
not ( n9740 , n9739 );
nand ( n9741 , n9738 , n3932 , n9740 );
nand ( n9742 , n202 , n9741 );
nand ( n9743 , n9733 , n9737 , n9742 );
or ( n9744 , n202 , n3842 );
not ( n9745 , n202 );
nand ( n9746 , n9745 , n3892 );
nand ( n9747 , n9744 , n3939 , n9746 );
nand ( n9748 , n203 , n9747 );
not ( n9749 , n202 );
not ( n9750 , n201 );
not ( n9751 , n3985 );
or ( n9752 , n9750 , n9751 );
not ( n9753 , n3833 );
nand ( n9754 , n201 , n9753 );
nand ( n9755 , n9752 , n9754 );
nand ( n9756 , n9749 , n9755 );
nand ( n9757 , n201 , n8285 );
nand ( n9758 , n9757 , n9538 );
nand ( n9759 , n3759 , n9672 );
not ( n9760 , n8375 );
not ( n9761 , n9760 );
or ( n9762 , n9761 , n3899 );
not ( n9763 , n3806 );
nand ( n9764 , n3989 , n9763 , n9569 );
nand ( n9765 , n202 , n9764 );
nand ( n9766 , n9759 , n9762 , n9765 );
or ( n9767 , n9758 , n9766 );
not ( n9768 , n203 );
nand ( n9769 , n9767 , n9768 );
nand ( n9770 , n9748 , n9756 , n9769 );
or ( n9771 , n9743 , n9770 );
nand ( n9772 , n9771 , n204 );
nand ( n9773 , n9695 , n9732 , n9772 );
not ( n9774 , n9773 );
not ( n9775 , n9774 );
or ( n9776 , n9659 , n9775 );
not ( n9777 , n9731 );
not ( n9778 , n9694 );
nand ( n9779 , n9777 , n9778 , n9772 );
not ( n9780 , n9779 );
not ( n9781 , n9657 );
buf ( n9782 , n9781 );
not ( n9783 , n9782 );
or ( n9784 , n9780 , n9783 );
nand ( n9785 , n9776 , n9784 );
and ( n9786 , n9516 , n9785 );
not ( n9787 , n9516 );
not ( n9788 , n9773 );
not ( n9789 , n9658 );
and ( n9790 , n9788 , n9789 );
and ( n9791 , n9779 , n9658 );
nor ( n9792 , n9790 , n9791 );
not ( n9793 , n9792 );
and ( n9794 , n9787 , n9793 );
nor ( n9795 , n9786 , n9794 );
not ( n9796 , n9795 );
nand ( n9797 , n9251 , n9796 );
nand ( n9798 , n9250 , n9795 );
nand ( n9799 , n9797 , n2352 , n9798 );
nand ( n9800 , n9121 , n9799 );
xnor ( n9801 , n390 , n391 );
or ( n9802 , n2352 , n9801 );
not ( n9803 , n390 );
not ( n9804 , n4298 );
or ( n9805 , n9803 , n9804 );
not ( n9806 , n4297 );
or ( n9807 , n390 , n9806 );
nand ( n9808 , n9805 , n9807 );
not ( n9809 , n9808 );
not ( n9810 , n4217 );
nand ( n9811 , n9810 , n154 );
not ( n9812 , n9811 );
nand ( n9813 , n158 , n9812 );
not ( n9814 , n9813 );
not ( n9815 , n9814 );
not ( n9816 , n158 );
not ( n9817 , n9816 );
not ( n9818 , n4221 );
or ( n9819 , n9817 , n9818 );
not ( n9820 , n154 );
nor ( n9821 , n156 , n157 );
nand ( n9822 , n9820 , n9821 );
not ( n9823 , n9822 );
nand ( n9824 , n4226 , n9823 );
nand ( n9825 , n9819 , n9824 );
not ( n9826 , n9825 );
nand ( n9827 , n159 , n4123 );
not ( n9828 , n159 );
not ( n9829 , n4119 );
nand ( n9830 , n154 , n9829 );
not ( n9831 , n9830 );
not ( n9832 , n158 );
nand ( n9833 , n9831 , n9832 );
nand ( n9834 , n4208 , n9833 );
nand ( n9835 , n9828 , n9834 );
nand ( n9836 , n9826 , n9827 , n9835 );
not ( n9837 , n159 );
not ( n9838 , n154 );
nand ( n9839 , n4078 , n9838 );
not ( n9840 , n9839 );
nand ( n9841 , n9837 , n9840 );
not ( n9842 , n9830 );
nand ( n9843 , n9842 , n158 );
nand ( n9844 , n9841 , n4138 , n9843 );
not ( n9845 , n9822 );
not ( n9846 , n4256 );
not ( n9847 , n158 );
nand ( n9848 , n9846 , n9847 );
not ( n9849 , n9848 );
or ( n9850 , n9845 , n9849 );
nand ( n9851 , n9850 , n159 );
nand ( n9852 , n4249 , n9851 );
nor ( n9853 , n9844 , n9852 );
and ( n9854 , n160 , n9853 );
not ( n9855 , n160 );
not ( n9856 , n158 );
nor ( n9857 , n154 , n4191 );
nand ( n9858 , n9856 , n9857 );
not ( n9859 , n4070 );
nand ( n9860 , n9859 , n4057 );
and ( n9861 , n4196 , n9860 );
and ( n9862 , n159 , n154 , n4066 );
nor ( n9863 , n9861 , n9862 );
and ( n9864 , n9858 , n9863 );
not ( n9865 , n159 );
and ( n9866 , n158 , n9865 );
nand ( n9867 , n9866 , n4080 );
and ( n9868 , n9864 , n4085 , n9867 );
and ( n9869 , n9855 , n9868 );
nor ( n9870 , n9854 , n9869 );
or ( n9871 , n9836 , n9870 );
nand ( n9872 , n9871 , n4144 );
not ( n9873 , n159 );
not ( n9874 , n158 );
nand ( n9875 , n9874 , n4285 );
nand ( n9876 , n9875 , n4182 , n4193 );
not ( n9877 , n9876 );
or ( n9878 , n9873 , n9877 );
nand ( n9879 , n9878 , n4041 );
not ( n9880 , n9879 );
not ( n9881 , n158 );
not ( n9882 , n154 );
nor ( n9883 , n9882 , n4057 );
nand ( n9884 , n9881 , n9883 );
and ( n9885 , n9884 , n4079 );
not ( n9886 , n158 );
not ( n9887 , n4031 );
nand ( n9888 , n9886 , n9887 );
nor ( n9889 , n159 , n9888 );
not ( n9890 , n4048 );
not ( n9891 , n9890 );
nor ( n9892 , n159 , n9891 );
nor ( n9893 , n9889 , n9892 );
nand ( n9894 , n9880 , n9885 , n9893 );
nand ( n9895 , n9894 , n160 );
not ( n9896 , n158 );
not ( n9897 , n4255 );
nor ( n9898 , n154 , n9897 );
not ( n9899 , n9898 );
nor ( n9900 , n9896 , n9899 );
not ( n9901 , n9900 );
not ( n9902 , n158 );
not ( n9903 , n4163 );
nand ( n9904 , n9902 , n9903 );
nand ( n9905 , n159 , n4137 );
and ( n9906 , n9904 , n9905 );
not ( n9907 , n9866 );
not ( n9908 , n4217 );
not ( n9909 , n9908 );
or ( n9910 , n9907 , n9909 );
not ( n9911 , n4039 );
nand ( n9912 , n4148 , n9911 );
nand ( n9913 , n9910 , n9912 );
not ( n9914 , n157 );
nand ( n9915 , n9914 , n156 );
nor ( n9916 , n154 , n9915 );
nand ( n9917 , n159 , n9916 );
not ( n9918 , n4157 );
nand ( n9919 , n9918 , n4042 );
not ( n9920 , n4136 );
nand ( n9921 , n4064 , n9920 );
nand ( n9922 , n9917 , n9919 , n9921 );
nor ( n9923 , n9913 , n9922 );
nand ( n9924 , n9906 , n4201 , n9923 );
nand ( n9925 , n9924 , n4054 );
nand ( n9926 , n9895 , n9901 , n9925 );
not ( n9927 , n154 );
not ( n9928 , n4281 );
not ( n9929 , n9908 );
nand ( n9930 , n9928 , n9929 );
not ( n9931 , n9930 );
or ( n9932 , n9927 , n9931 );
not ( n9933 , n154 );
not ( n9934 , n4088 );
nand ( n9935 , n9934 , n158 );
nor ( n9936 , n9933 , n9935 );
not ( n9937 , n9936 );
nand ( n9938 , n9932 , n9937 );
and ( n9939 , n159 , n9938 );
not ( n9940 , n159 );
not ( n9941 , n4119 );
nand ( n9942 , n158 , n9941 );
not ( n9943 , n4079 );
not ( n9944 , n158 );
nand ( n9945 , n9943 , n9944 );
nand ( n9946 , n9858 , n9942 , n9945 );
and ( n9947 , n9940 , n9946 );
nor ( n9948 , n9939 , n9947 );
not ( n9949 , n9948 );
or ( n9950 , n9926 , n9949 );
nand ( n9951 , n9950 , n161 );
nand ( n9952 , n9815 , n9872 , n9951 );
not ( n9953 , n9952 );
not ( n9954 , n160 );
not ( n9955 , n4148 );
nor ( n9956 , n155 , n156 );
nand ( n9957 , n154 , n9956 );
nand ( n9958 , n9957 , n4093 , n9839 );
not ( n9959 , n9958 );
or ( n9960 , n9955 , n9959 );
not ( n9961 , n9918 );
not ( n9962 , n4129 );
or ( n9963 , n9961 , n9962 );
nand ( n9964 , n9963 , n4041 );
nand ( n9965 , n159 , n9964 );
nand ( n9966 , n9960 , n9965 );
not ( n9967 , n9966 );
not ( n9968 , n159 );
not ( n9969 , n4238 );
nand ( n9970 , n9968 , n9969 );
nand ( n9971 , n9967 , n4081 , n9970 );
not ( n9972 , n9971 );
or ( n9973 , n9954 , n9972 );
not ( n9974 , n4073 );
not ( n9975 , n159 );
nand ( n9976 , n9974 , n4054 , n9975 );
nand ( n9977 , n9973 , n9976 );
not ( n9978 , n4054 );
not ( n9979 , n159 );
not ( n9980 , n4086 );
or ( n9981 , n9979 , n9980 );
nand ( n9982 , n4198 , n4221 );
nand ( n9983 , n9981 , n9982 );
not ( n9984 , n9983 );
or ( n9985 , n9978 , n9984 );
not ( n9986 , n9921 );
nand ( n9987 , n159 , n9986 );
nand ( n9988 , n9985 , n9987 );
nor ( n9989 , n9977 , n9988 );
not ( n9990 , n4039 );
not ( n9991 , n154 );
nand ( n9992 , n9990 , n9991 );
not ( n9993 , n9992 );
nand ( n9994 , n4226 , n9993 );
nand ( n9995 , n9953 , n9989 , n9994 );
not ( n9996 , n9995 );
not ( n9997 , n161 );
nor ( n9998 , n4147 , n9928 );
or ( n9999 , n4242 , n9998 );
nand ( n10000 , n9999 , n160 );
not ( n10001 , n159 );
nand ( n10002 , n4206 , n4227 , n9957 );
nand ( n10003 , n10001 , n10002 );
not ( n10004 , n159 );
nand ( n10005 , n10004 , n4154 );
nor ( n10006 , n4232 , n9889 );
not ( n10007 , n4196 );
not ( n10008 , n9857 );
or ( n10009 , n10007 , n10008 );
nand ( n10010 , n10009 , n4288 );
not ( n10011 , n10010 );
nand ( n10012 , n10003 , n10005 , n10006 , n10011 );
nand ( n10013 , n4054 , n10012 );
not ( n10014 , n159 );
not ( n10015 , n158 );
nand ( n10016 , n10015 , n4072 );
not ( n10017 , n158 );
nand ( n10018 , n154 , n4285 );
not ( n10019 , n10018 );
nand ( n10020 , n10017 , n10019 );
nand ( n10021 , n10016 , n4257 , n10020 );
not ( n10022 , n10021 );
or ( n10023 , n10014 , n10022 );
and ( n10024 , n159 , n160 );
not ( n10025 , n158 );
not ( n10026 , n9887 );
or ( n10027 , n10025 , n10026 );
not ( n10028 , n154 );
nand ( n10029 , n10028 , n155 );
nand ( n10030 , n10027 , n10029 );
not ( n10031 , n10030 );
not ( n10032 , n158 );
nand ( n10033 , n10032 , n4066 );
nand ( n10034 , n10031 , n9957 , n10033 );
nand ( n10035 , n10024 , n10034 );
nand ( n10036 , n10023 , n10035 );
nor ( n10037 , n4225 , n4174 );
not ( n10038 , n159 );
not ( n10039 , n10038 );
not ( n10040 , n4232 );
or ( n10041 , n10039 , n10040 );
not ( n10042 , n9915 );
nand ( n10043 , n10042 , n4115 );
nand ( n10044 , n10041 , n10043 );
nor ( n10045 , n10036 , n10037 , n10044 );
nand ( n10046 , n10000 , n10013 , n10045 );
not ( n10047 , n10046 );
or ( n10048 , n9997 , n10047 );
not ( n10049 , n4236 );
not ( n10050 , n10049 );
not ( n10051 , n4123 );
nand ( n10052 , n10051 , n4220 );
or ( n10053 , n10019 , n10052 );
nand ( n10054 , n10053 , n158 );
not ( n10055 , n10054 );
or ( n10056 , n10050 , n10055 );
nor ( n10057 , n4054 , n159 );
nand ( n10058 , n10056 , n10057 );
nand ( n10059 , n10048 , n10058 );
not ( n10060 , n10059 );
not ( n10061 , n4054 );
not ( n10062 , n159 );
nand ( n10063 , n158 , n9857 );
not ( n10064 , n10063 );
nand ( n10065 , n10062 , n10064 );
not ( n10066 , n9884 );
not ( n10067 , n10066 );
not ( n10068 , n158 );
nand ( n10069 , n10068 , n9941 );
not ( n10070 , n10069 );
not ( n10071 , n158 );
nand ( n10072 , n10071 , n9916 );
not ( n10073 , n10072 );
or ( n10074 , n10070 , n10073 );
not ( n10075 , n159 );
nand ( n10076 , n10074 , n10075 );
nand ( n10077 , n10065 , n10067 , n10076 );
not ( n10078 , n10077 );
or ( n10079 , n10061 , n10078 );
nand ( n10080 , n4042 , n4255 );
not ( n10081 , n10080 );
not ( n10082 , n4176 );
or ( n10083 , n10081 , n10082 );
not ( n10084 , n159 );
nand ( n10085 , n10083 , n10084 );
nand ( n10086 , n10079 , n10085 );
and ( n10087 , n159 , n4054 );
not ( n10088 , n10087 );
not ( n10089 , n158 );
nand ( n10090 , n10089 , n4228 );
not ( n10091 , n158 );
nor ( n10092 , n10091 , n4048 );
not ( n10093 , n10092 );
nand ( n10094 , n10090 , n10093 , n4243 );
not ( n10095 , n10094 );
or ( n10096 , n10088 , n10095 );
not ( n10097 , n158 );
not ( n10098 , n10097 );
not ( n10099 , n4072 );
nand ( n10100 , n10099 , n4100 , n4108 );
not ( n10101 , n10100 );
or ( n10102 , n10098 , n10101 );
and ( n10103 , n4283 , n9992 );
nand ( n10104 , n10102 , n10103 );
nand ( n10105 , n10024 , n10104 );
nand ( n10106 , n10096 , n10105 );
nor ( n10107 , n10086 , n10106 );
or ( n10108 , n4225 , n4193 );
nand ( n10109 , n10108 , n4166 );
nand ( n10110 , n4054 , n10109 );
not ( n10111 , n9830 );
not ( n10112 , n154 );
nor ( n10113 , n10112 , n4235 );
not ( n10114 , n10113 );
not ( n10115 , n10114 );
or ( n10116 , n10111 , n10115 );
nand ( n10117 , n10116 , n4226 );
nand ( n10118 , n10110 , n10076 , n10117 );
not ( n10119 , n4048 );
not ( n10120 , n154 );
nand ( n10121 , n10119 , n10120 );
not ( n10122 , n10121 );
nand ( n10123 , n4226 , n10122 );
not ( n10124 , n159 );
not ( n10125 , n154 );
nand ( n10126 , n10124 , n157 , n10125 );
not ( n10127 , n10126 );
not ( n10128 , n4059 );
nand ( n10129 , n10128 , n158 );
not ( n10130 , n10129 );
or ( n10131 , n10127 , n10130 );
nand ( n10132 , n10131 , n4054 );
and ( n10133 , n10123 , n10132 );
not ( n10134 , n4085 );
not ( n10135 , n4259 );
or ( n10136 , n10134 , n10135 );
not ( n10137 , n159 );
nand ( n10138 , n10136 , n10137 );
nand ( n10139 , n158 , n4183 );
not ( n10140 , n158 );
nand ( n10141 , n10140 , n4149 );
and ( n10142 , n10139 , n10141 );
not ( n10143 , n4197 );
nand ( n10144 , n10143 , n4268 );
nand ( n10145 , n4074 , n4064 );
not ( n10146 , n10145 );
not ( n10147 , n4217 );
nand ( n10148 , n10147 , n158 );
not ( n10149 , n10148 );
or ( n10150 , n10146 , n10149 );
not ( n10151 , n159 );
nand ( n10152 , n10150 , n10151 );
nand ( n10153 , n10142 , n10144 , n10152 );
nand ( n10154 , n160 , n10153 );
nand ( n10155 , n10133 , n10138 , n10154 );
or ( n10156 , n10118 , n10155 );
nand ( n10157 , n10156 , n4144 );
nand ( n10158 , n10060 , n10107 , n10157 );
not ( n10159 , n10158 );
not ( n10160 , n10159 );
and ( n10161 , n9996 , n10160 );
not ( n10162 , n9996 );
and ( n10163 , n10060 , n10107 , n10157 );
buf ( n10164 , n10163 );
and ( n10165 , n10162 , n10164 );
nor ( n10166 , n10161 , n10165 );
not ( n10167 , n10166 );
and ( n10168 , n9809 , n10167 );
and ( n10169 , n9808 , n10166 );
nor ( n10170 , n10168 , n10169 );
not ( n10171 , n10170 );
not ( n10172 , n169 );
not ( n10173 , n5393 );
or ( n10174 , n10172 , n10173 );
nand ( n10175 , n167 , n5482 );
not ( n10176 , n10175 );
not ( n10177 , n5512 );
or ( n10178 , n10176 , n10177 );
not ( n10179 , n169 );
nand ( n10180 , n10178 , n10179 );
nand ( n10181 , n10174 , n10180 );
not ( n10182 , n169 );
nor ( n10183 , n10182 , n167 );
not ( n10184 , n10183 );
not ( n10185 , n166 );
nand ( n10186 , n10185 , n5276 );
buf ( n10187 , n5235 );
nand ( n10188 , n10186 , n10187 , n5465 );
not ( n10189 , n10188 );
or ( n10190 , n10184 , n10189 );
not ( n10191 , n5539 );
not ( n10192 , n5314 );
nand ( n10193 , n10191 , n10192 );
nand ( n10194 , n10190 , n10193 );
nor ( n10195 , n10181 , n10194 );
or ( n10196 , n167 , n5573 );
or ( n10197 , n5373 , n5274 );
nand ( n10198 , n10197 , n5311 );
nand ( n10199 , n169 , n10198 );
nand ( n10200 , n10196 , n10199 );
not ( n10201 , n10200 );
not ( n10202 , n167 );
not ( n10203 , n166 );
not ( n10204 , n10203 );
not ( n10205 , n5594 );
or ( n10206 , n10204 , n10205 );
nand ( n10207 , n10206 , n5495 );
not ( n10208 , n10207 );
or ( n10209 , n10202 , n10208 );
not ( n10210 , n169 );
not ( n10211 , n5451 );
not ( n10212 , n5310 );
or ( n10213 , n10211 , n10212 );
not ( n10214 , n166 );
or ( n10215 , n10214 , n5318 );
nand ( n10216 , n10213 , n10215 );
nand ( n10217 , n10210 , n10216 );
nand ( n10218 , n10209 , n10217 );
not ( n10219 , n10218 );
nand ( n10220 , n10195 , n10201 , n10219 );
and ( n10221 , n10220 , n5449 );
not ( n10222 , n167 );
nand ( n10223 , n10222 , n5400 );
and ( n10224 , n10175 , n10223 );
not ( n10225 , n166 );
nor ( n10226 , n10224 , n10225 );
nor ( n10227 , n10221 , n10226 );
not ( n10228 , n5599 );
not ( n10229 , n10228 );
nand ( n10230 , n10229 , n167 );
not ( n10231 , n167 );
nor ( n10232 , n10231 , n5632 );
not ( n10233 , n10232 );
not ( n10234 , n5466 );
and ( n10235 , n10230 , n10233 , n10234 );
not ( n10236 , n167 );
nand ( n10237 , n5272 , n5556 );
nand ( n10238 , n166 , n10237 );
not ( n10239 , n5314 );
nand ( n10240 , n10239 , n5303 );
nand ( n10241 , n10238 , n5440 , n10240 );
nand ( n10242 , n10236 , n10241 );
nand ( n10243 , n10235 , n5489 , n10242 );
nand ( n10244 , n169 , n10243 );
not ( n10245 , n169 );
and ( n10246 , n5549 , n10193 );
not ( n10247 , n167 );
not ( n10248 , n166 );
nand ( n10249 , n10248 , n5557 );
not ( n10250 , n5329 );
not ( n10251 , n10250 );
not ( n10252 , n5388 );
nand ( n10253 , n10252 , n166 );
nand ( n10254 , n10249 , n10251 , n10253 );
nand ( n10255 , n10247 , n10254 );
not ( n10256 , n5613 );
nor ( n10257 , n166 , n5539 );
not ( n10258 , n10257 );
or ( n10259 , n5338 , n10239 );
nand ( n10260 , n10259 , n5339 );
nand ( n10261 , n5649 , n10256 , n10258 , n10260 );
nand ( n10262 , n167 , n10261 );
nand ( n10263 , n10246 , n10255 , n10262 );
nand ( n10264 , n10245 , n10263 );
not ( n10265 , n169 );
nand ( n10266 , n166 , n5644 );
and ( n10267 , n10266 , n5369 );
nand ( n10268 , n5220 , n5254 );
not ( n10269 , n10268 );
nand ( n10270 , n167 , n10269 );
not ( n10271 , n5458 );
not ( n10272 , n5360 );
or ( n10273 , n10271 , n10272 );
not ( n10274 , n167 );
nand ( n10275 , n10273 , n10274 );
nand ( n10276 , n10267 , n10270 , n10275 );
not ( n10277 , n10276 );
or ( n10278 , n10265 , n10277 );
not ( n10279 , n167 );
nand ( n10280 , n166 , n5457 );
not ( n10281 , n10280 );
not ( n10282 , n10281 );
nand ( n10283 , n5284 , n10282 , n10240 );
nand ( n10284 , n10279 , n10283 );
nand ( n10285 , n10278 , n10284 );
not ( n10286 , n167 );
not ( n10287 , n166 );
nor ( n10288 , n10287 , n5417 );
nand ( n10289 , n10286 , n10288 );
nand ( n10290 , n5353 , n10289 );
not ( n10291 , n167 );
nand ( n10292 , n10291 , n5521 );
not ( n10293 , n5422 );
nand ( n10294 , n166 , n10293 );
nand ( n10295 , n10292 , n10294 , n5462 );
nor ( n10296 , n10290 , n10295 );
or ( n10297 , n169 , n10296 );
and ( n10298 , n5220 , n5561 );
not ( n10299 , n163 );
and ( n10300 , n10299 , n5367 );
nor ( n10301 , n10298 , n10300 );
nand ( n10302 , n10301 , n5388 , n5436 );
nand ( n10303 , n167 , n10302 );
nand ( n10304 , n10297 , n10303 );
or ( n10305 , n10285 , n10304 );
nand ( n10306 , n10305 , n170 );
and ( n10307 , n10227 , n10244 , n10264 , n10306 );
and ( n10308 , n4847 , n10307 );
not ( n10309 , n4847 );
nand ( n10310 , n10227 , n10244 , n10264 , n10306 );
and ( n10311 , n10309 , n10310 );
nor ( n10312 , n10308 , n10311 );
not ( n10313 , n10312 );
not ( n10314 , n10313 );
or ( n10315 , n4310 , n4422 );
nand ( n10316 , n4330 , n10315 );
nor ( n10317 , n149 , n150 );
not ( n10318 , n10317 );
nor ( n10319 , n146 , n147 );
nand ( n10320 , n148 , n10319 );
not ( n10321 , n4326 );
not ( n10322 , n148 );
nand ( n10323 , n10321 , n10322 );
not ( n10324 , n10323 );
not ( n10325 , n10324 );
nand ( n10326 , n10320 , n4363 , n10325 );
not ( n10327 , n10326 );
or ( n10328 , n10318 , n10327 );
not ( n10329 , n148 );
nand ( n10330 , n10329 , n150 );
not ( n10331 , n10330 );
not ( n10332 , n10331 );
or ( n10333 , n4464 , n10332 );
nand ( n10334 , n10333 , n4399 );
nand ( n10335 , n149 , n10334 );
nand ( n10336 , n10328 , n10335 );
or ( n10337 , n10316 , n10336 );
nand ( n10338 , n10337 , n152 );
nand ( n10339 , n148 , n4454 );
not ( n10340 , n10339 );
nand ( n10341 , n150 , n10340 );
not ( n10342 , n4564 );
nand ( n10343 , n149 , n10342 );
and ( n10344 , n10341 , n10343 );
not ( n10345 , n149 );
nand ( n10346 , n10345 , n4532 );
nor ( n10347 , n10346 , n4322 );
not ( n10348 , n10347 );
not ( n10349 , n4463 );
not ( n10350 , n148 );
nand ( n10351 , n10350 , n4398 );
not ( n10352 , n10351 );
not ( n10353 , n10352 );
not ( n10354 , n10353 );
nand ( n10355 , n10349 , n10354 );
nand ( n10356 , n4480 , n4456 );
not ( n10357 , n10356 );
nand ( n10358 , n149 , n4385 );
not ( n10359 , n10358 );
or ( n10360 , n10357 , n10359 );
nand ( n10361 , n10360 , n4532 );
nand ( n10362 , n10348 , n10355 , n10361 );
not ( n10363 , n10362 );
and ( n10364 , n10338 , n10344 , n10363 );
not ( n10365 , n148 );
nand ( n10366 , n4419 , n4453 );
not ( n10367 , n10366 );
or ( n10368 , n10365 , n10367 );
not ( n10369 , n148 );
not ( n10370 , n4368 );
nand ( n10371 , n150 , n10370 );
or ( n10372 , n10369 , n10371 );
nand ( n10373 , n10368 , n10372 );
and ( n10374 , n149 , n10373 );
not ( n10375 , n149 );
not ( n10376 , n4328 );
not ( n10377 , n150 );
nand ( n10378 , n10376 , n10377 );
not ( n10379 , n10378 );
not ( n10380 , n10379 );
not ( n10381 , n148 );
nand ( n10382 , n10381 , n4432 );
nor ( n10383 , n150 , n10382 );
not ( n10384 , n10383 );
not ( n10385 , n4344 );
nand ( n10386 , n150 , n10385 );
nand ( n10387 , n10380 , n10384 , n10386 );
and ( n10388 , n10375 , n10387 );
nor ( n10389 , n10374 , n10388 );
not ( n10390 , n146 );
nand ( n10391 , n10390 , n147 );
or ( n10392 , n150 , n10391 );
nand ( n10393 , n10392 , n4326 , n4481 );
and ( n10394 , n149 , n10393 );
not ( n10395 , n4399 );
nor ( n10396 , n10394 , n10395 );
not ( n10397 , n10396 );
not ( n10398 , n149 );
not ( n10399 , n4361 );
not ( n10400 , n10399 );
nor ( n10401 , n150 , n10400 );
nand ( n10402 , n10398 , n10401 );
not ( n10403 , n149 );
not ( n10404 , n146 );
nor ( n10405 , n147 , n151 );
nand ( n10406 , n10403 , n10404 , n10405 );
and ( n10407 , n10402 , n10406 );
not ( n10408 , n150 );
not ( n10409 , n148 );
nor ( n10410 , n10409 , n4305 );
nand ( n10411 , n10408 , n10410 );
not ( n10412 , n4329 );
and ( n10413 , n10407 , n10411 , n10412 );
not ( n10414 , n10413 );
or ( n10415 , n10397 , n10414 );
nand ( n10416 , n10415 , n152 );
not ( n10417 , n4473 );
nand ( n10418 , n10331 , n10417 );
not ( n10419 , n4544 );
nand ( n10420 , n150 , n4454 );
not ( n10421 , n10420 );
or ( n10422 , n10419 , n10421 );
not ( n10423 , n149 );
nand ( n10424 , n10422 , n10423 );
not ( n10425 , n150 );
nand ( n10426 , n10425 , n4514 );
nand ( n10427 , n10424 , n10426 );
not ( n10428 , n10427 );
nand ( n10429 , n10428 , n4474 , n4564 );
nand ( n10430 , n149 , n4353 );
not ( n10431 , n151 );
nand ( n10432 , n10431 , n147 );
nor ( n10433 , n148 , n10432 );
nand ( n10434 , n149 , n10433 );
nor ( n10435 , n148 , n150 );
not ( n10436 , n10435 );
or ( n10437 , n4464 , n10436 );
nand ( n10438 , n10430 , n10434 , n10437 );
or ( n10439 , n10429 , n10438 );
nand ( n10440 , n10439 , n4532 );
nand ( n10441 , n10389 , n10416 , n10418 , n10440 );
and ( n10442 , n153 , n10441 );
not ( n10443 , n153 );
not ( n10444 , n149 );
nor ( n10445 , n10444 , n4349 );
not ( n10446 , n149 );
nand ( n10447 , n10446 , n10324 );
nand ( n10448 , n148 , n10385 );
not ( n10449 , n10448 );
nand ( n10450 , n150 , n10449 );
nand ( n10451 , n10447 , n4354 , n10450 );
not ( n10452 , n148 );
nand ( n10453 , n10452 , n10405 );
not ( n10454 , n10453 );
not ( n10455 , n150 );
nand ( n10456 , n10455 , n4535 );
not ( n10457 , n10456 );
or ( n10458 , n10454 , n10457 );
nand ( n10459 , n10458 , n149 );
nand ( n10460 , n4438 , n10459 );
nor ( n10461 , n10451 , n10460 );
or ( n10462 , n10461 , n4532 );
not ( n10463 , n150 );
nand ( n10464 , n10463 , n4456 );
nand ( n10465 , n10462 , n10464 );
nor ( n10466 , n10445 , n10465 );
not ( n10467 , n4462 );
nor ( n10468 , n10467 , n10453 );
not ( n10469 , n4310 );
and ( n10470 , n10469 , n4329 );
not ( n10471 , n149 );
not ( n10472 , n10471 );
not ( n10473 , n4312 );
and ( n10474 , n10472 , n10473 );
nor ( n10475 , n10474 , n10383 );
not ( n10476 , n4320 );
not ( n10477 , n4305 );
or ( n10478 , n10476 , n10477 );
nand ( n10479 , n10478 , n4480 );
nand ( n10480 , n10475 , n4384 , n10479 );
nor ( n10481 , n10470 , n10480 );
or ( n10482 , n10481 , n152 );
not ( n10483 , n149 );
nor ( n10484 , n150 , n10448 );
nor ( n10485 , n4477 , n10484 );
not ( n10486 , n10485 );
nand ( n10487 , n10483 , n10486 );
nand ( n10488 , n10482 , n10487 );
nor ( n10489 , n10468 , n10488 );
nand ( n10490 , n10466 , n10489 );
and ( n10491 , n10443 , n10490 );
nor ( n10492 , n10442 , n10491 );
nand ( n10493 , n10364 , n10492 );
not ( n10494 , n10493 );
not ( n10495 , n4405 );
not ( n10496 , n4382 );
not ( n10497 , n148 );
nand ( n10498 , n10496 , n10497 );
or ( n10499 , n4461 , n10498 );
not ( n10500 , n148 );
nand ( n10501 , n10500 , n151 );
not ( n10502 , n10501 );
not ( n10503 , n149 );
nand ( n10504 , n10502 , n10503 );
not ( n10505 , n10504 );
not ( n10506 , n4317 );
nand ( n10507 , n10506 , n150 );
not ( n10508 , n10507 );
or ( n10509 , n10505 , n10508 );
nand ( n10510 , n10509 , n4532 );
not ( n10511 , n150 );
nand ( n10512 , n10511 , n10385 );
not ( n10513 , n10512 );
not ( n10514 , n150 );
nand ( n10515 , n10514 , n10433 );
not ( n10516 , n10515 );
or ( n10517 , n10513 , n10516 );
not ( n10518 , n149 );
nand ( n10519 , n10517 , n10518 );
not ( n10520 , n10448 );
nand ( n10521 , n148 , n4374 );
not ( n10522 , n10521 );
or ( n10523 , n10520 , n10522 );
not ( n10524 , n4461 );
nand ( n10525 , n10523 , n10524 );
and ( n10526 , n10499 , n10510 , n10519 , n10525 );
not ( n10527 , n4384 );
not ( n10528 , n4536 );
or ( n10529 , n10527 , n10528 );
not ( n10530 , n149 );
nand ( n10531 , n10529 , n10530 );
not ( n10532 , n4460 );
not ( n10533 , n4482 );
or ( n10534 , n10532 , n10533 );
nand ( n10535 , n10534 , n4512 );
and ( n10536 , n4532 , n10535 );
not ( n10537 , n4532 );
not ( n10538 , n4326 );
nand ( n10539 , n10538 , n150 );
nand ( n10540 , n4480 , n4540 );
nand ( n10541 , n148 , n4340 );
not ( n10542 , n10541 );
not ( n10543 , n10420 );
or ( n10544 , n10542 , n10543 );
not ( n10545 , n149 );
nand ( n10546 , n10544 , n10545 );
nand ( n10547 , n10539 , n4525 , n10540 , n10546 );
and ( n10548 , n10537 , n10547 );
nor ( n10549 , n10536 , n10548 );
nand ( n10550 , n10526 , n10531 , n10549 );
not ( n10551 , n10550 );
or ( n10552 , n10495 , n10551 );
not ( n10553 , n150 );
nor ( n10554 , n148 , n4473 );
nand ( n10555 , n10553 , n10554 );
not ( n10556 , n10555 );
not ( n10557 , n4504 );
or ( n10558 , n10556 , n10557 );
not ( n10559 , n149 );
nand ( n10560 , n10558 , n10559 );
and ( n10561 , n149 , n4532 );
not ( n10562 , n150 );
nand ( n10563 , n10562 , n4467 );
not ( n10564 , n4391 );
nand ( n10565 , n10564 , n150 );
nand ( n10566 , n10563 , n10565 , n4444 );
nand ( n10567 , n10561 , n10566 );
not ( n10568 , n149 );
not ( n10569 , n150 );
nor ( n10570 , n10569 , n10382 );
nand ( n10571 , n10568 , n10570 );
nand ( n10572 , n10571 , n10411 , n10519 );
nand ( n10573 , n4532 , n10572 );
nand ( n10574 , n10560 , n10567 , n10573 );
not ( n10575 , n10574 );
nand ( n10576 , n10552 , n10575 );
not ( n10577 , n153 );
not ( n10578 , n10317 );
not ( n10579 , n4419 );
not ( n10580 , n10579 );
or ( n10581 , n10578 , n10580 );
nand ( n10582 , n10581 , n4444 );
nand ( n10583 , n152 , n10582 );
and ( n10584 , n4412 , n4556 );
nor ( n10585 , n149 , n4533 );
not ( n10586 , n10585 );
and ( n10587 , n10586 , n10402 );
not ( n10588 , n149 );
nand ( n10589 , n4409 , n4466 , n10320 );
and ( n10590 , n10588 , n10589 );
not ( n10591 , n10588 );
and ( n10592 , n10591 , n10383 );
nor ( n10593 , n10590 , n10592 );
nand ( n10594 , n10584 , n10587 , n10593 );
nand ( n10595 , n4532 , n10594 );
not ( n10596 , n149 );
not ( n10597 , n150 );
nand ( n10598 , n10597 , n4321 );
not ( n10599 , n4535 );
not ( n10600 , n150 );
not ( n10601 , n148 );
nor ( n10602 , n10601 , n10391 );
nand ( n10603 , n10600 , n10602 );
nand ( n10604 , n10598 , n10599 , n10603 );
not ( n10605 , n10604 );
or ( n10606 , n10596 , n10605 );
or ( n10607 , n149 , n4412 );
nand ( n10608 , n10606 , n10607 );
nor ( n10609 , n4461 , n4499 );
and ( n10610 , n149 , n152 );
not ( n10611 , n10610 );
not ( n10612 , n150 );
not ( n10613 , n10399 );
or ( n10614 , n10612 , n10613 );
not ( n10615 , n148 );
nand ( n10616 , n10615 , n146 );
nand ( n10617 , n10614 , n10616 );
not ( n10618 , n10617 );
not ( n10619 , n150 );
nand ( n10620 , n10619 , n4311 );
nand ( n10621 , n10618 , n10320 , n10620 );
not ( n10622 , n10621 );
or ( n10623 , n10611 , n10622 );
not ( n10624 , n10432 );
nand ( n10625 , n4336 , n10624 );
nand ( n10626 , n10623 , n10625 );
nor ( n10627 , n10608 , n10609 , n10626 );
nand ( n10628 , n10583 , n10595 , n10627 );
not ( n10629 , n10628 );
or ( n10630 , n10577 , n10629 );
not ( n10631 , n149 );
not ( n10632 , n150 );
nand ( n10633 , n4347 , n4455 );
nor ( n10634 , n10602 , n10633 );
or ( n10635 , n10632 , n10634 );
not ( n10636 , n4417 );
nand ( n10637 , n10635 , n10636 );
nand ( n10638 , n10631 , n10637 );
not ( n10639 , n10638 );
not ( n10640 , n150 );
not ( n10641 , n10640 );
not ( n10642 , n4321 );
nand ( n10643 , n10642 , n4365 , n4378 );
not ( n10644 , n10643 );
or ( n10645 , n10641 , n10644 );
and ( n10646 , n4562 , n10351 );
nand ( n10647 , n10645 , n10646 );
nand ( n10648 , n149 , n10647 );
not ( n10649 , n10648 );
or ( n10650 , n10639 , n10649 );
nand ( n10651 , n10650 , n152 );
nand ( n10652 , n10630 , n10651 );
nor ( n10653 , n10576 , n10652 );
buf ( n10654 , n10653 );
and ( n10655 , n10494 , n10654 );
not ( n10656 , n10494 );
nand ( n10657 , n4405 , n10550 );
nand ( n10658 , n153 , n10628 );
nand ( n10659 , n10657 , n10575 , n10651 , n10658 );
and ( n10660 , n10656 , n10659 );
nor ( n10661 , n10655 , n10660 );
not ( n10662 , n10661 );
or ( n10663 , n10314 , n10662 );
not ( n10664 , n10312 );
or ( n10665 , n10664 , n10661 );
nand ( n10666 , n10663 , n10665 );
nand ( n10667 , n10171 , n10666 );
not ( n10668 , n10666 );
nand ( n10669 , n10170 , n10668 );
nand ( n10670 , n10667 , n2352 , n10669 );
nand ( n10671 , n9802 , n10670 );
not ( n10672 , n169 );
not ( n10673 , n167 );
not ( n10674 , n10673 );
nand ( n10675 , n5645 , n5259 , n5549 );
not ( n10676 , n10675 );
or ( n10677 , n10674 , n10676 );
not ( n10678 , n167 );
and ( n10679 , n10678 , n10257 );
not ( n10680 , n10679 );
nand ( n10681 , n10677 , n10680 );
not ( n10682 , n10681 );
not ( n10683 , n5455 );
nand ( n10684 , n166 , n10683 );
not ( n10685 , n5453 );
nand ( n10686 , n166 , n10685 );
nand ( n10687 , n10686 , n5291 , n10253 );
nand ( n10688 , n167 , n10687 );
nand ( n10689 , n10682 , n10684 , n5465 , n10688 );
and ( n10690 , n10672 , n10689 );
not ( n10691 , n10672 );
not ( n10692 , n167 );
not ( n10693 , n5255 );
not ( n10694 , n10693 );
or ( n10695 , n5366 , n10694 );
nand ( n10696 , n10695 , n5650 );
nand ( n10697 , n10692 , n10696 );
not ( n10698 , n167 );
not ( n10699 , n5438 );
nand ( n10700 , n10698 , n10699 );
nand ( n10701 , n10697 , n10251 , n10700 );
and ( n10702 , n10691 , n10701 );
nor ( n10703 , n10690 , n10702 );
nand ( n10704 , n165 , n5244 );
not ( n10705 , n5229 );
nand ( n10706 , n10704 , n10705 , n5541 );
and ( n10707 , n5502 , n10706 );
nand ( n10708 , n5372 , n5310 );
not ( n10709 , n10708 );
nor ( n10710 , n10707 , n10709 );
not ( n10711 , n10193 );
not ( n10712 , n10239 );
nor ( n10713 , n10712 , n5250 );
nor ( n10714 , n10711 , n10713 );
not ( n10715 , n167 );
or ( n10716 , n10715 , n5318 );
not ( n10717 , n167 );
not ( n10718 , n168 );
not ( n10719 , n5367 );
or ( n10720 , n10718 , n10719 );
nand ( n10721 , n10720 , n5455 );
nand ( n10722 , n10717 , n10721 );
not ( n10723 , n167 );
nand ( n10724 , n164 , n5210 );
not ( n10725 , n10724 );
nand ( n10726 , n10723 , n5294 , n10725 );
nand ( n10727 , n10716 , n10722 , n10726 );
and ( n10728 , n169 , n10727 );
not ( n10729 , n169 );
not ( n10730 , n167 );
and ( n10731 , n10730 , n5319 );
not ( n10732 , n10730 );
not ( n10733 , n5295 );
and ( n10734 , n10732 , n10733 );
nor ( n10735 , n10731 , n10734 );
not ( n10736 , n167 );
not ( n10737 , n5487 );
nand ( n10738 , n10736 , n10737 );
nand ( n10739 , n5311 , n10270 );
nand ( n10740 , n5353 , n5530 , n10258 );
nor ( n10741 , n10739 , n10740 );
nand ( n10742 , n10735 , n10738 , n10741 );
and ( n10743 , n10729 , n10742 );
nor ( n10744 , n10728 , n10743 );
nand ( n10745 , n10710 , n10714 , n10744 );
and ( n10746 , n170 , n10745 );
not ( n10747 , n5518 );
or ( n10748 , n166 , n10747 );
not ( n10749 , n10737 );
nand ( n10750 , n10748 , n10749 );
and ( n10751 , n5379 , n10750 );
not ( n10752 , n5631 );
and ( n10753 , n5272 , n10752 );
not ( n10754 , n167 );
nor ( n10755 , n10753 , n10754 , n10712 );
nor ( n10756 , n10751 , n10755 );
nand ( n10757 , n169 , n5502 , n5400 );
and ( n10758 , n5467 , n10757 );
nand ( n10759 , n5502 , n10737 );
not ( n10760 , n167 );
not ( n10761 , n10266 );
nand ( n10762 , n10760 , n10761 );
and ( n10763 , n10759 , n10187 , n10762 );
not ( n10764 , n10763 );
not ( n10765 , n169 );
or ( n10766 , n5324 , n5411 );
nand ( n10767 , n10766 , n5291 );
and ( n10768 , n10765 , n10767 );
not ( n10769 , n10765 );
not ( n10770 , n167 );
not ( n10771 , n166 );
or ( n10772 , n10771 , n5351 );
not ( n10773 , n5556 );
nand ( n10774 , n166 , n10773 );
nand ( n10775 , n5406 , n10772 , n10774 );
nand ( n10776 , n10770 , n10775 );
not ( n10777 , n5589 );
not ( n10778 , n10280 );
or ( n10779 , n10777 , n10778 );
nand ( n10780 , n10779 , n167 );
nand ( n10781 , n10776 , n5570 , n10780 );
and ( n10782 , n10769 , n10781 );
nor ( n10783 , n10768 , n10782 );
not ( n10784 , n10783 );
or ( n10785 , n10764 , n10784 );
nand ( n10786 , n10785 , n5449 );
nand ( n10787 , n10756 , n10758 , n10786 );
nor ( n10788 , n10746 , n10787 );
nand ( n10789 , n10703 , n10788 );
not ( n10790 , n10789 );
not ( n10791 , n5665 );
or ( n10792 , n10790 , n10791 );
not ( n10793 , n10789 );
not ( n10794 , n5670 );
nand ( n10795 , n10793 , n10794 );
nand ( n10796 , n10792 , n10795 );
not ( n10797 , n5197 );
not ( n10798 , n5476 );
and ( n10799 , n10797 , n10798 );
nor ( n10800 , n5385 , n5475 );
and ( n10801 , n5197 , n10800 );
nor ( n10802 , n10799 , n10801 );
not ( n10803 , n10802 );
and ( n10804 , n10796 , n10803 );
not ( n10805 , n10796 );
and ( n10806 , n10805 , n10802 );
nor ( n10807 , n10804 , n10806 );
not ( n10808 , n10807 );
nand ( n10809 , n157 , n4044 );
and ( n10810 , n10809 , n4241 );
not ( n10811 , n159 );
nor ( n10812 , n10810 , n10811 );
not ( n10813 , n10812 );
not ( n10814 , n159 );
not ( n10815 , n4089 );
not ( n10816 , n4115 );
or ( n10817 , n10815 , n10816 );
nand ( n10818 , n10817 , n9992 );
nand ( n10819 , n10814 , n10818 );
not ( n10820 , n159 );
not ( n10821 , n4222 );
or ( n10822 , n10820 , n10821 );
not ( n10823 , n159 );
nand ( n10824 , n10823 , n9843 );
nand ( n10825 , n10822 , n10824 );
nand ( n10826 , n10819 , n4272 , n10825 );
not ( n10827 , n10826 );
and ( n10828 , n10813 , n10827 );
nor ( n10829 , n10828 , n4054 );
not ( n10830 , n10829 );
not ( n10831 , n159 );
nand ( n10832 , n10831 , n9900 );
not ( n10833 , n159 );
not ( n10834 , n155 );
not ( n10835 , n4115 );
or ( n10836 , n10834 , n10835 );
nand ( n10837 , n10836 , n9957 );
and ( n10838 , n10833 , n10837 );
and ( n10839 , n159 , n9903 );
nor ( n10840 , n10838 , n10839 );
nand ( n10841 , n10832 , n10840 );
nand ( n10842 , n160 , n10841 );
nand ( n10843 , n4044 , n4281 );
not ( n10844 , n9941 );
nand ( n10845 , n10114 , n10844 , n9811 );
nand ( n10846 , n4226 , n10845 );
nand ( n10847 , n10842 , n10843 , n10846 );
and ( n10848 , n4073 , n10072 );
not ( n10849 , n159 );
nand ( n10850 , n10849 , n4149 );
nand ( n10851 , n10848 , n4276 , n10850 );
not ( n10852 , n9888 );
and ( n10853 , n159 , n10852 );
not ( n10854 , n4201 );
nor ( n10855 , n10853 , n10854 );
not ( n10856 , n159 );
not ( n10857 , n9904 );
nand ( n10858 , n10856 , n10857 );
nand ( n10859 , n10855 , n4092 , n10858 );
or ( n10860 , n10851 , n10859 );
nand ( n10861 , n10860 , n4054 );
nand ( n10862 , n4198 , n4154 );
nand ( n10863 , n10861 , n10862 , n4152 , n161 );
or ( n10864 , n10847 , n10863 );
nor ( n10865 , n161 , n4080 );
and ( n10866 , n159 , n4242 );
nor ( n10867 , n159 , n4110 );
nand ( n10868 , n10042 , n9866 );
and ( n10869 , n9884 , n10868 );
nor ( n10870 , n10869 , n160 );
nor ( n10871 , n10866 , n10867 , n10870 );
nand ( n10872 , n158 , n4173 );
and ( n10873 , n158 , n4070 );
not ( n10874 , n10873 );
and ( n10875 , n10872 , n10874 , n9822 );
nor ( n10876 , n10875 , n159 );
not ( n10877 , n10876 );
not ( n10878 , n10139 );
not ( n10879 , n10878 );
not ( n10880 , n10033 );
not ( n10881 , n4036 );
or ( n10882 , n10880 , n10881 );
nand ( n10883 , n10882 , n159 );
nand ( n10884 , n10877 , n10879 , n10883 );
nand ( n10885 , n160 , n10884 );
nand ( n10886 , n10865 , n10871 , n10885 );
nand ( n10887 , n10864 , n10886 );
not ( n10888 , n4054 );
not ( n10889 , n9957 );
and ( n10890 , n158 , n10889 );
nand ( n10891 , n4148 , n4107 );
not ( n10892 , n10891 );
nor ( n10893 , n10890 , n4185 , n10892 );
and ( n10894 , n158 , n9956 );
or ( n10895 , n10894 , n10066 , n4264 );
nand ( n10896 , n10895 , n159 );
not ( n10897 , n4259 );
or ( n10898 , n10897 , n9936 , n4109 );
not ( n10899 , n159 );
nand ( n10900 , n10898 , n10899 );
nand ( n10901 , n10893 , n10896 , n10900 );
not ( n10902 , n10901 );
or ( n10903 , n10888 , n10902 );
not ( n10904 , n9970 );
and ( n10905 , n4191 , n4235 );
not ( n10906 , n154 );
nand ( n10907 , n10906 , n159 );
nor ( n10908 , n10905 , n158 , n10907 );
nor ( n10909 , n10904 , n10908 );
nand ( n10910 , n10903 , n10909 );
not ( n10911 , n10910 );
nand ( n10912 , n10830 , n10887 , n10911 );
not ( n10913 , n10912 );
not ( n10914 , n10913 );
and ( n10915 , n10466 , n10489 );
nor ( n10916 , n10915 , n153 );
not ( n10917 , n10916 );
nand ( n10918 , n10416 , n10418 , n10440 );
not ( n10919 , n10389 );
or ( n10920 , n10918 , n10919 );
nand ( n10921 , n10920 , n153 );
nand ( n10922 , n10917 , n10364 , n10921 );
not ( n10923 , n10922 );
not ( n10924 , n10923 );
or ( n10925 , n10914 , n10924 );
not ( n10926 , n10912 );
not ( n10927 , n10926 );
not ( n10928 , n10927 );
or ( n10929 , n10928 , n10923 );
nand ( n10930 , n10925 , n10929 );
and ( n10931 , n10160 , n338 );
not ( n10932 , n10160 );
not ( n10933 , n338 );
and ( n10934 , n10932 , n10933 );
nor ( n10935 , n10931 , n10934 );
not ( n10936 , n10935 );
and ( n10937 , n10930 , n10936 );
not ( n10938 , n10930 );
and ( n10939 , n10938 , n10935 );
nor ( n10940 , n10937 , n10939 );
not ( n10941 , n10940 );
or ( n10942 , n10808 , n10941 );
nand ( n10943 , n10942 , n2352 );
nor ( n10944 , n10940 , n10807 );
or ( n10945 , n10943 , n10944 );
and ( n10946 , n339 , n10933 );
not ( n10947 , n339 );
and ( n10948 , n10947 , n338 );
nor ( n10949 , n10946 , n10948 );
or ( n10950 , n2352 , n10949 );
nand ( n10951 , n10945 , n10950 );
not ( n10952 , n8929 );
not ( n10953 , n10952 );
not ( n10954 , n10953 );
xor ( n10955 , n359 , n9063 );
not ( n10956 , n10955 );
or ( n10957 , n10954 , n10956 );
not ( n10958 , n10952 );
or ( n10959 , n10958 , n10955 );
nand ( n10960 , n10957 , n10959 );
not ( n10961 , n202 );
not ( n10962 , n8418 );
and ( n10963 , n10961 , n10962 );
not ( n10964 , n4004 );
not ( n10965 , n202 );
nand ( n10966 , n10965 , n8288 );
not ( n10967 , n10966 );
nor ( n10968 , n10963 , n10964 , n10967 );
not ( n10969 , n10968 );
not ( n10970 , n203 );
not ( n10971 , n10970 );
not ( n10972 , n3898 );
not ( n10973 , n9636 );
and ( n10974 , n10972 , n10973 );
nor ( n10975 , n10974 , n3864 );
not ( n10976 , n3868 );
nor ( n10977 , n8424 , n3763 );
not ( n10978 , n10977 );
nand ( n10979 , n10978 , n3909 );
not ( n10980 , n10979 );
or ( n10981 , n10976 , n10980 );
nand ( n10982 , n10981 , n202 );
not ( n10983 , n202 );
not ( n10984 , n201 );
nand ( n10985 , n10984 , n3912 );
not ( n10986 , n3806 );
nand ( n10987 , n10985 , n10986 , n8412 );
nand ( n10988 , n10983 , n10987 );
nand ( n10989 , n10975 , n10982 , n10988 );
not ( n10990 , n10989 );
or ( n10991 , n10971 , n10990 );
nand ( n10992 , n3999 , n8411 );
not ( n10993 , n202 );
not ( n10994 , n8312 );
nand ( n10995 , n10993 , n10994 );
nand ( n10996 , n201 , n3893 );
nand ( n10997 , n10992 , n10995 , n10996 );
nand ( n10998 , n203 , n10997 );
nand ( n10999 , n10991 , n10998 );
nor ( n11000 , n10969 , n10999 );
not ( n11001 , n202 );
nand ( n11002 , n11001 , n3813 );
and ( n11003 , n10995 , n11002 );
not ( n11004 , n203 );
or ( n11005 , n3898 , n3954 );
or ( n11006 , n3998 , n3891 );
nand ( n11007 , n11005 , n11006 );
nand ( n11008 , n11004 , n11007 );
nand ( n11009 , n199 , n3890 );
not ( n11010 , n11009 );
nand ( n11011 , n11010 , n3904 );
not ( n11012 , n203 );
not ( n11013 , n3909 );
not ( n11014 , n3857 );
or ( n11015 , n11013 , n11014 );
nand ( n11016 , n11015 , n8403 );
nand ( n11017 , n11012 , n11016 );
and ( n11018 , n11008 , n11011 , n11017 );
nand ( n11019 , n11003 , n11018 );
not ( n11020 , n203 );
nand ( n11021 , n201 , n3976 );
not ( n11022 , n3802 );
nand ( n11023 , n11021 , n11022 , n3965 , n9617 );
not ( n11024 , n202 );
not ( n11025 , n201 );
nand ( n11026 , n11025 , n3971 );
not ( n11027 , n3755 );
nand ( n11028 , n11026 , n11027 , n9572 );
nand ( n11029 , n11024 , n11028 );
not ( n11030 , n3771 );
not ( n11031 , n8311 );
not ( n11032 , n9569 );
or ( n11033 , n11031 , n11032 );
nand ( n11034 , n11033 , n202 );
nand ( n11035 , n11029 , n11030 , n11034 );
nor ( n11036 , n11023 , n11035 );
or ( n11037 , n11020 , n11036 );
nand ( n11038 , n8379 , n9679 );
and ( n11039 , n202 , n11038 );
not ( n11040 , n201 );
not ( n11041 , n3890 );
nor ( n11042 , n11041 , n199 );
not ( n11043 , n11042 );
or ( n11044 , n11040 , n11043 );
nand ( n11045 , n11044 , n11021 );
and ( n11046 , n202 , n11045 );
nor ( n11047 , n11039 , n11046 );
nand ( n11048 , n11037 , n11047 , n3894 );
or ( n11049 , n11019 , n11048 );
nand ( n11050 , n11049 , n4008 );
not ( n11051 , n203 );
and ( n11052 , n9757 , n3910 );
nand ( n11053 , n11052 , n3932 , n3874 );
not ( n11054 , n11053 );
or ( n11055 , n11051 , n11054 );
not ( n11056 , n3868 );
nand ( n11057 , n202 , n11056 );
nand ( n11058 , n11055 , n11057 );
not ( n11059 , n11058 );
nand ( n11060 , n198 , n9672 );
nand ( n11061 , n11060 , n11009 , n3954 );
nand ( n11062 , n3880 , n11061 );
nand ( n11063 , n3999 , n3765 );
not ( n11064 , n9536 );
not ( n11065 , n3973 );
or ( n11066 , n11064 , n11065 );
not ( n11067 , n202 );
nand ( n11068 , n11066 , n11067 );
and ( n11069 , n11062 , n11063 , n11068 );
not ( n11070 , n203 );
not ( n11071 , n11070 );
not ( n11072 , n202 );
not ( n11073 , n11072 );
not ( n11074 , n8273 );
or ( n11075 , n11073 , n11074 );
or ( n11076 , n8332 , n8305 );
nand ( n11077 , n11076 , n202 );
nand ( n11078 , n11075 , n11077 );
nor ( n11079 , n9696 , n11078 );
not ( n11080 , n9576 );
nand ( n11081 , n11079 , n11080 , n3868 );
not ( n11082 , n11081 );
or ( n11083 , n11071 , n11082 );
not ( n11084 , n202 );
nand ( n11085 , n11084 , n3806 );
nand ( n11086 , n11083 , n11085 );
not ( n11087 , n11086 );
nand ( n11088 , n9672 , n3790 );
nand ( n11089 , n11059 , n11069 , n11087 , n11088 );
nand ( n11090 , n204 , n11089 );
nand ( n11091 , n11000 , n11050 , n11090 );
not ( n11092 , n11091 );
not ( n11093 , n3275 );
nor ( n11094 , n185 , n3341 );
not ( n11095 , n3013 );
nand ( n11096 , n184 , n8805 );
and ( n11097 , n3438 , n11096 );
nand ( n11098 , n185 , n3278 );
not ( n11099 , n185 );
nand ( n11100 , n11099 , n3124 );
nand ( n11101 , n11097 , n11098 , n11100 );
not ( n11102 , n11101 );
or ( n11103 , n11095 , n11102 );
nand ( n11104 , n11103 , n3246 );
nor ( n11105 , n11094 , n11104 );
not ( n11106 , n186 );
not ( n11107 , n3296 );
nand ( n11108 , n11107 , n185 );
not ( n11109 , n11108 );
not ( n11110 , n3235 );
nand ( n11111 , n11110 , n184 );
not ( n11112 , n11111 );
nor ( n11113 , n11109 , n11112 );
not ( n11114 , n3439 );
nand ( n11115 , n11114 , n3347 );
not ( n11116 , n185 );
not ( n11117 , n184 );
nand ( n11118 , n11117 , n3054 );
nand ( n11119 , n11118 , n3071 , n3176 );
nand ( n11120 , n11116 , n11119 );
nand ( n11121 , n11113 , n11115 , n11120 );
not ( n11122 , n11121 );
or ( n11123 , n11106 , n11122 );
not ( n11124 , n3326 );
not ( n11125 , n184 );
nand ( n11126 , n11124 , n11125 );
not ( n11127 , n11126 );
not ( n11128 , n3386 );
or ( n11129 , n11127 , n11128 );
nand ( n11130 , n11129 , n185 );
nand ( n11131 , n11123 , n11130 );
not ( n11132 , n11131 );
nand ( n11133 , n11105 , n11132 );
not ( n11134 , n11133 );
or ( n11135 , n11093 , n11134 );
nand ( n11136 , n185 , n3239 );
nand ( n11137 , n185 , n3397 );
and ( n11138 , n11136 , n11137 , n3178 );
not ( n11139 , n185 );
not ( n11140 , n184 );
nand ( n11141 , n3088 , n3002 );
not ( n11142 , n11141 );
or ( n11143 , n11140 , n11142 );
nand ( n11144 , n11143 , n8821 , n3221 );
nand ( n11145 , n11139 , n11144 );
nand ( n11146 , n11138 , n3319 , n11145 );
nand ( n11147 , n186 , n11146 );
nand ( n11148 , n11135 , n11147 );
not ( n11149 , n3013 );
and ( n11150 , n3432 , n3246 );
not ( n11151 , n185 );
or ( n11152 , n184 , n3345 );
nand ( n11153 , n11152 , n8828 , n9130 );
nand ( n11154 , n11151 , n11153 );
nand ( n11155 , n3293 , n9215 );
nand ( n11156 , n3253 , n3415 , n9207 );
or ( n11157 , n11155 , n11156 );
nand ( n11158 , n11157 , n185 );
nand ( n11159 , n11150 , n11154 , n11158 );
not ( n11160 , n11159 );
or ( n11161 , n11149 , n11160 );
not ( n11162 , n185 );
nand ( n11163 , n11162 , n3180 );
and ( n11164 , n11163 , n8834 , n3041 );
nand ( n11165 , n184 , n3306 );
nand ( n11166 , n185 , n8792 );
nand ( n11167 , n3013 , n11164 , n11165 , n11166 );
not ( n11168 , n11167 );
nand ( n11169 , n185 , n3133 );
not ( n11170 , n8861 );
not ( n11171 , n3143 );
or ( n11172 , n11170 , n11171 );
not ( n11173 , n185 );
nand ( n11174 , n11172 , n11173 );
nand ( n11175 , n11169 , n11174 );
not ( n11176 , n11175 );
nand ( n11177 , n186 , n11176 , n3216 , n8882 );
not ( n11178 , n11177 );
or ( n11179 , n11168 , n11178 );
nand ( n11180 , n183 , n3146 );
and ( n11181 , n11180 , n3023 );
not ( n11182 , n185 );
nor ( n11183 , n11181 , n11182 );
not ( n11184 , n185 );
not ( n11185 , n11184 );
nand ( n11186 , n3221 , n9135 , n8863 );
not ( n11187 , n11186 );
or ( n11188 , n11185 , n11187 );
not ( n11189 , n3350 );
or ( n11190 , n183 , n11189 );
nand ( n11191 , n11190 , n3222 );
nand ( n11192 , n185 , n11191 );
nand ( n11193 , n11188 , n11192 );
nor ( n11194 , n11183 , n11193 );
nand ( n11195 , n11179 , n11194 );
nand ( n11196 , n187 , n11195 );
nand ( n11197 , n11161 , n11196 );
nor ( n11198 , n11148 , n11197 );
not ( n11199 , n185 );
nand ( n11200 , n184 , n8895 );
not ( n11201 , n11200 );
and ( n11202 , n11199 , n11201 );
and ( n11203 , n3258 , n3278 );
nor ( n11204 , n11202 , n11203 );
nand ( n11205 , n11198 , n11204 );
not ( n11206 , n11205 );
not ( n11207 , n8609 );
or ( n11208 , n11206 , n11207 );
not ( n11209 , n11205 );
nand ( n11210 , n11209 , n8608 );
nand ( n11211 , n11208 , n11210 );
and ( n11212 , n11092 , n11211 );
not ( n11213 , n11092 );
not ( n11214 , n11211 );
and ( n11215 , n11213 , n11214 );
nor ( n11216 , n11212 , n11215 );
nor ( n11217 , n10960 , n11216 );
not ( n11218 , n10960 );
not ( n11219 , n11216 );
or ( n11220 , n11218 , n11219 );
nand ( n11221 , n11220 , n2352 );
or ( n11222 , n11217 , n11221 );
xnor ( n11223 , n359 , n360 );
or ( n11224 , n2352 , n11223 );
nand ( n11225 , n11222 , n11224 );
not ( n11226 , n371 );
and ( n11227 , n372 , n11226 );
not ( n11228 , n372 );
and ( n11229 , n11228 , n371 );
nor ( n11230 , n11227 , n11229 );
or ( n11231 , n2352 , n11230 );
not ( n11232 , n11226 );
not ( n11233 , n7089 );
or ( n11234 , n11232 , n11233 );
or ( n11235 , n7107 , n11226 );
nand ( n11236 , n11234 , n11235 );
not ( n11237 , n11236 );
not ( n11238 , n6569 );
nor ( n11239 , n6543 , n6785 );
nor ( n11240 , n11238 , n11239 );
not ( n11241 , n140 );
nand ( n11242 , n11241 , n142 );
or ( n11243 , n6662 , n11242 );
nand ( n11244 , n11243 , n6645 );
nand ( n11245 , n141 , n11244 );
nor ( n11246 , n141 , n142 );
nor ( n11247 , n138 , n139 );
nand ( n11248 , n140 , n11247 );
not ( n11249 , n6787 );
nor ( n11250 , n140 , n11249 );
not ( n11251 , n11250 );
nand ( n11252 , n6623 , n11248 , n11251 );
nand ( n11253 , n11246 , n11252 );
and ( n11254 , n11240 , n11245 , n11253 );
not ( n11255 , n144 );
nor ( n11256 , n11254 , n11255 );
not ( n11257 , n142 );
nand ( n11258 , n140 , n6656 );
nor ( n11259 , n11257 , n11258 );
not ( n11260 , n11259 );
not ( n11261 , n141 );
or ( n11262 , n11261 , n6708 );
nand ( n11263 , n11260 , n11262 );
not ( n11264 , n6661 );
nor ( n11265 , n140 , n6749 );
nand ( n11266 , n11264 , n11265 );
not ( n11267 , n6559 );
nor ( n11268 , n141 , n144 );
nand ( n11269 , n11267 , n11268 );
not ( n11270 , n144 );
not ( n11271 , n141 );
not ( n11272 , n6610 );
or ( n11273 , n11271 , n11272 );
nand ( n11274 , n6795 , n6658 );
nand ( n11275 , n11273 , n11274 );
nand ( n11276 , n11270 , n11275 );
nand ( n11277 , n11266 , n11269 , n11276 );
nor ( n11278 , n11256 , n11263 , n11277 );
not ( n11279 , n140 );
not ( n11280 , n6655 );
not ( n11281 , n11280 );
nand ( n11282 , n6696 , n11281 );
not ( n11283 , n11282 );
or ( n11284 , n11279 , n11283 );
not ( n11285 , n6561 );
nand ( n11286 , n11285 , n142 );
not ( n11287 , n11286 );
nand ( n11288 , n11287 , n140 );
nand ( n11289 , n11284 , n11288 );
and ( n11290 , n141 , n11289 );
not ( n11291 , n141 );
not ( n11292 , n6565 );
not ( n11293 , n142 );
nand ( n11294 , n11292 , n11293 );
not ( n11295 , n11294 );
not ( n11296 , n11295 );
not ( n11297 , n140 );
nand ( n11298 , n11297 , n6736 );
nor ( n11299 , n142 , n11298 );
not ( n11300 , n11299 );
not ( n11301 , n6584 );
nand ( n11302 , n142 , n11301 );
nand ( n11303 , n11296 , n11300 , n11302 );
and ( n11304 , n11291 , n11303 );
nor ( n11305 , n11290 , n11304 );
not ( n11306 , n141 );
not ( n11307 , n142 );
not ( n11308 , n6704 );
nand ( n11309 , n11307 , n11308 );
nand ( n11310 , n11309 , n6797 , n11249 );
not ( n11311 , n11310 );
or ( n11312 , n11306 , n11311 );
nand ( n11313 , n11312 , n6645 );
not ( n11314 , n11313 );
not ( n11315 , n142 );
not ( n11316 , n140 );
nor ( n11317 , n11316 , n6539 );
nand ( n11318 , n11315 , n11317 );
and ( n11319 , n11318 , n6567 );
not ( n11320 , n141 );
nor ( n11321 , n142 , n6621 );
nand ( n11322 , n11320 , n11321 );
not ( n11323 , n141 );
nand ( n11324 , n11323 , n6635 );
and ( n11325 , n11322 , n11324 );
nand ( n11326 , n11314 , n11319 , n11325 );
nand ( n11327 , n144 , n11326 );
not ( n11328 , n11242 );
nand ( n11329 , n11328 , n6701 );
or ( n11330 , n6662 , n6640 );
not ( n11331 , n141 );
not ( n11332 , n140 );
not ( n11333 , n138 );
nor ( n11334 , n11333 , n143 );
nand ( n11335 , n11332 , n11334 );
or ( n11336 , n11331 , n11335 );
nand ( n11337 , n141 , n6591 );
nand ( n11338 , n11330 , n11336 , n11337 );
not ( n11339 , n142 );
nor ( n11340 , n140 , n143 );
nand ( n11341 , n11339 , n11340 );
not ( n11342 , n11341 );
nand ( n11343 , n6669 , n11342 );
not ( n11344 , n6688 );
nand ( n11345 , n142 , n11280 );
not ( n11346 , n11345 );
or ( n11347 , n11344 , n11346 );
not ( n11348 , n141 );
nand ( n11349 , n11347 , n11348 );
nand ( n11350 , n11343 , n11349 );
not ( n11351 , n11350 );
nand ( n11352 , n11351 , n6801 , n6708 );
or ( n11353 , n11338 , n11352 );
not ( n11354 , n144 );
nand ( n11355 , n11353 , n11354 );
nand ( n11356 , n11305 , n11327 , n11329 , n11355 );
and ( n11357 , n137 , n11356 );
not ( n11358 , n137 );
not ( n11359 , n140 );
nor ( n11360 , n138 , n143 );
nand ( n11361 , n11359 , n11360 );
not ( n11362 , n11361 );
nand ( n11363 , n11264 , n11362 );
not ( n11364 , n141 );
not ( n11365 , n6584 );
nand ( n11366 , n11365 , n140 );
not ( n11367 , n11366 );
not ( n11368 , n142 );
nand ( n11369 , n11367 , n11368 );
nand ( n11370 , n6802 , n11369 );
nand ( n11371 , n11364 , n11370 );
not ( n11372 , n6566 );
nor ( n11373 , n11372 , n6543 );
not ( n11374 , n141 );
nor ( n11375 , n11374 , n6548 );
nor ( n11376 , n11375 , n11299 );
not ( n11377 , n6539 );
not ( n11378 , n6556 );
or ( n11379 , n11377 , n11378 );
nand ( n11380 , n11379 , n6795 );
nand ( n11381 , n11376 , n6777 , n11380 );
or ( n11382 , n11373 , n11381 );
not ( n11383 , n144 );
nand ( n11384 , n11382 , n11383 );
and ( n11385 , n11363 , n11371 , n11384 );
not ( n11386 , n6587 );
nand ( n11387 , n141 , n11386 );
not ( n11388 , n142 );
nand ( n11389 , n11388 , n6658 );
not ( n11390 , n141 );
nand ( n11391 , n11390 , n11250 );
not ( n11392 , n11366 );
nand ( n11393 , n11392 , n142 );
nand ( n11394 , n11391 , n6592 , n11393 );
not ( n11395 , n11361 );
not ( n11396 , n142 );
not ( n11397 , n6672 );
nand ( n11398 , n11396 , n11397 );
not ( n11399 , n11398 );
or ( n11400 , n11395 , n11399 );
nand ( n11401 , n11400 , n141 );
nand ( n11402 , n6742 , n11401 );
or ( n11403 , n11394 , n11402 );
nand ( n11404 , n11403 , n144 );
nand ( n11405 , n11385 , n11387 , n11389 , n11404 );
and ( n11406 , n11358 , n11405 );
nor ( n11407 , n11357 , n11406 );
nand ( n11408 , n11278 , n11407 );
not ( n11409 , n11408 );
not ( n11410 , n6808 );
not ( n11411 , n6777 );
not ( n11412 , n6674 );
or ( n11413 , n11411 , n11412 );
not ( n11414 , n141 );
nand ( n11415 , n11413 , n11414 );
not ( n11416 , n11415 );
not ( n11417 , n11416 );
not ( n11418 , n142 );
nand ( n11419 , n11418 , n11301 );
not ( n11420 , n11419 );
not ( n11421 , n11335 );
not ( n11422 , n142 );
nand ( n11423 , n11421 , n11422 );
not ( n11424 , n11423 );
or ( n11425 , n11420 , n11424 );
not ( n11426 , n141 );
nand ( n11427 , n11425 , n11426 );
not ( n11428 , n11366 );
and ( n11429 , n140 , n6599 );
not ( n11430 , n11429 );
not ( n11431 , n11430 );
or ( n11432 , n11428 , n11431 );
nand ( n11433 , n11432 , n11264 );
nand ( n11434 , n11427 , n11433 );
not ( n11435 , n144 );
not ( n11436 , n11435 );
not ( n11437 , n140 );
nand ( n11438 , n11437 , n143 );
or ( n11439 , n141 , n11438 );
nand ( n11440 , n142 , n6553 );
nand ( n11441 , n11439 , n11440 );
not ( n11442 , n11441 );
or ( n11443 , n11436 , n11442 );
not ( n11444 , n6605 );
not ( n11445 , n11444 );
not ( n11446 , n140 );
nand ( n11447 , n11445 , n11446 );
not ( n11448 , n11447 );
nand ( n11449 , n11448 , n11264 );
nand ( n11450 , n11443 , n11449 );
nor ( n11451 , n11434 , n11450 );
not ( n11452 , n6788 );
nand ( n11453 , n142 , n11452 );
nand ( n11454 , n6795 , n6684 );
nand ( n11455 , n140 , n6579 );
not ( n11456 , n11455 );
not ( n11457 , n11345 );
or ( n11458 , n11456 , n11457 );
not ( n11459 , n141 );
nand ( n11460 , n11458 , n11459 );
nand ( n11461 , n11453 , n6751 , n11454 , n11460 );
and ( n11462 , n144 , n11461 );
not ( n11463 , n144 );
not ( n11464 , n11264 );
not ( n11465 , n6798 );
or ( n11466 , n11464 , n11465 );
nand ( n11467 , n11466 , n6762 );
and ( n11468 , n11463 , n11467 );
nor ( n11469 , n11462 , n11468 );
nand ( n11470 , n11417 , n11451 , n11469 );
not ( n11471 , n11470 );
or ( n11472 , n11410 , n11471 );
not ( n11473 , n6723 );
not ( n11474 , n140 );
nor ( n11475 , n11474 , n6704 );
nand ( n11476 , n6587 , n6657 );
or ( n11477 , n11475 , n11476 );
nand ( n11478 , n11477 , n142 );
not ( n11479 , n11478 );
or ( n11480 , n11473 , n11479 );
not ( n11481 , n141 );
nand ( n11482 , n11480 , n11481 );
not ( n11483 , n11482 );
not ( n11484 , n142 );
not ( n11485 , n11484 );
nand ( n11486 , n6558 , n6626 , n6602 );
not ( n11487 , n11486 );
or ( n11488 , n11485 , n11487 );
not ( n11489 , n11265 );
and ( n11490 , n6702 , n11489 );
nand ( n11491 , n11488 , n11490 );
nand ( n11492 , n141 , n11491 );
not ( n11493 , n11492 );
or ( n11494 , n11483 , n11493 );
nand ( n11495 , n11494 , n144 );
nand ( n11496 , n11472 , n11495 );
not ( n11497 , n11496 );
and ( n11498 , n141 , n144 );
not ( n11499 , n6669 );
not ( n11500 , n140 );
and ( n11501 , n11499 , n11500 );
and ( n11502 , n142 , n6622 );
nor ( n11503 , n11501 , n11502 );
not ( n11504 , n142 );
not ( n11505 , n6546 );
and ( n11506 , n11504 , n11505 );
not ( n11507 , n11506 );
nand ( n11508 , n11503 , n11248 , n11507 );
nand ( n11509 , n11498 , n11508 );
not ( n11510 , n11509 );
not ( n11511 , n141 );
not ( n11512 , n11511 );
not ( n11513 , n6719 );
or ( n11514 , n11512 , n11513 );
or ( n11515 , n6661 , n6772 );
nand ( n11516 , n11514 , n11515 );
nor ( n11517 , n11510 , n11516 );
not ( n11518 , n144 );
not ( n11519 , n11246 );
nor ( n11520 , n11519 , n6696 );
nor ( n11521 , n6732 , n11520 );
or ( n11522 , n11518 , n11521 );
not ( n11523 , n142 );
nand ( n11524 , n11523 , n6557 );
not ( n11525 , n142 );
nand ( n11526 , n11525 , n11475 );
nand ( n11527 , n11524 , n6672 , n11526 );
nand ( n11528 , n141 , n11527 );
nand ( n11529 , n11522 , n11528 );
not ( n11530 , n11529 );
nand ( n11531 , n6575 , n11334 );
and ( n11532 , n6718 , n6706 );
not ( n11533 , n141 );
not ( n11534 , n6700 );
nand ( n11535 , n11533 , n11534 );
and ( n11536 , n11535 , n11322 );
not ( n11537 , n141 );
nand ( n11538 , n6716 , n6664 , n11248 );
and ( n11539 , n11537 , n11538 );
not ( n11540 , n11537 );
and ( n11541 , n11540 , n11299 );
nor ( n11542 , n11539 , n11541 );
nand ( n11543 , n11532 , n11536 , n11542 );
not ( n11544 , n144 );
nand ( n11545 , n11543 , n11544 );
nand ( n11546 , n11517 , n11530 , n11531 , n11545 );
and ( n11547 , n137 , n11546 );
nand ( n11548 , n6641 , n11534 );
not ( n11549 , n11548 );
not ( n11550 , n6779 );
or ( n11551 , n11549 , n11550 );
not ( n11552 , n141 );
nand ( n11553 , n11551 , n11552 );
not ( n11554 , n144 );
and ( n11555 , n141 , n11554 );
not ( n11556 , n142 );
not ( n11557 , n6664 );
nand ( n11558 , n11556 , n11557 );
not ( n11559 , n6635 );
not ( n11560 , n11559 );
nand ( n11561 , n11560 , n142 );
nand ( n11562 , n11558 , n11561 , n6733 );
nand ( n11563 , n11555 , n11562 );
not ( n11564 , n144 );
not ( n11565 , n141 );
not ( n11566 , n11298 );
nand ( n11567 , n11565 , n142 , n11566 );
nand ( n11568 , n11567 , n11318 , n11427 );
nand ( n11569 , n11564 , n11568 );
nand ( n11570 , n11553 , n11563 , n11569 );
nor ( n11571 , n11547 , n11570 );
nand ( n11572 , n11497 , n11571 );
buf ( n11573 , n11572 );
and ( n11574 , n11409 , n11573 );
not ( n11575 , n11409 );
nand ( n11576 , n6808 , n11470 );
not ( n11577 , n11570 );
nand ( n11578 , n137 , n11546 );
and ( n11579 , n11495 , n11576 , n11577 , n11578 );
not ( n11580 , n11579 );
not ( n11581 , n11580 );
and ( n11582 , n11575 , n11581 );
nor ( n11583 , n11574 , n11582 );
not ( n11584 , n11583 );
and ( n11585 , n11237 , n11584 );
and ( n11586 , n11236 , n11583 );
nor ( n11587 , n11585 , n11586 );
not ( n11588 , n11587 );
not ( n11589 , n117 );
not ( n11590 , n11589 );
and ( n11591 , n116 , n7376 );
nand ( n11592 , n115 , n11591 );
nand ( n11593 , n7556 , n11592 , n7581 );
not ( n11594 , n11593 );
or ( n11595 , n11590 , n11594 );
not ( n11596 , n7346 );
nor ( n11597 , n116 , n117 );
nand ( n11598 , n11596 , n11597 );
nand ( n11599 , n11595 , n11598 );
nor ( n11600 , n112 , n114 );
nand ( n11601 , n115 , n11600 );
not ( n11602 , n11601 );
nand ( n11603 , n116 , n11602 );
nand ( n11604 , n116 , n11600 );
not ( n11605 , n116 );
not ( n11606 , n112 );
nor ( n11607 , n11606 , n113 );
nand ( n11608 , n115 , n11607 );
not ( n11609 , n11608 );
nand ( n11610 , n11605 , n11609 );
not ( n11611 , n11610 );
not ( n11612 , n11611 );
nand ( n11613 , n11604 , n11612 , n7588 );
nand ( n11614 , n117 , n11613 );
nand ( n11615 , n11603 , n7382 , n11614 );
nor ( n11616 , n11599 , n11615 );
or ( n11617 , n118 , n11616 );
and ( n11618 , n117 , n118 );
not ( n11619 , n116 );
not ( n11620 , n11619 );
nor ( n11621 , n113 , n115 );
not ( n11622 , n11621 );
or ( n11623 , n11620 , n11622 );
not ( n11624 , n7441 );
nand ( n11625 , n11623 , n11624 );
nand ( n11626 , n11618 , n11625 );
nand ( n11627 , n11617 , n11626 );
not ( n11628 , n117 );
nand ( n11629 , n11628 , n7446 );
not ( n11630 , n7451 );
not ( n11631 , n7476 );
not ( n11632 , n11631 );
or ( n11633 , n11630 , n11632 );
nand ( n11634 , n11633 , n117 , n7349 );
nand ( n11635 , n11629 , n11634 );
nor ( n11636 , n11627 , n11635 );
not ( n11637 , n7376 );
not ( n11638 , n11637 );
nand ( n11639 , n7512 , n11638 );
not ( n11640 , n7333 );
not ( n11641 , n115 );
nand ( n11642 , n11640 , n11641 );
not ( n11643 , n11642 );
not ( n11644 , n11643 );
and ( n11645 , n11639 , n11644 );
or ( n11646 , n117 , n11645 );
nand ( n11647 , n115 , n7456 );
not ( n11648 , n11647 );
nand ( n11649 , n11648 , n116 );
or ( n11650 , n117 , n11649 );
nand ( n11651 , n11646 , n11650 , n7593 );
and ( n11652 , n118 , n11651 );
not ( n11653 , n117 );
nand ( n11654 , n116 , n118 );
not ( n11655 , n7490 );
nor ( n11656 , n11653 , n11654 , n11655 );
nor ( n11657 , n11652 , n11656 );
not ( n11658 , n118 );
nand ( n11659 , n112 , n113 );
or ( n11660 , n11659 , n7484 );
not ( n11661 , n11611 );
nand ( n11662 , n11660 , n11661 );
and ( n11663 , n11658 , n11662 );
not ( n11664 , n11658 );
not ( n11665 , n117 );
not ( n11666 , n112 );
nand ( n11667 , n11666 , n113 );
nor ( n11668 , n115 , n11667 );
not ( n11669 , n11668 );
nand ( n11670 , n116 , n7400 );
not ( n11671 , n7542 );
nand ( n11672 , n11671 , n116 );
nand ( n11673 , n11669 , n11670 , n11672 );
nand ( n11674 , n11665 , n11673 );
nand ( n11675 , n116 , n7371 );
not ( n11676 , n116 );
nand ( n11677 , n11676 , n7343 );
not ( n11678 , n11677 );
not ( n11679 , n7519 );
or ( n11680 , n11678 , n11679 );
nand ( n11681 , n11680 , n117 );
nand ( n11682 , n11674 , n11675 , n11681 );
and ( n11683 , n11664 , n11682 );
nor ( n11684 , n11663 , n11683 );
not ( n11685 , n7478 );
not ( n11686 , n11624 );
nand ( n11687 , n11685 , n11686 );
not ( n11688 , n117 );
nand ( n11689 , n11688 , n7557 );
nand ( n11690 , n11684 , n11687 , n7375 , n11689 );
and ( n11691 , n7325 , n11690 );
not ( n11692 , n7325 );
not ( n11693 , n118 );
not ( n11694 , n117 );
not ( n11695 , n116 );
not ( n11696 , n115 );
nand ( n11697 , n11696 , n7356 );
nor ( n11698 , n11695 , n11697 );
nand ( n11699 , n11694 , n11698 );
not ( n11700 , n117 );
not ( n11701 , n114 );
not ( n11702 , n7510 );
or ( n11703 , n11701 , n11702 );
nand ( n11704 , n11703 , n11601 );
and ( n11705 , n11700 , n11704 );
not ( n11706 , n11700 );
and ( n11707 , n11706 , n7418 );
nor ( n11708 , n11705 , n11707 );
nand ( n11709 , n11699 , n11708 );
not ( n11710 , n11709 );
or ( n11711 , n11693 , n11710 );
buf ( n11712 , n7456 );
not ( n11713 , n11712 );
not ( n11714 , n7488 );
not ( n11715 , n11714 );
nand ( n11716 , n115 , n11715 );
not ( n11717 , n7344 );
not ( n11718 , n11717 );
not ( n11719 , n115 );
nor ( n11720 , n11718 , n11719 );
not ( n11721 , n11720 );
nand ( n11722 , n11713 , n11716 , n11721 );
nand ( n11723 , n11685 , n11722 );
nand ( n11724 , n11711 , n11723 );
not ( n11725 , n11724 );
not ( n11726 , n7350 );
not ( n11727 , n7613 );
nor ( n11728 , n11726 , n11727 );
nand ( n11729 , n117 , n7426 );
nor ( n11730 , n116 , n7360 );
and ( n11731 , n117 , n11730 );
not ( n11732 , n117 );
not ( n11733 , n116 );
nand ( n11734 , n11733 , n7418 );
not ( n11735 , n11734 );
and ( n11736 , n11732 , n11735 );
or ( n11737 , n11731 , n11736 );
not ( n11738 , n7335 );
not ( n11739 , n117 );
nand ( n11740 , n11738 , n11739 );
and ( n11741 , n7359 , n7552 );
not ( n11742 , n116 );
nor ( n11743 , n115 , n11659 );
nand ( n11744 , n11742 , n11743 );
and ( n11745 , n11744 , n7598 );
nand ( n11746 , n11740 , n11741 , n7544 , n11745 );
or ( n11747 , n11737 , n11746 );
not ( n11748 , n118 );
nand ( n11749 , n11747 , n11748 );
nand ( n11750 , n11725 , n11728 , n11729 , n11749 );
and ( n11751 , n11692 , n11750 );
nor ( n11752 , n11691 , n11751 );
and ( n11753 , n11636 , n11657 , n11752 );
not ( n11754 , n11753 );
nand ( n11755 , n8154 , n8245 );
not ( n11756 , n11755 );
not ( n11757 , n11756 );
or ( n11758 , n11754 , n11757 );
or ( n11759 , n11753 , n11756 );
nand ( n11760 , n11758 , n11759 );
not ( n11761 , n117 );
not ( n11762 , n116 );
not ( n11763 , n115 );
nand ( n11764 , n11763 , n7389 );
nor ( n11765 , n11762 , n11764 );
nand ( n11766 , n11761 , n11765 );
not ( n11767 , n11744 );
not ( n11768 , n116 );
nand ( n11769 , n11768 , n11712 );
not ( n11770 , n11769 );
or ( n11771 , n11767 , n11770 );
not ( n11772 , n117 );
nand ( n11773 , n11771 , n11772 );
and ( n11774 , n11766 , n11612 , n11773 );
nor ( n11775 , n11774 , n118 );
not ( n11776 , n11775 );
not ( n11777 , n118 );
and ( n11778 , n117 , n11777 );
not ( n11779 , n11778 );
not ( n11780 , n7432 );
not ( n11781 , n116 );
nand ( n11782 , n11780 , n11781 );
not ( n11783 , n7406 );
nand ( n11784 , n11783 , n116 );
nand ( n11785 , n11782 , n11784 , n7442 );
not ( n11786 , n11785 );
or ( n11787 , n11779 , n11786 );
nand ( n11788 , n7348 , n7356 );
not ( n11789 , n11788 );
not ( n11790 , n7410 );
or ( n11791 , n11789 , n11790 );
not ( n11792 , n117 );
nand ( n11793 , n11791 , n11792 );
nand ( n11794 , n11787 , n11793 );
not ( n11795 , n11794 );
not ( n11796 , n117 );
not ( n11797 , n116 );
not ( n11798 , n11797 );
not ( n11799 , n7543 );
nand ( n11800 , n11799 , n7556 , n7567 );
not ( n11801 , n11800 );
or ( n11802 , n11798 , n11801 );
nor ( n11803 , n7608 , n11643 );
nand ( n11804 , n11802 , n11803 );
not ( n11805 , n11804 );
or ( n11806 , n11796 , n11805 );
not ( n11807 , n114 );
nand ( n11808 , n11807 , n115 , n112 );
not ( n11809 , n11808 );
not ( n11810 , n11809 );
nand ( n11811 , n11631 , n11810 , n11655 , n7457 );
nand ( n11812 , n7485 , n11811 );
nand ( n11813 , n11806 , n11812 );
nand ( n11814 , n118 , n11813 );
nand ( n11815 , n11776 , n11795 , n11814 );
not ( n11816 , n11815 );
not ( n11817 , n11685 );
not ( n11818 , n7402 );
or ( n11819 , n11817 , n11818 );
not ( n11820 , n117 );
and ( n11821 , n11820 , n7473 );
not ( n11822 , n11820 );
not ( n11823 , n116 );
nand ( n11824 , n11823 , n7543 );
not ( n11825 , n116 );
nand ( n11826 , n11825 , n11809 );
nand ( n11827 , n11824 , n7579 , n11826 );
and ( n11828 , n11822 , n11827 );
nor ( n11829 , n11821 , n11828 );
nand ( n11830 , n11819 , n11829 );
not ( n11831 , n11830 );
not ( n11832 , n7442 );
not ( n11833 , n7501 );
not ( n11834 , n11833 );
nand ( n11835 , n11597 , n11834 );
not ( n11836 , n11835 );
or ( n11837 , n11832 , n11836 );
nand ( n11838 , n11837 , n118 );
not ( n11839 , n118 );
nor ( n11840 , n7473 , n7604 );
not ( n11841 , n117 );
not ( n11842 , n7357 );
nand ( n11843 , n11841 , n11842 );
not ( n11844 , n117 );
nand ( n11845 , n11844 , n11730 );
and ( n11846 , n11843 , n11845 );
nor ( n11847 , n116 , n11764 );
and ( n11848 , n117 , n11847 );
not ( n11849 , n117 );
nand ( n11850 , n11601 , n7432 , n7362 );
and ( n11851 , n11849 , n11850 );
nor ( n11852 , n11848 , n11851 );
nand ( n11853 , n11840 , n11846 , n11852 );
nand ( n11854 , n11839 , n11853 );
not ( n11855 , n114 );
not ( n11856 , n11855 );
not ( n11857 , n115 );
and ( n11858 , n11856 , n11857 );
not ( n11859 , n7360 );
and ( n11860 , n116 , n11859 );
nor ( n11861 , n11858 , n11860 );
nand ( n11862 , n11861 , n11677 , n11601 );
and ( n11863 , n11618 , n11862 );
nor ( n11864 , n11659 , n7509 );
nor ( n11865 , n11863 , n11864 );
nand ( n11866 , n11831 , n11838 , n11854 , n11865 );
nand ( n11867 , n119 , n11866 );
not ( n11868 , n11647 );
not ( n11869 , n11720 );
not ( n11870 , n11869 );
or ( n11871 , n11868 , n11870 );
nand ( n11872 , n11871 , n11685 );
nor ( n11873 , n7478 , n7390 );
or ( n11874 , n7415 , n11873 );
not ( n11875 , n118 );
nand ( n11876 , n11874 , n11875 );
and ( n11877 , n11773 , n11872 , n11876 );
not ( n11878 , n7336 );
not ( n11879 , n117 );
not ( n11880 , n11855 );
not ( n11881 , n7468 );
or ( n11882 , n11880 , n11881 );
nand ( n11883 , n116 , n7488 );
nand ( n11884 , n11882 , n11883 );
and ( n11885 , n11879 , n11884 );
nor ( n11886 , n7387 , n7585 );
nor ( n11887 , n11885 , n11886 );
nand ( n11888 , n11878 , n11887 , n11675 );
and ( n11889 , n118 , n11888 );
not ( n11890 , n118 );
not ( n11891 , n117 );
not ( n11892 , n11891 );
not ( n11893 , n11621 );
or ( n11894 , n11892 , n11893 );
not ( n11895 , n116 );
nor ( n11896 , n11895 , n7532 );
not ( n11897 , n11896 );
nand ( n11898 , n11894 , n11897 );
and ( n11899 , n11890 , n11898 );
nor ( n11900 , n11889 , n11899 );
not ( n11901 , n115 );
and ( n11902 , n11901 , n7407 );
nand ( n11903 , n11685 , n11902 );
not ( n11904 , n7409 );
not ( n11905 , n11904 );
not ( n11906 , n7581 );
or ( n11907 , n11905 , n11906 );
not ( n11908 , n117 );
nand ( n11909 , n11907 , n11908 );
nand ( n11910 , n11877 , n11900 , n11903 , n11909 );
nand ( n11911 , n11910 , n7325 );
nand ( n11912 , n11816 , n11867 , n11911 );
buf ( n11913 , n11912 );
not ( n11914 , n6796 );
not ( n11915 , n6676 );
and ( n11916 , n11914 , n11915 );
not ( n11917 , n141 );
nor ( n11918 , n11916 , n11917 , n6640 );
nor ( n11919 , n11239 , n11918 );
or ( n11920 , n142 , n11438 );
not ( n11921 , n6731 );
not ( n11922 , n11921 );
nand ( n11923 , n11920 , n11922 );
nand ( n11924 , n11498 , n11923 );
not ( n11925 , n144 );
not ( n11926 , n11248 );
nand ( n11927 , n142 , n11926 );
nand ( n11928 , n11246 , n6676 );
and ( n11929 , n11927 , n6785 , n11928 );
not ( n11930 , n11247 );
not ( n11931 , n11930 );
nand ( n11932 , n142 , n11931 );
nand ( n11933 , n11932 , n11318 , n6690 );
nand ( n11934 , n141 , n11933 );
not ( n11935 , n141 );
nand ( n11936 , n6602 , n11288 , n6674 );
nand ( n11937 , n11935 , n11936 );
nand ( n11938 , n11929 , n11934 , n11937 );
nand ( n11939 , n11925 , n11938 );
and ( n11940 , n11919 , n11924 , n11939 );
not ( n11941 , n141 );
not ( n11942 , n11941 );
nand ( n11943 , n6562 , n6575 );
nand ( n11944 , n11943 , n11489 , n11393 );
not ( n11945 , n11944 );
or ( n11946 , n11942 , n11945 );
not ( n11947 , n6688 );
not ( n11948 , n11947 );
nand ( n11949 , n11946 , n11948 );
and ( n11950 , n11949 , n144 );
not ( n11951 , n11498 );
nor ( n11952 , n11951 , n6659 );
nor ( n11953 , n11950 , n11952 );
not ( n11954 , n11922 );
nand ( n11955 , n11264 , n11954 );
not ( n11956 , n6567 );
not ( n11957 , n11956 );
not ( n11958 , n141 );
not ( n11959 , n6604 );
nand ( n11960 , n11958 , n11959 );
nand ( n11961 , n11955 , n11957 , n11960 );
not ( n11962 , n141 );
not ( n11963 , n6556 );
nand ( n11964 , n142 , n11963 );
nand ( n11965 , n142 , n6771 );
nand ( n11966 , n11361 , n11964 , n11965 );
nand ( n11967 , n11962 , n11966 );
not ( n11968 , n11507 );
not ( n11969 , n6647 );
or ( n11970 , n11968 , n11969 );
nand ( n11971 , n11970 , n141 );
and ( n11972 , n11967 , n11453 , n11971 );
and ( n11973 , n144 , n11972 );
not ( n11974 , n144 );
and ( n11975 , n6544 , n11334 );
not ( n11976 , n11318 );
nor ( n11977 , n11975 , n11976 );
and ( n11978 , n11974 , n11977 );
nor ( n11979 , n11973 , n11978 );
or ( n11980 , n11961 , n11979 );
nand ( n11981 , n11980 , n6808 );
not ( n11982 , n144 );
not ( n11983 , n11982 );
not ( n11984 , n141 );
nand ( n11985 , n11984 , n11921 );
not ( n11986 , n6559 );
nor ( n11987 , n11986 , n6616 );
nand ( n11988 , n11423 , n6695 );
not ( n11989 , n141 );
and ( n11990 , n11989 , n11343 );
not ( n11991 , n11321 );
and ( n11992 , n11991 , n141 );
nor ( n11993 , n11990 , n11992 );
nor ( n11994 , n11988 , n11993 );
nand ( n11995 , n6801 , n11985 , n11987 , n11994 );
not ( n11996 , n11995 );
or ( n11997 , n11983 , n11996 );
and ( n11998 , n6795 , n6701 );
nor ( n11999 , n11998 , n6678 );
not ( n12000 , n141 );
or ( n12001 , n12000 , n6764 );
not ( n12002 , n141 );
or ( n12003 , n6669 , n6574 );
nand ( n12004 , n12003 , n11248 );
nand ( n12005 , n12002 , n12004 );
not ( n12006 , n141 );
not ( n12007 , n138 );
nor ( n12008 , n12007 , n11242 );
nand ( n12009 , n12006 , n6622 , n12008 );
nand ( n12010 , n12001 , n12005 , n12009 );
nand ( n12011 , n144 , n12010 );
and ( n12012 , n11999 , n6698 , n12011 );
nand ( n12013 , n11997 , n12012 );
not ( n12014 , n11301 );
and ( n12015 , n11430 , n12014 , n11258 );
nor ( n12016 , n12015 , n6661 );
or ( n12017 , n12013 , n12016 );
nand ( n12018 , n12017 , n137 );
nand ( n12019 , n11940 , n11953 , n11981 , n12018 );
not ( n12020 , n12019 );
and ( n12021 , n11913 , n12020 );
not ( n12022 , n11913 );
buf ( n12023 , n12019 );
and ( n12024 , n12022 , n12023 );
nor ( n12025 , n12021 , n12024 );
and ( n12026 , n11760 , n12025 );
not ( n12027 , n11760 );
not ( n12028 , n12025 );
and ( n12029 , n12027 , n12028 );
nor ( n12030 , n12026 , n12029 );
not ( n12031 , n12030 );
nand ( n12032 , n11588 , n12031 );
nand ( n12033 , n11587 , n12030 );
nand ( n12034 , n12032 , n2352 , n12033 );
nand ( n12035 , n11231 , n12034 );
xnor ( n12036 , n382 , n383 );
or ( n12037 , n2352 , n12036 );
not ( n12038 , n9996 );
and ( n12039 , n382 , n12038 );
not ( n12040 , n382 );
and ( n12041 , n12040 , n9996 );
nor ( n12042 , n12039 , n12041 );
not ( n12043 , n12042 );
not ( n12044 , n10493 );
not ( n12045 , n12044 );
not ( n12046 , n5197 );
and ( n12047 , n12045 , n12046 );
and ( n12048 , n10923 , n5205 );
nor ( n12049 , n12047 , n12048 );
not ( n12050 , n12049 );
and ( n12051 , n12043 , n12050 );
and ( n12052 , n12042 , n12049 );
nor ( n12053 , n12051 , n12052 );
not ( n12054 , n12053 );
not ( n12055 , n10796 );
not ( n12056 , n177 );
not ( n12057 , n4898 );
not ( n12058 , n4836 );
or ( n12059 , n12057 , n12058 );
nand ( n12060 , n12059 , n5017 );
and ( n12061 , n12056 , n12060 );
not ( n12062 , n12056 );
not ( n12063 , n176 );
nand ( n12064 , n172 , n4700 );
not ( n12065 , n4593 );
nand ( n12066 , n172 , n12065 );
nand ( n12067 , n5128 , n12064 , n12066 );
nand ( n12068 , n12063 , n12067 );
not ( n12069 , n4889 );
not ( n12070 , n4750 );
or ( n12071 , n12069 , n12070 );
nand ( n12072 , n12071 , n176 );
nand ( n12073 , n12068 , n4957 , n12072 );
and ( n12074 , n12062 , n12073 );
nor ( n12075 , n12061 , n12074 );
nand ( n12076 , n4982 , n4665 );
not ( n12077 , n176 );
not ( n12078 , n172 );
nor ( n12079 , n12078 , n4732 );
nand ( n12080 , n12077 , n12079 );
nand ( n12081 , n12075 , n12076 , n4706 , n12080 );
and ( n12082 , n4765 , n12081 );
not ( n12083 , n4869 );
nand ( n12084 , n172 , n12083 );
nand ( n12085 , n4906 , n4587 );
and ( n12086 , n12084 , n4668 , n12085 );
not ( n12087 , n176 );
not ( n12088 , n4733 );
nand ( n12089 , n5070 , n12088 , n4579 );
and ( n12090 , n12087 , n12089 );
not ( n12091 , n12087 );
not ( n12092 , n4868 );
not ( n12093 , n12092 );
nand ( n12094 , n172 , n12093 );
nand ( n12095 , n12094 , n5017 , n4608 );
and ( n12096 , n12091 , n12095 );
nor ( n12097 , n12090 , n12096 );
and ( n12098 , n12086 , n12097 );
nor ( n12099 , n12098 , n177 );
nor ( n12100 , n12082 , n12099 );
not ( n12101 , n12100 );
and ( n12102 , n4629 , n4588 );
nand ( n12103 , n176 , n4809 );
not ( n12104 , n177 );
not ( n12105 , n4618 );
not ( n12106 , n12105 );
not ( n12107 , n4813 );
nand ( n12108 , n4904 , n12107 );
and ( n12109 , n12108 , n4714 , n4929 );
not ( n12110 , n176 );
nor ( n12111 , n12110 , n4864 );
nor ( n12112 , n4702 , n12111 );
nor ( n12113 , n176 , n4664 );
nor ( n12114 , n4772 , n12113 );
nand ( n12115 , n12106 , n12109 , n12112 , n12114 );
nand ( n12116 , n12104 , n12115 );
nand ( n12117 , n12102 , n12103 , n12116 );
not ( n12118 , n177 );
not ( n12119 , n176 );
nand ( n12120 , n12119 , n5063 );
and ( n12121 , n176 , n4814 );
not ( n12122 , n176 );
not ( n12123 , n174 );
or ( n12124 , n12123 , n4739 );
nand ( n12125 , n12124 , n4869 );
and ( n12126 , n12122 , n12125 );
nor ( n12127 , n12121 , n12126 );
nand ( n12128 , n12120 , n12127 );
not ( n12129 , n12128 );
or ( n12130 , n12118 , n12129 );
not ( n12131 , n5084 );
nand ( n12132 , n173 , n5072 );
nand ( n12133 , n4979 , n12131 , n12132 );
nand ( n12134 , n4982 , n12133 );
nand ( n12135 , n12130 , n12134 );
nor ( n12136 , n12117 , n12135 );
or ( n12137 , n12136 , n4765 );
or ( n12138 , n172 , n4944 );
nand ( n12139 , n12138 , n4664 );
and ( n12140 , n4879 , n12139 );
and ( n12141 , n4646 , n5034 );
not ( n12142 , n176 );
nor ( n12143 , n12141 , n12142 , n4581 );
nor ( n12144 , n12140 , n12143 );
and ( n12145 , n172 , n177 );
nand ( n12146 , n176 , n12145 , n4842 );
and ( n12147 , n5183 , n12146 );
or ( n12148 , n176 , n5153 );
nand ( n12149 , n4899 , n5066 );
not ( n12150 , n12149 );
not ( n12151 , n5027 );
or ( n12152 , n12150 , n12151 );
not ( n12153 , n176 );
nand ( n12154 , n12152 , n12153 );
nand ( n12155 , n12148 , n12154 , n4601 );
nand ( n12156 , n177 , n12155 );
and ( n12157 , n12144 , n12147 , n12156 );
nand ( n12158 , n12137 , n12157 );
nor ( n12159 , n12101 , n12158 );
not ( n12160 , n12159 );
not ( n12161 , n5040 );
not ( n12162 , n12161 );
and ( n12163 , n12160 , n12162 );
not ( n12164 , n5040 );
and ( n12165 , n12159 , n12164 );
nor ( n12166 , n12163 , n12165 );
not ( n12167 , n12166 );
not ( n12168 , n12167 );
and ( n12169 , n12055 , n12168 );
and ( n12170 , n12167 , n10796 );
nor ( n12171 , n12169 , n12170 );
not ( n12172 , n12171 );
nand ( n12173 , n12054 , n12172 );
nand ( n12174 , n12053 , n12171 );
nand ( n12175 , n12173 , n2352 , n12174 );
nand ( n12176 , n12037 , n12175 );
xnor ( n12177 , n384 , n385 );
or ( n12178 , n2352 , n12177 );
not ( n12179 , n9836 );
not ( n12180 , n9870 );
nand ( n12181 , n12179 , n12180 );
and ( n12182 , n4144 , n12181 );
not ( n12183 , n4144 );
nand ( n12184 , n9948 , n9895 , n9901 , n9925 );
and ( n12185 , n12183 , n12184 );
nor ( n12186 , n12182 , n12185 );
nand ( n12187 , n12186 , n9994 , n9815 , n9989 );
and ( n12188 , n384 , n12187 );
not ( n12189 , n384 );
not ( n12190 , n12187 );
and ( n12191 , n12189 , n12190 );
nor ( n12192 , n12188 , n12191 );
not ( n12193 , n12192 );
not ( n12194 , n10661 );
and ( n12195 , n12193 , n12194 );
and ( n12196 , n12192 , n10661 );
nor ( n12197 , n12195 , n12196 );
not ( n12198 , n12197 );
not ( n12199 , n10315 );
not ( n12200 , n4433 );
not ( n12201 , n12200 );
not ( n12202 , n4415 );
not ( n12203 , n12202 );
and ( n12204 , n12201 , n12203 );
not ( n12205 , n149 );
not ( n12206 , n4393 );
nor ( n12207 , n12204 , n12205 , n12206 );
nor ( n12208 , n12199 , n12207 );
or ( n12209 , n150 , n10501 );
nand ( n12210 , n12209 , n4442 );
nand ( n12211 , n10610 , n12210 );
not ( n12212 , n149 );
not ( n12213 , n12212 );
nand ( n12214 , n10370 , n4336 );
nand ( n12215 , n12214 , n10353 , n10450 );
not ( n12216 , n12215 );
or ( n12217 , n12213 , n12216 );
nand ( n12218 , n12217 , n4546 );
nand ( n12219 , n152 , n12218 );
and ( n12220 , n12208 , n12211 , n12219 );
not ( n12221 , n4457 );
nand ( n12222 , n12221 , n10610 );
or ( n12223 , n4463 , n4442 );
not ( n12224 , n4488 );
not ( n12225 , n12224 );
not ( n12226 , n4380 );
not ( n12227 , n149 );
nand ( n12228 , n12226 , n12227 );
nand ( n12229 , n12223 , n12225 , n12228 );
and ( n12230 , n10469 , n10624 );
not ( n12231 , n10411 );
nor ( n12232 , n12230 , n12231 );
and ( n12233 , n4532 , n12232 );
not ( n12234 , n4532 );
not ( n12235 , n149 );
not ( n12236 , n150 );
nor ( n12237 , n12236 , n4320 );
not ( n12238 , n12237 );
nand ( n12239 , n150 , n4498 );
nand ( n12240 , n10453 , n12238 , n12239 );
nand ( n12241 , n12235 , n12240 );
not ( n12242 , n10620 );
not ( n12243 , n4400 );
or ( n12244 , n12242 , n12243 );
nand ( n12245 , n12244 , n149 );
and ( n12246 , n12241 , n10539 , n12245 );
and ( n12247 , n12234 , n12246 );
nor ( n12248 , n12233 , n12247 );
or ( n12249 , n12229 , n12248 );
nand ( n12250 , n12249 , n4405 );
not ( n12251 , n153 );
and ( n12252 , n10521 , n4344 , n10339 );
nor ( n12253 , n12252 , n4461 );
not ( n12254 , n12253 );
nand ( n12255 , n4480 , n10417 );
nand ( n12256 , n12255 , n4509 );
not ( n12257 , n152 );
nand ( n12258 , n146 , n4335 );
not ( n12259 , n12258 );
not ( n12260 , n10320 );
or ( n12261 , n12259 , n12260 );
not ( n12262 , n149 );
nand ( n12263 , n12261 , n12262 );
nand ( n12264 , n149 , n4514 );
nand ( n12265 , n10331 , n10585 );
nand ( n12266 , n12263 , n12264 , n12265 );
not ( n12267 , n12266 );
or ( n12268 , n12257 , n12267 );
nand ( n12269 , n12268 , n4566 );
nor ( n12270 , n12256 , n12269 );
not ( n12271 , n4559 );
nor ( n12272 , n149 , n4442 );
nor ( n12273 , n12271 , n12272 );
not ( n12274 , n149 );
not ( n12275 , n10401 );
or ( n12276 , n12274 , n12275 );
nand ( n12277 , n12276 , n4322 );
nand ( n12278 , n10317 , n4514 );
nand ( n12279 , n12278 , n4370 , n10515 );
nor ( n12280 , n12277 , n12279 );
nand ( n12281 , n12273 , n4474 , n12280 );
nand ( n12282 , n4532 , n12281 );
nand ( n12283 , n12254 , n12270 , n12282 );
not ( n12284 , n12283 );
or ( n12285 , n12251 , n12284 );
not ( n12286 , n10320 );
nand ( n12287 , n150 , n12286 );
nand ( n12288 , n10317 , n12202 );
and ( n12289 , n12287 , n4422 , n12288 );
nand ( n12290 , n150 , n10319 );
nand ( n12291 , n12290 , n10411 , n4548 );
nand ( n12292 , n149 , n12291 );
not ( n12293 , n149 );
nand ( n12294 , n4378 , n10372 , n4536 );
nand ( n12295 , n12293 , n12294 );
nand ( n12296 , n12289 , n12292 , n12295 );
nand ( n12297 , n4532 , n12296 );
nand ( n12298 , n12285 , n12297 );
not ( n12299 , n12298 );
nand ( n12300 , n12220 , n12222 , n12250 , n12299 );
not ( n12301 , n12300 );
not ( n12302 , n12166 );
not ( n12303 , n12302 );
or ( n12304 , n12301 , n12303 );
not ( n12305 , n12300 );
nand ( n12306 , n12305 , n12166 );
nand ( n12307 , n12304 , n12306 );
not ( n12308 , n10800 );
and ( n12309 , n12307 , n12308 );
not ( n12310 , n12307 );
and ( n12311 , n12310 , n10800 );
nor ( n12312 , n12309 , n12311 );
not ( n12313 , n12312 );
nand ( n12314 , n12198 , n12313 );
nand ( n12315 , n12197 , n12312 );
nand ( n12316 , n12314 , n2352 , n12315 );
nand ( n12317 , n12178 , n12316 );
not ( n12318 , n342 );
not ( n12319 , n194 );
and ( n12320 , n191 , n2955 );
not ( n12321 , n12320 );
nand ( n12322 , n193 , n2444 );
nand ( n12323 , n12321 , n12322 );
not ( n12324 , n193 );
not ( n12325 , n12324 );
not ( n12326 , n191 );
nand ( n12327 , n12326 , n2452 );
nand ( n12328 , n2589 , n12327 , n2787 );
not ( n12329 , n12328 );
or ( n12330 , n12325 , n12329 );
nand ( n12331 , n2561 , n2912 );
nand ( n12332 , n12330 , n12331 );
nor ( n12333 , n12323 , n12332 );
or ( n12334 , n12319 , n12333 );
nor ( n12335 , n2586 , n2817 );
not ( n12336 , n194 );
not ( n12337 , n12336 );
and ( n12338 , n2585 , n2444 );
and ( n12339 , n193 , n2510 );
nor ( n12340 , n12338 , n12339 );
not ( n12341 , n191 );
nor ( n12342 , n12341 , n2475 );
not ( n12343 , n12342 );
nand ( n12344 , n12340 , n2915 , n12343 );
not ( n12345 , n12344 );
or ( n12346 , n12337 , n12345 );
nand ( n12347 , n12346 , n2756 );
nor ( n12348 , n12335 , n12347 );
not ( n12349 , n191 );
not ( n12350 , n12349 );
not ( n12351 , n2978 );
or ( n12352 , n12350 , n12351 );
nand ( n12353 , n12352 , n2851 );
nand ( n12354 , n193 , n12353 );
nand ( n12355 , n12334 , n12348 , n12354 );
nand ( n12356 , n12355 , n2364 );
not ( n12357 , n193 );
not ( n12358 , n2567 );
nand ( n12359 , n2635 , n12358 , n2709 );
and ( n12360 , n12357 , n12359 );
or ( n12361 , n188 , n2781 );
not ( n12362 , n2711 );
nand ( n12363 , n12361 , n12362 );
and ( n12364 , n193 , n12363 );
not ( n12365 , n2376 );
not ( n12366 , n2771 );
not ( n12367 , n12366 );
or ( n12368 , n12365 , n12367 );
nand ( n12369 , n12368 , n2571 );
and ( n12370 , n193 , n12369 );
nor ( n12371 , n12360 , n12364 , n12370 );
not ( n12372 , n12371 );
not ( n12373 , n194 );
nand ( n12374 , n191 , n2872 );
not ( n12375 , n12374 );
nor ( n12376 , n12375 , n2666 );
not ( n12377 , n193 );
nand ( n12378 , n12377 , n2526 );
nand ( n12379 , n193 , n8956 );
nand ( n12380 , n12376 , n12378 , n9030 , n12379 );
and ( n12381 , n12373 , n12380 );
not ( n12382 , n12373 );
not ( n12383 , n193 );
not ( n12384 , n2634 );
nand ( n12385 , n12384 , n2811 );
and ( n12386 , n12383 , n12385 );
nand ( n12387 , n193 , n2804 );
not ( n12388 , n12387 );
nor ( n12389 , n12386 , n12388 );
nand ( n12390 , n12389 , n2716 , n2534 );
and ( n12391 , n12382 , n12390 );
nor ( n12392 , n12381 , n12391 );
not ( n12393 , n12392 );
or ( n12394 , n12372 , n12393 );
nand ( n12395 , n12394 , n195 );
not ( n12396 , n193 );
nand ( n12397 , n191 , n2380 );
not ( n12398 , n12397 );
and ( n12399 , n12396 , n12398 );
and ( n12400 , n2472 , n2512 );
nor ( n12401 , n12399 , n12400 );
nand ( n12402 , n193 , n2974 );
not ( n12403 , n193 );
nor ( n12404 , n12403 , n2828 );
not ( n12405 , n12404 );
and ( n12406 , n12402 , n12405 , n2767 );
not ( n12407 , n193 );
nand ( n12408 , n2409 , n2670 );
nand ( n12409 , n191 , n12408 );
nand ( n12410 , n2709 , n9056 , n12409 );
nand ( n12411 , n12407 , n12410 );
nand ( n12412 , n12406 , n2845 , n12411 );
nand ( n12413 , n194 , n12412 );
not ( n12414 , n194 );
and ( n12415 , n2887 , n2756 );
not ( n12416 , n193 );
not ( n12417 , n191 );
nand ( n12418 , n12417 , n2901 );
nand ( n12419 , n12418 , n2436 , n2573 );
nand ( n12420 , n12416 , n12419 );
not ( n12421 , n2483 );
nand ( n12422 , n12421 , n2944 );
not ( n12423 , n2575 );
nand ( n12424 , n2382 , n12423 );
not ( n12425 , n12424 );
not ( n12426 , n2547 );
or ( n12427 , n12425 , n12426 );
nand ( n12428 , n12427 , n2633 );
or ( n12429 , n12422 , n12428 );
nand ( n12430 , n12429 , n193 );
nand ( n12431 , n12415 , n12420 , n12430 );
nand ( n12432 , n12414 , n12431 );
and ( n12433 , n12401 , n12413 , n12432 );
and ( n12434 , n12356 , n12395 , n12433 );
not ( n12435 , n12434 );
not ( n12436 , n12435 );
or ( n12437 , n12318 , n12436 );
buf ( n12438 , n12434 );
not ( n12439 , n12438 );
or ( n12440 , n342 , n12439 );
nand ( n12441 , n12437 , n12440 );
not ( n12442 , n12441 );
not ( n12443 , n11211 );
not ( n12444 , n12443 );
or ( n12445 , n12442 , n12444 );
or ( n12446 , n12441 , n12443 );
nand ( n12447 , n12445 , n12446 );
not ( n12448 , n12447 );
buf ( n12449 , n9512 );
not ( n12450 , n12449 );
not ( n12451 , n211 );
not ( n12452 , n209 );
or ( n12453 , n12452 , n3679 );
nand ( n12454 , n12453 , n8760 );
and ( n12455 , n12451 , n12454 );
and ( n12456 , n8636 , n3514 );
nor ( n12457 , n12455 , n12456 );
not ( n12458 , n211 );
not ( n12459 , n8511 );
not ( n12460 , n209 );
nand ( n12461 , n12459 , n12460 );
nand ( n12462 , n3641 , n9448 , n8703 );
nand ( n12463 , n9303 , n12462 );
nand ( n12464 , n12461 , n8474 , n12463 );
not ( n12465 , n12464 );
or ( n12466 , n12458 , n12465 );
or ( n12467 , n3708 , n8440 );
nand ( n12468 , n12467 , n8457 );
nand ( n12469 , n3717 , n12468 );
nand ( n12470 , n12466 , n12469 );
not ( n12471 , n12470 );
and ( n12472 , n12457 , n12471 );
or ( n12473 , n8617 , n8463 );
not ( n12474 , n3469 );
or ( n12475 , n3579 , n8667 );
nand ( n12476 , n209 , n3588 );
nand ( n12477 , n12475 , n12476 );
not ( n12478 , n12477 );
not ( n12479 , n209 );
not ( n12480 , n12479 );
nand ( n12481 , n8556 , n3703 );
not ( n12482 , n12481 );
or ( n12483 , n12480 , n12482 );
not ( n12484 , n210 );
nand ( n12485 , n12484 , n8605 );
nand ( n12486 , n12483 , n12485 );
not ( n12487 , n12486 );
not ( n12488 , n211 );
nand ( n12489 , n209 , n208 , n3582 );
not ( n12490 , n3499 );
not ( n12491 , n3668 );
or ( n12492 , n12490 , n12491 );
nand ( n12493 , n12492 , n8561 );
nand ( n12494 , n12489 , n12493 );
nor ( n12495 , n9451 , n12494 );
not ( n12496 , n8568 );
not ( n12497 , n12496 );
nand ( n12498 , n12497 , n8604 );
nand ( n12499 , n12495 , n8581 , n12498 );
and ( n12500 , n12488 , n12499 );
not ( n12501 , n12488 );
nor ( n12502 , n8443 , n3521 );
not ( n12503 , n209 );
nand ( n12504 , n12503 , n3555 );
not ( n12505 , n8667 );
not ( n12506 , n8652 );
or ( n12507 , n12505 , n12506 );
nand ( n12508 , n12507 , n209 );
nand ( n12509 , n12502 , n12504 , n8503 , n12508 );
and ( n12510 , n12501 , n12509 );
nor ( n12511 , n12500 , n12510 );
nand ( n12512 , n12478 , n12487 , n12511 );
not ( n12513 , n12512 );
or ( n12514 , n12474 , n12513 );
nand ( n12515 , n12514 , n3606 );
not ( n12516 , n211 );
not ( n12517 , n3529 );
not ( n12518 , n3674 );
or ( n12519 , n12517 , n12518 );
not ( n12520 , n209 );
nand ( n12521 , n12519 , n12520 );
nand ( n12522 , n12516 , n12521 );
and ( n12523 , n3585 , n9306 );
nand ( n12524 , n209 , n8736 );
and ( n12525 , n12524 , n8554 , n9328 );
nand ( n12526 , n3687 , n12523 , n12525 );
or ( n12527 , n12522 , n12526 );
and ( n12528 , n8569 , n9455 );
and ( n12529 , n9428 , n8456 );
not ( n12530 , n209 );
not ( n12531 , n210 );
not ( n12532 , n207 );
nor ( n12533 , n12532 , n205 );
nand ( n12534 , n12531 , n12533 );
nand ( n12535 , n12534 , n8565 , n8558 );
not ( n12536 , n12535 );
or ( n12537 , n12530 , n12536 );
nand ( n12538 , n12537 , n211 );
not ( n12539 , n12538 );
nand ( n12540 , n12528 , n12529 , n3739 , n12539 );
nand ( n12541 , n12527 , n12540 );
not ( n12542 , n208 );
or ( n12543 , n8630 , n12542 );
nand ( n12544 , n12543 , n3546 );
nand ( n12545 , n209 , n12544 );
not ( n12546 , n209 );
not ( n12547 , n12546 );
not ( n12548 , n9451 );
nand ( n12549 , n12548 , n9253 , n3594 );
not ( n12550 , n12549 );
or ( n12551 , n12547 , n12550 );
nand ( n12552 , n12551 , n8759 );
not ( n12553 , n12552 );
nand ( n12554 , n12541 , n12545 , n12553 );
nand ( n12555 , n212 , n12554 );
not ( n12556 , n12555 );
nor ( n12557 , n12515 , n12556 );
and ( n12558 , n12472 , n12473 , n3744 , n12557 );
not ( n12559 , n12558 );
or ( n12560 , n12450 , n12559 );
not ( n12561 , n9513 );
nand ( n12562 , n3469 , n12512 );
and ( n12563 , n3744 , n12555 , n3606 , n12562 );
and ( n12564 , n12472 , n12473 , n12563 );
or ( n12565 , n12561 , n12564 );
nand ( n12566 , n12560 , n12565 );
not ( n12567 , n12566 );
not ( n12568 , n3910 );
nand ( n12569 , n12568 , n202 );
and ( n12570 , n11063 , n12569 );
or ( n12571 , n203 , n12570 );
not ( n12572 , n9672 );
or ( n12573 , n3842 , n12572 );
nand ( n12574 , n12573 , n3995 );
and ( n12575 , n3825 , n12574 );
and ( n12576 , n202 , n3848 );
nor ( n12577 , n12575 , n12576 );
and ( n12578 , n3906 , n8300 );
nand ( n12579 , n3948 , n3900 );
nor ( n12580 , n12578 , n12579 );
nand ( n12581 , n12571 , n12577 , n12580 );
not ( n12582 , n12581 );
not ( n12583 , n202 );
not ( n12584 , n201 );
not ( n12585 , n3886 );
nand ( n12586 , n12584 , n12585 );
not ( n12587 , n3769 );
nand ( n12588 , n12586 , n12587 , n8364 );
not ( n12589 , n12588 );
or ( n12590 , n12583 , n12589 );
nand ( n12591 , n12590 , n9630 );
not ( n12592 , n12591 );
and ( n12593 , n3995 , n8312 );
and ( n12594 , n9578 , n9746 );
nand ( n12595 , n12592 , n203 , n12593 , n12594 );
not ( n12596 , n203 );
not ( n12597 , n202 );
nor ( n12598 , n12597 , n9536 );
nor ( n12599 , n8369 , n12598 );
not ( n12600 , n3801 );
not ( n12601 , n3915 );
or ( n12602 , n12600 , n12601 );
not ( n12603 , n202 );
nand ( n12604 , n12602 , n12603 );
nand ( n12605 , n12599 , n12604 );
not ( n12606 , n12605 );
and ( n12607 , n9662 , n3865 );
nor ( n12608 , n3873 , n9677 );
nand ( n12609 , n12596 , n12606 , n12607 , n12608 );
nand ( n12610 , n12595 , n12609 );
not ( n12611 , n202 );
not ( n12612 , n9580 );
nand ( n12613 , n12612 , n9721 , n3932 );
nand ( n12614 , n12611 , n12613 );
or ( n12615 , n3758 , n10977 );
nand ( n12616 , n12615 , n3756 );
nand ( n12617 , n202 , n12616 );
nand ( n12618 , n12610 , n12614 , n11088 , n12617 );
and ( n12619 , n204 , n12618 );
not ( n12620 , n204 );
not ( n12621 , n203 );
not ( n12622 , n12621 );
not ( n12623 , n8304 );
nand ( n12624 , n202 , n12623 );
not ( n12625 , n3811 );
not ( n12626 , n3911 );
or ( n12627 , n12625 , n12626 );
nand ( n12628 , n12627 , n3999 );
nand ( n12629 , n12624 , n12628 );
nor ( n12630 , n8336 , n12629 );
not ( n12631 , n3929 );
nand ( n12632 , n3904 , n12631 );
nand ( n12633 , n12630 , n12612 , n12632 );
not ( n12634 , n12633 );
or ( n12635 , n12622 , n12634 );
nand ( n12636 , n202 , n3925 );
nand ( n12637 , n12635 , n12636 );
not ( n12638 , n12637 );
not ( n12639 , n11043 );
nand ( n12640 , n3897 , n12639 );
not ( n12641 , n202 );
not ( n12642 , n12641 );
nand ( n12643 , n8348 , n3868 );
not ( n12644 , n12643 );
or ( n12645 , n12642 , n12644 );
not ( n12646 , n201 );
nand ( n12647 , n12646 , n3765 );
nand ( n12648 , n12645 , n12647 );
not ( n12649 , n12648 );
not ( n12650 , n201 );
not ( n12651 , n12650 );
not ( n12652 , n8411 );
or ( n12653 , n12651 , n12652 );
nand ( n12654 , n12653 , n11043 );
nand ( n12655 , n202 , n12654 );
not ( n12656 , n202 );
nand ( n12657 , n12656 , n3771 );
nand ( n12658 , n12655 , n3820 , n12657 );
nand ( n12659 , n8274 , n8403 );
or ( n12660 , n12658 , n12659 );
nand ( n12661 , n12660 , n203 );
nand ( n12662 , n12638 , n12640 , n12649 , n12661 );
and ( n12663 , n12620 , n12662 );
nor ( n12664 , n12619 , n12663 );
not ( n12665 , n9761 );
nand ( n12666 , n8279 , n9583 , n11030 );
nand ( n12667 , n12665 , n12666 );
not ( n12668 , n8396 );
not ( n12669 , n202 );
nand ( n12670 , n12668 , n12669 );
nand ( n12671 , n12667 , n8314 , n12670 );
nand ( n12672 , n203 , n12671 );
nand ( n12673 , n12582 , n12664 , n12672 );
not ( n12674 , n12673 );
and ( n12675 , n12674 , n9658 );
not ( n12676 , n12674 );
not ( n12677 , n9658 );
and ( n12678 , n12676 , n12677 );
nor ( n12679 , n12675 , n12678 );
not ( n12680 , n12679 );
or ( n12681 , n12567 , n12680 );
or ( n12682 , n12566 , n12679 );
nand ( n12683 , n12681 , n12682 );
not ( n12684 , n12683 );
nor ( n12685 , n12448 , n12684 );
or ( n12686 , n12447 , n12683 );
nand ( n12687 , n12686 , n2352 );
or ( n12688 , n12685 , n12687 );
xnor ( n12689 , n342 , n343 );
or ( n12690 , n2352 , n12689 );
nand ( n12691 , n12688 , n12690 );
not ( n12692 , n10664 );
not ( n12693 , n290 );
not ( n12694 , n161 );
not ( n12695 , n159 );
not ( n12696 , n9833 );
not ( n12697 , n12696 );
or ( n12698 , n12695 , n12697 );
nand ( n12699 , n12698 , n9901 );
not ( n12700 , n160 );
not ( n12701 , n4086 );
not ( n12702 , n154 );
nor ( n12703 , n12702 , n4106 );
nand ( n12704 , n158 , n12703 );
nand ( n12705 , n158 , n4091 );
nand ( n12706 , n12701 , n9945 , n12704 , n12705 );
not ( n12707 , n12706 );
or ( n12708 , n12700 , n12707 );
not ( n12709 , n159 );
not ( n12710 , n9916 );
nand ( n12711 , n12710 , n4283 , n4036 );
nand ( n12712 , n12709 , n12711 );
nand ( n12713 , n12708 , n12712 );
nor ( n12714 , n12699 , n12713 );
not ( n12715 , n10850 );
not ( n12716 , n9982 );
nor ( n12717 , n12715 , n12716 );
not ( n12718 , n156 );
or ( n12719 , n12718 , n4131 );
nand ( n12720 , n154 , n9821 );
not ( n12721 , n154 );
nand ( n12722 , n12721 , n9956 );
nand ( n12723 , n12719 , n12720 , n12722 );
nand ( n12724 , n10057 , n12723 );
and ( n12725 , n4174 , n4067 );
not ( n12726 , n159 );
nor ( n12727 , n12725 , n12726 );
not ( n12728 , n159 );
nand ( n12729 , n12728 , n4137 );
and ( n12730 , n4283 , n10005 );
nand ( n12731 , n12729 , n9833 , n12730 );
or ( n12732 , n12727 , n12731 );
nand ( n12733 , n12732 , n4054 );
nand ( n12734 , n12714 , n12717 , n12724 , n12733 );
not ( n12735 , n12734 );
or ( n12736 , n12694 , n12735 );
and ( n12737 , n4226 , n10019 );
not ( n12738 , n9904 );
not ( n12739 , n12738 );
not ( n12740 , n12739 );
nor ( n12741 , n12737 , n12740 );
not ( n12742 , n9833 );
nand ( n12743 , n4115 , n9930 );
not ( n12744 , n12743 );
or ( n12745 , n12742 , n12744 );
nand ( n12746 , n12745 , n159 );
not ( n12747 , n159 );
or ( n12748 , n158 , n4059 );
nand ( n12749 , n12748 , n4241 , n4259 );
nand ( n12750 , n12747 , n12749 );
nand ( n12751 , n12741 , n12746 , n12750 );
nand ( n12752 , n4054 , n12751 );
nand ( n12753 , n12736 , n12752 );
not ( n12754 , n159 );
and ( n12755 , n158 , n9823 );
nor ( n12756 , n12755 , n9903 );
not ( n12757 , n158 );
not ( n12758 , n9883 );
nor ( n12759 , n12757 , n12758 );
not ( n12760 , n12759 );
nor ( n12761 , n158 , n9811 );
not ( n12762 , n12761 );
nand ( n12763 , n12756 , n12760 , n12762 );
not ( n12764 , n12763 );
or ( n12765 , n12754 , n12764 );
not ( n12766 , n159 );
nand ( n12767 , n12766 , n4080 );
nand ( n12768 , n12765 , n12767 );
nor ( n12769 , n159 , n9992 );
not ( n12770 , n12769 );
not ( n12771 , n9866 );
nor ( n12772 , n12771 , n12720 );
nor ( n12773 , n10122 , n12772 );
not ( n12774 , n160 );
not ( n12775 , n158 );
not ( n12776 , n12775 );
not ( n12777 , n4099 );
or ( n12778 , n12776 , n12777 );
not ( n12779 , n12722 );
nand ( n12780 , n4226 , n12779 );
nand ( n12781 , n12778 , n12780 );
not ( n12782 , n12781 );
nor ( n12783 , n158 , n4122 );
nor ( n12784 , n4197 , n9891 );
nor ( n12785 , n12783 , n12784 );
nand ( n12786 , n12774 , n12782 , n12785 );
not ( n12787 , n159 );
not ( n12788 , n12787 );
not ( n12789 , n158 );
not ( n12790 , n4034 );
nand ( n12791 , n12789 , n12790 );
nand ( n12792 , n12791 , n9935 , n10020 );
not ( n12793 , n12792 );
or ( n12794 , n12788 , n12793 );
nand ( n12795 , n12794 , n4272 );
not ( n12796 , n12795 );
not ( n12797 , n4062 );
not ( n12798 , n12797 );
not ( n12799 , n4257 );
or ( n12800 , n12798 , n12799 );
nand ( n12801 , n12800 , n159 );
nor ( n12802 , n12759 , n10092 );
and ( n12803 , n12802 , n9839 , n10080 );
nand ( n12804 , n12796 , n12801 , n160 , n12803 );
nand ( n12805 , n12786 , n12804 );
nand ( n12806 , n12770 , n12773 , n12805 );
nor ( n12807 , n12768 , n12806 );
or ( n12808 , n161 , n12807 );
not ( n12809 , n10867 );
not ( n12810 , n158 );
not ( n12811 , n10122 );
or ( n12812 , n12810 , n12811 );
nand ( n12813 , n12812 , n12767 );
nand ( n12814 , n160 , n12813 );
nand ( n12815 , n12809 , n12814 );
not ( n12816 , n9848 );
nand ( n12817 , n10024 , n12816 );
not ( n12818 , n12704 );
nand ( n12819 , n159 , n12818 );
nand ( n12820 , n12817 , n9912 , n12819 );
nor ( n12821 , n12815 , n12820 );
nand ( n12822 , n12808 , n12821 );
nor ( n12823 , n12753 , n12822 );
xnor ( n12824 , n12693 , n12823 );
not ( n12825 , n177 );
not ( n12826 , n12825 );
not ( n12827 , n5098 );
not ( n12828 , n12827 );
not ( n12829 , n5035 );
nand ( n12830 , n12829 , n4982 );
not ( n12831 , n4899 );
not ( n12832 , n5075 );
or ( n12833 , n12831 , n12832 );
nand ( n12834 , n12833 , n5122 );
nand ( n12835 , n176 , n12834 );
nand ( n12836 , n12828 , n12830 , n12835 );
not ( n12837 , n12836 );
or ( n12838 , n12826 , n12837 );
or ( n12839 , n172 , n4690 );
nand ( n12840 , n12839 , n4664 , n4579 );
nand ( n12841 , n5166 , n12840 );
nand ( n12842 , n12838 , n12841 );
not ( n12843 , n12842 );
not ( n12844 , n177 );
nand ( n12845 , n4795 , n4684 );
and ( n12846 , n176 , n12845 );
not ( n12847 , n176 );
and ( n12848 , n12847 , n4759 );
nor ( n12849 , n12846 , n12848 );
nand ( n12850 , n4614 , n5122 , n4857 , n12849 );
and ( n12851 , n12844 , n12850 );
not ( n12852 , n176 );
or ( n12853 , n12852 , n5122 );
not ( n12854 , n177 );
nor ( n12855 , n12854 , n176 );
not ( n12856 , n12855 );
or ( n12857 , n4622 , n4755 );
nand ( n12858 , n173 , n5127 );
not ( n12859 , n173 );
nand ( n12860 , n12859 , n4868 );
nand ( n12861 , n12857 , n12858 , n12860 );
not ( n12862 , n12861 );
or ( n12863 , n12856 , n12862 );
not ( n12864 , n12113 );
nand ( n12865 , n12863 , n12864 );
not ( n12866 , n12865 );
and ( n12867 , n5062 , n5193 );
nand ( n12868 , n12853 , n12866 , n12867 );
nor ( n12869 , n12851 , n12868 );
not ( n12870 , n5093 );
nand ( n12871 , n4614 , n4750 );
not ( n12872 , n12871 );
not ( n12873 , n12872 );
or ( n12874 , n12870 , n12873 );
not ( n12875 , n176 );
nand ( n12876 , n12874 , n12875 );
nand ( n12877 , n172 , n4713 );
not ( n12878 , n12877 );
nor ( n12879 , n12878 , n4719 );
not ( n12880 , n12879 );
not ( n12881 , n172 );
nor ( n12882 , n12881 , n4979 );
nor ( n12883 , n5087 , n12882 );
not ( n12884 , n12883 );
or ( n12885 , n12880 , n12884 );
nand ( n12886 , n12885 , n177 );
nand ( n12887 , n12869 , n12876 , n12886 );
nand ( n12888 , n178 , n12887 );
not ( n12889 , n4982 );
not ( n12890 , n4979 );
not ( n12891 , n12890 );
nor ( n12892 , n12889 , n12891 );
not ( n12893 , n12892 );
not ( n12894 , n176 );
not ( n12895 , n4601 );
nand ( n12896 , n12894 , n12895 );
nand ( n12897 , n12893 , n12896 , n12080 );
not ( n12898 , n177 );
not ( n12899 , n176 );
nand ( n12900 , n12899 , n4707 );
not ( n12901 , n4658 );
nand ( n12902 , n172 , n12901 );
and ( n12903 , n12900 , n12902 );
or ( n12904 , n12898 , n12903 );
or ( n12905 , n4878 , n5157 );
nand ( n12906 , n12904 , n12905 );
nor ( n12907 , n12897 , n12906 );
not ( n12908 , n176 );
not ( n12909 , n4814 );
nand ( n12910 , n172 , n5129 );
not ( n12911 , n5014 );
nand ( n12912 , n12911 , n172 );
nand ( n12913 , n4899 , n5072 );
nand ( n12914 , n12909 , n12910 , n12912 , n12913 );
not ( n12915 , n12914 );
or ( n12916 , n12908 , n12915 );
nand ( n12917 , n12916 , n12900 );
not ( n12918 , n12858 );
nand ( n12919 , n12918 , n4836 );
not ( n12920 , n176 );
nand ( n12921 , n12920 , n5028 );
and ( n12922 , n12919 , n12921 );
not ( n12923 , n12901 );
not ( n12924 , n177 );
not ( n12925 , n12860 );
nand ( n12926 , n12925 , n4828 );
not ( n12927 , n172 );
not ( n12928 , n4635 );
nand ( n12929 , n12927 , n12928 );
not ( n12930 , n4655 );
nand ( n12931 , n12930 , n4776 );
nand ( n12932 , n12926 , n12929 , n4651 , n12931 );
and ( n12933 , n12924 , n12932 );
not ( n12934 , n12924 );
nand ( n12935 , n4601 , n5003 );
nand ( n12936 , n12912 , n4994 );
nor ( n12937 , n12935 , n12936 );
not ( n12938 , n4694 );
not ( n12939 , n4577 );
or ( n12940 , n12938 , n12939 );
nand ( n12941 , n12940 , n176 );
nand ( n12942 , n5150 , n12941 );
not ( n12943 , n12942 );
not ( n12944 , n176 );
not ( n12945 , n172 );
nand ( n12946 , n12945 , n4749 );
nand ( n12947 , n12946 , n5067 , n4915 );
nand ( n12948 , n12944 , n12947 );
nand ( n12949 , n12937 , n12943 , n12948 );
and ( n12950 , n12934 , n12949 );
nor ( n12951 , n12933 , n12950 );
nand ( n12952 , n12922 , n12923 , n12951 );
or ( n12953 , n12917 , n12952 );
nand ( n12954 , n12953 , n4765 );
and ( n12955 , n12843 , n12888 , n12907 , n12954 );
not ( n12956 , n12955 );
not ( n12957 , n150 );
nand ( n12958 , n12957 , n4318 );
and ( n12959 , n12958 , n4442 , n4536 );
nor ( n12960 , n12959 , n10346 );
not ( n12961 , n12960 );
not ( n12962 , n150 );
nor ( n12963 , n12962 , n10521 );
not ( n12964 , n12963 );
not ( n12965 , n12964 );
nand ( n12966 , n12965 , n149 );
not ( n12967 , n149 );
not ( n12968 , n4546 );
nand ( n12969 , n12967 , n12968 );
not ( n12970 , n10456 );
nand ( n12971 , n12970 , n10610 );
and ( n12972 , n12969 , n12228 , n12971 );
not ( n12973 , n150 );
not ( n12974 , n10498 );
not ( n12975 , n12974 );
or ( n12976 , n12973 , n12975 );
not ( n12977 , n149 );
nand ( n12978 , n12977 , n12224 );
nand ( n12979 , n12976 , n12978 );
and ( n12980 , n152 , n12979 );
not ( n12981 , n152 );
and ( n12982 , n4462 , n10602 );
not ( n12983 , n10426 );
nor ( n12984 , n12982 , n12983 );
not ( n12985 , n4336 );
not ( n12986 , n10366 );
or ( n12987 , n12985 , n12986 );
not ( n12988 , n10484 );
nand ( n12989 , n12987 , n12988 );
nand ( n12990 , n149 , n12989 );
nand ( n12991 , n12984 , n12990 );
and ( n12992 , n12981 , n12991 );
nor ( n12993 , n12980 , n12992 );
and ( n12994 , n12966 , n12972 , n12993 );
nand ( n12995 , n150 , n4369 );
nand ( n12996 , n12995 , n10378 );
not ( n12997 , n12963 );
nand ( n12998 , n12997 , n4386 );
nor ( n12999 , n12996 , n12998 );
or ( n13000 , n4532 , n12999 );
nand ( n13001 , n149 , n10484 );
and ( n13002 , n4562 , n4400 );
not ( n13003 , n13002 );
or ( n13004 , n10433 , n13003 );
not ( n13005 , n149 );
nand ( n13006 , n13004 , n13005 );
nand ( n13007 , n13000 , n13001 , n13006 );
not ( n13008 , n150 );
not ( n13009 , n4312 );
not ( n13010 , n13009 );
or ( n13011 , n13008 , n13010 );
nand ( n13012 , n13011 , n4499 );
and ( n13013 , n149 , n13012 );
not ( n13014 , n149 );
and ( n13015 , n13014 , n4353 );
nor ( n13016 , n13013 , n13015 );
nand ( n13017 , n4562 , n12988 , n10586 , n13016 );
nand ( n13018 , n4532 , n13017 );
not ( n13019 , n12272 );
nor ( n13020 , n4532 , n149 );
not ( n13021 , n10330 );
nand ( n13022 , n147 , n13021 );
nand ( n13023 , n148 , n10405 );
not ( n13024 , n148 );
nand ( n13025 , n13024 , n10319 );
nand ( n13026 , n13022 , n13023 , n13025 );
nand ( n13027 , n13020 , n13026 );
and ( n13028 , n13019 , n13027 );
and ( n13029 , n13028 , n153 , n10418 , n10356 );
nand ( n13030 , n13018 , n13029 );
or ( n13031 , n13007 , n13030 );
not ( n13032 , n150 );
and ( n13033 , n13032 , n4563 );
nor ( n13034 , n4461 , n13025 );
nor ( n13035 , n13033 , n13034 );
nand ( n13036 , n4480 , n4511 );
nand ( n13037 , n4532 , n13035 , n4438 , n13036 );
not ( n13038 , n13037 );
nand ( n13039 , n150 , n10410 );
and ( n13040 , n4546 , n10565 , n13039 , n10555 );
not ( n13041 , n149 );
or ( n13042 , n150 , n4363 );
nand ( n13043 , n13042 , n10371 , n10603 );
and ( n13044 , n13041 , n13043 );
not ( n13045 , n4307 );
not ( n13046 , n10599 );
or ( n13047 , n13045 , n13046 );
nand ( n13048 , n13047 , n149 );
nand ( n13049 , n10325 , n13048 );
nor ( n13050 , n13044 , n13049 );
nand ( n13051 , n152 , n13040 , n13050 );
not ( n13052 , n13051 );
or ( n13053 , n13038 , n13052 );
not ( n13054 , n149 );
not ( n13055 , n150 );
or ( n13056 , n13055 , n10453 );
not ( n13057 , n4514 );
nand ( n13058 , n13056 , n13057 );
nand ( n13059 , n4336 , n4454 );
nand ( n13060 , n13039 , n13059 );
nor ( n13061 , n13058 , n13060 );
nor ( n13062 , n13054 , n13061 );
nor ( n13063 , n153 , n13062 );
not ( n13064 , n12975 );
nor ( n13065 , n4310 , n13023 );
nor ( n13066 , n13064 , n13065 );
not ( n13067 , n149 );
nand ( n13068 , n13067 , n10352 );
and ( n13069 , n13063 , n13066 , n12978 , n13068 );
nand ( n13070 , n13053 , n13069 );
nand ( n13071 , n13031 , n13070 );
nand ( n13072 , n12961 , n12994 , n13071 );
not ( n13073 , n13072 );
not ( n13074 , n13073 );
or ( n13075 , n12956 , n13074 );
not ( n13076 , n12955 );
nand ( n13077 , n13076 , n13072 );
nand ( n13078 , n13075 , n13077 );
and ( n13079 , n12824 , n13078 );
not ( n13080 , n12824 );
not ( n13081 , n13078 );
and ( n13082 , n13080 , n13081 );
nor ( n13083 , n13079 , n13082 );
not ( n13084 , n13083 );
nor ( n13085 , n12692 , n13084 );
or ( n13086 , n10664 , n13083 );
nand ( n13087 , n13086 , n2352 );
or ( n13088 , n13085 , n13087 );
and ( n13089 , n291 , n12693 );
not ( n13090 , n291 );
and ( n13091 , n13090 , n290 );
nor ( n13092 , n13089 , n13091 );
or ( n13093 , n2352 , n13092 );
nand ( n13094 , n13088 , n13093 );
not ( n13095 , n75 );
and ( n13096 , n76 , n13095 );
not ( n13097 , n76 );
and ( n13098 , n13097 , n75 );
nor ( n13099 , n13096 , n13098 );
or ( n13100 , n2352 , n13099 );
not ( n13101 , n7 );
not ( n13102 , n13101 );
nor ( n13103 , n3 , n1016 );
not ( n13104 , n1365 );
nor ( n13105 , n13103 , n13104 );
nand ( n13106 , n13105 , n1409 , n1138 );
not ( n13107 , n13106 );
or ( n13108 , n13102 , n13107 );
not ( n13109 , n3 );
nand ( n13110 , n13109 , n13104 );
nand ( n13111 , n13108 , n13110 );
nor ( n13112 , n13111 , n1393 );
not ( n13113 , n2331 );
nand ( n13114 , n7 , n13113 );
or ( n13115 , n1398 , n2295 , n1073 );
nand ( n13116 , n13115 , n7 );
nand ( n13117 , n13116 , n1270 , n2326 );
nand ( n13118 , n8 , n13117 );
not ( n13119 , n3 );
or ( n13120 , n1136 , n13119 , n999 );
nand ( n13121 , n13120 , n1138 );
or ( n13122 , n3 , n1237 );
or ( n13123 , n7 , n1064 );
nand ( n13124 , n13122 , n13123 , n1066 );
or ( n13125 , n13121 , n13124 );
nand ( n13126 , n13125 , n992 );
nand ( n13127 , n13112 , n13114 , n13118 , n13126 );
and ( n13128 , n9 , n13127 );
not ( n13129 , n9 );
not ( n13130 , n2274 );
nor ( n13131 , n13130 , n1253 );
nand ( n13132 , n7 , n1104 );
not ( n13133 , n1024 );
not ( n13134 , n1039 );
nor ( n13135 , n13133 , n13134 );
or ( n13136 , n2282 , n13135 );
not ( n13137 , n7 );
nand ( n13138 , n13136 , n13137 );
and ( n13139 , n13131 , n13132 , n2221 , n13138 );
or ( n13140 , n13139 , n8 );
not ( n13141 , n2221 );
not ( n13142 , n1086 );
or ( n13143 , n13141 , n13142 );
not ( n13144 , n7 );
nand ( n13145 , n13143 , n13144 );
nand ( n13146 , n13140 , n13145 );
not ( n13147 , n13146 );
not ( n13148 , n8 );
and ( n13149 , n1343 , n2301 );
not ( n13150 , n1121 );
not ( n13151 , n13150 );
not ( n13152 , n1303 );
or ( n13153 , n13151 , n13152 );
nand ( n13154 , n13153 , n7 );
nand ( n13155 , n1136 , n1115 );
not ( n13156 , n13155 );
not ( n13157 , n3 );
not ( n13158 , n1397 );
or ( n13159 , n13157 , n13158 );
not ( n13160 , n3 );
not ( n13161 , n1063 );
nand ( n13162 , n13160 , n13161 );
nand ( n13163 , n13159 , n13162 );
not ( n13164 , n13163 );
or ( n13165 , n13156 , n13164 );
not ( n13166 , n7 );
nand ( n13167 , n13165 , n13166 );
nand ( n13168 , n1291 , n13149 , n13154 , n13167 );
not ( n13169 , n13168 );
or ( n13170 , n13148 , n13169 );
nand ( n13171 , n13170 , n997 );
not ( n13172 , n13171 );
nand ( n13173 , n3 , n13104 );
not ( n13174 , n13173 );
nand ( n13175 , n7 , n13174 );
not ( n13176 , n3 );
not ( n13177 , n13176 );
not ( n13178 , n1350 );
or ( n13179 , n13177 , n13178 );
not ( n13180 , n1147 );
not ( n13181 , n3 );
nand ( n13182 , n13180 , n13181 );
nand ( n13183 , n13179 , n13182 );
nand ( n13184 , n7 , n13183 );
nand ( n13185 , n13147 , n13172 , n13175 , n13184 );
and ( n13186 , n13129 , n13185 );
nor ( n13187 , n13128 , n13186 );
not ( n13188 , n7 );
nand ( n13189 , n1030 , n1359 , n1262 );
nand ( n13190 , n13188 , n13189 );
not ( n13191 , n1255 );
not ( n13192 , n13174 );
nand ( n13193 , n13190 , n13191 , n13192 );
nand ( n13194 , n992 , n13193 );
or ( n13195 , n3 , n1059 );
nand ( n13196 , n13195 , n997 , n1183 );
nand ( n13197 , n1285 , n13196 );
and ( n13198 , n13197 , n1256 , n1352 );
nand ( n13199 , n1136 , n1051 );
not ( n13200 , n2253 );
not ( n13201 , n3 );
nand ( n13202 , n13201 , n1456 );
not ( n13203 , n1351 );
and ( n13204 , n13199 , n13200 , n13202 , n13203 );
or ( n13205 , n7 , n13204 );
not ( n13206 , n1164 );
not ( n13207 , n1290 );
or ( n13208 , n13206 , n13207 );
nand ( n13209 , n13205 , n13208 );
and ( n13210 , n13209 , n8 );
not ( n13211 , n1393 );
not ( n13212 , n1461 );
not ( n13213 , n1270 );
or ( n13214 , n13212 , n13213 );
nand ( n13215 , n13214 , n3 );
nand ( n13216 , n13211 , n13215 );
and ( n13217 , n1425 , n13216 );
nor ( n13218 , n13210 , n13217 );
nand ( n13219 , n13187 , n13194 , n13198 , n13218 );
not ( n13220 , n13219 );
and ( n13221 , n13220 , n9101 );
not ( n13222 , n13220 );
and ( n13223 , n13222 , n9104 );
nor ( n13224 , n13221 , n13223 );
not ( n13225 , n13095 );
not ( n13226 , n16 );
or ( n13227 , n13226 , n771 );
nand ( n13228 , n5784 , n803 , n13227 );
not ( n13229 , n16 );
not ( n13230 , n13229 );
nand ( n13231 , n846 , n813 );
nand ( n13232 , n5757 , n13231 );
not ( n13233 , n13232 );
or ( n13234 , n13230 , n13233 );
nand ( n13235 , n13234 , n5794 );
nor ( n13236 , n13228 , n13235 );
or ( n13237 , n17 , n13236 );
not ( n13238 , n923 );
nand ( n13239 , n13238 , n744 );
nand ( n13240 , n13237 , n13239 );
not ( n13241 , n13240 );
not ( n13242 , n17 );
nand ( n13243 , n5848 , n5706 );
not ( n13244 , n13243 );
not ( n13245 , n12 );
nand ( n13246 , n13245 , n5791 );
not ( n13247 , n13 );
not ( n13248 , n5903 );
or ( n13249 , n13247 , n13248 );
not ( n13250 , n13 );
not ( n13251 , n914 );
nand ( n13252 , n13250 , n13251 );
nand ( n13253 , n13249 , n13252 );
nand ( n13254 , n13246 , n13253 );
not ( n13255 , n16 );
and ( n13256 , n13254 , n13255 );
not ( n13257 , n969 );
nand ( n13258 , n13257 , n5873 );
and ( n13259 , n16 , n13258 );
nor ( n13260 , n13256 , n13259 );
nand ( n13261 , n13244 , n13260 , n5887 );
not ( n13262 , n13261 );
or ( n13263 , n13242 , n13262 );
not ( n13264 , n13 );
not ( n13265 , n13264 );
nor ( n13266 , n11 , n12 );
not ( n13267 , n13266 );
or ( n13268 , n13265 , n13267 );
or ( n13269 , n13 , n5928 );
nand ( n13270 , n13268 , n13269 );
and ( n13271 , n16 , n13270 );
not ( n13272 , n941 );
nor ( n13273 , n13271 , n13272 );
nand ( n13274 , n13263 , n13273 );
not ( n13275 , n13274 );
or ( n13276 , n16 , n5794 );
not ( n13277 , n16 );
and ( n13278 , n13 , n5754 );
not ( n13279 , n13278 );
or ( n13280 , n13277 , n13279 );
nand ( n13281 , n13241 , n13275 , n13276 , n13280 );
and ( n13282 , n13281 , n841 );
not ( n13283 , n5783 );
nand ( n13284 , n5702 , n13283 , n5755 , n884 );
not ( n13285 , n16 );
and ( n13286 , n13284 , n13285 );
not ( n13287 , n5901 );
not ( n13288 , n13287 );
not ( n13289 , n13288 );
not ( n13290 , n13289 );
nor ( n13291 , n13286 , n13290 );
not ( n13292 , n17 );
nand ( n13293 , n878 , n5697 , n5903 );
nand ( n13294 , n16 , n13293 );
nand ( n13295 , n13294 , n816 , n854 );
not ( n13296 , n13295 );
or ( n13297 , n13292 , n13296 );
nand ( n13298 , n16 , n5815 );
nand ( n13299 , n13297 , n13298 );
nor ( n13300 , n16 , n915 );
nor ( n13301 , n916 , n13300 );
not ( n13302 , n13 );
and ( n13303 , n13302 , n842 );
and ( n13304 , n796 , n5682 );
nor ( n13305 , n13303 , n13304 );
and ( n13306 , n13301 , n884 , n13305 );
nor ( n13307 , n13306 , n17 );
nor ( n13308 , n13 , n5755 );
nor ( n13309 , n13299 , n13307 , n13308 );
and ( n13310 , n13291 , n13309 );
nor ( n13311 , n13310 , n841 );
nor ( n13312 , n13282 , n13311 );
nand ( n13313 , n782 , n977 );
or ( n13314 , n13 , n5973 );
not ( n13315 , n12 );
nand ( n13316 , n13315 , n977 );
nand ( n13317 , n13314 , n13316 );
not ( n13318 , n861 );
not ( n13319 , n12 );
nand ( n13320 , n13318 , n13319 );
not ( n13321 , n13320 );
or ( n13322 , n13317 , n13321 , n5776 );
not ( n13323 , n16 );
nand ( n13324 , n13322 , n13323 );
and ( n13325 , n13313 , n13324 );
nor ( n13326 , n13325 , n793 );
not ( n13327 , n13 );
nand ( n13328 , n13327 , n5980 );
not ( n13329 , n894 );
nand ( n13330 , n13328 , n941 , n13329 );
and ( n13331 , n5881 , n13330 );
not ( n13332 , n5884 );
not ( n13333 , n815 );
not ( n13334 , n13333 );
or ( n13335 , n13332 , n13334 );
nand ( n13336 , n13335 , n13 );
nand ( n13337 , n13287 , n13336 );
and ( n13338 , n13337 , n5839 );
nor ( n13339 , n13331 , n13338 );
not ( n13340 , n16 );
not ( n13341 , n13340 );
nand ( n13342 , n5897 , n5911 , n830 );
not ( n13343 , n13342 );
or ( n13344 , n13341 , n13343 );
nor ( n13345 , n806 , n13278 );
nand ( n13346 , n13344 , n13345 );
nand ( n13347 , n793 , n13346 );
nand ( n13348 , n13339 , n13347 , n807 , n5932 );
nor ( n13349 , n13326 , n13348 );
nand ( n13350 , n13312 , n13349 );
not ( n13351 , n13350 );
not ( n13352 , n13351 );
and ( n13353 , n13225 , n13352 );
not ( n13354 , n13350 );
and ( n13355 , n13095 , n13354 );
nor ( n13356 , n13353 , n13355 );
not ( n13357 , n13356 );
and ( n13358 , n13224 , n13357 );
not ( n13359 , n13224 );
and ( n13360 , n13359 , n13356 );
nor ( n13361 , n13358 , n13360 );
not ( n13362 , n13361 );
nand ( n13363 , n25 , n6252 );
nor ( n13364 , n23 , n1914 );
not ( n13365 , n13364 );
nand ( n13366 , n13365 , n6215 );
nand ( n13367 , n6279 , n1813 );
or ( n13368 , n13366 , n13367 );
not ( n13369 , n25 );
nand ( n13370 , n13368 , n13369 );
nand ( n13371 , n13363 , n6406 , n13370 );
not ( n13372 , n13371 );
not ( n13373 , n26 );
not ( n13374 , n25 );
and ( n13375 , n13374 , n1968 );
and ( n13376 , n1940 , n6197 );
nor ( n13377 , n13375 , n13376 );
not ( n13378 , n23 );
nand ( n13379 , n13378 , n1829 );
and ( n13380 , n1969 , n1813 );
nand ( n13381 , n13377 , n13379 , n13380 );
nand ( n13382 , n13373 , n13381 );
not ( n13383 , n6410 );
not ( n13384 , n1780 );
nand ( n13385 , n13383 , n6211 , n13384 );
and ( n13386 , n1987 , n13385 );
not ( n13387 , n23 );
and ( n13388 , n13387 , n6280 );
nor ( n13389 , n13386 , n13388 );
nand ( n13390 , n13372 , n13382 , n13389 );
and ( n13391 , n1875 , n1827 );
not ( n13392 , n26 );
nor ( n13393 , n13391 , n13392 );
or ( n13394 , n13390 , n13393 );
nand ( n13395 , n13394 , n19 );
not ( n13396 , n26 );
nor ( n13397 , n13396 , n25 );
not ( n13398 , n6452 );
not ( n13399 , n6164 );
not ( n13400 , n23 );
nand ( n13401 , n13400 , n6354 );
not ( n13402 , n6363 );
nand ( n13403 , n13398 , n13399 , n13401 , n13402 );
and ( n13404 , n13397 , n13403 );
not ( n13405 , n23 );
or ( n13406 , n13405 , n6350 );
nand ( n13407 , n13406 , n6406 , n1877 );
and ( n13408 , n1987 , n13407 );
nor ( n13409 , n13404 , n13408 );
not ( n13410 , n1975 );
nand ( n13411 , n6370 , n1934 , n1998 );
not ( n13412 , n13411 );
or ( n13413 , n13410 , n13412 );
nand ( n13414 , n26 , n1768 , n1785 );
nand ( n13415 , n13413 , n13414 );
not ( n13416 , n23 );
nand ( n13417 , n13416 , n6333 );
not ( n13418 , n1922 );
not ( n13419 , n1845 );
and ( n13420 , n13417 , n13418 , n13419 );
not ( n13421 , n6462 );
nor ( n13422 , n13420 , n13421 );
not ( n13423 , n1941 );
nand ( n13424 , n1940 , n6163 );
not ( n13425 , n13424 );
or ( n13426 , n13423 , n13425 );
not ( n13427 , n26 );
nand ( n13428 , n13426 , n13427 );
not ( n13429 , n1985 );
nand ( n13430 , n13428 , n13429 , n6364 );
nor ( n13431 , n13415 , n13422 , n13430 );
not ( n13432 , n13424 );
nand ( n13433 , n25 , n13432 );
not ( n13434 , n23 );
not ( n13435 , n13434 );
nor ( n13436 , n21 , n22 );
not ( n13437 , n13436 );
or ( n13438 , n13435 , n13437 );
not ( n13439 , n23 );
nand ( n13440 , n13439 , n1785 );
nand ( n13441 , n13438 , n13440 );
nand ( n13442 , n25 , n13441 );
and ( n13443 , n13418 , n13433 , n13442 );
not ( n13444 , n26 );
not ( n13445 , n25 );
or ( n13446 , n13445 , n1894 );
nand ( n13447 , n13446 , n6300 );
and ( n13448 , n13444 , n13447 );
not ( n13449 , n13444 );
not ( n13450 , n22 );
nand ( n13451 , n13450 , n1859 );
not ( n13452 , n13451 );
and ( n13453 , n23 , n6410 );
not ( n13454 , n23 );
and ( n13455 , n13454 , n6245 );
nor ( n13456 , n13453 , n13455 );
not ( n13457 , n13456 );
or ( n13458 , n13452 , n13457 );
not ( n13459 , n25 );
nand ( n13460 , n13458 , n13459 );
not ( n13461 , n6219 );
nor ( n13462 , n6444 , n13461 );
nand ( n13463 , n13460 , n6465 , n13462 );
and ( n13464 , n13449 , n13463 );
nor ( n13465 , n13448 , n13464 );
nand ( n13466 , n13443 , n13465 );
not ( n13467 , n26 );
not ( n13468 , n6277 );
nand ( n13469 , n6275 , n1893 );
not ( n13470 , n13469 );
or ( n13471 , n13468 , n13470 );
not ( n13472 , n25 );
nand ( n13473 , n13471 , n13472 );
not ( n13474 , n1982 );
nand ( n13475 , n13473 , n6170 , n13474 );
nand ( n13476 , n13467 , n13475 );
not ( n13477 , n6392 );
or ( n13478 , n1899 , n13477 );
nand ( n13479 , n13478 , n1987 );
not ( n13480 , n6170 );
not ( n13481 , n1956 );
or ( n13482 , n13480 , n13481 );
not ( n13483 , n25 );
nand ( n13484 , n13482 , n13483 );
nand ( n13485 , n13476 , n13479 , n13484 );
or ( n13486 , n13466 , n13485 );
nand ( n13487 , n13486 , n1853 );
nand ( n13488 , n13395 , n13409 , n13431 , n13487 );
not ( n13489 , n13488 );
not ( n13490 , n13489 );
not ( n13491 , n1673 );
not ( n13492 , n31 );
not ( n13493 , n13492 );
nand ( n13494 , n2158 , n1749 );
not ( n13495 , n13494 );
or ( n13496 , n13493 , n13495 );
nand ( n13497 , n1629 , n1497 );
not ( n13498 , n13497 );
not ( n13499 , n32 );
nand ( n13500 , n13498 , n13499 );
nand ( n13501 , n13496 , n13500 );
not ( n13502 , n33 );
nand ( n13503 , n13501 , n13502 );
not ( n13504 , n31 );
not ( n13505 , n27 );
nand ( n13506 , n13505 , n1611 );
not ( n13507 , n13506 );
nand ( n13508 , n13504 , n13507 );
and ( n13509 , n6023 , n13508 );
nand ( n13510 , n6022 , n13509 );
not ( n13511 , n32 );
and ( n13512 , n13510 , n13511 );
not ( n13513 , n1615 );
not ( n13514 , n13513 );
or ( n13515 , n31 , n13514 );
nand ( n13516 , n13515 , n1710 );
and ( n13517 , n2188 , n13516 );
nor ( n13518 , n13512 , n13517 );
nand ( n13519 , n1698 , n1735 );
nand ( n13520 , n32 , n6072 , n13519 );
not ( n13521 , n32 );
or ( n13522 , n13521 , n2171 );
nand ( n13523 , n1733 , n1608 );
not ( n13524 , n1498 );
nand ( n13525 , n13522 , n13523 , n13524 );
nand ( n13526 , n1701 , n1629 );
nand ( n13527 , n1714 , n13526 );
or ( n13528 , n13525 , n13527 );
nand ( n13529 , n13528 , n33 );
nand ( n13530 , n13503 , n13518 , n13520 , n13529 );
not ( n13531 , n13530 );
or ( n13532 , n13491 , n13531 );
not ( n13533 , n33 );
nand ( n13534 , n1515 , n1521 );
not ( n13535 , n32 );
not ( n13536 , n31 );
nand ( n13537 , n13536 , n2068 );
nand ( n13538 , n13537 , n2115 , n1548 );
nand ( n13539 , n13535 , n13538 );
nand ( n13540 , n13534 , n1495 , n13539 );
and ( n13541 , n13533 , n13540 );
not ( n13542 , n1677 );
not ( n13543 , n13542 );
not ( n13544 , n31 );
nand ( n13545 , n13544 , n2039 );
not ( n13546 , n13545 );
nor ( n13547 , n13543 , n13546 );
nor ( n13548 , n2125 , n1532 );
nand ( n13549 , n32 , n13548 );
not ( n13550 , n32 );
not ( n13551 , n1617 );
nand ( n13552 , n13550 , n13551 );
not ( n13553 , n6039 );
and ( n13554 , n13549 , n13552 , n13553 );
and ( n13555 , n13547 , n13554 );
not ( n13556 , n33 );
nor ( n13557 , n13555 , n13556 );
nor ( n13558 , n13541 , n13557 );
nand ( n13559 , n13532 , n13558 );
not ( n13560 , n13559 );
not ( n13561 , n32 );
not ( n13562 , n13526 );
nand ( n13563 , n13561 , n13562 );
not ( n13564 , n2198 );
nand ( n13565 , n32 , n13564 );
not ( n13566 , n6043 );
not ( n13567 , n1546 );
or ( n13568 , n13566 , n13567 );
nand ( n13569 , n13568 , n2188 );
and ( n13570 , n13563 , n13565 , n13569 );
and ( n13571 , n1553 , n1727 );
not ( n13572 , n32 );
not ( n13573 , n2126 );
nand ( n13574 , n13573 , n1652 );
nand ( n13575 , n13572 , n13574 );
nand ( n13576 , n2056 , n6022 );
not ( n13577 , n27 );
nor ( n13578 , n13577 , n1517 );
and ( n13579 , n31 , n13578 );
not ( n13580 , n13579 );
nand ( n13581 , n1607 , n13580 );
or ( n13582 , n13576 , n13581 );
nand ( n13583 , n13582 , n32 );
nand ( n13584 , n13571 , n13575 , n13583 );
not ( n13585 , n32 );
nand ( n13586 , n13585 , n6042 );
nand ( n13587 , n13586 , n1534 , n5998 );
nand ( n13588 , n33 , n13587 );
not ( n13589 , n32 );
not ( n13590 , n31 );
nor ( n13591 , n27 , n29 );
not ( n13592 , n13591 );
or ( n13593 , n13590 , n13592 );
nand ( n13594 , n13593 , n1700 );
nand ( n13595 , n13589 , n13594 );
nand ( n13596 , n31 , n1589 );
nand ( n13597 , n13596 , n1574 );
nand ( n13598 , n1540 , n6072 );
not ( n13599 , n2166 );
nand ( n13600 , n1608 , n13599 );
not ( n13601 , n31 );
nand ( n13602 , n13601 , n2064 , n1704 );
nand ( n13603 , n13602 , n1582 , n2142 );
nand ( n13604 , n32 , n13603 );
nand ( n13605 , n13598 , n13600 , n13604 );
or ( n13606 , n13597 , n13605 );
not ( n13607 , n33 );
nand ( n13608 , n13606 , n13607 );
nand ( n13609 , n13588 , n13595 , n13608 );
or ( n13610 , n13584 , n13609 );
nand ( n13611 , n13610 , n34 );
and ( n13612 , n13560 , n13570 , n13611 );
buf ( n13613 , n13612 );
not ( n13614 , n13613 );
or ( n13615 , n13490 , n13614 );
buf ( n13616 , n13488 );
not ( n13617 , n13616 );
or ( n13618 , n13613 , n13617 );
nand ( n13619 , n13615 , n13618 );
not ( n13620 , n9 );
or ( n13621 , n7 , n1037 );
and ( n13622 , n13621 , n2283 , n1116 );
nor ( n13623 , n13622 , n992 );
not ( n13624 , n7 );
not ( n13625 , n1359 );
nor ( n13626 , n13625 , n1220 );
nand ( n13627 , n13626 , n1086 , n13173 );
not ( n13628 , n13627 );
or ( n13629 , n13624 , n13628 );
not ( n13630 , n1181 );
not ( n13631 , n1453 );
or ( n13632 , n13630 , n13631 );
not ( n13633 , n7 );
nand ( n13634 , n13632 , n13633 );
nand ( n13635 , n13629 , n13634 );
nor ( n13636 , n13623 , n13635 );
not ( n13637 , n13103 );
nand ( n13638 , n3 , n1222 );
and ( n13639 , n13637 , n13638 );
not ( n13640 , n2245 );
nand ( n13641 , n3 , n13640 );
and ( n13642 , n13641 , n1306 );
not ( n13643 , n6 );
nand ( n13644 , n13643 , n1050 );
not ( n13645 , n1042 );
nand ( n13646 , n1229 , n13645 );
nand ( n13647 , n1293 , n1373 , n13182 );
nand ( n13648 , n7 , n13647 );
nand ( n13649 , n13642 , n13644 , n13646 , n13648 );
and ( n13650 , n992 , n13649 );
nand ( n13651 , n3 , n1350 );
and ( n13652 , n2297 , n13651 );
nor ( n13653 , n13652 , n7 );
nor ( n13654 , n13650 , n13653 );
nand ( n13655 , n13636 , n13639 , n13654 );
not ( n13656 , n13655 );
or ( n13657 , n13620 , n13656 );
and ( n13658 , n7 , n1278 );
not ( n13659 , n7 );
nand ( n13660 , n4 , n2295 );
and ( n13661 , n13659 , n13660 );
or ( n13662 , n13658 , n13661 );
nand ( n13663 , n13657 , n13662 );
nand ( n13664 , n1277 , n1290 );
nor ( n13665 , n1392 , n1057 );
and ( n13666 , n7 , n13665 );
not ( n13667 , n7 );
and ( n13668 , n13667 , n1123 );
nor ( n13669 , n13666 , n13668 );
not ( n13670 , n2317 );
nand ( n13671 , n13664 , n13669 , n1012 , n13670 );
nand ( n13672 , n8 , n13671 );
not ( n13673 , n7 );
not ( n13674 , n3 );
nand ( n13675 , n13674 , n1056 );
nand ( n13676 , n13675 , n1416 , n2279 );
and ( n13677 , n13673 , n13676 );
not ( n13678 , n13673 );
nand ( n13679 , n1040 , n2278 );
and ( n13680 , n13678 , n13679 );
nor ( n13681 , n13677 , n13680 );
nand ( n13682 , n13681 , n13175 , n2270 );
nand ( n13683 , n992 , n13682 );
not ( n13684 , n7 );
not ( n13685 , n13684 );
not ( n13686 , n13155 );
not ( n13687 , n3 );
nand ( n13688 , n13686 , n13687 );
nand ( n13689 , n13688 , n1079 , n1086 );
not ( n13690 , n13689 );
or ( n13691 , n13685 , n13690 );
not ( n13692 , n2214 );
nand ( n13693 , n1447 , n13692 );
nand ( n13694 , n13693 , n7 , n1050 );
nand ( n13695 , n13691 , n13694 );
nand ( n13696 , n1097 , n1229 );
nand ( n13697 , n13696 , n1433 , n13660 );
not ( n13698 , n13697 );
not ( n13699 , n1343 );
nand ( n13700 , n7 , n13699 );
not ( n13701 , n2265 );
nand ( n13702 , n13698 , n13700 , n13701 );
nand ( n13703 , n8 , n13702 );
or ( n13704 , n3 , n1120 );
nand ( n13705 , n13704 , n1096 );
nand ( n13706 , n1285 , n13705 );
not ( n13707 , n3 );
not ( n13708 , n13707 );
not ( n13709 , n1326 );
or ( n13710 , n13708 , n13709 );
nand ( n13711 , n1164 , n1152 );
nand ( n13712 , n13710 , n13711 );
nand ( n13713 , n992 , n13712 );
nand ( n13714 , n13703 , n13706 , n13713 );
or ( n13715 , n13695 , n13714 );
nand ( n13716 , n13715 , n1133 );
nand ( n13717 , n13672 , n13683 , n13716 );
nor ( n13718 , n13663 , n13717 );
xor ( n13719 , n13718 , n2209 );
and ( n13720 , n13619 , n13719 );
not ( n13721 , n13619 );
not ( n13722 , n13719 );
and ( n13723 , n13721 , n13722 );
nor ( n13724 , n13720 , n13723 );
not ( n13725 , n13724 );
nand ( n13726 , n13362 , n13725 );
nand ( n13727 , n13361 , n13724 );
nand ( n13728 , n13726 , n2352 , n13727 );
nand ( n13729 , n13100 , n13728 );
not ( n13730 , n5989 );
not ( n13731 , n86 );
and ( n13732 , n13730 , n13731 );
not ( n13733 , n13730 );
and ( n13734 , n13733 , n86 );
nor ( n13735 , n13732 , n13734 );
not ( n13736 , n992 );
and ( n13737 , n1375 , n2279 );
not ( n13738 , n7 );
not ( n13739 , n3 );
nand ( n13740 , n13739 , n1398 );
not ( n13741 , n2330 );
nand ( n13742 , n13740 , n13741 , n2221 );
nand ( n13743 , n13738 , n13742 );
nand ( n13744 , n1457 , n13200 );
nand ( n13745 , n2278 , n1343 , n1044 );
or ( n13746 , n13744 , n13745 );
nand ( n13747 , n13746 , n7 );
nand ( n13748 , n13737 , n13743 , n13747 );
not ( n13749 , n13748 );
or ( n13750 , n13736 , n13749 );
not ( n13751 , n7 );
nand ( n13752 , n13751 , n2290 );
nand ( n13753 , n13750 , n13752 );
not ( n13754 , n13753 );
nand ( n13755 , n1170 , n1288 );
not ( n13756 , n1416 );
nand ( n13757 , n7 , n13756 );
nand ( n13758 , n7 , n1319 );
and ( n13759 , n13757 , n13758 , n13638 );
not ( n13760 , n7 );
not ( n13761 , n3 );
nand ( n13762 , n1072 , n1447 );
not ( n13763 , n13762 );
or ( n13764 , n13761 , n13763 );
nand ( n13765 , n13764 , n1201 , n13664 );
nand ( n13766 , n13760 , n13765 );
nand ( n13767 , n13759 , n1295 , n13766 );
nand ( n13768 , n8 , n13767 );
and ( n13769 , n13755 , n13768 );
not ( n13770 , n8 );
and ( n13771 , n1179 , n1018 );
nand ( n13772 , n1159 , n1381 );
not ( n13773 , n7 );
not ( n13774 , n3 );
not ( n13775 , n1096 );
nand ( n13776 , n13774 , n13775 );
nand ( n13777 , n1221 , n1215 , n13776 );
nand ( n13778 , n13773 , n13777 );
nand ( n13779 , n13771 , n13772 , n13778 );
not ( n13780 , n13779 );
or ( n13781 , n13770 , n13780 );
not ( n13782 , n3 );
not ( n13783 , n13782 );
not ( n13784 , n1448 );
or ( n13785 , n13783 , n13784 );
nand ( n13786 , n13785 , n1280 );
nand ( n13787 , n7 , n13786 );
nand ( n13788 , n13781 , n13787 );
not ( n13789 , n13788 );
not ( n13790 , n7 );
not ( n13791 , n13211 );
and ( n13792 , n13790 , n13791 );
nand ( n13793 , n3 , n2265 );
nand ( n13794 , n7 , n1288 );
not ( n13795 , n7 );
nand ( n13796 , n13795 , n13103 );
nand ( n13797 , n13793 , n1384 , n13794 , n13796 );
and ( n13798 , n13797 , n992 );
nor ( n13799 , n13792 , n13798 );
nand ( n13800 , n13789 , n1133 , n2279 , n13799 );
not ( n13801 , n8 );
not ( n13802 , n1262 );
nor ( n13803 , n13802 , n2317 );
not ( n13804 , n1231 );
not ( n13805 , n1042 );
or ( n13806 , n13804 , n13805 );
not ( n13807 , n7 );
nand ( n13808 , n13806 , n13807 );
nand ( n13809 , n13803 , n2247 , n13808 );
not ( n13810 , n13809 );
or ( n13811 , n13801 , n13810 );
not ( n13812 , n7 );
nand ( n13813 , n13664 , n1105 , n2301 );
nand ( n13814 , n13812 , n13813 );
nand ( n13815 , n13811 , n13814 );
not ( n13816 , n13815 );
and ( n13817 , n1136 , n1401 );
and ( n13818 , n1114 , n2324 );
nor ( n13819 , n13817 , n13818 );
not ( n13820 , n1194 );
nand ( n13821 , n13819 , n1142 , n13820 );
nand ( n13822 , n7 , n13821 );
not ( n13823 , n1248 );
nand ( n13824 , n13823 , n13711 );
not ( n13825 , n7 );
nand ( n13826 , n13825 , n1358 );
not ( n13827 , n1120 );
nand ( n13828 , n3 , n13827 );
nand ( n13829 , n13826 , n13828 , n1217 );
or ( n13830 , n13824 , n13829 );
nand ( n13831 , n13830 , n992 );
nand ( n13832 , n13816 , n9 , n13822 , n13831 );
nand ( n13833 , n13800 , n13832 );
nand ( n13834 , n13754 , n13769 , n13833 );
and ( n13835 , n13834 , n987 );
not ( n13836 , n13834 );
and ( n13837 , n13836 , n986 );
nor ( n13838 , n13835 , n13837 );
xor ( n13839 , n13735 , n13838 );
not ( n13840 , n13839 );
not ( n13841 , n26 );
not ( n13842 , n13841 );
not ( n13843 , n6276 );
nor ( n13844 , n13843 , n6178 );
not ( n13845 , n25 );
not ( n13846 , n23 );
nand ( n13847 , n13846 , n6410 );
not ( n13848 , n6252 );
nand ( n13849 , n13847 , n13848 , n6170 );
nand ( n13850 , n13845 , n13849 );
nor ( n13851 , n6444 , n6302 );
nand ( n13852 , n13851 , n13399 , n6355 , n1941 );
nand ( n13853 , n25 , n13852 );
nand ( n13854 , n13844 , n13850 , n13853 );
not ( n13855 , n13854 );
or ( n13856 , n13842 , n13855 );
not ( n13857 , n1814 );
or ( n13858 , n25 , n13857 );
nand ( n13859 , n25 , n6349 );
nand ( n13860 , n13858 , n13859 );
nand ( n13861 , n23 , n13860 );
nand ( n13862 , n13856 , n13861 );
not ( n13863 , n13862 );
not ( n13864 , n6342 );
nand ( n13865 , n13864 , n25 );
nor ( n13866 , n1799 , n6235 );
not ( n13867 , n13866 );
and ( n13868 , n13865 , n13867 , n1868 );
not ( n13869 , n25 );
nand ( n13870 , n6206 , n1779 );
nand ( n13871 , n23 , n13870 );
not ( n13872 , n1784 );
nand ( n13873 , n13872 , n6275 );
nand ( n13874 , n13871 , n1839 , n13873 );
nand ( n13875 , n13869 , n13874 );
nand ( n13876 , n13868 , n6331 , n13875 );
nand ( n13877 , n26 , n13876 );
not ( n13878 , n26 );
not ( n13879 , n13878 );
not ( n13880 , n1858 );
not ( n13881 , n1984 );
or ( n13882 , n13880 , n13881 );
not ( n13883 , n25 );
nand ( n13884 , n13882 , n13883 );
and ( n13885 , n6268 , n6191 , n1998 , n13884 );
not ( n13886 , n13885 );
and ( n13887 , n13879 , n13886 );
not ( n13888 , n25 );
nand ( n13889 , n1894 , n6219 , n13873 );
and ( n13890 , n13888 , n13889 );
nor ( n13891 , n13887 , n13890 );
not ( n13892 , n21 );
and ( n13893 , n13892 , n1997 );
and ( n13894 , n1812 , n6414 );
nor ( n13895 , n13893 , n13894 );
nand ( n13896 , n13895 , n1849 , n1834 );
nand ( n13897 , n25 , n13896 );
not ( n13898 , n1980 );
not ( n13899 , n25 );
not ( n13900 , n1774 );
nand ( n13901 , n13900 , n23 );
not ( n13902 , n13901 );
nand ( n13903 , n13899 , n13902 );
nand ( n13904 , n13898 , n13903 );
not ( n13905 , n25 );
nand ( n13906 , n13905 , n6369 );
not ( n13907 , n1789 );
nand ( n13908 , n23 , n13907 );
nand ( n13909 , n13906 , n13908 , n1865 );
or ( n13910 , n13904 , n13909 );
not ( n13911 , n26 );
nand ( n13912 , n13910 , n13911 );
nand ( n13913 , n13891 , n13897 , n13912 );
or ( n13914 , n13913 , n1853 );
or ( n13915 , n23 , n6311 );
nand ( n13916 , n13915 , n6456 );
and ( n13917 , n25 , n13916 );
not ( n13918 , n23 );
not ( n13919 , n1887 );
nand ( n13920 , n13918 , n13919 );
not ( n13921 , n1765 );
and ( n13922 , n13920 , n13921 , n6160 );
not ( n13923 , n13397 );
nor ( n13924 , n13922 , n13923 );
nor ( n13925 , n13917 , n13924 );
not ( n13926 , n25 );
not ( n13927 , n6406 );
nand ( n13928 , n13926 , n13927 );
nor ( n13929 , n1793 , n1889 );
nor ( n13930 , n1915 , n13929 );
and ( n13931 , n26 , n13930 );
not ( n13932 , n26 );
not ( n13933 , n1855 );
not ( n13934 , n13933 );
not ( n13935 , n1914 );
and ( n13936 , n13934 , n13935 );
not ( n13937 , n23 );
nor ( n13938 , n13937 , n1921 );
nor ( n13939 , n13936 , n13938 );
and ( n13940 , n13932 , n13939 );
nor ( n13941 , n13931 , n13940 );
nand ( n13942 , n26 , n1844 );
not ( n13943 , n13859 );
not ( n13944 , n6381 );
or ( n13945 , n13943 , n13944 );
not ( n13946 , n26 );
nand ( n13947 , n13945 , n13946 );
nand ( n13948 , n13942 , n6276 , n13947 );
nor ( n13949 , n13941 , n13948 , n19 );
nand ( n13950 , n13925 , n13928 , n13949 );
nand ( n13951 , n13914 , n13950 );
and ( n13952 , n13863 , n13877 , n13951 );
or ( n13953 , n28 , n6073 );
nand ( n13954 , n13953 , n6124 );
nand ( n13955 , n32 , n13954 );
or ( n13956 , n29 , n2125 );
nand ( n13957 , n13956 , n2158 );
and ( n13958 , n32 , n13957 );
not ( n13959 , n32 );
nand ( n13960 , n6076 , n1717 , n13545 );
and ( n13961 , n13959 , n13960 );
nor ( n13962 , n13958 , n13961 );
not ( n13963 , n33 );
not ( n13964 , n32 );
nand ( n13965 , n13964 , n2055 );
nand ( n13966 , n31 , n13513 );
and ( n13967 , n13965 , n13966 , n13500 );
nand ( n13968 , n13967 , n1569 , n6067 );
nand ( n13969 , n13963 , n13968 );
nand ( n13970 , n13542 , n6052 );
not ( n13971 , n6059 );
not ( n13972 , n2166 );
or ( n13973 , n13971 , n13972 );
not ( n13974 , n32 );
nand ( n13975 , n13973 , n13974 );
nand ( n13976 , n1590 , n13975 );
or ( n13977 , n13970 , n13976 );
nand ( n13978 , n13977 , n33 );
nand ( n13979 , n13955 , n13962 , n13969 , n13978 );
and ( n13980 , n34 , n13979 );
not ( n13981 , n34 );
not ( n13982 , n33 );
not ( n13983 , n31 );
nor ( n13984 , n13983 , n13524 );
not ( n13985 , n13984 );
and ( n13986 , n13985 , n2034 );
not ( n13987 , n32 );
and ( n13988 , n13987 , n1553 );
not ( n13989 , n13987 );
and ( n13990 , n13989 , n2091 );
or ( n13991 , n13988 , n13990 );
nand ( n13992 , n13986 , n13991 );
and ( n13993 , n13982 , n13992 );
nor ( n13994 , n32 , n2060 );
nor ( n13995 , n13993 , n13994 );
not ( n13996 , n31 );
not ( n13997 , n13996 );
not ( n13998 , n2130 );
or ( n13999 , n13997 , n13998 );
nand ( n14000 , n13999 , n2201 );
nand ( n14001 , n32 , n14000 );
nand ( n14002 , n6097 , n1592 );
not ( n14003 , n32 );
not ( n14004 , n14003 );
not ( n14005 , n31 );
not ( n14006 , n1710 );
nand ( n14007 , n14005 , n14006 );
nand ( n14008 , n14007 , n6002 , n1607 );
not ( n14009 , n14008 );
or ( n14010 , n14004 , n14009 );
nand ( n14011 , n2074 , n2027 );
nand ( n14012 , n14010 , n14011 );
or ( n14013 , n14002 , n14012 );
nand ( n14014 , n14013 , n33 );
nand ( n14015 , n13995 , n1548 , n14001 , n14014 );
and ( n14016 , n13981 , n14015 );
nor ( n14017 , n13980 , n14016 );
not ( n14018 , n33 );
and ( n14019 , n1630 , n1548 );
not ( n14020 , n32 );
not ( n14021 , n2077 );
not ( n14022 , n31 );
nand ( n14023 , n14021 , n14022 );
nand ( n14024 , n14023 , n1669 , n1624 );
nand ( n14025 , n14020 , n14024 );
buf ( n14026 , n2171 );
nand ( n14027 , n14026 , n2109 );
nand ( n14028 , n1546 , n1576 , n6036 );
or ( n14029 , n14027 , n14028 );
nand ( n14030 , n14029 , n32 );
nand ( n14031 , n14019 , n14025 , n14030 );
nand ( n14032 , n14018 , n14031 );
not ( n14033 , n33 );
not ( n14034 , n2115 );
and ( n14035 , n32 , n14034 );
nor ( n14036 , n1514 , n1519 );
nor ( n14037 , n14035 , n14036 );
or ( n14038 , n14033 , n14037 );
not ( n14039 , n6054 );
or ( n14040 , n1692 , n14039 );
nand ( n14041 , n14038 , n14040 );
not ( n14042 , n33 );
not ( n14043 , n32 );
not ( n14044 , n14043 );
nand ( n14045 , n1698 , n1732 );
nand ( n14046 , n31 , n14045 );
nand ( n14047 , n14046 , n6127 , n13545 );
not ( n14048 , n14047 );
or ( n14049 , n14044 , n14048 );
and ( n14050 , n2133 , n1727 );
nand ( n14051 , n14049 , n14050 );
not ( n14052 , n14051 );
or ( n14053 , n14042 , n14052 );
nand ( n14054 , n32 , n6042 , n1629 );
nand ( n14055 , n14053 , n14054 );
nor ( n14056 , n14041 , n14055 );
and ( n14057 , n14017 , n14032 , n14056 );
and ( n14058 , n13952 , n14057 );
not ( n14059 , n13952 );
nand ( n14060 , n14032 , n14056 );
not ( n14061 , n14060 );
nand ( n14062 , n14061 , n14017 );
buf ( n14063 , n14062 );
and ( n14064 , n14059 , n14063 );
nor ( n14065 , n14058 , n14064 );
not ( n14066 , n14065 );
not ( n14067 , n14066 );
nor ( n14068 , n6151 , n6481 );
not ( n14069 , n14068 );
not ( n14070 , n6473 );
nand ( n14071 , n14070 , n6151 );
nand ( n14072 , n14069 , n14071 );
not ( n14073 , n14072 );
or ( n14074 , n14067 , n14073 );
and ( n14075 , n13863 , n13877 , n13951 );
xor ( n14076 , n14062 , n14075 );
buf ( n14077 , n14076 );
or ( n14078 , n14077 , n14072 );
nand ( n14079 , n14074 , n14078 );
not ( n14080 , n14079 );
or ( n14081 , n13840 , n14080 );
nand ( n14082 , n14081 , n2352 );
nor ( n14083 , n13839 , n14079 );
or ( n14084 , n14082 , n14083 );
and ( n14085 , n87 , n13731 );
not ( n14086 , n87 );
and ( n14087 , n14086 , n86 );
nor ( n14088 , n14085 , n14087 );
or ( n14089 , n2352 , n14088 );
nand ( n14090 , n14084 , n14089 );
not ( n14091 , n78 );
not ( n14092 , n14091 );
not ( n14093 , n17 );
not ( n14094 , n893 );
and ( n14095 , n14094 , n931 );
nand ( n14096 , n833 , n5925 );
not ( n14097 , n16 );
not ( n14098 , n960 );
not ( n14099 , n13 );
nand ( n14100 , n14098 , n14099 );
nand ( n14101 , n14100 , n5722 , n789 );
nand ( n14102 , n14097 , n14101 );
nand ( n14103 , n14095 , n14096 , n14102 );
not ( n14104 , n14103 );
or ( n14105 , n14093 , n14104 );
or ( n14106 , n13 , n5948 );
nand ( n14107 , n14106 , n5861 );
nand ( n14108 , n16 , n14107 );
nand ( n14109 , n14105 , n14108 );
not ( n14110 , n13 );
nor ( n14111 , n14110 , n939 );
nor ( n14112 , n14111 , n5929 );
not ( n14113 , n14112 );
and ( n14114 , n16 , n5885 );
not ( n14115 , n16 );
and ( n14116 , n14115 , n5783 );
nor ( n14117 , n14114 , n14116 );
not ( n14118 , n14117 );
or ( n14119 , n14113 , n14118 );
nand ( n14120 , n14119 , n793 );
not ( n14121 , n16 );
nand ( n14122 , n14121 , n13288 );
nand ( n14123 , n14120 , n5749 , n14122 );
or ( n14124 , n14109 , n14123 );
nand ( n14125 , n14124 , n841 );
not ( n14126 , n14125 );
not ( n14127 , n14126 );
not ( n14128 , n10 );
not ( n14129 , n793 );
not ( n14130 , n795 );
nand ( n14131 , n14130 , n866 );
not ( n14132 , n14131 );
not ( n14133 , n16 );
nand ( n14134 , n14132 , n14133 );
not ( n14135 , n14134 );
not ( n14136 , n5896 );
nor ( n14137 , n16 , n14136 );
not ( n14138 , n13 );
nor ( n14139 , n14138 , n868 );
nor ( n14140 , n14135 , n14137 , n14139 );
nand ( n14141 , n14140 , n820 , n779 );
not ( n14142 , n14141 );
or ( n14143 , n14129 , n14142 );
not ( n14144 , n12 );
and ( n14145 , n14144 , n5907 );
not ( n14146 , n858 );
and ( n14147 , n755 , n14146 );
nor ( n14148 , n14145 , n14147 );
nand ( n14149 , n14148 , n902 , n844 );
nand ( n14150 , n16 , n14149 );
nand ( n14151 , n14143 , n14150 );
not ( n14152 , n14151 );
not ( n14153 , n16 );
not ( n14154 , n846 );
or ( n14155 , n14154 , n5928 );
nand ( n14156 , n14155 , n771 , n5706 );
nand ( n14157 , n14153 , n14156 );
and ( n14158 , n5718 , n830 );
not ( n14159 , n754 );
not ( n14160 , n5844 );
or ( n14161 , n14159 , n14160 );
not ( n14162 , n16 );
nand ( n14163 , n14161 , n14162 );
nand ( n14164 , n14158 , n5768 , n14163 );
nand ( n14165 , n17 , n14164 );
nand ( n14166 , n14152 , n14157 , n14165 );
not ( n14167 , n14166 );
or ( n14168 , n14128 , n14167 );
not ( n14169 , n16 );
and ( n14170 , n14169 , n5811 );
and ( n14171 , n810 , n5885 );
nor ( n14172 , n14170 , n14171 );
nand ( n14173 , n14168 , n14172 );
not ( n14174 , n14173 );
and ( n14175 , n5803 , n5749 );
not ( n14176 , n16 );
or ( n14177 , n13 , n5903 );
nand ( n14178 , n14177 , n5814 , n5794 );
and ( n14179 , n14176 , n14178 );
not ( n14180 , n14176 );
nor ( n14181 , n5776 , n5745 );
not ( n14182 , n5848 );
not ( n14183 , n5974 );
nand ( n14184 , n14183 , n805 );
nor ( n14185 , n14182 , n14184 );
nand ( n14186 , n14181 , n14185 );
and ( n14187 , n14180 , n14186 );
nor ( n14188 , n14179 , n14187 );
nand ( n14189 , n14175 , n14188 );
nand ( n14190 , n14189 , n793 );
nand ( n14191 , n16 , n5962 );
nand ( n14192 , n810 , n5774 );
nand ( n14193 , n13 , n790 );
and ( n14194 , n14191 , n14192 , n14193 );
not ( n14195 , n16 );
not ( n14196 , n13 );
nand ( n14197 , n876 , n5693 );
not ( n14198 , n14197 );
or ( n14199 , n14196 , n14198 );
nand ( n14200 , n14199 , n850 , n14155 );
and ( n14201 , n14195 , n14200 );
not ( n14202 , n5890 );
nor ( n14203 , n14201 , n14202 );
nand ( n14204 , n14194 , n14203 );
nand ( n14205 , n17 , n14204 );
nand ( n14206 , n14127 , n14174 , n14190 , n14205 );
not ( n14207 , n14206 );
not ( n14208 , n14207 );
and ( n14209 , n14092 , n14208 );
not ( n14210 , n14206 );
and ( n14211 , n14091 , n14210 );
nor ( n14212 , n14209 , n14211 );
and ( n14213 , n13800 , n13832 );
nor ( n14214 , n14213 , n13753 );
nand ( n14215 , n13769 , n14214 );
not ( n14216 , n14215 );
not ( n14217 , n14216 );
not ( n14218 , n14057 );
and ( n14219 , n14217 , n14218 );
not ( n14220 , n14215 );
and ( n14221 , n14220 , n14057 );
nor ( n14222 , n14219 , n14221 );
xor ( n14223 , n14212 , n14222 );
not ( n14224 , n14223 );
not ( n14225 , n14072 );
not ( n14226 , n2209 );
not ( n14227 , n14226 );
not ( n14228 , n6145 );
not ( n14229 , n14228 );
and ( n14230 , n14227 , n14229 );
and ( n14231 , n14226 , n14228 );
nor ( n14232 , n14230 , n14231 );
not ( n14233 , n14232 );
or ( n14234 , n14225 , n14233 );
or ( n14235 , n14232 , n14072 );
nand ( n14236 , n14234 , n14235 );
not ( n14237 , n14236 );
nor ( n14238 , n14224 , n14237 );
or ( n14239 , n14236 , n14223 );
nand ( n14240 , n14239 , n2352 );
or ( n14241 , n14238 , n14240 );
and ( n14242 , n92 , n14091 );
not ( n14243 , n92 );
and ( n14244 , n14243 , n78 );
nor ( n14245 , n14242 , n14244 );
or ( n14246 , n2352 , n14245 );
nand ( n14247 , n14241 , n14246 );
not ( n14248 , n13219 );
not ( n14249 , n10 );
not ( n14250 , n853 );
not ( n14251 , n5945 );
and ( n14252 , n14250 , n14251 );
nor ( n14253 , n14252 , n16 );
not ( n14254 , n16 );
not ( n14255 , n5897 );
nor ( n14256 , n14255 , n13278 );
nand ( n14257 , n789 , n926 , n14256 );
not ( n14258 , n14257 );
or ( n14259 , n14254 , n14258 );
nand ( n14260 , n14259 , n13283 );
nor ( n14261 , n14253 , n14260 );
or ( n14262 , n16 , n765 );
not ( n14263 , n978 );
nand ( n14264 , n14262 , n5757 , n14263 );
and ( n14265 , n17 , n14264 );
not ( n14266 , n16 );
not ( n14267 , n13 );
not ( n14268 , n13266 );
or ( n14269 , n14267 , n14268 );
nand ( n14270 , n14269 , n5695 );
and ( n14271 , n14266 , n14270 );
nor ( n14272 , n14265 , n14271 );
not ( n14273 , n5766 );
nand ( n14274 , n13 , n14273 );
nand ( n14275 , n14274 , n5770 );
nand ( n14276 , n13 , n834 );
not ( n14277 , n5844 );
nand ( n14278 , n14277 , n744 );
nand ( n14279 , n13269 , n5720 , n5954 );
nand ( n14280 , n16 , n14279 );
nand ( n14281 , n14276 , n14278 , n14280 );
or ( n14282 , n14275 , n14281 );
nand ( n14283 , n14282 , n793 );
nand ( n14284 , n14261 , n14272 , n14193 , n14283 );
not ( n14285 , n14284 );
or ( n14286 , n14249 , n14285 );
not ( n14287 , n846 );
not ( n14288 , n931 );
not ( n14289 , n14288 );
or ( n14290 , n14287 , n14289 );
not ( n14291 , n932 );
or ( n14292 , n14291 , n5745 );
nand ( n14293 , n14292 , n16 );
not ( n14294 , n16 );
not ( n14295 , n13 );
nand ( n14296 , n14295 , n802 );
nand ( n14297 , n14296 , n5963 , n5749 );
nand ( n14298 , n14294 , n14297 );
nand ( n14299 , n13280 , n5740 , n14293 , n14298 );
nand ( n14300 , n793 , n14299 );
nand ( n14301 , n14290 , n14300 );
or ( n14302 , n13 , n868 );
nand ( n14303 , n14302 , n960 );
nand ( n14304 , n5881 , n14303 );
nand ( n14305 , n5693 , n5831 );
nand ( n14306 , n16 , n929 , n14305 );
not ( n14307 , n921 );
nand ( n14308 , n846 , n5791 );
not ( n14309 , n14308 );
or ( n14310 , n14307 , n14309 );
not ( n14311 , n16 );
nand ( n14312 , n14310 , n14311 );
and ( n14313 , n14306 , n13239 , n14312 );
nand ( n14314 , n12 , n11 , n13 );
nor ( n14315 , n5731 , n14314 );
not ( n14316 , n14315 );
nand ( n14317 , n16 , n14182 );
and ( n14318 , n877 , n743 );
nand ( n14319 , n939 , n5704 );
nor ( n14320 , n14318 , n14319 );
nand ( n14321 , n14316 , n14317 , n14320 );
and ( n14322 , n17 , n14321 );
not ( n14323 , n17 );
not ( n14324 , n13 );
not ( n14325 , n14324 );
nand ( n14326 , n902 , n5810 );
not ( n14327 , n14326 );
or ( n14328 , n14325 , n14327 );
nand ( n14329 , n14328 , n14134 );
and ( n14330 , n14323 , n14329 );
nor ( n14331 , n14322 , n14330 );
nand ( n14332 , n14304 , n14313 , n14331 );
nand ( n14333 , n841 , n14332 );
not ( n14334 , n16 );
and ( n14335 , n14334 , n971 );
not ( n14336 , n14334 );
nor ( n14337 , n13 , n5757 );
and ( n14338 , n14336 , n14337 );
nor ( n14339 , n14335 , n14338 );
not ( n14340 , n936 );
nand ( n14341 , n14155 , n14339 , n14340 , n5718 );
nand ( n14342 , n17 , n14341 );
not ( n14343 , n16 );
nand ( n14344 , n14343 , n14315 );
nand ( n14345 , n14333 , n14342 , n14344 );
nor ( n14346 , n14301 , n14345 );
nand ( n14347 , n14286 , n14346 );
not ( n14348 , n14347 );
and ( n14349 , n14248 , n14348 );
not ( n14350 , n14248 );
and ( n14351 , n14350 , n14347 );
nor ( n14352 , n14349 , n14351 );
and ( n14353 , n71 , n5989 );
not ( n14354 , n71 );
not ( n14355 , n5989 );
and ( n14356 , n14354 , n14355 );
nor ( n14357 , n14353 , n14356 );
and ( n14358 , n14352 , n14357 );
not ( n14359 , n14352 );
not ( n14360 , n14357 );
and ( n14361 , n14359 , n14360 );
nor ( n14362 , n14358 , n14361 );
not ( n14363 , n14362 );
nand ( n14364 , n23 , n13436 );
and ( n14365 , n6208 , n14364 );
nor ( n14366 , n14365 , n25 );
not ( n14367 , n14366 );
not ( n14368 , n1825 );
not ( n14369 , n6314 );
or ( n14370 , n14368 , n14369 );
not ( n14371 , n25 );
nand ( n14372 , n14370 , n14371 );
nand ( n14373 , n6370 , n13424 );
not ( n14374 , n14373 );
nand ( n14375 , n6160 , n1956 , n14374 );
nand ( n14376 , n25 , n14375 );
nand ( n14377 , n14367 , n14372 , n14376 );
and ( n14378 , n13365 , n1868 );
or ( n14379 , n25 , n1916 );
not ( n14380 , n1907 );
nand ( n14381 , n14379 , n6277 , n14380 );
nand ( n14382 , n26 , n14381 );
nor ( n14383 , n13933 , n1984 );
not ( n14384 , n25 );
nand ( n14385 , n6317 , n6187 , n13440 );
not ( n14386 , n14385 );
or ( n14387 , n14384 , n14386 );
nand ( n14388 , n1783 , n1960 );
nand ( n14389 , n23 , n6267 );
and ( n14390 , n14388 , n14389 , n6270 );
nand ( n14391 , n14387 , n14390 );
or ( n14392 , n14383 , n14391 );
not ( n14393 , n26 );
nand ( n14394 , n14392 , n14393 );
nand ( n14395 , n14378 , n14382 , n14394 );
nor ( n14396 , n14377 , n14395 );
or ( n14397 , n14396 , n1853 );
and ( n14398 , n25 , n6453 );
not ( n14399 , n25 );
nand ( n14400 , n22 , n6210 );
and ( n14401 , n14399 , n14400 );
or ( n14402 , n14398 , n14401 );
nand ( n14403 , n14397 , n14402 );
not ( n14404 , n25 );
not ( n14405 , n14404 );
not ( n14406 , n23 );
not ( n14407 , n13451 );
nand ( n14408 , n14406 , n14407 );
nand ( n14409 , n14408 , n1953 , n1956 );
not ( n14410 , n14409 );
or ( n14411 , n14405 , n14410 );
nand ( n14412 , n6206 , n6235 );
nand ( n14413 , n14412 , n25 , n1960 );
nand ( n14414 , n14411 , n14413 );
not ( n14415 , n1799 );
not ( n14416 , n6294 );
and ( n14417 , n14415 , n14416 );
not ( n14418 , n6217 );
nor ( n14419 , n14417 , n14418 );
not ( n14420 , n14419 );
nand ( n14421 , n1888 , n1855 );
and ( n14422 , n14421 , n1921 , n14400 );
not ( n14423 , n14422 );
or ( n14424 , n14420 , n14423 );
nand ( n14425 , n14424 , n26 );
or ( n14426 , n23 , n1789 );
nand ( n14427 , n14426 , n1887 );
nand ( n14428 , n6462 , n14427 );
not ( n14429 , n26 );
not ( n14430 , n23 );
not ( n14431 , n14430 );
nand ( n14432 , n1836 , n1813 );
not ( n14433 , n14432 );
or ( n14434 , n14431 , n14433 );
nand ( n14435 , n14434 , n13903 );
nand ( n14436 , n14429 , n14435 );
nand ( n14437 , n14425 , n14428 , n14436 );
or ( n14438 , n14414 , n14437 );
nand ( n14439 , n14438 , n1853 );
not ( n14440 , n26 );
and ( n14441 , n13433 , n6296 );
or ( n14442 , n1919 , n6302 );
nand ( n14443 , n14442 , n25 );
not ( n14444 , n25 );
not ( n14445 , n23 );
nand ( n14446 , n14445 , n1933 );
nand ( n14447 , n14446 , n6342 , n6276 );
nand ( n14448 , n14444 , n14447 );
nand ( n14449 , n14441 , n14443 , n14448 );
nand ( n14450 , n14440 , n14449 );
not ( n14451 , n1944 );
not ( n14452 , n6192 );
nand ( n14453 , n1997 , n1933 );
and ( n14454 , n25 , n14453 );
not ( n14455 , n25 );
and ( n14456 , n14455 , n1900 );
or ( n14457 , n14454 , n14456 );
nand ( n14458 , n14451 , n14452 , n13873 , n14457 );
nand ( n14459 , n26 , n14458 );
nand ( n14460 , n14439 , n14450 , n14459 );
nor ( n14461 , n14403 , n14460 );
not ( n14462 , n14461 );
not ( n14463 , n6473 );
not ( n14464 , n14463 );
or ( n14465 , n14462 , n14464 );
nor ( n14466 , n14403 , n14460 );
buf ( n14467 , n14466 );
or ( n14468 , n14467 , n14070 );
nand ( n14469 , n14465 , n14468 );
not ( n14470 , n14469 );
not ( n14471 , n31 );
nand ( n14472 , n14471 , n1661 );
not ( n14473 , n14472 );
not ( n14474 , n1534 );
or ( n14475 , n14473 , n14474 );
not ( n14476 , n32 );
nand ( n14477 , n14475 , n14476 );
nand ( n14478 , n14477 , n1624 );
nand ( n14479 , n32 , n6075 );
nand ( n14480 , n14479 , n6083 , n1554 );
or ( n14481 , n14478 , n14480 );
not ( n14482 , n33 );
nand ( n14483 , n14481 , n14482 );
not ( n14484 , n1562 );
not ( n14485 , n14484 );
not ( n14486 , n1624 );
not ( n14487 , n6022 );
or ( n14488 , n14486 , n14487 );
not ( n14489 , n32 );
nand ( n14490 , n14488 , n14489 );
nand ( n14491 , n14485 , n14490 );
not ( n14492 , n14491 );
not ( n14493 , n2192 );
nand ( n14494 , n14026 , n1717 );
nor ( n14495 , n14493 , n14494 );
not ( n14496 , n14495 );
not ( n14497 , n1616 );
nand ( n14498 , n14497 , n2013 );
and ( n14499 , n32 , n14498 );
not ( n14500 , n32 );
and ( n14501 , n31 , n2077 );
not ( n14502 , n31 );
and ( n14503 , n14502 , n1588 );
or ( n14504 , n14501 , n14503 );
nand ( n14505 , n13506 , n14504 );
and ( n14506 , n14500 , n14505 );
nor ( n14507 , n14499 , n14506 );
not ( n14508 , n14507 );
or ( n14509 , n14496 , n14508 );
nand ( n14510 , n14509 , n33 );
nand ( n14511 , n14483 , n14492 , n13534 , n14510 );
not ( n14512 , n31 );
nand ( n14513 , n14512 , n13591 );
and ( n14514 , n14513 , n13602 );
not ( n14515 , n32 );
nor ( n14516 , n14514 , n14515 );
or ( n14517 , n14511 , n14516 );
nand ( n14518 , n14517 , n1673 );
not ( n14519 , n33 );
not ( n14520 , n14519 );
nand ( n14521 , n1635 , n1749 );
not ( n14522 , n14521 );
not ( n14523 , n31 );
nand ( n14524 , n14523 , n6131 );
not ( n14525 , n1634 );
not ( n14526 , n14525 );
not ( n14527 , n32 );
nand ( n14528 , n14526 , n14527 );
not ( n14529 , n1572 );
nand ( n14530 , n1629 , n14529 );
nand ( n14531 , n14522 , n14524 , n14528 , n14530 );
not ( n14532 , n14531 );
or ( n14533 , n14520 , n14532 );
not ( n14534 , n32 );
nand ( n14535 , n1712 , n1522 , n1553 , n1749 );
nand ( n14536 , n14534 , n14535 );
nand ( n14537 , n14533 , n14536 );
not ( n14538 , n14537 );
not ( n14539 , n1669 );
nand ( n14540 , n32 , n14539 );
not ( n14541 , n33 );
nand ( n14542 , n2077 , n1702 , n2101 );
nand ( n14543 , n32 , n14542 );
nand ( n14544 , n14543 , n6088 , n1654 );
not ( n14545 , n14544 );
or ( n14546 , n14541 , n14545 );
not ( n14547 , n31 );
not ( n14548 , n1522 );
nand ( n14549 , n14547 , n14548 );
nand ( n14550 , n14546 , n14549 );
not ( n14551 , n14550 );
nand ( n14552 , n14538 , n2060 , n14540 , n14551 );
nand ( n14553 , n34 , n14552 );
not ( n14554 , n33 );
not ( n14555 , n14554 );
not ( n14556 , n32 );
not ( n14557 , n14556 );
nand ( n14558 , n2056 , n2069 , n6052 );
not ( n14559 , n14558 );
or ( n14560 , n14557 , n14559 );
and ( n14561 , n6036 , n13580 );
nand ( n14562 , n14560 , n14561 );
not ( n14563 , n14562 );
or ( n14564 , n14555 , n14563 );
or ( n14565 , n31 , n6012 );
nand ( n14566 , n14565 , n14485 , n6101 );
nand ( n14567 , n2188 , n14566 );
nand ( n14568 , n14564 , n14567 );
not ( n14569 , n14568 );
not ( n14570 , n2060 );
not ( n14571 , n2091 );
not ( n14572 , n6088 );
or ( n14573 , n14571 , n14572 );
nand ( n14574 , n14573 , n31 );
not ( n14575 , n14574 );
or ( n14576 , n14570 , n14575 );
nand ( n14577 , n14576 , n1739 );
not ( n14578 , n32 );
not ( n14579 , n31 );
nand ( n14580 , n14579 , n2108 );
and ( n14581 , n14580 , n1576 );
not ( n14582 , n2039 );
nand ( n14583 , n14581 , n1493 , n14582 );
and ( n14584 , n33 , n14578 , n14583 );
not ( n14585 , n1751 );
nor ( n14586 , n14585 , n5998 );
nor ( n14587 , n14584 , n14586 );
and ( n14588 , n14577 , n14587 , n6085 , n2040 );
nand ( n14589 , n14518 , n14553 , n14569 , n14588 );
not ( n14590 , n14589 );
not ( n14591 , n14590 );
not ( n14592 , n13616 );
and ( n14593 , n14591 , n14592 );
not ( n14594 , n14589 );
and ( n14595 , n14594 , n13616 );
nor ( n14596 , n14593 , n14595 );
not ( n14597 , n14596 );
not ( n14598 , n14597 );
or ( n14599 , n14470 , n14598 );
not ( n14600 , n14589 );
not ( n14601 , n14600 );
not ( n14602 , n13489 );
and ( n14603 , n14601 , n14602 );
and ( n14604 , n14594 , n13489 );
nor ( n14605 , n14603 , n14604 );
not ( n14606 , n14605 );
not ( n14607 , n14461 );
not ( n14608 , n6473 );
and ( n14609 , n14607 , n14608 );
not ( n14610 , n6481 );
and ( n14611 , n14610 , n14461 );
nor ( n14612 , n14609 , n14611 );
not ( n14613 , n14612 );
nand ( n14614 , n14606 , n14613 );
nand ( n14615 , n14599 , n14614 );
not ( n14616 , n14615 );
nor ( n14617 , n14363 , n14616 );
or ( n14618 , n14615 , n14362 );
nand ( n14619 , n14618 , n2352 );
or ( n14620 , n14617 , n14619 );
xnor ( n14621 , n71 , n72 );
or ( n14622 , n2352 , n14621 );
nand ( n14623 , n14620 , n14622 );
xnor ( n14624 , n93 , n94 );
or ( n14625 , n2352 , n14624 );
nor ( n14626 , n13584 , n13609 );
or ( n14627 , n14626 , n1673 );
nand ( n14628 , n14627 , n13570 );
not ( n14629 , n14628 );
not ( n14630 , n13559 );
nand ( n14631 , n14629 , n14630 );
not ( n14632 , n14631 );
nor ( n14633 , n13663 , n13717 );
not ( n14634 , n14633 );
and ( n14635 , n14632 , n14634 );
and ( n14636 , n14633 , n14631 );
nor ( n14637 , n14635 , n14636 );
or ( n14638 , n14637 , n14469 );
nand ( n14639 , n14637 , n14612 );
nand ( n14640 , n14638 , n14639 );
not ( n14641 , n5989 );
not ( n14642 , n14641 );
xor ( n14643 , n93 , n14642 );
not ( n14644 , n14643 );
and ( n14645 , n14640 , n14644 );
not ( n14646 , n14640 );
and ( n14647 , n14646 , n14643 );
nor ( n14648 , n14645 , n14647 );
nand ( n14649 , n14648 , n2352 );
nand ( n14650 , n14625 , n14649 );
not ( n14651 , n69 );
and ( n14652 , n97 , n14651 );
not ( n14653 , n97 );
and ( n14654 , n14653 , n69 );
nor ( n14655 , n14652 , n14654 );
or ( n14656 , n2352 , n14655 );
not ( n14657 , n14248 );
not ( n14658 , n14590 );
and ( n14659 , n14657 , n14658 );
buf ( n14660 , n13219 );
not ( n14661 , n14660 );
and ( n14662 , n14661 , n14594 );
nor ( n14663 , n14659 , n14662 );
not ( n14664 , n14651 );
not ( n14665 , n13350 );
not ( n14666 , n14665 );
and ( n14667 , n14664 , n14666 );
and ( n14668 , n14651 , n13354 );
nor ( n14669 , n14667 , n14668 );
not ( n14670 , n14669 );
and ( n14671 , n14663 , n14670 );
not ( n14672 , n14663 );
and ( n14673 , n14672 , n14669 );
nor ( n14674 , n14671 , n14673 );
not ( n14675 , n14674 );
not ( n14676 , n13613 );
not ( n14677 , n2210 );
and ( n14678 , n14676 , n14677 );
and ( n14679 , n13613 , n2340 );
nor ( n14680 , n14678 , n14679 );
and ( n14681 , n14680 , n14469 );
not ( n14682 , n14680 );
and ( n14683 , n14682 , n14613 );
nor ( n14684 , n14681 , n14683 );
not ( n14685 , n14684 );
nand ( n14686 , n14675 , n14685 );
nand ( n14687 , n14684 , n14674 );
nand ( n14688 , n14686 , n2352 , n14687 );
nand ( n14689 , n14656 , n14688 );
not ( n14690 , n232 );
and ( n14691 , n233 , n14690 );
not ( n14692 , n233 );
and ( n14693 , n14692 , n232 );
nor ( n14694 , n14691 , n14693 );
or ( n14695 , n2352 , n14694 );
not ( n14696 , n4406 );
and ( n14697 , n4471 , n4531 , n4571 , n14696 );
and ( n14698 , n9996 , n14697 );
not ( n14699 , n9996 );
not ( n14700 , n4572 );
not ( n14701 , n14700 );
and ( n14702 , n14699 , n14701 );
nor ( n14703 , n14698 , n14702 );
not ( n14704 , n14690 );
not ( n14705 , n10164 );
or ( n14706 , n14704 , n14705 );
buf ( n14707 , n10163 );
or ( n14708 , n14707 , n14690 );
nand ( n14709 , n14706 , n14708 );
not ( n14710 , n14709 );
and ( n14711 , n14703 , n14710 );
not ( n14712 , n14703 );
and ( n14713 , n14712 , n14709 );
nor ( n14714 , n14711 , n14713 );
not ( n14715 , n14714 );
not ( n14716 , n10313 );
not ( n14717 , n5673 );
or ( n14718 , n14716 , n14717 );
or ( n14719 , n10313 , n5673 );
nand ( n14720 , n14718 , n14719 );
not ( n14721 , n14720 );
nand ( n14722 , n14715 , n14721 );
nand ( n14723 , n14714 , n14720 );
nand ( n14724 , n14722 , n2352 , n14723 );
nand ( n14725 , n14695 , n14724 );
not ( n14726 , n242 );
and ( n14727 , n243 , n14726 );
not ( n14728 , n243 );
and ( n14729 , n14728 , n242 );
nor ( n14730 , n14727 , n14729 );
or ( n14731 , n2352 , n14730 );
nand ( n14732 , n12299 , n12222 , n12250 , n12220 );
not ( n14733 , n14732 );
not ( n14734 , n14733 );
not ( n14735 , n4054 );
not ( n14736 , n159 );
not ( n14737 , n4086 );
nand ( n14738 , n10129 , n10148 , n14737 );
nand ( n14739 , n14736 , n14738 );
not ( n14740 , n9986 );
nand ( n14741 , n14739 , n14740 , n12704 );
not ( n14742 , n14741 );
or ( n14743 , n14735 , n14742 );
not ( n14744 , n10087 );
not ( n14745 , n158 );
not ( n14746 , n9928 );
nand ( n14747 , n14745 , n14746 );
nand ( n14748 , n14747 , n12739 , n9833 );
not ( n14749 , n14748 );
or ( n14750 , n14744 , n14749 );
and ( n14751 , n9987 , n10123 );
nand ( n14752 , n14750 , n14751 );
not ( n14753 , n160 );
not ( n14754 , n159 );
not ( n14755 , n14754 );
nor ( n14756 , n9898 , n4275 );
not ( n14757 , n158 );
nand ( n14758 , n14757 , n4287 );
nand ( n14759 , n14756 , n14758 , n10121 );
not ( n14760 , n14759 );
or ( n14761 , n14755 , n14760 );
nand ( n14762 , n9866 , n4049 );
nand ( n14763 , n14761 , n14762 );
not ( n14764 , n14763 );
or ( n14765 , n14753 , n14764 );
not ( n14766 , n10141 );
not ( n14767 , n14766 );
not ( n14768 , n14767 );
not ( n14769 , n4227 );
not ( n14770 , n9992 );
or ( n14771 , n14769 , n14770 );
nand ( n14772 , n14771 , n158 );
not ( n14773 , n14772 );
or ( n14774 , n14768 , n14773 );
nand ( n14775 , n14774 , n10024 );
nand ( n14776 , n14765 , n14775 );
nor ( n14777 , n14752 , n14776 );
nand ( n14778 , n14743 , n14777 );
not ( n14779 , n14778 );
nand ( n14780 , n9937 , n4220 );
nand ( n14781 , n4064 , n10042 );
not ( n14782 , n9935 );
not ( n14783 , n159 );
nand ( n14784 , n14782 , n14783 );
not ( n14785 , n158 );
not ( n14786 , n9839 );
nand ( n14787 , n14785 , n14786 );
nand ( n14788 , n14781 , n14784 , n14787 );
nor ( n14789 , n14780 , n14788 );
or ( n14790 , n160 , n14789 );
nand ( n14791 , n14790 , n14767 );
not ( n14792 , n14791 );
or ( n14793 , n4268 , n10873 , n9857 );
nand ( n14794 , n14793 , n159 );
nand ( n14795 , n14794 , n9992 , n9843 );
nand ( n14796 , n160 , n14795 );
not ( n14797 , n159 );
or ( n14798 , n14797 , n4272 );
not ( n14799 , n159 );
not ( n14800 , n14799 );
nor ( n14801 , n10878 , n10113 );
not ( n14802 , n158 );
nand ( n14803 , n14802 , n4154 );
nand ( n14804 , n14801 , n14803 , n4220 );
not ( n14805 , n14804 );
or ( n14806 , n14800 , n14805 );
not ( n14807 , n158 );
nand ( n14808 , n14807 , n10113 );
nand ( n14809 , n14806 , n14808 );
not ( n14810 , n14809 );
nand ( n14811 , n14792 , n14796 , n14798 , n14810 );
nand ( n14812 , n161 , n14811 );
nand ( n14813 , n10862 , n9813 );
not ( n14814 , n4264 );
not ( n14815 , n4041 );
nand ( n14816 , n159 , n14815 );
not ( n14817 , n4043 );
nand ( n14818 , n14817 , n9911 );
not ( n14819 , n14818 );
or ( n14820 , n9812 , n14819 );
not ( n14821 , n159 );
nand ( n14822 , n14820 , n14821 );
nand ( n14823 , n14814 , n14816 , n14822 );
nor ( n14824 , n14813 , n14823 );
or ( n14825 , n160 , n14824 );
nand ( n14826 , n4148 , n4080 );
and ( n14827 , n12819 , n14826 );
nand ( n14828 , n14825 , n14827 );
not ( n14829 , n12722 );
and ( n14830 , n158 , n4268 );
not ( n14831 , n158 );
and ( n14832 , n14831 , n4089 );
nor ( n14833 , n14830 , n14832 );
not ( n14834 , n14833 );
or ( n14835 , n14829 , n14834 );
not ( n14836 , n159 );
nand ( n14837 , n14835 , n14836 );
not ( n14838 , n12758 );
not ( n14839 , n10069 );
or ( n14840 , n14838 , n14839 );
nand ( n14841 , n14840 , n159 );
and ( n14842 , n4036 , n10093 );
nand ( n14843 , n14837 , n14841 , n4283 , n14842 );
nand ( n14844 , n160 , n14843 );
not ( n14845 , n159 );
nand ( n14846 , n14845 , n4264 );
not ( n14847 , n157 );
nand ( n14848 , n14847 , n14817 );
not ( n14849 , n158 );
nand ( n14850 , n14849 , n9890 );
nand ( n14851 , n14848 , n14850 );
and ( n14852 , n159 , n14851 );
nor ( n14853 , n14852 , n12738 );
nand ( n14854 , n14844 , n14846 , n14853 );
or ( n14855 , n14828 , n14854 );
nand ( n14856 , n14855 , n4144 );
nand ( n14857 , n14779 , n14812 , n14856 );
not ( n14858 , n14857 );
not ( n14859 , n14858 );
or ( n14860 , n14734 , n14859 );
not ( n14861 , n14732 );
not ( n14862 , n14778 );
nand ( n14863 , n14862 , n14812 , n14856 );
not ( n14864 , n14863 );
or ( n14865 , n14861 , n14864 );
nand ( n14866 , n14860 , n14865 );
and ( n14867 , n14866 , n242 );
not ( n14868 , n14866 );
and ( n14869 , n14868 , n14726 );
nor ( n14870 , n14867 , n14869 );
not ( n14871 , n14870 );
not ( n14872 , n5339 );
or ( n14873 , n166 , n14872 );
nor ( n14874 , n166 , n5318 );
not ( n14875 , n14874 );
not ( n14876 , n5396 );
not ( n14877 , n14876 );
not ( n14878 , n14877 );
nand ( n14879 , n14873 , n14875 , n14878 );
nand ( n14880 , n5478 , n14879 );
not ( n14881 , n166 );
or ( n14882 , n14881 , n5605 );
nand ( n14883 , n14882 , n5573 , n5473 );
nand ( n14884 , n5379 , n14883 );
and ( n14885 , n14880 , n14884 );
not ( n14886 , n167 );
not ( n14887 , n14886 );
not ( n14888 , n10251 );
and ( n14889 , n14887 , n14888 );
nand ( n14890 , n5570 , n5541 );
nor ( n14891 , n166 , n5216 );
not ( n14892 , n14891 );
nand ( n14893 , n14892 , n5374 );
nor ( n14894 , n14890 , n14893 );
or ( n14895 , n167 , n14894 );
or ( n14896 , n166 , n5541 );
nand ( n14897 , n14895 , n14896 );
nor ( n14898 , n14889 , n14897 );
not ( n14899 , n14898 );
not ( n14900 , n5650 );
not ( n14901 , n5438 );
or ( n14902 , n14900 , n14901 );
nand ( n14903 , n14902 , n169 );
not ( n14904 , n5223 );
not ( n14905 , n10772 );
or ( n14906 , n14904 , n14905 , n5557 );
nand ( n14907 , n14906 , n5379 );
nand ( n14908 , n14903 , n14907 );
not ( n14909 , n5400 );
nand ( n14910 , n5259 , n14909 );
not ( n14911 , n166 );
not ( n14912 , n14911 );
not ( n14913 , n5434 );
or ( n14914 , n14912 , n14913 );
not ( n14915 , n167 );
not ( n14916 , n5257 );
and ( n14917 , n14915 , n14916 );
and ( n14918 , n5338 , n5596 );
nor ( n14919 , n14917 , n14918 );
nand ( n14920 , n14914 , n14919 );
nor ( n14921 , n14910 , n14920 );
or ( n14922 , n169 , n14921 );
nand ( n14923 , n14922 , n5573 );
nor ( n14924 , n14908 , n14923 );
not ( n14925 , n14924 );
or ( n14926 , n14899 , n14925 );
nand ( n14927 , n14926 , n170 );
not ( n14928 , n5303 );
nor ( n14929 , n5411 , n14928 );
and ( n14930 , n169 , n14929 );
not ( n14931 , n169 );
nor ( n14932 , n5337 , n5539 );
not ( n14933 , n14932 );
nand ( n14934 , n5340 , n14933 );
and ( n14935 , n14931 , n14934 );
nor ( n14936 , n14930 , n14935 );
nand ( n14937 , n5522 , n5332 , n5369 );
nand ( n14938 , n5355 , n14937 );
nand ( n14939 , n5220 , n5310 );
not ( n14940 , n166 );
not ( n14941 , n5611 );
nand ( n14942 , n14940 , n14941 );
nand ( n14943 , n14939 , n14942 , n10258 , n5504 );
nand ( n14944 , n10183 , n14943 );
and ( n14945 , n14936 , n14938 , n14944 );
and ( n14946 , n14945 , n5361 , n5506 );
not ( n14947 , n169 );
not ( n14948 , n14947 );
not ( n14949 , n167 );
or ( n14950 , n14949 , n5284 );
nand ( n14951 , n14950 , n10708 );
not ( n14952 , n14951 );
or ( n14953 , n14948 , n14952 );
not ( n14954 , n166 );
not ( n14955 , n14954 );
nor ( n14956 , n163 , n165 );
not ( n14957 , n14956 );
or ( n14958 , n14955 , n14957 );
not ( n14959 , n166 );
nand ( n14960 , n14959 , n5484 );
nand ( n14961 , n14958 , n14960 );
nand ( n14962 , n167 , n14961 );
nand ( n14963 , n14953 , n14962 );
not ( n14964 , n14963 );
not ( n14965 , n10253 );
not ( n14966 , n5237 );
or ( n14967 , n14965 , n14966 );
not ( n14968 , n167 );
nand ( n14969 , n14967 , n14968 );
and ( n14970 , n14964 , n14875 , n14969 );
not ( n14971 , n169 );
not ( n14972 , n14971 );
not ( n14973 , n10704 );
not ( n14974 , n166 );
nand ( n14975 , n14974 , n5472 );
not ( n14976 , n14975 );
or ( n14977 , n14973 , n14976 );
not ( n14978 , n167 );
nand ( n14979 , n14977 , n14978 );
nand ( n14980 , n14979 , n10253 , n5357 );
not ( n14981 , n14980 );
or ( n14982 , n14972 , n14981 );
nand ( n14983 , n167 , n14932 );
nand ( n14984 , n14982 , n14983 );
not ( n14985 , n14984 );
not ( n14986 , n169 );
not ( n14987 , n165 );
nand ( n14988 , n14987 , n10685 );
not ( n14989 , n14988 );
and ( n14990 , n166 , n5557 );
not ( n14991 , n166 );
and ( n14992 , n14991 , n10693 );
nor ( n14993 , n14990 , n14992 );
not ( n14994 , n14993 );
or ( n14995 , n14989 , n14994 );
not ( n14996 , n167 );
nand ( n14997 , n14995 , n14996 );
not ( n14998 , n5649 );
nor ( n14999 , n14998 , n10281 );
nand ( n15000 , n14997 , n5485 , n14999 );
not ( n15001 , n15000 );
or ( n15002 , n14986 , n15001 );
not ( n15003 , n5290 );
not ( n15004 , n15003 );
not ( n15005 , n5533 );
or ( n15006 , n15004 , n15005 );
nand ( n15007 , n15006 , n5379 );
nand ( n15008 , n15002 , n15007 );
not ( n15009 , n15008 );
nand ( n15010 , n14970 , n14985 , n15009 );
nand ( n15011 , n5449 , n15010 );
nand ( n15012 , n14885 , n14927 , n14946 , n15011 );
not ( n15013 , n15012 );
not ( n15014 , n15013 );
or ( n15015 , n12135 , n12117 );
nand ( n15016 , n15015 , n178 );
and ( n15017 , n12100 , n12157 , n15016 );
and ( n15018 , n10793 , n15017 );
not ( n15019 , n10793 );
not ( n15020 , n15017 );
and ( n15021 , n15019 , n15020 );
nor ( n15022 , n15018 , n15021 );
not ( n15023 , n15022 );
not ( n15024 , n15023 );
or ( n15025 , n15014 , n15024 );
not ( n15026 , n15013 );
nand ( n15027 , n15026 , n15022 );
nand ( n15028 , n15025 , n15027 );
not ( n15029 , n15028 );
nand ( n15030 , n14871 , n15029 );
nand ( n15031 , n14870 , n15028 );
nand ( n15032 , n15030 , n2352 , n15031 );
nand ( n15033 , n14731 , n15032 );
not ( n15034 , n250 );
not ( n15035 , n7317 );
not ( n15036 , n15035 );
or ( n15037 , n15034 , n15036 );
not ( n15038 , n7317 );
or ( n15039 , n250 , n15038 );
nand ( n15040 , n15037 , n15039 );
not ( n15041 , n142 );
nand ( n15042 , n15041 , n11429 );
nand ( n15043 , n6757 , n11430 );
nand ( n15044 , n11453 , n6657 );
or ( n15045 , n15043 , n15044 );
not ( n15046 , n141 );
nand ( n15047 , n15045 , n15046 );
nand ( n15048 , n6751 , n15042 , n15047 );
not ( n15049 , n15048 );
nand ( n15050 , n141 , n11947 );
not ( n15051 , n144 );
nand ( n15052 , n142 , n140 , n11334 );
and ( n15053 , n15052 , n6657 );
or ( n15054 , n141 , n11286 );
not ( n15055 , n142 );
nand ( n15056 , n15055 , n11250 );
nand ( n15057 , n15053 , n11288 , n15054 , n15056 );
and ( n15058 , n15051 , n15057 );
nand ( n15059 , n11298 , n11964 , n6685 );
nand ( n15060 , n141 , n15059 );
and ( n15061 , n15060 , n11489 , n11393 );
not ( n15062 , n144 );
nor ( n15063 , n15061 , n15062 );
nor ( n15064 , n15058 , n15063 );
nand ( n15065 , n137 , n15049 , n15050 , n15064 );
not ( n15066 , n11341 );
nand ( n15067 , n6588 , n11506 );
not ( n15068 , n15067 );
or ( n15069 , n15066 , n15068 );
nand ( n15070 , n15069 , n141 );
and ( n15071 , n6808 , n15070 );
nand ( n15072 , n142 , n11429 );
not ( n15073 , n15072 );
nand ( n15074 , n15073 , n141 );
nand ( n15075 , n6702 , n6647 );
not ( n15076 , n15075 );
not ( n15077 , n11317 );
not ( n15078 , n15077 );
not ( n15079 , n11419 );
or ( n15080 , n15078 , n15079 );
nand ( n15081 , n15080 , n141 );
not ( n15082 , n140 );
nand ( n15083 , n15082 , n11247 );
not ( n15084 , n15083 );
not ( n15085 , n142 );
and ( n15086 , n15085 , n6562 );
not ( n15087 , n15085 );
and ( n15088 , n15087 , n6684 );
nor ( n15089 , n15086 , n15088 );
not ( n15090 , n15089 );
or ( n15091 , n15084 , n15090 );
not ( n15092 , n141 );
nand ( n15093 , n15091 , n15092 );
nand ( n15094 , n11561 , n15076 , n15081 , n15093 );
and ( n15095 , n144 , n15094 );
not ( n15096 , n11343 );
nor ( n15097 , n15095 , n15096 );
not ( n15098 , n6690 );
not ( n15099 , n11294 );
or ( n15100 , n15098 , n15099 );
not ( n15101 , n141 );
nand ( n15102 , n15100 , n15101 );
not ( n15103 , n15102 );
nor ( n15104 , n11998 , n11259 );
nand ( n15105 , n141 , n6644 );
not ( n15106 , n140 );
nor ( n15107 , n15106 , n11281 );
nor ( n15108 , n6640 , n6749 );
or ( n15109 , n15107 , n15108 );
not ( n15110 , n141 );
nand ( n15111 , n15109 , n15110 );
and ( n15112 , n15105 , n6690 , n15111 );
and ( n15113 , n15104 , n15112 );
nor ( n15114 , n15113 , n144 );
nor ( n15115 , n15103 , n15114 );
nand ( n15116 , n15071 , n15074 , n15097 , n15115 );
nand ( n15117 , n15065 , n15116 );
not ( n15118 , n11555 );
or ( n15119 , n142 , n6696 );
nand ( n15120 , n15119 , n11343 , n11369 );
not ( n15121 , n15120 );
or ( n15122 , n15118 , n15121 );
nand ( n15123 , n15122 , n11262 );
not ( n15124 , n6751 );
not ( n15125 , n6664 );
not ( n15126 , n11489 );
or ( n15127 , n15125 , n15126 );
nand ( n15128 , n15127 , n142 );
not ( n15129 , n15128 );
or ( n15130 , n15124 , n15129 );
nand ( n15131 , n15130 , n11498 );
not ( n15132 , n11447 );
not ( n15133 , n142 );
not ( n15134 , n15133 );
not ( n15135 , n6705 );
or ( n15136 , n15134 , n15135 );
nand ( n15137 , n15136 , n6695 );
not ( n15138 , n140 );
and ( n15139 , n15138 , n11534 );
nor ( n15140 , n15132 , n15137 , n15139 );
or ( n15141 , n141 , n15140 );
not ( n15142 , n11559 );
nand ( n15143 , n6544 , n15142 );
nand ( n15144 , n15141 , n15143 );
nand ( n15145 , n144 , n15144 );
nand ( n15146 , n11449 , n15131 , n15145 );
nor ( n15147 , n15123 , n15146 );
not ( n15148 , n144 );
not ( n15149 , n141 );
not ( n15150 , n15149 );
nand ( n15151 , n11440 , n11345 , n6611 );
not ( n15152 , n15151 );
or ( n15153 , n15150 , n15152 );
and ( n15154 , n6708 , n15072 );
nand ( n15155 , n15153 , n15154 );
nand ( n15156 , n15148 , n15155 );
nand ( n15157 , n15117 , n15147 , n15156 );
not ( n15158 , n15157 );
not ( n15159 , n134 );
not ( n15160 , n132 );
not ( n15161 , n15160 );
not ( n15162 , n7290 );
or ( n15163 , n15161 , n15162 );
not ( n15164 , n133 );
nand ( n15165 , n15164 , n6840 , n6987 );
nand ( n15166 , n15163 , n15165 );
nand ( n15167 , n15159 , n15166 );
or ( n15168 , n6968 , n6863 );
not ( n15169 , n133 );
or ( n15170 , n15169 , n7309 );
not ( n15171 , n6989 );
not ( n15172 , n15171 );
not ( n15173 , n15172 );
nand ( n15174 , n15168 , n15170 , n15173 );
not ( n15175 , n7203 );
not ( n15176 , n6876 );
not ( n15177 , n15176 );
nor ( n15178 , n15177 , n6839 );
or ( n15179 , n15174 , n15175 , n15178 );
nand ( n15180 , n15179 , n134 );
not ( n15181 , n133 );
nor ( n15182 , n128 , n129 );
not ( n15183 , n15182 );
not ( n15184 , n15183 );
buf ( n15185 , n7013 );
nand ( n15186 , n15184 , n15185 );
nand ( n15187 , n6934 , n15186 );
and ( n15188 , n15181 , n15187 );
not ( n15189 , n7178 );
not ( n15190 , n6951 );
not ( n15191 , n15190 );
or ( n15192 , n132 , n15191 );
nand ( n15193 , n15192 , n6967 );
not ( n15194 , n15193 );
or ( n15195 , n15189 , n15194 );
not ( n15196 , n6887 );
not ( n15197 , n15196 );
nand ( n15198 , n6864 , n15197 );
nand ( n15199 , n15195 , n15198 );
not ( n15200 , n7284 );
not ( n15201 , n15200 );
and ( n15202 , n7169 , n15201 );
not ( n15203 , n132 );
not ( n15204 , n131 );
nand ( n15205 , n15204 , n133 );
nor ( n15206 , n15202 , n15203 , n15205 );
nor ( n15207 , n15188 , n15199 , n15206 );
and ( n15208 , n15167 , n15180 , n15207 );
nor ( n15209 , n15208 , n135 );
not ( n15210 , n15209 );
not ( n15211 , n130 );
nand ( n15212 , n15211 , n15185 );
not ( n15213 , n15212 );
not ( n15214 , n6869 );
not ( n15215 , n15214 );
nand ( n15216 , n15213 , n133 , n15215 );
not ( n15217 , n6996 );
buf ( n15218 , n6820 );
nand ( n15219 , n15185 , n15218 );
not ( n15220 , n133 );
not ( n15221 , n6954 );
and ( n15222 , n15220 , n15221 );
not ( n15223 , n15220 );
nor ( n15224 , n132 , n6913 );
and ( n15225 , n15223 , n15224 );
nor ( n15226 , n15222 , n15225 );
not ( n15227 , n7305 );
nand ( n15228 , n15227 , n132 );
nand ( n15229 , n15217 , n15219 , n15226 , n15228 );
nand ( n15230 , n134 , n15229 );
nand ( n15231 , n15216 , n15230 );
not ( n15232 , n133 );
not ( n15233 , n15232 );
not ( n15234 , n15178 );
or ( n15235 , n15233 , n15234 );
not ( n15236 , n134 );
nand ( n15237 , n15185 , n6916 );
nand ( n15238 , n7014 , n15237 );
and ( n15239 , n133 , n15238 );
not ( n15240 , n133 );
not ( n15241 , n132 );
nand ( n15242 , n15241 , n7004 );
nand ( n15243 , n15185 , n15200 );
nand ( n15244 , n15242 , n7259 , n15243 );
and ( n15245 , n15240 , n15244 );
nor ( n15246 , n15239 , n15245 );
not ( n15247 , n7129 );
nand ( n15248 , n132 , n15247 );
not ( n15249 , n15248 );
nand ( n15250 , n15249 , n133 );
not ( n15251 , n133 );
nand ( n15252 , n15251 , n6983 );
nand ( n15253 , n15246 , n15250 , n15252 );
nand ( n15254 , n15236 , n15253 );
nand ( n15255 , n15235 , n15254 );
nor ( n15256 , n15231 , n15255 );
not ( n15257 , n133 );
not ( n15258 , n15257 );
or ( n15259 , n130 , n6872 );
nand ( n15260 , n132 , n7229 );
nand ( n15261 , n15259 , n15260 );
not ( n15262 , n15261 );
or ( n15263 , n15258 , n15262 );
nor ( n15264 , n131 , n6922 );
nand ( n15265 , n132 , n15264 );
nand ( n15266 , n15265 , n7121 );
nand ( n15267 , n6817 , n6873 );
not ( n15268 , n6865 );
nand ( n15269 , n15268 , n7302 );
not ( n15270 , n7153 );
not ( n15271 , n15270 );
not ( n15272 , n132 );
nand ( n15273 , n15272 , n15218 );
nand ( n15274 , n15271 , n7220 , n15273 );
nand ( n15275 , n133 , n15274 );
nand ( n15276 , n15267 , n15269 , n15275 );
or ( n15277 , n15266 , n15276 );
not ( n15278 , n134 );
nand ( n15279 , n15277 , n15278 );
nand ( n15280 , n15263 , n15279 );
not ( n15281 , n132 );
not ( n15282 , n6980 );
nand ( n15283 , n15281 , n15282 );
and ( n15284 , n15283 , n6891 );
or ( n15285 , n133 , n15214 );
nand ( n15286 , n15285 , n6913 , n6958 );
nand ( n15287 , n134 , n15286 );
not ( n15288 , n133 );
nand ( n15289 , n15288 , n7038 , n7209 );
not ( n15290 , n6890 );
and ( n15291 , n133 , n7139 , n15290 );
buf ( n15292 , n15248 );
nand ( n15293 , n15291 , n6929 , n15292 );
nand ( n15294 , n15289 , n15293 );
nand ( n15295 , n15284 , n15287 , n15294 );
or ( n15296 , n15280 , n15295 );
nand ( n15297 , n15296 , n135 );
nand ( n15298 , n15210 , n15256 , n15297 );
not ( n15299 , n15298 );
and ( n15300 , n15158 , n15299 );
not ( n15301 , n15158 );
not ( n15302 , n15299 );
and ( n15303 , n15301 , n15302 );
nor ( n15304 , n15300 , n15303 );
xnor ( n15305 , n15040 , n15304 );
not ( n15306 , n15305 );
not ( n15307 , n7735 );
nor ( n15308 , n8007 , n15307 );
or ( n15309 , n121 , n15308 );
not ( n15310 , n7685 );
nand ( n15311 , n15309 , n15310 );
nand ( n15312 , n126 , n15311 );
not ( n15313 , n7948 );
or ( n15314 , n121 , n7695 );
nand ( n15315 , n15314 , n8186 );
nand ( n15316 , n15313 , n15315 );
not ( n15317 , n126 );
not ( n15318 , n124 );
nor ( n15319 , n15318 , n123 );
nand ( n15320 , n15319 , n121 );
nor ( n15321 , n7642 , n15320 );
not ( n15322 , n15321 );
not ( n15323 , n7755 );
nand ( n15324 , n15323 , n7813 );
and ( n15325 , n15324 , n7811 , n8058 );
nand ( n15326 , n7992 , n7814 );
nand ( n15327 , n15322 , n15325 , n15326 );
nand ( n15328 , n15317 , n15327 );
nand ( n15329 , n15312 , n15316 , n15328 );
not ( n15330 , n120 );
not ( n15331 , n15330 );
not ( n15332 , n121 );
not ( n15333 , n8060 );
nand ( n15334 , n15332 , n15333 );
nand ( n15335 , n15334 , n8158 , n8160 );
not ( n15336 , n15335 );
or ( n15337 , n15331 , n15336 );
nand ( n15338 , n7797 , n7975 );
nand ( n15339 , n15338 , n120 , n8175 );
nand ( n15340 , n15337 , n15339 );
or ( n15341 , n15329 , n15340 );
nand ( n15342 , n15341 , n7748 );
not ( n15343 , n120 );
nand ( n15344 , n121 , n122 );
nor ( n15345 , n125 , n15344 );
nand ( n15346 , n15345 , n7681 );
or ( n15347 , n15343 , n15346 );
nand ( n15348 , n8175 , n8066 );
and ( n15349 , n15347 , n15348 );
not ( n15350 , n15349 );
not ( n15351 , n7634 );
nand ( n15352 , n15351 , n7874 );
nand ( n15353 , n8204 , n15352 );
and ( n15354 , n120 , n15353 );
not ( n15355 , n120 );
not ( n15356 , n121 );
not ( n15357 , n8165 );
nand ( n15358 , n15356 , n15357 );
nand ( n15359 , n15358 , n7834 , n7863 );
and ( n15360 , n15355 , n15359 );
nor ( n15361 , n15354 , n15360 );
not ( n15362 , n15361 );
or ( n15363 , n15350 , n15362 );
nand ( n15364 , n15363 , n126 );
not ( n15365 , n120 );
not ( n15366 , n7941 );
or ( n15367 , n15365 , n15366 );
or ( n15368 , n120 , n15321 );
nand ( n15369 , n15367 , n15368 );
nand ( n15370 , n15342 , n15364 , n15369 );
not ( n15371 , n15370 );
not ( n15372 , n127 );
not ( n15373 , n120 );
not ( n15374 , n15373 );
nand ( n15375 , n7647 , n8092 );
not ( n15376 , n15375 );
or ( n15377 , n15374 , n15376 );
not ( n15378 , n120 );
not ( n15379 , n121 );
nor ( n15380 , n124 , n125 );
not ( n15381 , n15380 );
or ( n15382 , n15379 , n15381 );
not ( n15383 , n123 );
nor ( n15384 , n15383 , n122 );
nand ( n15385 , n121 , n15384 );
nand ( n15386 , n15382 , n15385 );
and ( n15387 , n15378 , n15386 );
not ( n15388 , n15378 );
nand ( n15389 , n8017 , n15346 );
not ( n15390 , n15389 );
nand ( n15391 , n15390 , n8228 , n8160 );
and ( n15392 , n15388 , n15391 );
nor ( n15393 , n15387 , n15392 );
nand ( n15394 , n15377 , n15393 );
not ( n15395 , n15394 );
nor ( n15396 , n121 , n7759 );
not ( n15397 , n15396 );
and ( n15398 , n15397 , n7841 );
nand ( n15399 , n7813 , n7824 );
nand ( n15400 , n7642 , n121 , n7659 );
nand ( n15401 , n121 , n7717 );
and ( n15402 , n15400 , n15401 , n7930 );
not ( n15403 , n7860 );
not ( n15404 , n121 );
not ( n15405 , n7668 );
nand ( n15406 , n15404 , n15405 );
nand ( n15407 , n125 , n7661 );
nand ( n15408 , n15403 , n15406 , n15407 );
nand ( n15409 , n120 , n15408 );
nand ( n15410 , n15399 , n15402 , n15409 );
and ( n15411 , n126 , n15410 );
not ( n15412 , n126 );
or ( n15413 , n120 , n7739 );
nand ( n15414 , n125 , n15357 );
nand ( n15415 , n15413 , n8182 , n15414 );
and ( n15416 , n15412 , n15415 );
nor ( n15417 , n15411 , n15416 );
nand ( n15418 , n15395 , n15398 , n15417 );
not ( n15419 , n15418 );
or ( n15420 , n15372 , n15419 );
not ( n15421 , n120 );
and ( n15422 , n15421 , n7921 );
not ( n15423 , n15421 );
nand ( n15424 , n7670 , n15357 );
and ( n15425 , n15423 , n15424 );
nor ( n15426 , n15422 , n15425 );
nor ( n15427 , n15426 , n8235 );
not ( n15428 , n8215 );
nand ( n15429 , n15427 , n7723 , n15428 );
not ( n15430 , n126 );
nand ( n15431 , n15429 , n15430 );
nand ( n15432 , n15420 , n15431 );
not ( n15433 , n15432 );
nand ( n15434 , n15371 , n15433 );
not ( n15435 , n8100 );
and ( n15436 , n15434 , n15435 );
not ( n15437 , n15434 );
not ( n15438 , n8099 );
not ( n15439 , n15438 );
not ( n15440 , n15439 );
and ( n15441 , n15437 , n15440 );
nor ( n15442 , n15436 , n15441 );
not ( n15443 , n15442 );
not ( n15444 , n7748 );
nor ( n15445 , n7897 , n8226 );
not ( n15446 , n15445 );
not ( n15447 , n15414 );
not ( n15448 , n121 );
nand ( n15449 , n15448 , n8101 );
not ( n15450 , n15449 );
or ( n15451 , n15447 , n15450 );
not ( n15452 , n120 );
nand ( n15453 , n15451 , n15452 );
not ( n15454 , n15453 );
or ( n15455 , n15446 , n15454 );
nand ( n15456 , n15455 , n126 );
not ( n15457 , n8160 );
not ( n15458 , n7898 );
or ( n15459 , n15457 , n15458 );
not ( n15460 , n120 );
nand ( n15461 , n15459 , n15460 );
not ( n15462 , n120 );
not ( n15463 , n7663 );
or ( n15464 , n15462 , n15463 );
nand ( n15465 , n7751 , n7814 );
nand ( n15466 , n15464 , n15465 );
nand ( n15467 , n126 , n15466 );
and ( n15468 , n15461 , n15467 );
not ( n15469 , n7924 );
or ( n15470 , n7692 , n15469 );
nand ( n15471 , n15470 , n8050 );
nand ( n15472 , n8200 , n15471 );
not ( n15473 , n120 );
not ( n15474 , n121 );
not ( n15475 , n15474 );
not ( n15476 , n15380 );
or ( n15477 , n15475 , n15476 );
nand ( n15478 , n15477 , n15406 );
not ( n15479 , n15478 );
or ( n15480 , n15473 , n15479 );
nand ( n15481 , n15480 , n15347 );
nor ( n15482 , n15472 , n15481 );
not ( n15483 , n126 );
not ( n15484 , n8060 );
not ( n15485 , n121 );
not ( n15486 , n7624 );
and ( n15487 , n15485 , n15486 );
not ( n15488 , n15485 );
and ( n15489 , n15488 , n7891 );
nor ( n15490 , n15487 , n15489 );
not ( n15491 , n15490 );
or ( n15492 , n15484 , n15491 );
not ( n15493 , n120 );
nand ( n15494 , n15492 , n15493 );
not ( n15495 , n7868 );
nor ( n15496 , n15495 , n7655 );
nand ( n15497 , n15494 , n7954 , n15496 );
nand ( n15498 , n15483 , n15497 );
nand ( n15499 , n15456 , n15468 , n15482 , n15498 );
not ( n15500 , n15499 );
or ( n15501 , n15444 , n15500 );
not ( n15502 , n126 );
and ( n15503 , n15502 , n7972 , n8181 );
nand ( n15504 , n15346 , n8212 );
and ( n15505 , n126 , n15504 );
nor ( n15506 , n15503 , n15505 );
not ( n15507 , n8017 );
not ( n15508 , n8029 );
nor ( n15509 , n15507 , n15508 );
nand ( n15510 , n7671 , n15509 );
nand ( n15511 , n8223 , n15510 );
not ( n15512 , n8229 );
and ( n15513 , n15506 , n15511 , n15512 , n7995 );
nand ( n15514 , n15501 , n15513 );
not ( n15515 , n15514 );
or ( n15516 , n7869 , n7928 );
or ( n15517 , n120 , n8170 );
nand ( n15518 , n15516 , n15517 , n8171 );
not ( n15519 , n8160 );
or ( n15520 , n15518 , n7736 , n15519 );
nand ( n15521 , n15520 , n126 );
not ( n15522 , n120 );
not ( n15523 , n8006 );
nand ( n15524 , n15523 , n15397 , n8036 , n7737 );
nand ( n15525 , n15522 , n15524 );
not ( n15526 , n7891 );
nand ( n15527 , n15526 , n7916 , n15320 );
and ( n15528 , n8050 , n15527 );
not ( n15529 , n7896 );
and ( n15530 , n120 , n15529 );
nor ( n15531 , n15528 , n15530 );
or ( n15532 , n121 , n15523 );
not ( n15533 , n7790 );
not ( n15534 , n7965 );
not ( n15535 , n7898 );
or ( n15536 , n15534 , n15535 );
not ( n15537 , n126 );
nand ( n15538 , n15536 , n15537 );
and ( n15539 , n15532 , n15533 , n15538 );
nand ( n15540 , n15521 , n15525 , n15531 , n15539 );
nand ( n15541 , n127 , n15540 );
not ( n15542 , n121 );
nand ( n15543 , n15542 , n7874 );
not ( n15544 , n7850 );
and ( n15545 , n15543 , n8200 , n15544 );
not ( n15546 , n15545 );
not ( n15547 , n7948 );
and ( n15548 , n15546 , n15547 );
not ( n15549 , n121 );
and ( n15550 , n15549 , n7885 );
nor ( n15551 , n15550 , n7880 );
not ( n15552 , n7994 );
not ( n15553 , n15552 );
not ( n15554 , n15553 );
not ( n15555 , n15403 );
not ( n15556 , n15555 );
and ( n15557 , n15551 , n15554 , n15556 );
nor ( n15558 , n15557 , n7819 );
nor ( n15559 , n15548 , n15558 );
not ( n15560 , n121 );
or ( n15561 , n15560 , n7950 );
nand ( n15562 , n15561 , n15533 , n8102 );
nand ( n15563 , n8050 , n15562 );
nand ( n15564 , n15515 , n15541 , n15559 , n15563 );
not ( n15565 , n15564 );
not ( n15566 , n7338 );
not ( n15567 , n15566 );
not ( n15568 , n7432 );
not ( n15569 , n11643 );
not ( n15570 , n15569 );
or ( n15571 , n15568 , n15570 );
nand ( n15572 , n15571 , n116 );
not ( n15573 , n15572 );
or ( n15574 , n15567 , n15573 );
nand ( n15575 , n15574 , n11618 );
not ( n15576 , n7406 );
not ( n15577 , n117 );
nand ( n15578 , n15576 , n15577 );
or ( n15579 , n11654 , n15578 );
not ( n15580 , n7610 );
nand ( n15581 , n117 , n15580 );
and ( n15582 , n15579 , n11903 , n15581 );
not ( n15583 , n11778 );
not ( n15584 , n116 );
nand ( n15585 , n15584 , n11834 );
not ( n15586 , n11735 );
not ( n15587 , n11647 );
not ( n15588 , n116 );
nand ( n15589 , n15587 , n15588 );
nand ( n15590 , n15585 , n15586 , n15589 );
not ( n15591 , n15590 );
or ( n15592 , n15583 , n15591 );
not ( n15593 , n117 );
not ( n15594 , n116 );
nand ( n15595 , n15594 , n7602 );
and ( n15596 , n11697 , n15595 );
not ( n15597 , n7599 );
not ( n15598 , n11902 );
nand ( n15599 , n15596 , n15597 , n15598 );
nand ( n15600 , n118 , n15593 , n15599 );
nand ( n15601 , n15592 , n15600 );
not ( n15602 , n15601 );
nand ( n15603 , n15575 , n15582 , n15602 );
not ( n15604 , n15603 );
not ( n15605 , n7589 );
not ( n15606 , n116 );
not ( n15607 , n7374 );
nand ( n15608 , n15606 , n15607 );
not ( n15609 , n15608 );
not ( n15610 , n15609 );
not ( n15611 , n15610 );
or ( n15612 , n15605 , n15611 );
not ( n15613 , n117 );
nand ( n15614 , n15612 , n15613 );
not ( n15615 , n11721 );
nand ( n15616 , n11685 , n15615 );
not ( n15617 , n115 );
nand ( n15618 , n15617 , n113 );
not ( n15619 , n15618 );
not ( n15620 , n116 );
nand ( n15621 , n15619 , n15620 );
not ( n15622 , n15621 );
not ( n15623 , n116 );
nand ( n15624 , n15623 , n7407 );
not ( n15625 , n15624 );
or ( n15626 , n15622 , n15625 );
nand ( n15627 , n15626 , n117 );
and ( n15628 , n15616 , n15586 , n15627 );
not ( n15629 , n118 );
nand ( n15630 , n117 , n7522 );
not ( n15631 , n11714 );
nand ( n15632 , n7468 , n15631 );
and ( n15633 , n15630 , n15632 , n11729 );
not ( n15634 , n11716 );
not ( n15635 , n11642 );
not ( n15636 , n116 );
nand ( n15637 , n15635 , n15636 );
not ( n15638 , n15637 );
or ( n15639 , n15634 , n15638 );
not ( n15640 , n117 );
nand ( n15641 , n15639 , n15640 );
nand ( n15642 , n15633 , n7589 , n15641 );
nand ( n15643 , n15629 , n15642 );
not ( n15644 , n11608 );
not ( n15645 , n15644 );
nand ( n15646 , n15645 , n11769 );
and ( n15647 , n117 , n15646 );
not ( n15648 , n117 );
not ( n15649 , n115 );
nand ( n15650 , n15649 , n11600 );
and ( n15651 , n116 , n7585 );
not ( n15652 , n116 );
and ( n15653 , n15652 , n11637 );
or ( n15654 , n15651 , n15653 );
nand ( n15655 , n15650 , n15654 );
and ( n15656 , n15648 , n15655 );
nor ( n15657 , n15647 , n15656 );
and ( n15658 , n7609 , n7519 );
nand ( n15659 , n15657 , n11784 , n15658 );
nand ( n15660 , n118 , n15659 );
nand ( n15661 , n15614 , n15628 , n15643 , n15660 );
and ( n15662 , n7325 , n15661 );
not ( n15663 , n7325 );
not ( n15664 , n118 );
not ( n15665 , n15664 );
not ( n15666 , n11659 );
nand ( n15667 , n15666 , n7468 );
and ( n15668 , n15667 , n11655 , n11592 );
not ( n15669 , n11591 );
not ( n15670 , n15669 );
not ( n15671 , n117 );
nand ( n15672 , n15670 , n15671 );
not ( n15673 , n116 );
not ( n15674 , n115 );
nand ( n15675 , n15674 , n7371 );
not ( n15676 , n15675 );
nand ( n15677 , n15673 , n15676 );
nand ( n15678 , n15668 , n15672 , n15677 );
not ( n15679 , n15678 );
or ( n15680 , n15665 , n15679 );
nand ( n15681 , n15680 , n15566 );
not ( n15682 , n15681 );
nand ( n15683 , n7585 , n11672 , n11764 );
nand ( n15684 , n117 , n15683 );
nand ( n15685 , n15684 , n15569 , n11649 );
nand ( n15686 , n118 , n15685 );
not ( n15687 , n7593 );
nand ( n15688 , n117 , n15687 );
not ( n15689 , n117 );
not ( n15690 , n7426 );
nand ( n15691 , n11721 , n11655 , n15690 , n11675 );
and ( n15692 , n15689 , n15691 );
nor ( n15693 , n116 , n11721 );
nor ( n15694 , n15692 , n15693 );
nand ( n15695 , n15682 , n15686 , n15688 , n15694 );
and ( n15696 , n15663 , n15695 );
nor ( n15697 , n15662 , n15696 );
not ( n15698 , n118 );
not ( n15699 , n7561 );
and ( n15700 , n11883 , n11897 );
not ( n15701 , n15700 );
or ( n15702 , n15699 , n15701 );
not ( n15703 , n117 );
nand ( n15704 , n15702 , n15703 );
nand ( n15705 , n116 , n11720 );
not ( n15706 , n15705 );
not ( n15707 , n15706 );
not ( n15708 , n15580 );
nand ( n15709 , n15704 , n15707 , n15708 );
nand ( n15710 , n15698 , n15709 );
nand ( n15711 , n15604 , n15697 , n15710 );
not ( n15712 , n15711 );
not ( n15713 , n15712 );
and ( n15714 , n15565 , n15713 );
not ( n15715 , n15565 );
and ( n15716 , n15715 , n15712 );
nor ( n15717 , n15714 , n15716 );
not ( n15718 , n15717 );
not ( n15719 , n15718 );
or ( n15720 , n15443 , n15719 );
not ( n15721 , n15434 );
not ( n15722 , n15439 );
and ( n15723 , n15721 , n15722 );
not ( n15724 , n15340 );
nand ( n15725 , n15724 , n15328 , n15316 , n15312 );
and ( n15726 , n7748 , n15725 );
not ( n15727 , n15364 );
nor ( n15728 , n15726 , n15727 );
nand ( n15729 , n127 , n15418 );
nand ( n15730 , n15369 , n15728 , n15431 , n15729 );
and ( n15731 , n15730 , n15435 );
nor ( n15732 , n15723 , n15731 );
not ( n15733 , n15732 );
and ( n15734 , n15565 , n15712 );
not ( n15735 , n15565 );
and ( n15736 , n15735 , n15713 );
nor ( n15737 , n15734 , n15736 );
not ( n15738 , n15737 );
nand ( n15739 , n15733 , n15738 );
nand ( n15740 , n15720 , n15739 );
not ( n15741 , n15740 );
nor ( n15742 , n15306 , n15741 );
or ( n15743 , n15740 , n15305 );
nand ( n15744 , n15743 , n2352 );
or ( n15745 , n15742 , n15744 );
xnor ( n15746 , n250 , n251 );
or ( n15747 , n2352 , n15746 );
nand ( n15748 , n15745 , n15747 );
not ( n15749 , n10240 );
not ( n15750 , n167 );
and ( n15751 , n15750 , n5291 );
not ( n15752 , n15750 );
nand ( n15753 , n5367 , n5244 );
and ( n15754 , n15752 , n15753 );
nor ( n15755 , n15751 , n15754 );
nor ( n15756 , n15749 , n15755 );
and ( n15757 , n15756 , n5343 , n10266 );
not ( n15758 , n169 );
nor ( n15759 , n15757 , n15758 );
not ( n15760 , n15759 );
not ( n15761 , n169 );
or ( n15762 , n5315 , n10713 );
nand ( n15763 , n15762 , n167 );
not ( n15764 , n167 );
not ( n15765 , n5331 );
or ( n15766 , n166 , n15765 );
nand ( n15767 , n15766 , n10228 , n10193 );
nand ( n15768 , n15764 , n15767 );
nand ( n15769 , n14983 , n10726 , n15763 , n15768 );
nand ( n15770 , n15761 , n15769 );
not ( n15771 , n167 );
not ( n15772 , n15771 );
not ( n15773 , n166 );
not ( n15774 , n14988 );
nand ( n15775 , n15773 , n15774 );
nand ( n15776 , n15775 , n5230 , n5237 );
not ( n15777 , n15776 );
or ( n15778 , n15772 , n15777 );
nand ( n15779 , n5556 , n10752 );
nand ( n15780 , n15779 , n167 , n5210 );
nand ( n15781 , n15778 , n15780 );
nand ( n15782 , n5222 , n5451 );
and ( n15783 , n15782 , n5318 , n5589 );
nand ( n15784 , n165 , n14905 );
nand ( n15785 , n167 , n14998 );
nand ( n15786 , n15783 , n15784 , n15785 );
nand ( n15787 , n169 , n15786 );
or ( n15788 , n166 , n5422 );
nand ( n15789 , n15788 , n5277 );
nand ( n15790 , n5478 , n15789 );
not ( n15791 , n169 );
not ( n15792 , n166 );
not ( n15793 , n15792 );
not ( n15794 , n5634 );
or ( n15795 , n15793 , n15794 );
nand ( n15796 , n15795 , n10289 );
nand ( n15797 , n15791 , n15796 );
nand ( n15798 , n15787 , n15790 , n15797 );
or ( n15799 , n15781 , n15798 );
nand ( n15800 , n15799 , n5449 );
nand ( n15801 , n15760 , n15770 , n15800 );
not ( n15802 , n15801 );
not ( n15803 , n167 );
not ( n15804 , n15803 );
not ( n15805 , n15784 );
or ( n15806 , n15804 , n15805 );
not ( n15807 , n167 );
or ( n15808 , n15807 , n5493 );
nand ( n15809 , n15806 , n15808 );
not ( n15810 , n169 );
or ( n15811 , n167 , n5312 );
nand ( n15812 , n15811 , n10704 , n5304 );
not ( n15813 , n15812 );
or ( n15814 , n15810 , n15813 );
and ( n15815 , n166 , n14956 );
not ( n15816 , n10774 );
nor ( n15817 , n15815 , n15816 );
or ( n15818 , n167 , n15817 );
nand ( n15819 , n15814 , n15818 );
not ( n15820 , n15819 );
nand ( n15821 , n15820 , n14892 , n10234 );
nand ( n15822 , n5441 , n5487 , n14960 );
nand ( n15823 , n167 , n15822 );
not ( n15824 , n15823 );
not ( n15825 , n10268 );
nand ( n15826 , n15825 , n166 );
nand ( n15827 , n15826 , n5530 );
nor ( n15828 , n164 , n5211 );
not ( n15829 , n5451 );
nor ( n15830 , n15829 , n5360 );
nor ( n15831 , n15824 , n15827 , n15828 , n15830 );
or ( n15832 , n169 , n15831 );
not ( n15833 , n5395 );
not ( n15834 , n5597 );
or ( n15835 , n15833 , n15834 );
not ( n15836 , n167 );
nand ( n15837 , n15835 , n15836 );
nand ( n15838 , n5522 , n14933 );
not ( n15839 , n15838 );
nand ( n15840 , n5465 , n5237 , n15839 );
nand ( n15841 , n167 , n15840 );
nand ( n15842 , n15832 , n15837 , n15841 );
or ( n15843 , n15821 , n15842 );
nand ( n15844 , n15843 , n170 );
and ( n15845 , n15802 , n15809 , n15844 );
not ( n15846 , n15845 );
not ( n15847 , n10794 );
and ( n15848 , n15846 , n15847 );
and ( n15849 , n15802 , n15809 , n15844 );
and ( n15850 , n15849 , n5671 );
nor ( n15851 , n15848 , n15850 );
not ( n15852 , n15851 );
not ( n15853 , n4959 );
not ( n15854 , n4805 );
not ( n15855 , n5168 );
or ( n15856 , n15854 , n15855 );
nand ( n15857 , n15856 , n172 );
not ( n15858 , n15857 );
or ( n15859 , n15853 , n15858 );
nand ( n15860 , n15859 , n4879 );
not ( n15861 , n5056 );
nand ( n15862 , n15861 , n12145 );
and ( n15863 , n15862 , n5115 , n4921 );
not ( n15864 , n172 );
nand ( n15865 , n15864 , n4628 );
nand ( n15866 , n15865 , n5098 , n5122 );
nand ( n15867 , n5006 , n15866 );
not ( n15868 , n176 );
not ( n15869 , n172 );
nand ( n15870 , n15869 , n4632 );
not ( n15871 , n5061 );
not ( n15872 , n12901 );
nand ( n15873 , n15870 , n4618 , n15871 , n15872 );
nand ( n15874 , n177 , n15868 , n15873 );
and ( n15875 , n15867 , n15874 );
nand ( n15876 , n15860 , n15863 , n15875 );
not ( n15877 , n15876 );
not ( n15878 , n177 );
not ( n15879 , n176 );
not ( n15880 , n15879 );
nand ( n15881 , n4949 , n4967 , n4720 );
not ( n15882 , n15881 );
or ( n15883 , n15880 , n15882 );
not ( n15884 , n12882 );
and ( n15885 , n4637 , n15884 );
nand ( n15886 , n15883 , n15885 );
nand ( n15887 , n15878 , n15886 );
not ( n15888 , n177 );
not ( n15889 , n15888 );
not ( n15890 , n172 );
not ( n15891 , n5150 );
nand ( n15892 , n15890 , n15891 );
not ( n15893 , n5067 );
not ( n15894 , n176 );
nand ( n15895 , n15893 , n15894 );
nand ( n15896 , n4680 , n4898 );
nor ( n15897 , n5069 , n4842 );
nand ( n15898 , n15892 , n15895 , n15896 , n15897 );
not ( n15899 , n15898 );
or ( n15900 , n15889 , n15899 );
nand ( n15901 , n15900 , n4959 );
not ( n15902 , n15901 );
not ( n15903 , n4859 );
nand ( n15904 , n4595 , n12064 , n15903 );
nand ( n15905 , n176 , n15904 );
nand ( n15906 , n15905 , n5168 , n5153 );
nand ( n15907 , n177 , n15906 );
nand ( n15908 , n176 , n12895 );
not ( n15909 , n176 );
not ( n15910 , n4809 );
not ( n15911 , n12890 );
nand ( n15912 , n4957 , n15910 , n15911 , n4843 );
and ( n15913 , n15909 , n15912 );
nor ( n15914 , n172 , n15911 );
nor ( n15915 , n15913 , n15914 );
nand ( n15916 , n15902 , n15907 , n15908 , n15915 );
and ( n15917 , n178 , n15916 );
not ( n15918 , n178 );
not ( n15919 , n176 );
nor ( n15920 , n171 , n173 );
not ( n15921 , n15920 );
or ( n15922 , n172 , n15921 );
not ( n15923 , n172 );
nand ( n15924 , n15923 , n4717 );
nand ( n15925 , n15922 , n15924 );
not ( n15926 , n15925 );
or ( n15927 , n15919 , n15926 );
not ( n15928 , n4608 );
not ( n15929 , n5088 );
or ( n15930 , n15928 , n15929 );
not ( n15931 , n176 );
nand ( n15932 , n15930 , n15931 );
nand ( n15933 , n15927 , n15932 );
not ( n15934 , n15933 );
not ( n15935 , n177 );
nand ( n15936 , n176 , n4747 );
and ( n15937 , n15936 , n5113 , n12103 );
not ( n15938 , n12132 );
not ( n15939 , n172 );
not ( n15940 , n5027 );
nand ( n15941 , n15939 , n15940 );
not ( n15942 , n15941 );
or ( n15943 , n15938 , n15942 );
not ( n15944 , n176 );
nand ( n15945 , n15943 , n15944 );
nand ( n15946 , n15935 , n15937 , n4608 , n15945 );
not ( n15947 , n12860 );
not ( n15948 , n172 );
not ( n15949 , n4595 );
or ( n15950 , n15948 , n15949 );
not ( n15951 , n172 );
not ( n15952 , n5066 );
nand ( n15953 , n15951 , n15952 );
nand ( n15954 , n15950 , n15953 );
not ( n15955 , n15954 );
or ( n15956 , n15947 , n15955 );
not ( n15957 , n176 );
nand ( n15958 , n15956 , n15957 );
not ( n15959 , n5003 );
nor ( n15960 , n15959 , n12871 );
not ( n15961 , n5014 );
not ( n15962 , n4925 );
or ( n15963 , n15961 , n15962 );
nand ( n15964 , n15963 , n176 );
nand ( n15965 , n15958 , n15960 , n15964 , n177 );
nand ( n15966 , n15946 , n15965 );
nor ( n15967 , n12827 , n12892 );
nand ( n15968 , n15934 , n15966 , n15967 );
and ( n15969 , n15918 , n15968 );
nor ( n15970 , n15917 , n15969 );
nand ( n15971 , n15877 , n15887 , n15970 );
not ( n15972 , n15971 );
nand ( n15973 , n14885 , n14927 , n14946 , n15011 );
not ( n15974 , n15973 );
not ( n15975 , n15974 );
and ( n15976 , n15972 , n15975 );
and ( n15977 , n15971 , n15013 );
nor ( n15978 , n15976 , n15977 );
not ( n15979 , n15978 );
nand ( n15980 , n15852 , n15979 );
not ( n15981 , n15845 );
not ( n15982 , n5665 );
and ( n15983 , n15981 , n15982 );
and ( n15984 , n15849 , n5665 );
nor ( n15985 , n15983 , n15984 );
not ( n15986 , n15985 );
not ( n15987 , n15876 );
nand ( n15988 , n15987 , n15970 , n15887 );
not ( n15989 , n15988 );
not ( n15990 , n15989 );
not ( n15991 , n15974 );
and ( n15992 , n15990 , n15991 );
not ( n15993 , n15971 );
and ( n15994 , n15993 , n15013 );
nor ( n15995 , n15992 , n15994 );
not ( n15996 , n15995 );
nand ( n15997 , n15986 , n15996 );
and ( n15998 , n15980 , n15997 );
not ( n15999 , n258 );
not ( n16000 , n15999 );
not ( n16001 , n10164 );
or ( n16002 , n16000 , n16001 );
or ( n16003 , n15999 , n14707 );
nand ( n16004 , n16002 , n16003 );
not ( n16005 , n14848 );
not ( n16006 , n9918 );
not ( n16007 , n16006 );
nand ( n16008 , n16005 , n159 , n16007 );
not ( n16009 , n159 );
and ( n16010 , n16009 , n10066 );
not ( n16011 , n16009 );
and ( n16012 , n16011 , n12761 );
nor ( n16013 , n16010 , n16012 );
nand ( n16014 , n4050 , n16013 , n9905 , n4110 );
nand ( n16015 , n160 , n16014 );
not ( n16016 , n159 );
nor ( n16017 , n9859 , n4063 );
nand ( n16018 , n16016 , n16017 );
nand ( n16019 , n12819 , n10832 );
not ( n16020 , n159 );
not ( n16021 , n16020 );
not ( n16022 , n158 );
not ( n16023 , n9929 );
nand ( n16024 , n16022 , n16023 );
not ( n16025 , n4232 );
nand ( n16026 , n16024 , n16025 , n4152 );
not ( n16027 , n16026 );
or ( n16028 , n16021 , n16027 );
not ( n16029 , n9919 );
not ( n16030 , n10843 );
or ( n16031 , n16029 , n16030 );
nand ( n16032 , n16031 , n159 );
nand ( n16033 , n16028 , n16032 );
or ( n16034 , n16019 , n16033 );
nand ( n16035 , n16034 , n4054 );
nand ( n16036 , n16008 , n16015 , n16018 , n16035 );
not ( n16037 , n16036 );
not ( n16038 , n4054 );
not ( n16039 , n158 );
not ( n16040 , n16039 );
not ( n16041 , n10052 );
or ( n16042 , n16040 , n16041 );
not ( n16043 , n4068 );
nand ( n16044 , n16042 , n16043 );
not ( n16045 , n16044 );
or ( n16046 , n16038 , n16045 );
not ( n16047 , n10033 );
nor ( n16048 , n16047 , n16017 );
nand ( n16049 , n4192 , n4148 );
not ( n16050 , n4283 );
nand ( n16051 , n159 , n16050 );
nand ( n16052 , n16048 , n16049 , n4163 , n16051 );
nand ( n16053 , n160 , n16052 );
not ( n16054 , n4172 );
not ( n16055 , n4235 );
or ( n16056 , n16054 , n16055 );
not ( n16057 , n158 );
nor ( n16058 , n16057 , n10907 );
nand ( n16059 , n16056 , n16058 );
and ( n16060 , n14826 , n16059 );
not ( n16061 , n159 );
nand ( n16062 , n9956 , n4044 );
nand ( n16063 , n9942 , n16062 );
and ( n16064 , n16061 , n16063 );
or ( n16065 , n158 , n4057 );
not ( n16066 , n4183 );
nand ( n16067 , n16065 , n16066 );
and ( n16068 , n10087 , n16067 );
nor ( n16069 , n16064 , n16068 );
and ( n16070 , n16053 , n16060 , n16069 );
nand ( n16071 , n16046 , n16070 );
nand ( n16072 , n4144 , n16071 );
not ( n16073 , n9969 );
not ( n16074 , n9830 );
not ( n16075 , n10043 );
or ( n16076 , n16074 , n16075 );
not ( n16077 , n159 );
nand ( n16078 , n16076 , n16077 );
nand ( n16079 , n16073 , n14803 , n16078 );
or ( n16080 , n159 , n16006 );
not ( n16081 , n9892 );
nand ( n16082 , n16080 , n9811 , n16081 );
and ( n16083 , n160 , n16082 );
not ( n16084 , n159 );
not ( n16085 , n4130 );
or ( n16086 , n157 , n16085 );
nand ( n16087 , n16086 , n10872 );
and ( n16088 , n16084 , n16087 );
nor ( n16089 , n16083 , n16088 );
and ( n16090 , n10129 , n4186 );
nand ( n16091 , n16090 , n9945 , n12704 );
nand ( n16092 , n159 , n16091 );
nand ( n16093 , n12705 , n10072 );
not ( n16094 , n156 );
nand ( n16095 , n16094 , n4130 );
nand ( n16096 , n4148 , n4099 );
nand ( n16097 , n4257 , n4241 , n14850 );
nand ( n16098 , n159 , n16097 );
nand ( n16099 , n16095 , n16096 , n16098 );
or ( n16100 , n16093 , n16099 );
nand ( n16101 , n16100 , n4054 );
nand ( n16102 , n16089 , n16092 , n16101 );
or ( n16103 , n16079 , n16102 );
nand ( n16104 , n16103 , n161 );
nand ( n16105 , n16037 , n16072 , n16104 );
not ( n16106 , n16105 );
not ( n16107 , n16106 );
nand ( n16108 , n12255 , n10341 );
not ( n16109 , n149 );
nor ( n16110 , n16109 , n4399 );
not ( n16111 , n16110 );
not ( n16112 , n10339 );
nand ( n16113 , n10435 , n4398 );
not ( n16114 , n16113 );
or ( n16115 , n16112 , n16114 );
not ( n16116 , n149 );
nand ( n16117 , n16115 , n16116 );
nand ( n16118 , n16111 , n4548 , n16117 );
nor ( n16119 , n16108 , n16118 );
or ( n16120 , n152 , n16119 );
nand ( n16121 , n16120 , n10426 );
not ( n16122 , n4548 );
not ( n16123 , n10378 );
or ( n16124 , n16122 , n16123 );
not ( n16125 , n149 );
nand ( n16126 , n16124 , n16125 );
not ( n16127 , n16126 );
not ( n16128 , n150 );
not ( n16129 , n16128 );
nor ( n16130 , n148 , n151 );
not ( n16131 , n16130 );
or ( n16132 , n16129 , n16131 );
not ( n16133 , n4391 );
not ( n16134 , n150 );
nand ( n16135 , n16133 , n16134 );
nand ( n16136 , n16132 , n16135 );
nand ( n16137 , n149 , n16136 );
nand ( n16138 , n10565 , n13002 );
not ( n16139 , n10410 );
not ( n16140 , n16139 );
not ( n16141 , n10512 );
or ( n16142 , n16140 , n16141 );
nand ( n16143 , n16142 , n149 );
not ( n16144 , n13025 );
not ( n16145 , n150 );
and ( n16146 , n16145 , n10370 );
not ( n16147 , n16145 );
and ( n16148 , n16147 , n4540 );
nor ( n16149 , n16146 , n16148 );
not ( n16150 , n16149 );
or ( n16151 , n16144 , n16150 );
not ( n16152 , n149 );
nand ( n16153 , n16151 , n16152 );
nand ( n16154 , n16143 , n16153 );
or ( n16155 , n16138 , n16154 );
nand ( n16156 , n16155 , n152 );
nand ( n16157 , n16137 , n12966 , n16156 );
nor ( n16158 , n16121 , n16127 , n16157 );
or ( n16159 , n153 , n16158 );
not ( n16160 , n149 );
not ( n16161 , n16160 );
nand ( n16162 , n10507 , n10420 , n4386 );
not ( n16163 , n16162 );
or ( n16164 , n16161 , n16163 );
and ( n16165 , n4564 , n12997 );
nand ( n16166 , n16164 , n16165 );
nand ( n16167 , n4532 , n16166 );
nand ( n16168 , n16159 , n16167 );
not ( n16169 , n16168 );
not ( n16170 , n153 );
not ( n16171 , n149 );
not ( n16172 , n16171 );
nand ( n16173 , n10539 , n10521 , n4520 , n4455 );
not ( n16174 , n16173 );
or ( n16175 , n16172 , n16174 );
and ( n16176 , n149 , n4545 );
not ( n16177 , n4525 );
nor ( n16178 , n16176 , n16177 );
nand ( n16179 , n16175 , n16178 );
not ( n16180 , n16179 );
not ( n16181 , n150 );
not ( n16182 , n10521 );
nand ( n16183 , n16181 , n16182 );
nand ( n16184 , n10382 , n12238 , n4541 );
nand ( n16185 , n149 , n16184 );
nand ( n16186 , n16185 , n10353 , n10450 );
nand ( n16187 , n152 , n16186 );
not ( n16188 , n150 );
not ( n16189 , n148 );
or ( n16190 , n16188 , n16189 , n10432 );
nand ( n16191 , n16190 , n4455 );
not ( n16192 , n10324 );
or ( n16193 , n150 , n16192 );
or ( n16194 , n149 , n10371 );
nand ( n16195 , n16193 , n16194 , n10372 );
or ( n16196 , n16191 , n16195 );
nand ( n16197 , n16196 , n4532 );
nand ( n16198 , n16180 , n16183 , n16187 , n16197 );
not ( n16199 , n16198 );
or ( n16200 , n16170 , n16199 );
not ( n16201 , n10561 );
or ( n16202 , n150 , n4419 );
nand ( n16203 , n16202 , n10426 , n12988 );
not ( n16204 , n16203 );
or ( n16205 , n16201 , n16204 );
nand ( n16206 , n16205 , n10343 );
not ( n16207 , n4525 );
not ( n16208 , n4466 );
not ( n16209 , n10351 );
or ( n16210 , n16208 , n16209 );
nand ( n16211 , n16210 , n150 );
not ( n16212 , n16211 );
or ( n16213 , n16207 , n16212 );
nand ( n16214 , n16213 , n10610 );
not ( n16215 , n149 );
not ( n16216 , n16215 );
not ( n16217 , n150 );
not ( n16218 , n4554 );
and ( n16219 , n16217 , n16218 );
nor ( n16220 , n16219 , n10554 );
nand ( n16221 , n16220 , n4559 , n10498 );
not ( n16222 , n16221 );
or ( n16223 , n16216 , n16222 );
nand ( n16224 , n10469 , n4511 );
nand ( n16225 , n16223 , n16224 );
nand ( n16226 , n152 , n16225 );
nand ( n16227 , n10499 , n16214 , n16226 );
nor ( n16228 , n16206 , n16227 );
nand ( n16229 , n16200 , n16228 );
not ( n16230 , n16229 );
nand ( n16231 , n16169 , n16230 );
not ( n16232 , n16231 );
and ( n16233 , n16107 , n16232 );
not ( n16234 , n16105 );
not ( n16235 , n16231 );
not ( n16236 , n16235 );
and ( n16237 , n16234 , n16236 );
nor ( n16238 , n16233 , n16237 );
and ( n16239 , n16004 , n16238 );
not ( n16240 , n16004 );
not ( n16241 , n16238 );
and ( n16242 , n16240 , n16241 );
nor ( n16243 , n16239 , n16242 );
not ( n16244 , n16243 );
nor ( n16245 , n15998 , n16244 );
nand ( n16246 , n15980 , n15997 );
or ( n16247 , n16243 , n16246 );
nand ( n16248 , n16247 , n2352 );
or ( n16249 , n16245 , n16248 );
and ( n16250 , n259 , n15999 );
not ( n16251 , n259 );
and ( n16252 , n16251 , n258 );
nor ( n16253 , n16250 , n16252 );
or ( n16254 , n2352 , n16253 );
nand ( n16255 , n16249 , n16254 );
not ( n16256 , n14697 );
not ( n16257 , n10654 );
and ( n16258 , n16256 , n16257 );
not ( n16259 , n10654 );
not ( n16260 , n16259 );
and ( n16261 , n14697 , n16260 );
nor ( n16262 , n16258 , n16261 );
not ( n16263 , n286 );
and ( n16264 , n4301 , n16263 );
not ( n16265 , n4301 );
and ( n16266 , n16265 , n286 );
nor ( n16267 , n16264 , n16266 );
and ( n16268 , n16262 , n16267 );
not ( n16269 , n16262 );
not ( n16270 , n16267 );
and ( n16271 , n16269 , n16270 );
nor ( n16272 , n16268 , n16271 );
not ( n16273 , n16272 );
not ( n16274 , n10307 );
not ( n16275 , n5205 );
and ( n16276 , n16274 , n16275 );
and ( n16277 , n10307 , n5205 );
nor ( n16278 , n16276 , n16277 );
not ( n16279 , n5042 );
and ( n16280 , n12044 , n16279 );
not ( n16281 , n12044 );
and ( n16282 , n16281 , n5200 );
nor ( n16283 , n16280 , n16282 );
not ( n16284 , n16283 );
and ( n16285 , n16278 , n16284 );
not ( n16286 , n16278 );
and ( n16287 , n16286 , n16283 );
nor ( n16288 , n16285 , n16287 );
not ( n16289 , n16288 );
nor ( n16290 , n16273 , n16289 );
or ( n16291 , n16272 , n16288 );
nand ( n16292 , n16291 , n2352 );
or ( n16293 , n16290 , n16292 );
and ( n16294 , n287 , n16263 );
not ( n16295 , n287 );
and ( n16296 , n16295 , n286 );
nor ( n16297 , n16294 , n16296 );
or ( n16298 , n2352 , n16297 );
nand ( n16299 , n16293 , n16298 );
not ( n16300 , n340 );
and ( n16301 , n341 , n16300 );
not ( n16302 , n341 );
and ( n16303 , n16302 , n340 );
nor ( n16304 , n16301 , n16303 );
or ( n16305 , n2352 , n16304 );
not ( n16306 , n3275 );
not ( n16307 , n9189 );
not ( n16308 , n16307 );
not ( n16309 , n8802 );
not ( n16310 , n8908 );
or ( n16311 , n16309 , n16310 );
nand ( n16312 , n16311 , n185 );
not ( n16313 , n185 );
not ( n16314 , n8850 );
nand ( n16315 , n16313 , n16314 );
and ( n16316 , n16315 , n3222 , n8821 );
nand ( n16317 , n16308 , n16312 , n16316 );
nand ( n16318 , n16317 , n186 );
nand ( n16319 , n8795 , n8792 );
and ( n16320 , n185 , n183 , n3081 );
and ( n16321 , n3047 , n3095 );
not ( n16322 , n3283 );
nor ( n16323 , n16321 , n16322 );
nor ( n16324 , n16320 , n16323 );
not ( n16325 , n184 );
not ( n16326 , n3376 );
nand ( n16327 , n16325 , n16326 );
nand ( n16328 , n16319 , n16324 , n16327 , n3427 );
nand ( n16329 , n3013 , n16328 );
not ( n16330 , n184 );
and ( n16331 , n16330 , n8895 );
and ( n16332 , n3258 , n8803 );
nor ( n16333 , n16331 , n16332 );
not ( n16334 , n185 );
not ( n16335 , n16334 );
nand ( n16336 , n11111 , n8781 );
not ( n16337 , n16336 );
or ( n16338 , n16335 , n16337 );
not ( n16339 , n185 );
or ( n16340 , n16339 , n3023 );
nand ( n16341 , n16338 , n16340 );
not ( n16342 , n16341 );
nand ( n16343 , n16318 , n16329 , n16333 , n16342 );
not ( n16344 , n16343 );
or ( n16345 , n16306 , n16344 );
not ( n16346 , n185 );
or ( n16347 , n16346 , n8882 );
nand ( n16348 , n16347 , n8896 );
nand ( n16349 , n3013 , n16348 );
nand ( n16350 , n16345 , n16349 );
not ( n16351 , n16350 );
nand ( n16352 , n9138 , n9208 );
or ( n16353 , n8768 , n11165 );
or ( n16354 , n3011 , n3417 );
not ( n16355 , n9218 );
not ( n16356 , n3176 );
nand ( n16357 , n16355 , n16356 );
and ( n16358 , n11166 , n16357 );
not ( n16359 , n16358 );
not ( n16360 , n185 );
or ( n16361 , n3112 , n3129 );
nand ( n16362 , n16361 , n9135 );
not ( n16363 , n16362 );
or ( n16364 , n16360 , n16363 );
nand ( n16365 , n8861 , n3276 , n8850 );
nand ( n16366 , n3092 , n16365 );
nand ( n16367 , n16364 , n16366 );
not ( n16368 , n16367 );
not ( n16369 , n16368 );
or ( n16370 , n16359 , n16369 );
nand ( n16371 , n16370 , n186 );
nand ( n16372 , n16353 , n16354 , n16371 );
nor ( n16373 , n16352 , n16372 );
not ( n16374 , n185 );
not ( n16375 , n184 );
nand ( n16376 , n16375 , n3290 );
nand ( n16377 , n16376 , n3439 , n3053 );
not ( n16378 , n16377 );
or ( n16379 , n16374 , n16378 );
nand ( n16380 , n16379 , n9135 );
not ( n16381 , n16380 );
and ( n16382 , n3213 , n3071 );
nand ( n16383 , n16381 , n16382 , n3301 , n3117 );
and ( n16384 , n186 , n16383 );
not ( n16385 , n186 );
not ( n16386 , n8858 );
nand ( n16387 , n16386 , n185 );
not ( n16388 , n8828 );
not ( n16389 , n3353 );
or ( n16390 , n16388 , n16389 );
not ( n16391 , n185 );
nand ( n16392 , n16390 , n16391 );
and ( n16393 , n3251 , n16387 , n16392 );
nor ( n16394 , n8776 , n3224 );
and ( n16395 , n16394 , n11108 , n9207 );
nand ( n16396 , n16393 , n16395 );
and ( n16397 , n16385 , n16396 );
nor ( n16398 , n16384 , n16397 );
not ( n16399 , n183 );
not ( n16400 , n8784 );
or ( n16401 , n16399 , n16400 );
nand ( n16402 , n16401 , n9182 );
nand ( n16403 , n185 , n16402 );
not ( n16404 , n16327 );
or ( n16405 , n16404 , n3075 );
not ( n16406 , n185 );
nand ( n16407 , n16405 , n16406 );
nand ( n16408 , n16398 , n16403 , n8894 , n16407 );
nand ( n16409 , n16408 , n187 );
nand ( n16410 , n16351 , n16373 , n16409 );
not ( n16411 , n16410 );
not ( n16412 , n16411 );
not ( n16413 , n12558 );
and ( n16414 , n16412 , n16413 );
and ( n16415 , n16411 , n12564 );
nor ( n16416 , n16414 , n16415 );
not ( n16417 , n2364 );
not ( n16418 , n191 );
not ( n16419 , n2418 );
nand ( n16420 , n16418 , n16419 );
and ( n16421 , n193 , n192 , n2474 );
and ( n16422 , n2412 , n2525 );
nor ( n16423 , n16422 , n2560 );
nor ( n16424 , n16421 , n16423 );
and ( n16425 , n16420 , n16424 );
not ( n16426 , n194 );
nand ( n16427 , n2504 , n8956 );
nand ( n16428 , n16425 , n16426 , n2531 , n16427 );
not ( n16429 , n9014 );
not ( n16430 , n8966 );
or ( n16431 , n16429 , n16430 );
nand ( n16432 , n16431 , n193 );
not ( n16433 , n194 );
not ( n16434 , n9056 );
nor ( n16435 , n16433 , n16434 );
not ( n16436 , n193 );
nand ( n16437 , n16436 , n2394 );
and ( n16438 , n16437 , n12362 , n2431 );
nand ( n16439 , n16432 , n16435 , n16438 );
nand ( n16440 , n16428 , n16439 );
not ( n16441 , n193 );
not ( n16442 , n2554 );
nor ( n16443 , n12320 , n16442 );
not ( n16444 , n16443 );
nand ( n16445 , n16441 , n16444 );
nand ( n16446 , n193 , n2572 );
not ( n16447 , n191 );
and ( n16448 , n16447 , n2380 );
and ( n16449 , n2472 , n9015 );
nor ( n16450 , n16448 , n16449 );
nand ( n16451 , n16440 , n16445 , n16446 , n16450 );
not ( n16452 , n16451 );
or ( n16453 , n16417 , n16452 );
not ( n16454 , n194 );
not ( n16455 , n193 );
not ( n16456 , n2534 );
not ( n16457 , n16456 );
or ( n16458 , n16455 , n16457 );
nand ( n16459 , n16458 , n8980 );
nand ( n16460 , n16454 , n16459 );
nand ( n16461 , n16453 , n16460 );
not ( n16462 , n16461 );
not ( n16463 , n2585 );
not ( n16464 , n2394 );
nand ( n16465 , n2956 , n12384 , n16464 );
not ( n16466 , n16465 );
or ( n16467 , n16463 , n16466 );
or ( n16468 , n2795 , n2781 );
not ( n16469 , n2567 );
nand ( n16470 , n16468 , n16469 );
nand ( n16471 , n193 , n16470 );
nand ( n16472 , n16467 , n16471 );
not ( n16473 , n16472 );
not ( n16474 , n2767 );
not ( n16475 , n193 );
nand ( n16476 , n16474 , n16475 );
nand ( n16477 , n16473 , n12379 , n16476 );
nand ( n16478 , n194 , n16477 );
not ( n16479 , n194 );
not ( n16480 , n193 );
and ( n16481 , n16479 , n16480 , n12375 );
nor ( n16482 , n16481 , n2470 );
not ( n16483 , n193 );
nand ( n16484 , n16420 , n2687 , n2789 );
nand ( n16485 , n16483 , n16484 );
not ( n16486 , n192 );
or ( n16487 , n8940 , n16486 );
nand ( n16488 , n16487 , n2373 );
and ( n16489 , n16488 , n193 );
nor ( n16490 , n16489 , n2735 );
not ( n16491 , n193 );
not ( n16492 , n191 );
not ( n16493 , n2489 );
nand ( n16494 , n16492 , n16493 );
nand ( n16495 , n16494 , n2391 , n2911 );
not ( n16496 , n16495 );
or ( n16497 , n16491 , n16496 );
nand ( n16498 , n16497 , n12358 );
not ( n16499 , n16498 );
not ( n16500 , n2588 );
nor ( n16501 , n16500 , n2721 );
nor ( n16502 , n2799 , n2951 );
nand ( n16503 , n194 , n16499 , n16501 , n16502 );
nand ( n16504 , n2740 , n2469 );
nand ( n16505 , n12322 , n8969 );
nor ( n16506 , n16504 , n16505 );
and ( n16507 , n2504 , n2528 );
and ( n16508 , n193 , n2807 );
nor ( n16509 , n16507 , n16508 );
nor ( n16510 , n2550 , n194 );
nand ( n16511 , n16506 , n2712 , n16509 , n16510 );
nand ( n16512 , n16503 , n16511 );
nand ( n16513 , n16485 , n16490 , n16512 );
nand ( n16514 , n195 , n16513 );
and ( n16515 , n16478 , n16482 , n16514 );
nand ( n16516 , n2472 , n2423 );
not ( n16517 , n2565 );
not ( n16518 , n16517 );
nand ( n16519 , n16462 , n16515 , n16516 , n16518 );
not ( n16520 , n16519 );
not ( n16521 , n16520 );
not ( n16522 , n16300 );
and ( n16523 , n16521 , n16522 );
not ( n16524 , n16461 );
nand ( n16525 , n16524 , n16515 , n16516 , n16518 );
not ( n16526 , n16525 );
and ( n16527 , n16526 , n16300 );
nor ( n16528 , n16523 , n16527 );
and ( n16529 , n16416 , n16528 );
not ( n16530 , n16416 );
not ( n16531 , n16528 );
and ( n16532 , n16530 , n16531 );
nor ( n16533 , n16529 , n16532 );
not ( n16534 , n16533 );
not ( n16535 , n211 );
not ( n16536 , n3561 );
not ( n16537 , n8604 );
or ( n16538 , n16536 , n16537 );
nand ( n16539 , n16538 , n9428 );
and ( n16540 , n16535 , n16539 );
not ( n16541 , n16535 );
not ( n16542 , n209 );
nand ( n16543 , n9358 , n3501 , n8667 );
nand ( n16544 , n16542 , n16543 );
not ( n16545 , n9278 );
not ( n16546 , n3643 );
or ( n16547 , n16545 , n16546 );
nand ( n16548 , n16547 , n209 );
nand ( n16549 , n16544 , n3483 , n16548 );
and ( n16550 , n16541 , n16549 );
nor ( n16551 , n16540 , n16550 );
not ( n16552 , n16551 );
nand ( n16553 , n8636 , n8621 );
not ( n16554 , n8473 );
nand ( n16555 , n16553 , n16554 , n8660 );
nor ( n16556 , n16552 , n16555 );
nor ( n16557 , n16556 , n212 );
not ( n16558 , n16557 );
or ( n16559 , n210 , n9407 );
not ( n16560 , n8621 );
nand ( n16561 , n16559 , n16560 );
and ( n16562 , n3717 , n16561 );
not ( n16563 , n3725 );
and ( n16564 , n8499 , n16563 );
not ( n16565 , n209 );
nor ( n16566 , n16564 , n16565 , n8454 );
nor ( n16567 , n16562 , n16566 );
and ( n16568 , n209 , n3741 , n8605 );
not ( n16569 , n12461 );
nor ( n16570 , n16568 , n16569 );
or ( n16571 , n209 , n3522 );
not ( n16572 , n209 );
not ( n16573 , n3543 );
not ( n16574 , n8673 );
or ( n16575 , n16573 , n16574 );
nand ( n16576 , n16575 , n3513 );
nand ( n16577 , n16572 , n16576 );
nand ( n16578 , n16571 , n16577 , n3529 );
nand ( n16579 , n211 , n16578 );
and ( n16580 , n16567 , n16570 , n16579 );
nand ( n16581 , n3610 , n3518 , n3480 );
and ( n16582 , n8636 , n16581 );
nor ( n16583 , n16582 , n8538 );
and ( n16584 , n3607 , n8531 );
not ( n16585 , n9318 );
not ( n16586 , n209 );
not ( n16587 , n205 );
or ( n16588 , n16587 , n8448 );
nand ( n16589 , n16588 , n9448 );
and ( n16590 , n16586 , n16589 );
and ( n16591 , n209 , n8670 );
nor ( n16592 , n16590 , n16591 );
not ( n16593 , n16592 );
or ( n16594 , n16585 , n16593 );
nand ( n16595 , n16594 , n211 );
not ( n16596 , n211 );
and ( n16597 , n209 , n8714 );
not ( n16598 , n209 );
and ( n16599 , n16598 , n3584 );
nor ( n16600 , n16597 , n16599 );
and ( n16601 , n8486 , n3726 );
and ( n16602 , n8463 , n8554 , n9348 );
nand ( n16603 , n16600 , n8749 , n16601 , n16602 );
nand ( n16604 , n16596 , n16603 );
nand ( n16605 , n16583 , n16584 , n16595 , n16604 );
nand ( n16606 , n212 , n16605 );
not ( n16607 , n209 );
not ( n16608 , n16607 );
nand ( n16609 , n8489 , n3546 , n8530 );
not ( n16610 , n16609 );
or ( n16611 , n16608 , n16610 );
nand ( n16612 , n9303 , n3725 );
nand ( n16613 , n16611 , n16612 );
nand ( n16614 , n210 , n3622 );
nand ( n16615 , n16614 , n9428 , n3589 );
nand ( n16616 , n209 , n16615 );
not ( n16617 , n9448 );
nand ( n16618 , n210 , n16617 );
nand ( n16619 , n16616 , n8509 , n16618 );
nor ( n16620 , n16613 , n16619 );
nor ( n16621 , n211 , n16620 );
not ( n16622 , n16621 );
nand ( n16623 , n16558 , n16580 , n16606 , n16622 );
not ( n16624 , n16623 );
not ( n16625 , n16624 );
not ( n16626 , n9509 );
and ( n16627 , n16625 , n16626 );
not ( n16628 , n16623 );
and ( n16629 , n9514 , n16628 );
nor ( n16630 , n16627 , n16629 );
not ( n16631 , n16630 );
not ( n16632 , n202 );
not ( n16633 , n3958 );
not ( n16634 , n16633 );
not ( n16635 , n3909 );
or ( n16636 , n16634 , n16635 );
nand ( n16637 , n16636 , n3814 );
nand ( n16638 , n16632 , n16637 );
not ( n16639 , n10962 );
not ( n16640 , n202 );
not ( n16641 , n3820 );
nand ( n16642 , n16640 , n16641 );
nand ( n16643 , n16638 , n16639 , n16642 );
and ( n16644 , n203 , n16643 );
not ( n16645 , n203 );
not ( n16646 , n202 );
not ( n16647 , n16646 );
nand ( n16648 , n9646 , n3756 , n8412 );
not ( n16649 , n16648 );
or ( n16650 , n16647 , n16649 );
not ( n16651 , n202 );
nand ( n16652 , n16651 , n3882 );
nand ( n16653 , n16650 , n16652 );
not ( n16654 , n16653 );
not ( n16655 , n9583 );
nand ( n16656 , n201 , n16655 );
nand ( n16657 , n201 , n3953 );
nand ( n16658 , n16657 , n9630 , n3926 );
nand ( n16659 , n202 , n16658 );
nand ( n16660 , n16654 , n16656 , n9738 , n16659 );
and ( n16661 , n16645 , n16660 );
nor ( n16662 , n16644 , n16661 );
not ( n16663 , n9549 );
or ( n16664 , n201 , n16663 );
nand ( n16665 , n16664 , n10986 );
and ( n16666 , n3825 , n16665 );
and ( n16667 , n8362 , n9725 );
not ( n16668 , n202 );
not ( n16669 , n8293 );
nor ( n16670 , n16667 , n16668 , n16669 );
nor ( n16671 , n16666 , n16670 );
nand ( n16672 , n203 , n3897 , n3765 );
and ( n16673 , n12670 , n16672 );
nand ( n16674 , n3897 , n3806 );
and ( n16675 , n16674 , n8312 , n10966 );
not ( n16676 , n203 );
not ( n16677 , n3778 );
not ( n16678 , n3904 );
or ( n16679 , n16677 , n16678 );
nand ( n16680 , n16679 , n9630 );
nand ( n16681 , n16676 , n16680 );
not ( n16682 , n9754 );
nor ( n16683 , n3830 , n11042 );
not ( n16684 , n16683 );
or ( n16685 , n16682 , n16684 );
not ( n16686 , n202 );
nand ( n16687 , n16685 , n16686 );
not ( n16688 , n9605 );
not ( n16689 , n3972 );
or ( n16690 , n16688 , n16689 );
nand ( n16691 , n16690 , n202 );
nand ( n16692 , n16687 , n3787 , n16691 );
nand ( n16693 , n203 , n16692 );
nand ( n16694 , n16675 , n16681 , n16693 );
nand ( n16695 , n4008 , n16694 );
nand ( n16696 , n16671 , n16673 , n16695 );
not ( n16697 , n16696 );
not ( n16698 , n203 );
and ( n16699 , n8370 , n11085 );
and ( n16700 , n8299 , n8286 );
and ( n16701 , n3969 , n3999 );
not ( n16702 , n202 );
not ( n16703 , n16702 );
not ( n16704 , n3864 );
or ( n16705 , n16703 , n16704 );
nand ( n16706 , n16705 , n9538 );
nor ( n16707 , n16701 , n16706 );
nand ( n16708 , n16699 , n3883 , n16700 , n16707 );
nand ( n16709 , n16698 , n16708 );
not ( n16710 , n16709 );
not ( n16711 , n3979 );
nand ( n16712 , n3939 , n16711 , n3795 );
nand ( n16713 , n3897 , n16712 );
nand ( n16714 , n8345 , n16713 );
not ( n16715 , n203 );
not ( n16716 , n202 );
or ( n16717 , n3889 , n3908 );
nand ( n16718 , n16717 , n9583 );
nand ( n16719 , n16716 , n16718 );
not ( n16720 , n8379 );
nand ( n16721 , n16720 , n202 );
nand ( n16722 , n16719 , n16721 , n9673 );
not ( n16723 , n16722 );
or ( n16724 , n16715 , n16723 );
and ( n16725 , n4000 , n8425 );
nand ( n16726 , n16724 , n16725 );
nor ( n16727 , n16714 , n16726 );
not ( n16728 , n16727 );
or ( n16729 , n16710 , n16728 );
nand ( n16730 , n16729 , n204 );
and ( n16731 , n16662 , n16697 , n16730 );
and ( n16732 , n9782 , n16731 );
not ( n16733 , n9782 );
not ( n16734 , n16730 );
nor ( n16735 , n16696 , n16734 );
nand ( n16736 , n16662 , n16735 );
and ( n16737 , n16733 , n16736 );
nor ( n16738 , n16732 , n16737 );
not ( n16739 , n16738 );
and ( n16740 , n16631 , n16739 );
and ( n16741 , n16630 , n16738 );
nor ( n16742 , n16740 , n16741 );
not ( n16743 , n16742 );
nand ( n16744 , n16534 , n16743 );
nand ( n16745 , n16533 , n16742 );
nand ( n16746 , n16744 , n2352 , n16745 );
nand ( n16747 , n16305 , n16746 );
not ( n16748 , n16525 );
not ( n16749 , n16748 );
not ( n16750 , n98 );
not ( n16751 , n16750 );
and ( n16752 , n16749 , n16751 );
not ( n16753 , n98 );
and ( n16754 , n16753 , n16526 );
nor ( n16755 , n16752 , n16754 );
not ( n16756 , n2364 );
not ( n16757 , n193 );
or ( n16758 , n16757 , n2845 );
nand ( n16759 , n16758 , n2589 , n8963 );
not ( n16760 , n194 );
not ( n16761 , n2676 );
not ( n16762 , n2635 );
or ( n16763 , n16761 , n16762 );
nand ( n16764 , n16763 , n193 );
not ( n16765 , n193 );
nand ( n16766 , n2414 , n2783 , n9014 );
nand ( n16767 , n16765 , n16766 );
nand ( n16768 , n16764 , n2453 , n16767 );
not ( n16769 , n16768 );
or ( n16770 , n16760 , n16769 );
not ( n16771 , n194 );
or ( n16772 , n2385 , n2503 );
nand ( n16773 , n16772 , n2720 );
nand ( n16774 , n16771 , n16773 );
nand ( n16775 , n16770 , n16774 );
nor ( n16776 , n16759 , n16775 );
not ( n16777 , n16776 );
or ( n16778 , n16756 , n16777 );
not ( n16779 , n2472 );
not ( n16780 , n2614 );
nand ( n16781 , n2451 , n16780 , n2563 );
not ( n16782 , n16781 );
or ( n16783 , n16779 , n16782 );
nand ( n16784 , n16783 , n2742 );
not ( n16785 , n16784 );
not ( n16786 , n2756 );
not ( n16787 , n2562 );
nor ( n16788 , n16786 , n16787 );
not ( n16789 , n2736 );
and ( n16790 , n193 , n2476 );
not ( n16791 , n193 );
or ( n16792 , n2894 , n2771 );
nand ( n16793 , n16792 , n2956 );
and ( n16794 , n16791 , n16793 );
nor ( n16795 , n16790 , n16794 );
not ( n16796 , n16795 );
or ( n16797 , n16789 , n16796 );
nand ( n16798 , n16797 , n194 );
nand ( n16799 , n16785 , n16788 , n16798 );
not ( n16800 , n16799 );
nand ( n16801 , n12374 , n2808 );
nor ( n16802 , n16801 , n2483 , n8974 );
not ( n16803 , n16802 );
not ( n16804 , n193 );
or ( n16805 , n16804 , n2950 );
nand ( n16806 , n16805 , n12322 );
not ( n16807 , n193 );
not ( n16808 , n16807 );
not ( n16809 , n2550 );
or ( n16810 , n16808 , n16809 );
nand ( n16811 , n16810 , n12387 );
nor ( n16812 , n16806 , n16811 );
not ( n16813 , n16812 );
or ( n16814 , n16803 , n16813 );
not ( n16815 , n194 );
nand ( n16816 , n16814 , n16815 );
nand ( n16817 , n16800 , n195 , n16816 );
nand ( n16818 , n16778 , n16817 );
not ( n16819 , n2599 );
or ( n16820 , n2376 , n16819 );
nand ( n16821 , n16820 , n2817 );
nand ( n16822 , n193 , n16821 );
not ( n16823 , n16822 );
not ( n16824 , n193 );
or ( n16825 , n2803 , n2771 );
nand ( n16826 , n16825 , n2424 );
nand ( n16827 , n16824 , n16826 );
not ( n16828 , n193 );
not ( n16829 , n12397 );
or ( n16830 , n16828 , n16829 );
not ( n16831 , n193 );
nand ( n16832 , n16831 , n2431 );
nand ( n16833 , n16830 , n16832 );
and ( n16834 , n16827 , n2436 , n16833 );
not ( n16835 , n16834 );
or ( n16836 , n16823 , n16835 );
nand ( n16837 , n16836 , n194 );
not ( n16838 , n194 );
not ( n16839 , n193 );
not ( n16840 , n16839 );
nand ( n16841 , n2714 , n2373 , n2887 );
not ( n16842 , n16841 );
or ( n16843 , n16840 , n16842 );
nor ( n16844 , n2586 , n2482 );
not ( n16845 , n16844 );
nand ( n16846 , n16843 , n16845 );
not ( n16847 , n16846 );
not ( n16848 , n191 );
nor ( n16849 , n16848 , n2956 );
not ( n16850 , n193 );
nand ( n16851 , n191 , n2625 );
nand ( n16852 , n16851 , n2720 , n2573 );
not ( n16853 , n16852 );
or ( n16854 , n16850 , n16853 );
nand ( n16855 , n16854 , n2787 );
nor ( n16856 , n16849 , n16855 );
nand ( n16857 , n16847 , n16856 );
and ( n16858 , n16838 , n16857 );
and ( n16859 , n2670 , n2482 );
nor ( n16860 , n16859 , n191 , n2700 );
not ( n16861 , n16860 );
nand ( n16862 , n16861 , n16476 );
nor ( n16863 , n16858 , n16862 );
and ( n16864 , n16818 , n16837 , n16863 );
buf ( n16865 , n16864 );
not ( n16866 , n2991 );
and ( n16867 , n16865 , n16866 );
not ( n16868 , n16865 );
and ( n16869 , n16868 , n2987 );
nor ( n16870 , n16867 , n16869 );
not ( n16871 , n16870 );
nand ( n16872 , n16755 , n16871 );
not ( n16873 , n16755 );
nand ( n16874 , n16873 , n16870 );
nand ( n16875 , n16872 , n16874 );
not ( n16876 , n16875 );
not ( n16877 , n3084 );
not ( n16878 , n8863 );
or ( n16879 , n16877 , n16878 );
nand ( n16880 , n16879 , n185 );
not ( n16881 , n9169 );
not ( n16882 , n185 );
nand ( n16883 , n8802 , n3097 , n3159 );
nand ( n16884 , n16882 , n16883 );
nand ( n16885 , n16880 , n16881 , n16884 );
nand ( n16886 , n186 , n16885 );
not ( n16887 , n185 );
or ( n16888 , n16887 , n3319 );
nand ( n16889 , n16886 , n8904 , n16888 );
not ( n16890 , n3013 );
or ( n16891 , n3137 , n9218 );
nand ( n16892 , n16891 , n3213 );
not ( n16893 , n16892 );
or ( n16894 , n16890 , n16893 );
not ( n16895 , n8792 );
nand ( n16896 , n16894 , n16895 );
or ( n16897 , n16889 , n16896 );
nand ( n16898 , n16897 , n3275 );
not ( n16899 , n181 );
not ( n16900 , n3220 );
or ( n16901 , n16899 , n16900 );
nand ( n16902 , n16901 , n3149 );
and ( n16903 , n3329 , n16902 );
and ( n16904 , n3088 , n3009 );
not ( n16905 , n3347 );
nor ( n16906 , n16904 , n183 , n16905 );
nor ( n16907 , n16903 , n16906 );
not ( n16908 , n11200 );
nand ( n16909 , n3329 , n16908 );
not ( n16910 , n185 );
not ( n16911 , n16910 );
nand ( n16912 , n183 , n9152 );
nand ( n16913 , n16912 , n3417 , n9189 );
not ( n16914 , n16913 );
or ( n16915 , n16911 , n16914 );
nand ( n16916 , n16915 , n8828 );
nand ( n16917 , n186 , n16916 );
and ( n16918 , n16907 , n16909 , n16357 , n16917 );
nand ( n16919 , n16898 , n16918 );
not ( n16920 , n16919 );
nand ( n16921 , n3314 , n3008 );
and ( n16922 , n3179 , n16921 );
not ( n16923 , n184 );
not ( n16924 , n3063 );
or ( n16925 , n16923 , n16924 );
nand ( n16926 , n16925 , n3213 , n9130 );
nand ( n16927 , n185 , n16926 );
not ( n16928 , n3276 );
nand ( n16929 , n16928 , n184 );
not ( n16930 , n185 );
nand ( n16931 , n3243 , n9182 , n3432 );
nand ( n16932 , n16930 , n16931 );
nand ( n16933 , n16922 , n16927 , n16929 , n16932 );
nand ( n16934 , n3013 , n16933 );
not ( n16935 , n3258 );
not ( n16936 , n9194 );
not ( n16937 , n3068 );
nand ( n16938 , n16936 , n16937 , n3115 );
not ( n16939 , n16938 );
or ( n16940 , n16935 , n16939 );
nand ( n16941 , n16940 , n3253 );
not ( n16942 , n16941 );
and ( n16943 , n9134 , n3246 );
not ( n16944 , n3300 );
not ( n16945 , n3283 );
or ( n16946 , n16944 , n16945 );
nand ( n16947 , n16946 , n11169 );
not ( n16948 , n185 );
not ( n16949 , n16948 );
not ( n16950 , n8776 );
or ( n16951 , n16949 , n16950 );
nand ( n16952 , n16951 , n9215 );
nor ( n16953 , n16947 , n16952 );
and ( n16954 , n11165 , n3139 );
nor ( n16955 , n11109 , n8886 );
nand ( n16956 , n16953 , n16954 , n16955 );
and ( n16957 , n3013 , n16956 );
not ( n16958 , n3013 );
nand ( n16959 , n185 , n8805 );
not ( n16960 , n185 );
not ( n16961 , n182 );
not ( n16962 , n3167 );
or ( n16963 , n16961 , n16962 );
nand ( n16964 , n16963 , n3276 );
nand ( n16965 , n16960 , n16964 );
nand ( n16966 , n3266 , n16959 , n16965 );
and ( n16967 , n16958 , n16966 );
nor ( n16968 , n16957 , n16967 );
nand ( n16969 , n16942 , n16943 , n16968 );
nand ( n16970 , n187 , n16969 );
and ( n16971 , n16920 , n16934 , n16970 );
not ( n16972 , n16971 );
not ( n16973 , n3460 );
or ( n16974 , n3336 , n3325 );
nand ( n16975 , n16974 , n187 );
not ( n16976 , n3408 );
not ( n16977 , n3420 );
or ( n16978 , n16976 , n16977 );
nand ( n16979 , n16978 , n186 );
nand ( n16980 , n16973 , n3393 , n16975 , n16979 );
not ( n16981 , n16980 );
buf ( n16982 , n16981 );
not ( n16983 , n16982 );
and ( n16984 , n16972 , n16983 );
not ( n16985 , n16971 );
not ( n16986 , n16985 );
not ( n16987 , n16980 );
not ( n16988 , n16987 );
not ( n16989 , n16988 );
and ( n16990 , n16986 , n16989 );
nor ( n16991 , n16984 , n16990 );
not ( n16992 , n12558 );
not ( n16993 , n12674 );
and ( n16994 , n16992 , n16993 );
and ( n16995 , n12558 , n12674 );
nor ( n16996 , n16994 , n16995 );
and ( n16997 , n16991 , n16996 );
not ( n16998 , n16991 );
not ( n16999 , n16996 );
and ( n17000 , n16998 , n16999 );
nor ( n17001 , n16997 , n17000 );
not ( n17002 , n17001 );
or ( n17003 , n16876 , n17002 );
nand ( n17004 , n17003 , n2352 );
nor ( n17005 , n16875 , n17001 );
or ( n17006 , n17004 , n17005 );
not ( n17007 , n98 );
and ( n17008 , n315 , n17007 );
not ( n17009 , n315 );
and ( n17010 , n17009 , n98 );
nor ( n17011 , n17008 , n17010 );
or ( n17012 , n2352 , n17011 );
nand ( n17013 , n17006 , n17012 );
not ( n17014 , n320 );
not ( n17015 , n4296 );
or ( n17016 , n17014 , n17015 );
not ( n17017 , n320 );
nand ( n17018 , n17017 , n4297 );
nand ( n17019 , n17016 , n17018 );
buf ( n17020 , n13072 );
xnor ( n17021 , n17019 , n17020 );
nand ( n17022 , n12888 , n12907 , n12954 );
nor ( n17023 , n12842 , n17022 );
not ( n17024 , n17023 );
not ( n17025 , n5449 );
not ( n17026 , n169 );
not ( n17027 , n5369 );
nor ( n17028 , n17027 , n14932 );
nand ( n17029 , n17028 , n15826 , n5237 );
not ( n17030 , n17029 );
or ( n17031 , n17026 , n17030 );
not ( n17032 , n5326 );
not ( n17033 , n14999 );
or ( n17034 , n17032 , n17033 );
not ( n17035 , n167 );
nand ( n17036 , n17034 , n17035 );
nand ( n17037 , n17031 , n17036 );
not ( n17038 , n169 );
not ( n17039 , n17038 );
or ( n17040 , n5594 , n10288 );
nand ( n17041 , n17040 , n167 );
not ( n17042 , n167 );
nand ( n17043 , n17042 , n5342 );
nor ( n17044 , n14998 , n5615 );
nand ( n17045 , n14876 , n17041 , n17043 , n17044 );
not ( n17046 , n17045 );
or ( n17047 , n17039 , n17046 );
not ( n17048 , n10183 );
nand ( n17049 , n165 , n5405 );
nand ( n17050 , n10724 , n17049 , n14988 );
not ( n17051 , n17050 );
or ( n17052 , n17048 , n17051 );
nand ( n17053 , n17052 , n10738 );
not ( n17054 , n167 );
not ( n17055 , n5396 );
or ( n17056 , n17054 , n17055 );
nor ( n17057 , n5217 , n5375 );
nand ( n17058 , n17056 , n17057 );
nor ( n17059 , n17053 , n17058 );
nand ( n17060 , n17047 , n17059 );
nor ( n17061 , n17037 , n17060 );
not ( n17062 , n17061 );
and ( n17063 , n17025 , n17062 );
not ( n17064 , n167 );
nand ( n17065 , n17064 , n10250 );
and ( n17066 , n17065 , n14983 , n10762 );
not ( n17067 , n169 );
not ( n17068 , n17067 );
not ( n17069 , n167 );
nand ( n17070 , n17069 , n5413 );
not ( n17071 , n17070 );
and ( n17072 , n17068 , n17071 );
not ( n17073 , n5372 );
not ( n17074 , n5548 );
or ( n17075 , n17073 , n17074 );
not ( n17076 , n166 );
or ( n17077 , n17076 , n5504 );
nand ( n17078 , n17075 , n17077 );
and ( n17079 , n169 , n17078 );
nor ( n17080 , n17072 , n17079 );
nand ( n17081 , n17066 , n17080 );
nor ( n17082 , n17063 , n17081 );
not ( n17083 , n169 );
and ( n17084 , n5502 , n5623 );
nor ( n17085 , n17084 , n14874 );
and ( n17086 , n5245 , n14872 );
nor ( n17087 , n17086 , n5366 );
or ( n17088 , n14877 , n17087 );
nand ( n17089 , n17088 , n167 );
not ( n17090 , n167 );
not ( n17091 , n166 );
nand ( n17092 , n17091 , n5521 );
nand ( n17093 , n17092 , n10749 , n5549 );
nand ( n17094 , n17090 , n17093 );
nand ( n17095 , n17085 , n17089 , n17094 );
nand ( n17096 , n17083 , n17095 );
not ( n17097 , n169 );
not ( n17098 , n5502 );
not ( n17099 , n15774 );
or ( n17100 , n17098 , n17099 );
nand ( n17101 , n5372 , n5303 );
nand ( n17102 , n17100 , n17101 );
and ( n17103 , n17097 , n17102 );
not ( n17104 , n166 );
or ( n17105 , n17104 , n5406 );
nand ( n17106 , n166 , n5290 );
nand ( n17107 , n17105 , n17106 );
and ( n17108 , n167 , n17107 );
nor ( n17109 , n17103 , n17108 );
not ( n17110 , n167 );
nand ( n17111 , n17110 , n5472 );
not ( n17112 , n17111 );
nor ( n17113 , n5505 , n17112 );
nand ( n17114 , n5318 , n15753 );
and ( n17115 , n167 , n17114 );
nor ( n17116 , n5411 , n17049 );
nor ( n17117 , n17115 , n17116 );
and ( n17118 , n17070 , n17109 , n17113 , n17117 );
not ( n17119 , n17118 );
not ( n17120 , n169 );
not ( n17121 , n5367 );
not ( n17122 , n14872 );
not ( n17123 , n17122 );
or ( n17124 , n17121 , n17123 );
nand ( n17125 , n17124 , n5440 );
and ( n17126 , n17120 , n17125 );
not ( n17127 , n17120 );
not ( n17128 , n167 );
not ( n17129 , n17128 );
not ( n17130 , n166 );
nand ( n17131 , n17130 , n5457 );
nand ( n17132 , n17131 , n5257 , n5624 );
not ( n17133 , n17132 );
or ( n17134 , n17129 , n17133 );
not ( n17135 , n17106 );
nor ( n17136 , n17135 , n5493 );
nand ( n17137 , n17134 , n17136 );
not ( n17138 , n17137 );
not ( n17139 , n10294 );
not ( n17140 , n5441 );
or ( n17141 , n17139 , n17140 );
nand ( n17142 , n17141 , n167 );
not ( n17143 , n5485 );
nor ( n17144 , n17143 , n10250 );
nand ( n17145 , n17138 , n17142 , n5459 , n17144 );
and ( n17146 , n17127 , n17145 );
nor ( n17147 , n17126 , n17146 );
not ( n17148 , n17147 );
or ( n17149 , n17119 , n17148 );
nand ( n17150 , n17149 , n5449 );
nand ( n17151 , n17082 , n17096 , n17150 );
not ( n17152 , n17151 );
and ( n17153 , n17024 , n17152 );
and ( n17154 , n17023 , n17151 );
nor ( n17155 , n17153 , n17154 );
not ( n17156 , n17155 );
and ( n17157 , n10310 , n17156 );
not ( n17158 , n10310 );
and ( n17159 , n17158 , n17155 );
nor ( n17160 , n17157 , n17159 );
nor ( n17161 , n17021 , n17160 );
not ( n17162 , n17021 );
not ( n17163 , n17160 );
or ( n17164 , n17162 , n17163 );
nand ( n17165 , n17164 , n2352 );
or ( n17166 , n17161 , n17165 );
xnor ( n17167 , n320 , n321 );
or ( n17168 , n2352 , n17167 );
nand ( n17169 , n17166 , n17168 );
not ( n17170 , n301 );
not ( n17171 , n17170 );
not ( n17172 , n7089 );
or ( n17173 , n17171 , n17172 );
or ( n17174 , n17170 , n7107 );
nand ( n17175 , n17173 , n17174 );
not ( n17176 , n17175 );
nand ( n17177 , n130 , n15185 );
and ( n17178 , n17177 , n15271 );
not ( n17179 , n133 );
nor ( n17180 , n17178 , n17179 );
not ( n17181 , n17180 );
not ( n17182 , n133 );
not ( n17183 , n6922 );
not ( n17184 , n17183 );
not ( n17185 , n7208 );
or ( n17186 , n17184 , n17185 );
nand ( n17187 , n17186 , n6908 );
nand ( n17188 , n17182 , n17187 );
not ( n17189 , n6880 );
not ( n17190 , n132 );
nand ( n17191 , n17189 , n17190 );
nand ( n17192 , n132 , n6833 );
and ( n17193 , n133 , n17192 );
not ( n17194 , n133 );
and ( n17195 , n17194 , n7068 );
or ( n17196 , n17193 , n17195 );
nand ( n17197 , n17188 , n17191 , n17196 );
not ( n17198 , n17197 );
and ( n17199 , n17181 , n17198 );
not ( n17200 , n134 );
nor ( n17201 , n17199 , n17200 );
not ( n17202 , n17201 );
not ( n17203 , n134 );
not ( n17204 , n17203 );
not ( n17205 , n6853 );
and ( n17206 , n132 , n17205 );
nand ( n17207 , n6862 , n15200 );
not ( n17208 , n17207 );
nor ( n17209 , n17206 , n6890 , n17208 );
nand ( n17210 , n132 , n15184 );
nand ( n17211 , n132 , n7047 );
nand ( n17212 , n17210 , n6954 , n17211 );
nand ( n17213 , n133 , n17212 );
not ( n17214 , n7305 );
not ( n17215 , n6924 );
not ( n17216 , n7145 );
or ( n17217 , n17214 , n17215 , n17216 );
not ( n17218 , n133 );
nand ( n17219 , n17217 , n17218 );
nand ( n17220 , n17209 , n17213 , n17219 );
not ( n17221 , n17220 );
or ( n17222 , n17204 , n17221 );
not ( n17223 , n6892 );
and ( n17224 , n6968 , n15201 );
nor ( n17225 , n17224 , n132 , n15205 );
nor ( n17226 , n17223 , n17225 );
nand ( n17227 , n17222 , n17226 );
not ( n17228 , n17227 );
not ( n17229 , n15197 );
not ( n17230 , n17229 );
nor ( n17231 , n135 , n17230 );
not ( n17232 , n133 );
nand ( n17233 , n132 , n15176 );
nand ( n17234 , n15260 , n17233 , n7028 );
nand ( n17235 , n17232 , n17234 );
not ( n17236 , n7203 );
nand ( n17237 , n132 , n6855 );
not ( n17238 , n17237 );
or ( n17239 , n17236 , n17238 );
nand ( n17240 , n17239 , n133 );
nand ( n17241 , n17235 , n7151 , n17240 );
nand ( n17242 , n134 , n17241 );
not ( n17243 , n15228 );
not ( n17244 , n133 );
nand ( n17245 , n17243 , n17244 );
not ( n17246 , n134 );
not ( n17247 , n7206 );
not ( n17248 , n7002 );
or ( n17249 , n17247 , n17248 );
nand ( n17250 , n17249 , n6954 );
and ( n17251 , n17246 , n17250 );
not ( n17252 , n15271 );
and ( n17253 , n6906 , n17252 );
nor ( n17254 , n17251 , n17253 );
nand ( n17255 , n17231 , n17242 , n17245 , n17254 );
not ( n17256 , n133 );
not ( n17257 , n7208 );
or ( n17258 , n6841 , n17257 );
not ( n17259 , n6852 );
nand ( n17260 , n17258 , n17259 );
and ( n17261 , n17256 , n17260 );
and ( n17262 , n133 , n15172 );
nor ( n17263 , n17261 , n17262 );
nand ( n17264 , n15252 , n17263 );
and ( n17265 , n134 , n17264 );
not ( n17266 , n6906 );
not ( n17267 , n6933 );
nand ( n17268 , n7129 , n17267 , n6913 );
not ( n17269 , n17268 );
or ( n17270 , n17266 , n17269 );
nand ( n17271 , n17270 , n15237 );
nor ( n17272 , n17265 , n17271 );
nand ( n17273 , n6827 , n15282 );
not ( n17274 , n134 );
not ( n17275 , n133 );
not ( n17276 , n6946 );
or ( n17277 , n17275 , n17276 );
nand ( n17278 , n17277 , n6999 );
not ( n17279 , n133 );
not ( n17280 , n17279 );
not ( n17281 , n6990 );
not ( n17282 , n17281 );
or ( n17283 , n17280 , n17282 );
nand ( n17284 , n133 , n15264 );
nand ( n17285 , n17283 , n17284 );
nor ( n17286 , n17278 , n17285 );
not ( n17287 , n6901 );
and ( n17288 , n17287 , n7121 );
not ( n17289 , n7127 );
not ( n17290 , n132 );
nand ( n17291 , n17289 , n17290 );
not ( n17292 , n133 );
nand ( n17293 , n17292 , n15270 );
nand ( n17294 , n17286 , n17288 , n17291 , n17293 );
and ( n17295 , n17274 , n17294 );
not ( n17296 , n15243 );
nor ( n17297 , n17295 , n17296 );
nand ( n17298 , n17272 , n135 , n17273 , n17297 );
nand ( n17299 , n17255 , n17298 );
nand ( n17300 , n17202 , n17228 , n17299 );
not ( n17301 , n17300 );
not ( n17302 , n17301 );
not ( n17303 , n7317 );
or ( n17304 , n17302 , n17303 );
not ( n17305 , n17201 );
nand ( n17306 , n17228 , n17305 , n17299 );
not ( n17307 , n17306 );
or ( n17308 , n17307 , n7317 );
nand ( n17309 , n17304 , n17308 );
not ( n17310 , n17309 );
or ( n17311 , n17176 , n17310 );
or ( n17312 , n17175 , n17309 );
nand ( n17313 , n17311 , n17312 );
not ( n17314 , n17313 );
not ( n17315 , n12019 );
buf ( n17316 , n11579 );
not ( n17317 , n17316 );
and ( n17318 , n17315 , n17317 );
not ( n17319 , n11580 );
and ( n17320 , n12023 , n17319 );
nor ( n17321 , n17318 , n17320 );
not ( n17322 , n17321 );
not ( n17323 , n11755 );
not ( n17324 , n17323 );
not ( n17325 , n7325 );
or ( n17326 , n116 , n11655 );
or ( n17327 , n7478 , n11669 );
nand ( n17328 , n17326 , n17327 );
not ( n17329 , n117 );
not ( n17330 , n17329 );
nand ( n17331 , n7364 , n15589 );
not ( n17332 , n17331 );
or ( n17333 , n17330 , n17332 );
nand ( n17334 , n117 , n7587 );
nand ( n17335 , n17333 , n17334 );
nor ( n17336 , n17328 , n17335 );
not ( n17337 , n11847 );
and ( n17338 , n117 , n115 , n7343 );
nor ( n17339 , n17338 , n118 );
not ( n17340 , n7531 );
and ( n17341 , n17340 , n7542 );
nor ( n17342 , n17341 , n7387 );
nor ( n17343 , n7409 , n17342 );
not ( n17344 , n7375 );
nand ( n17345 , n7485 , n17344 );
nand ( n17346 , n17337 , n17339 , n17343 , n17345 );
not ( n17347 , n11669 );
not ( n17348 , n116 );
not ( n17349 , n7579 );
nand ( n17350 , n17348 , n17349 );
not ( n17351 , n17350 );
or ( n17352 , n17347 , n17351 );
nand ( n17353 , n17352 , n117 );
not ( n17354 , n118 );
nor ( n17355 , n17354 , n7458 );
nor ( n17356 , n117 , n15675 );
nand ( n17357 , n7504 , n11649 );
nor ( n17358 , n17356 , n17357 );
nand ( n17359 , n17353 , n17355 , n17358 );
nand ( n17360 , n17346 , n17359 );
nand ( n17361 , n17336 , n17360 );
not ( n17362 , n17361 );
or ( n17363 , n17325 , n17362 );
not ( n17364 , n7431 );
not ( n17365 , n7498 );
or ( n17366 , n17364 , n17365 );
nand ( n17367 , n17366 , n7523 );
and ( n17368 , n11618 , n17367 );
nor ( n17369 , n117 , n118 );
not ( n17370 , n7544 );
and ( n17371 , n17369 , n17370 );
nor ( n17372 , n17368 , n17371 );
nand ( n17373 , n17363 , n17372 );
not ( n17374 , n17373 );
nand ( n17375 , n7562 , n11601 , n15675 );
nand ( n17376 , n11597 , n17375 );
nand ( n17377 , n17376 , n7546 , n11629 );
nand ( n17378 , n118 , n17377 );
not ( n17379 , n15569 );
nand ( n17380 , n11685 , n17379 );
and ( n17381 , n17380 , n15632 , n15581 );
not ( n17382 , n17381 );
nand ( n17383 , n11714 , n11833 );
nand ( n17384 , n115 , n17383 );
and ( n17385 , n11592 , n17384 );
not ( n17386 , n117 );
nor ( n17387 , n17385 , n17386 );
not ( n17388 , n17387 );
not ( n17389 , n117 );
not ( n17390 , n11847 );
nand ( n17391 , n116 , n11712 );
nand ( n17392 , n17390 , n17391 , n15608 );
nand ( n17393 , n17389 , n17392 );
nand ( n17394 , n11845 , n7521 );
not ( n17395 , n17394 );
nand ( n17396 , n11610 , n7374 );
not ( n17397 , n17396 );
not ( n17398 , n112 );
nor ( n17399 , n17398 , n116 , n114 );
nand ( n17400 , n7390 , n7370 );
or ( n17401 , n17399 , n17400 );
nand ( n17402 , n17401 , n117 );
nand ( n17403 , n17395 , n17397 , n15578 , n17402 );
nand ( n17404 , n118 , n17403 );
nand ( n17405 , n17388 , n17393 , n17404 );
not ( n17406 , n11883 );
not ( n17407 , n7591 );
or ( n17408 , n17406 , n17407 );
not ( n17409 , n117 );
nand ( n17410 , n17408 , n17409 );
nand ( n17411 , n17410 , n7610 , n7359 , n11734 );
nand ( n17412 , n117 , n7503 );
nand ( n17413 , n117 , n11743 );
nand ( n17414 , n7431 , n7348 );
nand ( n17415 , n17412 , n17413 , n17414 );
nor ( n17416 , n17411 , n17415 );
or ( n17417 , n118 , n17416 );
not ( n17418 , n11698 );
nand ( n17419 , n17417 , n17418 );
nor ( n17420 , n17405 , n17419 );
or ( n17421 , n17420 , n7325 );
not ( n17422 , n118 );
not ( n17423 , n117 );
not ( n17424 , n7561 );
not ( n17425 , n17424 );
or ( n17426 , n17423 , n17425 );
nand ( n17427 , n7388 , n7490 );
nand ( n17428 , n17426 , n17427 );
nand ( n17429 , n17422 , n17428 );
nand ( n17430 , n17421 , n17429 );
nor ( n17431 , n17382 , n17430 );
and ( n17432 , n17374 , n17378 , n17431 );
not ( n17433 , n17432 );
and ( n17434 , n17324 , n17433 );
and ( n17435 , n11756 , n17432 );
nor ( n17436 , n17434 , n17435 );
not ( n17437 , n17436 );
not ( n17438 , n17437 );
or ( n17439 , n17322 , n17438 );
or ( n17440 , n17321 , n17437 );
nand ( n17441 , n17439 , n17440 );
not ( n17442 , n17441 );
nor ( n17443 , n17314 , n17442 );
or ( n17444 , n17313 , n17441 );
nand ( n17445 , n17444 , n2352 );
or ( n17446 , n17443 , n17445 );
and ( n17447 , n302 , n17170 );
not ( n17448 , n302 );
and ( n17449 , n17448 , n301 );
nor ( n17450 , n17447 , n17449 );
or ( n17451 , n2352 , n17450 );
nand ( n17452 , n17446 , n17451 );
not ( n17453 , n1 );
xor ( n17454 , n332 , n333 );
not ( n17455 , n17454 );
or ( n17456 , n17453 , n17455 );
xnor ( n17457 , n332 , n15035 );
not ( n17458 , n144 );
or ( n17459 , n141 , n6662 );
nand ( n17460 , n17459 , n11258 , n11324 );
not ( n17461 , n17460 );
or ( n17462 , n17458 , n17461 );
not ( n17463 , n141 );
not ( n17464 , n142 );
not ( n17465 , n11340 );
or ( n17466 , n17464 , n17465 );
nand ( n17467 , n17466 , n11965 );
nand ( n17468 , n17463 , n17467 );
nand ( n17469 , n17462 , n17468 );
nand ( n17470 , n6757 , n6728 );
nor ( n17471 , n17469 , n17470 );
not ( n17472 , n11366 );
not ( n17473 , n11531 );
or ( n17474 , n17472 , n17473 );
not ( n17475 , n141 );
nand ( n17476 , n17474 , n17475 );
not ( n17477 , n11440 );
nor ( n17478 , n17477 , n6727 );
nand ( n17479 , n17478 , n11294 , n15072 );
nand ( n17480 , n141 , n17479 );
not ( n17481 , n6707 );
or ( n17482 , n17481 , n11519 );
nand ( n17483 , n6588 , n11328 );
and ( n17484 , n17483 , n11423 );
nand ( n17485 , n17482 , n17484 );
not ( n17486 , n141 );
nand ( n17487 , n15067 , n6731 , n6672 );
not ( n17488 , n17487 );
or ( n17489 , n17486 , n17488 );
nand ( n17490 , n142 , n6613 );
nand ( n17491 , n17489 , n17490 );
or ( n17492 , n17485 , n17491 );
not ( n17493 , n144 );
nand ( n17494 , n17492 , n17493 );
and ( n17495 , n17471 , n17476 , n17480 , n17494 );
or ( n17496 , n17495 , n6808 );
and ( n17497 , n141 , n11548 );
not ( n17498 , n141 );
not ( n17499 , n140 );
or ( n17500 , n17499 , n11964 );
and ( n17501 , n17498 , n17500 );
or ( n17502 , n17497 , n17501 );
nand ( n17503 , n17496 , n17502 );
nand ( n17504 , n11931 , n6641 );
and ( n17505 , n17504 , n11302 , n11294 );
or ( n17506 , n141 , n17505 );
nand ( n17507 , n6683 , n11915 );
nand ( n17508 , n17507 , n141 , n11328 );
nand ( n17509 , n17506 , n17508 );
nand ( n17510 , n6796 , n11246 );
and ( n17511 , n17510 , n6764 , n11507 );
nand ( n17512 , n11264 , n6701 );
nand ( n17513 , n17511 , n17500 , n17512 );
nand ( n17514 , n144 , n17513 );
or ( n17515 , n142 , n6539 );
nand ( n17516 , n17515 , n6788 );
nand ( n17517 , n11555 , n17516 );
not ( n17518 , n144 );
not ( n17519 , n142 );
not ( n17520 , n17519 );
not ( n17521 , n11476 );
or ( n17522 , n17520 , n17521 );
nand ( n17523 , n17522 , n6550 );
nand ( n17524 , n17518 , n17523 );
nand ( n17525 , n17514 , n17517 , n17524 );
or ( n17526 , n17509 , n17525 );
nand ( n17527 , n17526 , n6808 );
not ( n17528 , n144 );
not ( n17529 , n141 );
not ( n17530 , n142 );
not ( n17531 , n11281 );
nand ( n17532 , n17530 , n17531 );
nand ( n17533 , n17532 , n6720 , n6677 );
and ( n17534 , n17529 , n17533 );
not ( n17535 , n17529 );
nand ( n17536 , n11330 , n6698 );
and ( n17537 , n17535 , n17536 );
nor ( n17538 , n17534 , n17537 );
nand ( n17539 , n17538 , n15074 , n12009 );
nand ( n17540 , n17528 , n17539 );
not ( n17541 , n6642 );
nand ( n17542 , n6575 , n6656 );
and ( n17543 , n141 , n17542 );
not ( n17544 , n141 );
and ( n17545 , n17544 , n11318 );
nor ( n17546 , n17543 , n17545 );
nor ( n17547 , n17541 , n17546 );
not ( n17548 , n11959 );
nand ( n17549 , n17547 , n11337 , n17548 );
nand ( n17550 , n144 , n17549 );
nand ( n17551 , n17527 , n17540 , n17550 );
nor ( n17552 , n17503 , n17551 );
not ( n17553 , n17552 );
not ( n17554 , n17553 );
not ( n17555 , n15616 );
not ( n17556 , n117 );
not ( n17557 , n17556 );
not ( n17558 , n116 );
nand ( n17559 , n17558 , n11715 );
nand ( n17560 , n17559 , n7472 , n7350 );
not ( n17561 , n17560 );
or ( n17562 , n17557 , n17561 );
nand ( n17563 , n17562 , n11699 );
or ( n17564 , n17555 , n17563 );
not ( n17565 , n118 );
nand ( n17566 , n17564 , n17565 );
and ( n17567 , n117 , n11788 );
not ( n17568 , n117 );
not ( n17569 , n7542 );
nand ( n17570 , n7468 , n17569 );
and ( n17571 , n17568 , n17570 );
or ( n17572 , n17567 , n17571 );
not ( n17573 , n17414 );
not ( n17574 , n7613 );
or ( n17575 , n17573 , n17574 );
nand ( n17576 , n17575 , n11778 );
not ( n17577 , n7557 );
nand ( n17578 , n17577 , n7461 );
nor ( n17579 , n7511 , n11714 );
nand ( n17580 , n117 , n17579 );
not ( n17581 , n15645 );
nand ( n17582 , n17581 , n11597 );
nand ( n17583 , n17580 , n17582 , n17412 );
or ( n17584 , n17578 , n17583 );
nand ( n17585 , n17584 , n118 );
and ( n17586 , n17566 , n17572 , n17576 , n17585 );
not ( n17587 , n117 );
not ( n17588 , n116 );
not ( n17589 , n15650 );
nand ( n17590 , n17588 , n17589 );
nand ( n17591 , n17391 , n17590 , n15610 );
nand ( n17592 , n17587 , n17591 );
not ( n17593 , n118 );
not ( n17594 , n116 );
not ( n17595 , n17594 );
nand ( n17596 , n11655 , n7457 );
not ( n17597 , n17596 );
or ( n17598 , n17595 , n17597 );
nand ( n17599 , n17598 , n7540 );
nand ( n17600 , n17593 , n17599 );
nand ( n17601 , n7450 , n11631 );
nand ( n17602 , n117 , n7498 , n17601 );
not ( n17603 , n118 );
and ( n17604 , n11677 , n17570 );
nand ( n17605 , n11630 , n11597 );
nand ( n17606 , n117 , n7608 );
nand ( n17607 , n17604 , n17605 , n7419 , n17606 );
not ( n17608 , n17607 );
or ( n17609 , n17603 , n17608 );
or ( n17610 , n116 , n17340 );
nand ( n17611 , n17610 , n7370 );
nand ( n17612 , n11778 , n17611 );
nand ( n17613 , n17609 , n17612 );
not ( n17614 , n17613 );
nand ( n17615 , n17592 , n17600 , n17602 , n17614 );
nand ( n17616 , n7325 , n17615 );
not ( n17617 , n117 );
nand ( n17618 , n17617 , n7431 );
nand ( n17619 , n17618 , n11716 , n15578 );
nand ( n17620 , n118 , n17619 );
or ( n17621 , n11864 , n11648 );
not ( n17622 , n117 );
nand ( n17623 , n17621 , n17622 );
not ( n17624 , n7380 );
nor ( n17625 , n17624 , n11896 );
nand ( n17626 , n17625 , n15705 , n15608 );
nand ( n17627 , n117 , n17626 );
nand ( n17628 , n17620 , n17623 , n17627 );
not ( n17629 , n17628 );
not ( n17630 , n17629 );
not ( n17631 , n15690 );
nor ( n17632 , n17631 , n7446 );
not ( n17633 , n117 );
not ( n17634 , n116 );
or ( n17635 , n17634 , n15618 );
nand ( n17636 , n17635 , n11670 );
nand ( n17637 , n17633 , n17636 );
not ( n17638 , n7551 );
not ( n17639 , n17638 );
nand ( n17640 , n17639 , n116 );
nand ( n17641 , n11744 , n17640 );
nand ( n17642 , n7329 , n7498 );
not ( n17643 , n7567 );
nand ( n17644 , n11597 , n17643 );
nand ( n17645 , n15624 , n7579 , n7335 );
nand ( n17646 , n117 , n17645 );
nand ( n17647 , n17642 , n17644 , n17646 );
or ( n17648 , n17641 , n17647 );
not ( n17649 , n118 );
nand ( n17650 , n17648 , n17649 );
nand ( n17651 , n17632 , n17637 , n17650 );
or ( n17652 , n17630 , n17651 );
nand ( n17653 , n17652 , n119 );
and ( n17654 , n17586 , n17616 , n17653 );
not ( n17655 , n17654 );
and ( n17656 , n17554 , n17655 );
and ( n17657 , n17553 , n17654 );
nor ( n17658 , n17656 , n17657 );
or ( n17659 , n17658 , n15442 );
nand ( n17660 , n17658 , n15732 );
nand ( n17661 , n17659 , n17660 );
nor ( n17662 , n17457 , n17661 );
not ( n17663 , n17662 );
nand ( n17664 , n17457 , n17661 );
nand ( n17665 , n17663 , n17664 , n2352 );
nand ( n17666 , n17456 , n17665 );
and ( n17667 , n334 , n12187 );
not ( n17668 , n334 );
not ( n17669 , n12187 );
and ( n17670 , n17668 , n17669 );
nor ( n17671 , n17667 , n17670 );
not ( n17672 , n17671 );
not ( n17673 , n10913 );
not ( n17674 , n14707 );
and ( n17675 , n17673 , n17674 );
not ( n17676 , n10927 );
and ( n17677 , n17676 , n14707 );
nor ( n17678 , n17675 , n17677 );
not ( n17679 , n17678 );
or ( n17680 , n17672 , n17679 );
or ( n17681 , n17671 , n17678 );
nand ( n17682 , n17680 , n17681 );
not ( n17683 , n17682 );
not ( n17684 , n14861 );
not ( n17685 , n10659 );
not ( n17686 , n17685 );
not ( n17687 , n17686 );
or ( n17688 , n17684 , n17687 );
not ( n17689 , n17685 );
not ( n17690 , n12300 );
or ( n17691 , n17689 , n17690 );
nand ( n17692 , n17688 , n17691 );
not ( n17693 , n17692 );
not ( n17694 , n10802 );
or ( n17695 , n17693 , n17694 );
or ( n17696 , n17692 , n10802 );
nand ( n17697 , n17695 , n17696 );
not ( n17698 , n17697 );
nor ( n17699 , n17683 , n17698 );
or ( n17700 , n17697 , n17682 );
nand ( n17701 , n17700 , n2352 );
or ( n17702 , n17699 , n17701 );
xnor ( n17703 , n334 , n335 );
or ( n17704 , n2352 , n17703 );
nand ( n17705 , n17702 , n17704 );
not ( n17706 , n303 );
and ( n17707 , n304 , n17706 );
not ( n17708 , n304 );
and ( n17709 , n17708 , n303 );
nor ( n17710 , n17707 , n17709 );
or ( n17711 , n2352 , n17710 );
not ( n17712 , n17706 );
not ( n17713 , n134 );
nand ( n17714 , n17237 , n7185 );
not ( n17715 , n17714 );
not ( n17716 , n131 );
nand ( n17717 , n17716 , n15182 );
not ( n17718 , n17717 );
not ( n17719 , n132 );
and ( n17720 , n17719 , n17183 );
not ( n17721 , n17719 );
and ( n17722 , n17721 , n7170 );
nor ( n17723 , n17720 , n17722 );
not ( n17724 , n17723 );
or ( n17725 , n17718 , n17724 );
not ( n17726 , n133 );
nand ( n17727 , n17725 , n17726 );
not ( n17728 , n6952 );
not ( n17729 , n17728 );
not ( n17730 , n7118 );
or ( n17731 , n17729 , n17730 );
nand ( n17732 , n17731 , n133 );
nand ( n17733 , n17715 , n17727 , n17732 , n7309 );
not ( n17734 , n17733 );
or ( n17735 , n17713 , n17734 );
nand ( n17736 , n17735 , n15250 );
not ( n17737 , n17736 );
not ( n17738 , n6991 );
not ( n17739 , n15212 );
not ( n17740 , n15273 );
or ( n17741 , n17739 , n17740 );
nand ( n17742 , n17741 , n133 );
and ( n17743 , n15198 , n17738 , n17742 );
or ( n17744 , n133 , n17211 );
nand ( n17745 , n17273 , n6914 );
not ( n17746 , n133 );
or ( n17747 , n17746 , n6882 );
not ( n17748 , n6913 );
not ( n17749 , n6880 );
nand ( n17750 , n15185 , n17749 );
not ( n17751 , n17750 );
or ( n17752 , n17748 , n17751 );
not ( n17753 , n133 );
nand ( n17754 , n17752 , n17753 );
nand ( n17755 , n17747 , n17211 , n17754 );
or ( n17756 , n17745 , n17755 );
not ( n17757 , n134 );
nand ( n17758 , n17756 , n17757 );
nand ( n17759 , n17737 , n17743 , n17744 , n17758 );
nand ( n17760 , n7099 , n17759 );
not ( n17761 , n134 );
not ( n17762 , n133 );
not ( n17763 , n17762 );
nand ( n17764 , n7139 , n7163 , n6824 );
not ( n17765 , n17764 );
or ( n17766 , n17763 , n17765 );
and ( n17767 , n6846 , n15292 );
nand ( n17768 , n17766 , n17767 );
nand ( n17769 , n17761 , n17768 );
not ( n17770 , n7178 );
not ( n17771 , n132 );
not ( n17772 , n6917 );
nand ( n17773 , n17771 , n17772 );
nand ( n17774 , n17773 , n17738 , n7041 );
not ( n17775 , n17774 );
or ( n17776 , n17770 , n17775 );
not ( n17777 , n6847 );
nor ( n17778 , n17777 , n7135 );
nand ( n17779 , n17776 , n17778 );
not ( n17780 , n17779 );
buf ( n17781 , n7156 );
not ( n17782 , n17781 );
or ( n17783 , n7181 , n6909 );
nand ( n17784 , n17783 , n132 );
not ( n17785 , n17784 );
or ( n17786 , n17782 , n17785 );
nand ( n17787 , n17786 , n7195 );
not ( n17788 , n133 );
not ( n17789 , n17788 );
not ( n17790 , n6982 );
not ( n17791 , n17291 );
nor ( n17792 , n17790 , n17791 );
not ( n17793 , n132 );
not ( n17794 , n7243 );
nand ( n17795 , n17793 , n17794 );
nand ( n17796 , n17792 , n17795 , n7134 );
not ( n17797 , n17796 );
or ( n17798 , n17789 , n17797 );
nand ( n17799 , n7002 , n15218 );
nand ( n17800 , n17798 , n17799 );
nand ( n17801 , n134 , n17800 );
and ( n17802 , n17780 , n17787 , n17801 );
not ( n17803 , n134 );
not ( n17804 , n17803 );
nand ( n17805 , n6924 , n6832 );
not ( n17806 , n17805 );
not ( n17807 , n6923 );
or ( n17808 , n133 , n17807 );
not ( n17809 , n132 );
nand ( n17810 , n17809 , n7064 );
nand ( n17811 , n6840 , n7206 );
nand ( n17812 , n17806 , n17808 , n17810 , n17811 );
not ( n17813 , n17812 );
or ( n17814 , n17804 , n17813 );
nand ( n17815 , n17814 , n17781 );
not ( n17816 , n17815 );
not ( n17817 , n133 );
not ( n17818 , n17817 );
and ( n17819 , n7151 , n15283 );
not ( n17820 , n6833 );
nand ( n17821 , n17819 , n7129 , n17820 );
not ( n17822 , n17821 );
or ( n17823 , n17818 , n17822 );
not ( n17824 , n132 );
nand ( n17825 , n17824 , n15247 );
nand ( n17826 , n17823 , n17825 );
not ( n17827 , n17826 );
not ( n17828 , n133 );
or ( n17829 , n17828 , n17191 );
not ( n17830 , n6938 );
not ( n17831 , n7170 );
nand ( n17832 , n17830 , n17831 , n17233 );
nand ( n17833 , n133 , n17832 );
nand ( n17834 , n17833 , n6908 , n7068 );
nand ( n17835 , n134 , n17834 );
nand ( n17836 , n17816 , n17827 , n17829 , n17835 );
nand ( n17837 , n135 , n17836 );
nand ( n17838 , n17760 , n17769 , n17802 , n17837 );
not ( n17839 , n17838 );
not ( n17840 , n17839 );
or ( n17841 , n17712 , n17840 );
or ( n17842 , n17706 , n17839 );
nand ( n17843 , n17841 , n17842 );
and ( n17844 , n15158 , n17319 );
not ( n17845 , n15158 );
and ( n17846 , n17845 , n11573 );
nor ( n17847 , n17844 , n17846 );
and ( n17848 , n17843 , n17847 );
not ( n17849 , n17843 );
not ( n17850 , n17847 );
and ( n17851 , n17849 , n17850 );
nor ( n17852 , n17848 , n17851 );
not ( n17853 , n17852 );
not ( n17854 , n17586 );
not ( n17855 , n7325 );
not ( n17856 , n17615 );
or ( n17857 , n17855 , n17856 );
and ( n17858 , n17629 , n17632 , n17637 , n17650 );
or ( n17859 , n7325 , n17858 );
nand ( n17860 , n17857 , n17859 );
nor ( n17861 , n17854 , n17860 );
buf ( n17862 , n17861 );
not ( n17863 , n17862 );
not ( n17864 , n15565 );
or ( n17865 , n17863 , n17864 );
or ( n17866 , n17862 , n15565 );
nand ( n17867 , n17865 , n17866 );
nor ( n17868 , n17551 , n17503 );
not ( n17869 , n17868 );
and ( n17870 , n17869 , n11913 );
not ( n17871 , n17869 );
not ( n17872 , n11913 );
and ( n17873 , n17871 , n17872 );
nor ( n17874 , n17870 , n17873 );
and ( n17875 , n17867 , n17874 );
not ( n17876 , n17867 );
not ( n17877 , n17874 );
and ( n17878 , n17876 , n17877 );
nor ( n17879 , n17875 , n17878 );
not ( n17880 , n17879 );
nand ( n17881 , n17853 , n17880 );
nand ( n17882 , n17852 , n17879 );
nand ( n17883 , n17881 , n2352 , n17882 );
nand ( n17884 , n17711 , n17883 );
not ( n17885 , n309 );
and ( n17886 , n310 , n17885 );
not ( n17887 , n310 );
and ( n17888 , n17887 , n309 );
nor ( n17889 , n17886 , n17888 );
or ( n17890 , n2352 , n17889 );
not ( n17891 , n135 );
and ( n17892 , n17237 , n6882 , n15219 );
nor ( n17893 , n17892 , n133 );
not ( n17894 , n17893 );
or ( n17895 , n130 , n17257 );
nand ( n17896 , n17895 , n7046 );
nand ( n17897 , n133 , n17896 );
or ( n17898 , n128 , n6872 );
nand ( n17899 , n17898 , n7066 );
nand ( n17900 , n133 , n17899 );
not ( n17901 , n6856 );
not ( n17902 , n7303 );
or ( n17903 , n17901 , n17902 );
not ( n17904 , n133 );
nand ( n17905 , n17903 , n17904 );
nand ( n17906 , n17284 , n17905 );
not ( n17907 , n17906 );
nand ( n17908 , n17907 , n15228 , n6824 );
and ( n17909 , n134 , n17908 );
not ( n17910 , n6901 );
nand ( n17911 , n17910 , n15165 );
not ( n17912 , n133 );
nand ( n17913 , n17912 , n7138 );
nand ( n17914 , n132 , n15190 );
nand ( n17915 , n17913 , n17914 , n6888 );
nor ( n17916 , n17911 , n17915 );
nor ( n17917 , n134 , n17916 );
nor ( n17918 , n17909 , n17917 );
nand ( n17919 , n17894 , n17897 , n17900 , n17918 );
not ( n17920 , n17919 );
or ( n17921 , n17891 , n17920 );
not ( n17922 , n134 );
not ( n17923 , n17922 );
and ( n17924 , n6862 , n15282 );
and ( n17925 , n133 , n7181 );
nor ( n17926 , n17924 , n17925 );
not ( n17927 , n132 );
nor ( n17928 , n17927 , n15171 );
not ( n17929 , n17928 );
nand ( n17930 , n17926 , n7110 , n17929 );
not ( n17931 , n17930 );
or ( n17932 , n17923 , n17931 );
not ( n17933 , n132 );
not ( n17934 , n17933 );
not ( n17935 , n7231 );
or ( n17936 , n17934 , n17935 );
nand ( n17937 , n17936 , n7276 );
nand ( n17938 , n133 , n17937 );
nand ( n17939 , n17932 , n17938 );
not ( n17940 , n17939 );
or ( n17941 , n133 , n17781 );
nand ( n17942 , n6999 , n7036 );
not ( n17943 , n133 );
not ( n17944 , n17943 );
not ( n17945 , n132 );
nand ( n17946 , n17945 , n6966 );
nand ( n17947 , n17946 , n15196 , n15290 );
not ( n17948 , n17947 );
or ( n17949 , n17944 , n17948 );
not ( n17950 , n6970 );
nand ( n17951 , n17950 , n6827 );
nand ( n17952 , n17949 , n17951 );
or ( n17953 , n17942 , n17952 );
nand ( n17954 , n17953 , n134 );
nand ( n17955 , n17940 , n17941 , n15243 , n17954 );
and ( n17956 , n7099 , n17955 );
not ( n17957 , n133 );
not ( n17958 , n17192 );
and ( n17959 , n17957 , n17958 );
and ( n17960 , n6906 , n7181 );
nor ( n17961 , n17959 , n17960 );
not ( n17962 , n7189 );
not ( n17963 , n133 );
nand ( n17964 , n7169 , n6968 );
nand ( n17965 , n132 , n17964 );
nand ( n17966 , n17965 , n7072 , n15219 );
nand ( n17967 , n17963 , n17966 );
nand ( n17968 , n133 , n7258 );
nand ( n17969 , n133 , n7285 );
and ( n17970 , n17968 , n17969 , n6891 );
nand ( n17971 , n17962 , n17967 , n17970 );
and ( n17972 , n134 , n17971 );
not ( n17973 , n134 );
nand ( n17974 , n7145 , n15243 );
not ( n17975 , n17974 );
not ( n17976 , n133 );
not ( n17977 , n132 );
nand ( n17978 , n17977 , n7170 );
nand ( n17979 , n17978 , n17191 , n17211 );
nand ( n17980 , n17976 , n17979 );
not ( n17981 , n7244 );
or ( n17982 , n6840 , n7013 );
nand ( n17983 , n17982 , n6916 );
nand ( n17984 , n17981 , n17291 , n7309 , n17983 );
nand ( n17985 , n133 , n17984 );
nand ( n17986 , n17975 , n17980 , n17985 );
and ( n17987 , n17973 , n17986 );
nor ( n17988 , n17972 , n17987 );
nand ( n17989 , n17961 , n17988 );
nor ( n17990 , n17956 , n17989 );
nand ( n17991 , n17921 , n17990 );
not ( n17992 , n17991 );
not ( n17993 , n17992 );
not ( n17994 , n17885 );
and ( n17995 , n17993 , n17994 );
not ( n17996 , n17991 );
and ( n17997 , n17885 , n17996 );
nor ( n17998 , n17995 , n17997 );
not ( n17999 , n17998 );
not ( n18000 , n7317 );
not ( n18001 , n18000 );
not ( n18002 , n7107 );
or ( n18003 , n18001 , n18002 );
not ( n18004 , n7317 );
or ( n18005 , n18004 , n7107 );
nand ( n18006 , n18003 , n18005 );
not ( n18007 , n18006 );
or ( n18008 , n17999 , n18007 );
or ( n18009 , n17998 , n18006 );
nand ( n18010 , n18008 , n18009 );
not ( n18011 , n7912 );
not ( n18012 , n18011 );
not ( n18013 , n11583 );
not ( n18014 , n18013 );
or ( n18015 , n18012 , n18014 );
not ( n18016 , n7912 );
not ( n18017 , n11583 );
or ( n18018 , n18016 , n18017 );
nand ( n18019 , n18015 , n18018 );
or ( n18020 , n18010 , n18019 );
nand ( n18021 , n18010 , n18019 );
nand ( n18022 , n18020 , n18021 , n2352 );
nand ( n18023 , n17890 , n18022 );
not ( n18024 , n12753 );
not ( n18025 , n12822 );
nand ( n18026 , n18024 , n18025 );
xor ( n18027 , n326 , n18026 );
xnor ( n18028 , n18027 , n9806 );
not ( n18029 , n14700 );
not ( n18030 , n18029 );
not ( n18031 , n17156 );
or ( n18032 , n18030 , n18031 );
or ( n18033 , n18029 , n17156 );
nand ( n18034 , n18032 , n18033 );
nor ( n18035 , n18028 , n18034 );
not ( n18036 , n18028 );
not ( n18037 , n18034 );
or ( n18038 , n18036 , n18037 );
nand ( n18039 , n18038 , n2352 );
or ( n18040 , n18035 , n18039 );
xnor ( n18041 , n326 , n327 );
or ( n18042 , n2352 , n18041 );
nand ( n18043 , n18040 , n18042 );
not ( n18044 , n344 );
and ( n18045 , n345 , n18044 );
not ( n18046 , n345 );
and ( n18047 , n18046 , n344 );
nor ( n18048 , n18045 , n18047 );
or ( n18049 , n2352 , n18048 );
and ( n18050 , n15712 , n15158 );
not ( n18051 , n15712 );
and ( n18052 , n18051 , n15157 );
nor ( n18053 , n18050 , n18052 );
and ( n18054 , n17838 , n344 );
not ( n18055 , n17838 );
and ( n18056 , n18055 , n18044 );
nor ( n18057 , n18054 , n18056 );
and ( n18058 , n18053 , n18057 );
not ( n18059 , n18053 );
not ( n18060 , n18057 );
and ( n18061 , n18059 , n18060 );
nor ( n18062 , n18058 , n18061 );
not ( n18063 , n18062 );
not ( n18064 , n17862 );
not ( n18065 , n11913 );
not ( n18066 , n18065 );
or ( n18067 , n18064 , n18066 );
or ( n18068 , n17862 , n17872 );
nand ( n18069 , n18067 , n18068 );
and ( n18070 , n18069 , n15732 );
not ( n18071 , n18069 );
not ( n18072 , n15442 );
and ( n18073 , n18071 , n18072 );
nor ( n18074 , n18070 , n18073 );
not ( n18075 , n18074 );
nand ( n18076 , n18063 , n18075 );
nand ( n18077 , n18062 , n18074 );
nand ( n18078 , n18076 , n2352 , n18077 );
nand ( n18079 , n18049 , n18078 );
not ( n18080 , n2826 );
and ( n18081 , n9239 , n18080 );
not ( n18082 , n9239 );
buf ( n18083 , n2826 );
and ( n18084 , n18082 , n18083 );
nor ( n18085 , n18081 , n18084 );
not ( n18086 , n2991 );
and ( n18087 , n367 , n18086 );
not ( n18088 , n367 );
and ( n18089 , n18088 , n2987 );
nor ( n18090 , n18087 , n18089 );
and ( n18091 , n18085 , n18090 );
not ( n18092 , n18085 );
not ( n18093 , n18090 );
and ( n18094 , n18092 , n18093 );
nor ( n18095 , n18091 , n18094 );
not ( n18096 , n18095 );
not ( n18097 , n4015 );
or ( n18098 , n9785 , n18097 );
not ( n18099 , n4015 );
nand ( n18100 , n9792 , n18099 );
nand ( n18101 , n18098 , n18100 );
not ( n18102 , n18101 );
nor ( n18103 , n18096 , n18102 );
or ( n18104 , n18095 , n18101 );
nand ( n18105 , n18104 , n2352 );
or ( n18106 , n18103 , n18105 );
xnor ( n18107 , n367 , n368 );
or ( n18108 , n2352 , n18107 );
nand ( n18109 , n18106 , n18108 );
and ( n18110 , n105 , n18083 );
not ( n18111 , n105 );
and ( n18112 , n18111 , n18080 );
nor ( n18113 , n18110 , n18112 );
not ( n18114 , n18113 );
not ( n18115 , n9774 );
not ( n18116 , n9369 );
and ( n18117 , n18115 , n18116 );
not ( n18118 , n9779 );
and ( n18119 , n18118 , n9369 );
nor ( n18120 , n18117 , n18119 );
not ( n18121 , n18120 );
not ( n18122 , n16981 );
not ( n18123 , n2986 );
and ( n18124 , n18122 , n18123 );
not ( n18125 , n2985 );
and ( n18126 , n16982 , n18125 );
nor ( n18127 , n18124 , n18126 );
not ( n18128 , n18127 );
not ( n18129 , n18128 );
or ( n18130 , n18121 , n18129 );
not ( n18131 , n18120 );
nand ( n18132 , n18131 , n18127 );
nand ( n18133 , n18130 , n18132 );
not ( n18134 , n18133 );
nor ( n18135 , n18114 , n18134 );
or ( n18136 , n18113 , n18133 );
nand ( n18137 , n18136 , n2352 );
or ( n18138 , n18135 , n18137 );
not ( n18139 , n105 );
and ( n18140 , n375 , n18139 );
not ( n18141 , n375 );
and ( n18142 , n18141 , n105 );
nor ( n18143 , n18140 , n18142 );
or ( n18144 , n2352 , n18143 );
nand ( n18145 , n18138 , n18144 );
not ( n18146 , n376 );
and ( n18147 , n377 , n18146 );
not ( n18148 , n377 );
and ( n18149 , n18148 , n376 );
nor ( n18150 , n18147 , n18149 );
or ( n18151 , n2352 , n18150 );
and ( n18152 , n18146 , n2991 );
not ( n18153 , n18146 );
and ( n18154 , n18153 , n2986 );
or ( n18155 , n18152 , n18154 );
not ( n18156 , n18155 );
not ( n18157 , n11205 );
not ( n18158 , n18157 );
not ( n18159 , n16520 );
and ( n18160 , n18158 , n18159 );
not ( n18161 , n11148 );
nand ( n18162 , n3013 , n11159 );
nand ( n18163 , n18161 , n11204 , n18162 , n11196 );
not ( n18164 , n18163 );
and ( n18165 , n18164 , n16520 );
nor ( n18166 , n18160 , n18165 );
not ( n18167 , n18166 );
or ( n18168 , n18156 , n18167 );
or ( n18169 , n18155 , n18166 );
nand ( n18170 , n18168 , n18169 );
not ( n18171 , n18170 );
not ( n18172 , n18171 );
not ( n18173 , n8614 );
not ( n18174 , n12679 );
or ( n18175 , n18173 , n18174 );
or ( n18176 , n8614 , n12679 );
nand ( n18177 , n18175 , n18176 );
not ( n18178 , n18177 );
or ( n18179 , n18172 , n18178 );
not ( n18180 , n18177 );
and ( n18181 , n18170 , n18180 );
nor ( n18182 , n18181 , n1 );
nand ( n18183 , n18179 , n18182 );
nand ( n18184 , n18151 , n18183 );
not ( n18185 , n1 );
xor ( n18186 , n388 , n389 );
not ( n18187 , n18186 );
or ( n18188 , n18185 , n18187 );
xor ( n18189 , n388 , n18086 );
not ( n18190 , n18189 );
and ( n18191 , n9369 , n3273 );
not ( n18192 , n9369 );
and ( n18193 , n18192 , n3272 );
nor ( n18194 , n18191 , n18193 );
or ( n18195 , n18194 , n9785 );
nand ( n18196 , n18194 , n9792 );
nand ( n18197 , n18195 , n18196 );
not ( n18198 , n18197 );
or ( n18199 , n18190 , n18198 );
nor ( n18200 , n18189 , n18197 );
nor ( n18201 , n1 , n18200 );
nand ( n18202 , n18199 , n18201 );
nand ( n18203 , n18188 , n18202 );
not ( n18204 , n84 );
not ( n18205 , n18204 );
nand ( n18206 , n14174 , n14190 , n14205 , n14125 );
not ( n18207 , n18206 );
not ( n18208 , n18207 );
or ( n18209 , n18205 , n18208 );
not ( n18210 , n18206 );
or ( n18211 , n18204 , n18210 );
nand ( n18212 , n18209 , n18211 );
not ( n18213 , n18212 );
not ( n18214 , n13834 );
not ( n18215 , n9101 );
or ( n18216 , n18214 , n18215 );
not ( n18217 , n9101 );
nand ( n18218 , n14220 , n18217 );
nand ( n18219 , n18216 , n18218 );
not ( n18220 , n18219 );
or ( n18221 , n18213 , n18220 );
or ( n18222 , n18212 , n18219 );
nand ( n18223 , n18221 , n18222 );
not ( n18224 , n18223 );
not ( n18225 , n13952 );
not ( n18226 , n6150 );
and ( n18227 , n18225 , n18226 );
not ( n18228 , n13952 );
not ( n18229 , n18228 );
not ( n18230 , n6145 );
and ( n18231 , n18229 , n18230 );
nor ( n18232 , n18227 , n18231 );
not ( n18233 , n18232 );
not ( n18234 , n2209 );
not ( n18235 , n1276 );
and ( n18236 , n18234 , n18235 );
not ( n18237 , n5837 );
and ( n18238 , n2209 , n18237 );
nor ( n18239 , n18236 , n18238 );
not ( n18240 , n18239 );
and ( n18241 , n18233 , n18240 );
and ( n18242 , n18239 , n18232 );
nor ( n18243 , n18241 , n18242 );
not ( n18244 , n18243 );
nor ( n18245 , n18224 , n18244 );
or ( n18246 , n18223 , n18243 );
nand ( n18247 , n18246 , n2352 );
or ( n18248 , n18245 , n18247 );
and ( n18249 , n85 , n18204 );
not ( n18250 , n85 );
and ( n18251 , n18250 , n84 );
nor ( n18252 , n18249 , n18251 );
or ( n18253 , n2352 , n18252 );
nand ( n18254 , n18248 , n18253 );
and ( n18255 , n14348 , n77 );
not ( n18256 , n14348 );
not ( n18257 , n77 );
and ( n18258 , n18256 , n18257 );
or ( n18259 , n18255 , n18258 );
not ( n18260 , n2037 );
nand ( n18261 , n2048 , n2058 , n2081 );
or ( n18262 , n18260 , n18261 );
nand ( n18263 , n18262 , n1673 );
nand ( n18264 , n2207 , n18263 , n2151 );
not ( n18265 , n18264 );
not ( n18266 , n18265 );
not ( n18267 , n6472 );
not ( n18268 , n18267 );
and ( n18269 , n18266 , n18268 );
and ( n18270 , n18265 , n18267 );
nor ( n18271 , n18269 , n18270 );
not ( n18272 , n18271 );
xor ( n18273 , n14637 , n18272 );
nor ( n18274 , n18259 , n18273 );
not ( n18275 , n18259 );
not ( n18276 , n18273 );
or ( n18277 , n18275 , n18276 );
nand ( n18278 , n18277 , n2352 );
or ( n18279 , n18274 , n18278 );
and ( n18280 , n88 , n18257 );
not ( n18281 , n88 );
and ( n18282 , n18281 , n77 );
nor ( n18283 , n18280 , n18282 );
or ( n18284 , n2352 , n18283 );
nand ( n18285 , n18279 , n18284 );
xnor ( n18286 , n41 , n42 );
or ( n18287 , n2352 , n18286 );
not ( n18288 , n41 );
not ( n18289 , n1472 );
and ( n18290 , n18288 , n18289 );
and ( n18291 , n41 , n9101 );
nor ( n18292 , n18290 , n18291 );
not ( n18293 , n5839 );
and ( n18294 , n13 , n842 );
nand ( n18295 , n864 , n941 );
nor ( n18296 , n18294 , n18295 );
or ( n18297 , n18293 , n18296 );
not ( n18298 , n803 );
nand ( n18299 , n18298 , n16 );
nand ( n18300 , n833 , n977 );
and ( n18301 , n18299 , n18300 , n14155 );
nand ( n18302 , n18297 , n18301 , n881 );
not ( n18303 , n18302 );
not ( n18304 , n16 );
not ( n18305 , n18304 );
not ( n18306 , n12 );
or ( n18307 , n18306 , n5782 );
and ( n18308 , n929 , n14197 );
nor ( n18309 , n13 , n748 );
nor ( n18310 , n18308 , n18309 );
nand ( n18311 , n18307 , n18310 , n771 );
not ( n18312 , n18311 );
or ( n18313 , n18305 , n18312 );
not ( n18314 , n5803 );
not ( n18315 , n13 );
not ( n18316 , n18315 );
not ( n18317 , n855 );
or ( n18318 , n18316 , n18317 );
nand ( n18319 , n18318 , n970 );
and ( n18320 , n16 , n18319 );
nor ( n18321 , n16 , n13316 );
nor ( n18322 , n18320 , n18321 );
not ( n18323 , n18322 );
or ( n18324 , n18314 , n18323 );
nand ( n18325 , n18324 , n17 );
nand ( n18326 , n18313 , n18325 );
not ( n18327 , n18326 );
not ( n18328 , n14308 );
not ( n18329 , n13287 );
or ( n18330 , n18328 , n18329 );
nand ( n18331 , n18330 , n16 );
and ( n18332 , n13 , n879 );
not ( n18333 , n16 );
not ( n18334 , n14314 );
and ( n18335 , n18333 , n18334 );
nor ( n18336 , n18332 , n18335 );
not ( n18337 , n13 );
nand ( n18338 , n18337 , n14273 );
and ( n18339 , n18338 , n13320 , n14192 );
nand ( n18340 , n13289 , n18336 , n18339 );
nand ( n18341 , n793 , n18340 );
nand ( n18342 , n841 , n18327 , n18331 , n18341 );
not ( n18343 , n17 );
not ( n18344 , n12 );
nor ( n18345 , n18344 , n15 );
or ( n18346 , n18345 , n5791 );
nand ( n18347 , n18346 , n743 );
nand ( n18348 , n13231 , n5966 , n760 );
nand ( n18349 , n16 , n18348 );
nand ( n18350 , n18347 , n14256 , n18349 );
not ( n18351 , n18350 );
or ( n18352 , n18343 , n18351 );
not ( n18353 , n5956 );
or ( n18354 , n13321 , n18353 );
not ( n18355 , n16 );
nand ( n18356 , n18354 , n18355 );
nand ( n18357 , n18352 , n18356 );
not ( n18358 , n18357 );
not ( n18359 , n16 );
nand ( n18360 , n13316 , n844 , n895 );
not ( n18361 , n18360 );
or ( n18362 , n18359 , n18361 );
nand ( n18363 , n755 , n18345 );
not ( n18364 , n18363 );
nand ( n18365 , n18364 , n782 );
not ( n18366 , n14314 );
not ( n18367 , n801 );
or ( n18368 , n18366 , n18367 );
nand ( n18369 , n18368 , n16 );
nand ( n18370 , n18365 , n18369 );
not ( n18371 , n16 );
nand ( n18372 , n18371 , n815 );
nand ( n18373 , n18372 , n5722 , n5789 );
or ( n18374 , n18370 , n18373 );
nand ( n18375 , n18374 , n793 );
nand ( n18376 , n18362 , n18375 );
not ( n18377 , n18376 );
nand ( n18378 , n10 , n18358 , n18377 );
nand ( n18379 , n18342 , n18378 );
and ( n18380 , n17 , n5719 );
not ( n18381 , n17 );
and ( n18382 , n16 , n14111 );
nor ( n18383 , n18382 , n916 , n14291 );
not ( n18384 , n16 );
nand ( n18385 , n5722 , n5702 , n5757 );
nand ( n18386 , n18384 , n18385 );
nand ( n18387 , n18383 , n903 , n18386 );
and ( n18388 , n18381 , n18387 );
nor ( n18389 , n18380 , n18388 );
nand ( n18390 , n18303 , n18379 , n18389 );
not ( n18391 , n18390 );
not ( n18392 , n18391 );
not ( n18393 , n18392 );
not ( n18394 , n18393 );
and ( n18395 , n18292 , n18394 );
not ( n18396 , n18292 );
and ( n18397 , n18396 , n18393 );
nor ( n18398 , n18395 , n18397 );
not ( n18399 , n18398 );
and ( n18400 , n25 , n13938 );
nor ( n18401 , n18400 , n6175 , n1919 );
not ( n18402 , n25 );
nand ( n18403 , n1766 , n6215 , n6277 );
nand ( n18404 , n18402 , n18403 );
and ( n18405 , n18401 , n1850 , n18404 );
nor ( n18406 , n18405 , n26 );
not ( n18407 , n1987 );
nand ( n18408 , n23 , n1829 );
and ( n18409 , n18408 , n1786 , n13418 );
or ( n18410 , n18407 , n18409 );
nand ( n18411 , n25 , n1982 );
nand ( n18412 , n1794 , n1785 );
and ( n18413 , n18411 , n18412 , n13873 );
not ( n18414 , n1770 );
nand ( n18415 , n18410 , n18413 , n18414 );
nor ( n18416 , n18406 , n18415 );
not ( n18417 , n6193 );
nand ( n18418 , n26 , n18417 );
not ( n18419 , n14408 );
not ( n18420 , n6406 );
or ( n18421 , n18419 , n18420 );
nand ( n18422 , n18421 , n25 );
not ( n18423 , n25 );
not ( n18424 , n18423 );
not ( n18425 , n6363 );
or ( n18426 , n18424 , n18425 );
not ( n18427 , n6178 );
nand ( n18428 , n18426 , n18427 );
or ( n18429 , n23 , n1803 );
nand ( n18430 , n18429 , n1900 );
and ( n18431 , n25 , n18430 );
or ( n18432 , n18428 , n18431 );
nand ( n18433 , n18432 , n26 );
not ( n18434 , n25 );
and ( n18435 , n1960 , n13870 );
not ( n18436 , n23 );
not ( n18437 , n1860 );
and ( n18438 , n18436 , n18437 );
nor ( n18439 , n18435 , n18438 );
nand ( n18440 , n22 , n13364 );
nand ( n18441 , n18439 , n1894 , n18440 );
nand ( n18442 , n18434 , n18441 );
not ( n18443 , n13866 );
nand ( n18444 , n18443 , n13398 , n6406 , n6427 );
not ( n18445 , n6267 );
or ( n18446 , n23 , n18445 );
nand ( n18447 , n21 , n1940 );
or ( n18448 , n25 , n18447 );
nand ( n18449 , n18446 , n18448 );
or ( n18450 , n18444 , n18449 );
not ( n18451 , n26 );
nand ( n18452 , n18450 , n18451 );
nand ( n18453 , n18422 , n18433 , n18442 , n18452 );
and ( n18454 , n1853 , n18453 );
not ( n18455 , n1853 );
not ( n18456 , n1987 );
nand ( n18457 , n13469 , n1843 , n1861 );
not ( n18458 , n18457 );
or ( n18459 , n18456 , n18458 );
nand ( n18460 , n26 , n14373 );
nand ( n18461 , n18459 , n18460 );
not ( n18462 , n18447 );
or ( n18463 , n18462 , n1933 );
nand ( n18464 , n18463 , n6462 );
not ( n18465 , n6320 );
not ( n18466 , n13398 );
or ( n18467 , n18465 , n18466 );
not ( n18468 , n25 );
nand ( n18469 , n18467 , n18468 );
nand ( n18470 , n18464 , n18469 );
nor ( n18471 , n18461 , n18470 );
not ( n18472 , n1859 );
nand ( n18473 , n22 , n1783 );
nand ( n18474 , n18472 , n18473 );
nand ( n18475 , n26 , n1855 , n18474 );
not ( n18476 , n13402 );
not ( n18477 , n1846 );
or ( n18478 , n18476 , n18477 );
nand ( n18479 , n18478 , n25 );
nand ( n18480 , n18475 , n18479 );
not ( n18481 , n26 );
not ( n18482 , n18481 );
not ( n18483 , n1864 );
not ( n18484 , n25 );
nand ( n18485 , n18484 , n1876 );
nand ( n18486 , n22 , n1802 );
not ( n18487 , n18486 );
nand ( n18488 , n18487 , n1768 );
nand ( n18489 , n18483 , n18485 , n6165 , n18488 );
not ( n18490 , n18489 );
or ( n18491 , n18482 , n18490 );
nand ( n18492 , n18491 , n14451 );
nor ( n18493 , n18480 , n18492 );
nand ( n18494 , n18471 , n18493 );
and ( n18495 , n18455 , n18494 );
nor ( n18496 , n18454 , n18495 );
nand ( n18497 , n18416 , n18418 , n18496 );
not ( n18498 , n18497 );
not ( n18499 , n18498 );
not ( n18500 , n18499 );
not ( n18501 , n18500 );
not ( n18502 , n18272 );
and ( n18503 , n18501 , n18502 );
and ( n18504 , n18500 , n18272 );
nor ( n18505 , n18503 , n18504 );
not ( n18506 , n18505 );
nand ( n18507 , n18399 , n18506 );
nand ( n18508 , n18398 , n18505 );
nand ( n18509 , n18507 , n2352 , n18508 );
nand ( n18510 , n18287 , n18509 );
not ( n18511 , n81 );
and ( n18512 , n18511 , n14206 );
not ( n18513 , n18511 );
and ( n18514 , n18513 , n14207 );
nor ( n18515 , n18512 , n18514 );
and ( n18516 , n987 , n13730 );
not ( n18517 , n987 );
and ( n18518 , n18517 , n5989 );
nor ( n18519 , n18516 , n18518 );
xor ( n18520 , n18515 , n18519 );
not ( n18521 , n18520 );
not ( n18522 , n14066 );
or ( n18523 , n18522 , n1477 );
not ( n18524 , n14076 );
nand ( n18525 , n18524 , n1477 );
nand ( n18526 , n18523 , n18525 );
not ( n18527 , n18526 );
nor ( n18528 , n18521 , n18527 );
or ( n18529 , n18520 , n18526 );
nand ( n18530 , n18529 , n2352 );
or ( n18531 , n18528 , n18530 );
and ( n18532 , n82 , n18511 );
not ( n18533 , n82 );
and ( n18534 , n18533 , n81 );
nor ( n18535 , n18532 , n18534 );
or ( n18536 , n2352 , n18535 );
nand ( n18537 , n18531 , n18536 );
not ( n18538 , n215 );
and ( n18539 , n216 , n18538 );
not ( n18540 , n216 );
and ( n18541 , n18540 , n215 );
nor ( n18542 , n18539 , n18541 );
or ( n18543 , n2352 , n18542 );
not ( n18544 , n118 );
not ( n18545 , n11810 );
nand ( n18546 , n18545 , n11685 );
not ( n18547 , n15589 );
nand ( n18548 , n7512 , n17383 );
not ( n18549 , n18548 );
or ( n18550 , n18547 , n18549 );
nand ( n18551 , n18550 , n117 );
nand ( n18552 , n15586 , n18546 , n18551 );
and ( n18553 , n18544 , n18552 );
not ( n18554 , n117 );
nand ( n18555 , n18554 , n17344 );
nand ( n18556 , n116 , n11902 );
and ( n18557 , n18555 , n18556 );
not ( n18558 , n118 );
nor ( n18559 , n18557 , n18558 );
nor ( n18560 , n18553 , n18559 );
not ( n18561 , n118 );
nor ( n18562 , n15706 , n15609 );
nand ( n18563 , n18562 , n17640 , n7561 );
not ( n18564 , n18563 );
or ( n18565 , n18561 , n18564 );
not ( n18566 , n11743 );
not ( n18567 , n18566 );
not ( n18568 , n15658 );
or ( n18569 , n18567 , n18568 );
not ( n18570 , n117 );
nand ( n18571 , n18569 , n18570 );
nand ( n18572 , n18565 , n18571 );
not ( n18573 , n118 );
not ( n18574 , n18573 );
not ( n18575 , n7608 );
nand ( n18576 , n7401 , n7538 );
and ( n18577 , n117 , n18576 );
not ( n18578 , n117 );
and ( n18579 , n18578 , n7503 );
nor ( n18580 , n18577 , n18579 );
nand ( n18581 , n18575 , n11843 , n18580 , n15589 );
not ( n18582 , n18581 );
or ( n18583 , n18574 , n18582 );
nand ( n18584 , n112 , n7498 );
not ( n18585 , n11667 );
nand ( n18586 , n115 , n18585 );
nand ( n18587 , n18584 , n18586 , n15650 );
not ( n18588 , n117 );
nand ( n18589 , n18587 , n118 , n18588 );
nand ( n18590 , n11740 , n18589 );
not ( n18591 , n117 );
not ( n18592 , n15589 );
not ( n18593 , n18592 );
or ( n18594 , n18591 , n18593 );
and ( n18595 , n17418 , n17427 );
nand ( n18596 , n18594 , n18595 );
nor ( n18597 , n18590 , n18596 );
nand ( n18598 , n18583 , n18597 );
or ( n18599 , n18572 , n18598 );
nand ( n18600 , n18599 , n119 );
not ( n18601 , n117 );
nand ( n18602 , n18601 , n15687 );
nand ( n18603 , n18602 , n15616 , n11689 );
not ( n18604 , n17369 );
not ( n18605 , n116 );
nand ( n18606 , n18605 , n7533 );
nand ( n18607 , n18606 , n11624 , n7581 );
not ( n18608 , n18607 );
or ( n18609 , n18604 , n18608 );
not ( n18610 , n116 );
nand ( n18611 , n11618 , n18610 , n17349 );
nand ( n18612 , n18609 , n18611 );
nor ( n18613 , n18603 , n18612 );
nor ( n18614 , n7484 , n18586 );
not ( n18615 , n18614 );
nand ( n18616 , n18615 , n18555 );
nor ( n18617 , n117 , n11642 );
not ( n18618 , n18617 );
nand ( n18619 , n15598 , n18618 );
and ( n18620 , n116 , n11668 );
nor ( n18621 , n18620 , n7418 );
nand ( n18622 , n116 , n15644 );
not ( n18623 , n18622 );
nor ( n18624 , n18623 , n17579 );
and ( n18625 , n18621 , n18624 );
not ( n18626 , n117 );
nor ( n18627 , n18625 , n18626 );
nor ( n18628 , n18616 , n18619 , n18627 );
not ( n18629 , n18628 );
not ( n18630 , n118 );
not ( n18631 , n7592 );
and ( n18632 , n18622 , n18631 , n11784 , n11788 );
not ( n18633 , n117 );
not ( n18634 , n116 );
nand ( n18635 , n18634 , n7518 );
nand ( n18636 , n18635 , n15669 , n11826 );
nand ( n18637 , n18633 , n18636 );
not ( n18638 , n7535 );
not ( n18639 , n7579 );
or ( n18640 , n18638 , n18639 );
nand ( n18641 , n18640 , n117 );
nand ( n18642 , n18632 , n18637 , n15675 , n18641 );
or ( n18643 , n18630 , n18642 );
not ( n18644 , n118 );
not ( n18645 , n7407 );
nor ( n18646 , n18645 , n7387 );
nor ( n18647 , n18646 , n7458 );
not ( n18648 , n15650 );
nand ( n18649 , n18648 , n11685 );
not ( n18650 , n116 );
nand ( n18651 , n18650 , n17643 );
nand ( n18652 , n18644 , n18647 , n18649 , n18651 );
nand ( n18653 , n18643 , n18652 );
not ( n18654 , n18653 );
or ( n18655 , n18629 , n18654 );
nand ( n18656 , n18655 , n7325 );
and ( n18657 , n18560 , n18600 , n18613 , n18656 );
not ( n18658 , n18657 );
not ( n18659 , n127 );
and ( n18660 , n8209 , n15496 );
nor ( n18661 , n18660 , n120 );
not ( n18662 , n18661 );
nand ( n18663 , n7868 , n15544 );
not ( n18664 , n120 );
nand ( n18665 , n18664 , n7629 );
not ( n18666 , n8066 );
not ( n18667 , n7798 );
not ( n18668 , n18667 );
not ( n18669 , n7684 );
or ( n18670 , n18668 , n18669 );
nand ( n18671 , n18670 , n120 );
nand ( n18672 , n18665 , n18666 , n18671 );
or ( n18673 , n18663 , n18672 );
nand ( n18674 , n18673 , n126 );
nor ( n18675 , n120 , n15407 );
not ( n18676 , n15345 );
not ( n18677 , n125 );
nand ( n18678 , n18677 , n8135 );
and ( n18679 , n18676 , n8060 , n18678 );
nor ( n18680 , n18679 , n7819 );
nor ( n18681 , n18675 , n18680 );
not ( n18682 , n18681 );
not ( n18683 , n120 );
not ( n18684 , n7850 );
or ( n18685 , n18683 , n18684 );
nor ( n18686 , n8176 , n8239 );
nand ( n18687 , n18685 , n18686 );
nor ( n18688 , n18682 , n18687 );
nand ( n18689 , n15401 , n8160 );
nand ( n18690 , n15346 , n7671 );
or ( n18691 , n18689 , n18690 );
not ( n18692 , n126 );
nand ( n18693 , n18691 , n18692 );
nand ( n18694 , n18662 , n18674 , n18688 , n18693 );
not ( n18695 , n18694 );
or ( n18696 , n18659 , n18695 );
not ( n18697 , n120 );
and ( n18698 , n18697 , n15529 );
not ( n18699 , n8143 );
or ( n18700 , n126 , n18699 );
nand ( n18701 , n18700 , n15347 );
nor ( n18702 , n18698 , n18701 );
not ( n18703 , n120 );
nand ( n18704 , n18703 , n7722 );
not ( n18705 , n126 );
not ( n18706 , n121 );
not ( n18707 , n15552 );
not ( n18708 , n18707 );
or ( n18709 , n18706 , n18708 );
nand ( n18710 , n7751 , n15555 );
nand ( n18711 , n18709 , n18710 );
nand ( n18712 , n18705 , n18711 );
and ( n18713 , n18702 , n18704 , n18712 );
nand ( n18714 , n18696 , n18713 );
not ( n18715 , n18714 );
not ( n18716 , n120 );
not ( n18717 , n18716 );
nand ( n18718 , n7921 , n15407 , n7861 );
not ( n18719 , n18718 );
or ( n18720 , n18717 , n18719 );
nand ( n18721 , n18720 , n8200 );
not ( n18722 , n18721 );
not ( n18723 , n8148 );
or ( n18724 , n18723 , n7974 );
not ( n18725 , n15544 );
nand ( n18726 , n7635 , n8166 );
not ( n18727 , n18726 );
or ( n18728 , n18725 , n18727 );
nand ( n18729 , n18728 , n120 );
nand ( n18730 , n18722 , n18724 , n18729 );
nand ( n18731 , n126 , n18730 );
not ( n18732 , n126 );
or ( n18733 , n8004 , n8060 );
nand ( n18734 , n7751 , n8181 );
nand ( n18735 , n18733 , n18734 );
not ( n18736 , n18735 );
or ( n18737 , n18732 , n18736 );
not ( n18738 , n15352 );
not ( n18739 , n15544 );
or ( n18740 , n18738 , n18739 );
nand ( n18741 , n18740 , n126 );
nand ( n18742 , n18737 , n18741 );
not ( n18743 , n18742 );
not ( n18744 , n120 );
nand ( n18745 , n18744 , n8101 );
not ( n18746 , n7811 );
not ( n18747 , n15424 );
or ( n18748 , n18746 , n18747 );
nand ( n18749 , n18748 , n120 );
and ( n18750 , n18745 , n18749 );
not ( n18751 , n8017 );
nand ( n18752 , n121 , n8137 );
not ( n18753 , n18752 );
or ( n18754 , n18751 , n18753 );
nand ( n18755 , n18754 , n120 );
nor ( n18756 , n7971 , n18678 );
not ( n18757 , n18756 );
and ( n18758 , n18755 , n15552 , n18757 );
and ( n18759 , n18699 , n18750 , n18758 );
not ( n18760 , n126 );
nor ( n18761 , n7953 , n7895 );
not ( n18762 , n120 );
or ( n18763 , n121 , n7653 );
nand ( n18764 , n18763 , n8170 , n8085 );
nand ( n18765 , n18762 , n18764 );
nand ( n18766 , n18761 , n18765 , n8017 , n7941 );
not ( n18767 , n18766 );
or ( n18768 , n7696 , n15555 );
nand ( n18769 , n18768 , n120 );
nand ( n18770 , n18767 , n18769 , n8106 );
nand ( n18771 , n18760 , n18770 );
nand ( n18772 , n18743 , n18759 , n18771 );
nand ( n18773 , n7748 , n18772 );
nand ( n18774 , n18715 , n18731 , n18773 );
not ( n18775 , n18774 );
or ( n18776 , n18658 , n18775 );
not ( n18777 , n18657 );
not ( n18778 , n7748 );
not ( n18779 , n18772 );
or ( n18780 , n18778 , n18779 );
nand ( n18781 , n18780 , n18731 );
nor ( n18782 , n18714 , n18781 );
nand ( n18783 , n18777 , n18782 );
nand ( n18784 , n18776 , n18783 );
not ( n18785 , n18784 );
not ( n18786 , n18785 );
not ( n18787 , n118 );
nand ( n18788 , n117 , n7420 );
and ( n18789 , n18788 , n17414 , n11592 );
not ( n18790 , n117 );
nand ( n18791 , n11716 , n7375 , n11675 );
nand ( n18792 , n18790 , n18791 );
nand ( n18793 , n18789 , n17334 , n18792 );
and ( n18794 , n18787 , n18793 );
not ( n18795 , n117 );
or ( n18796 , n18795 , n15632 );
not ( n18797 , n18646 );
and ( n18798 , n18796 , n18797 , n17345 );
nand ( n18799 , n116 , n15676 );
not ( n18800 , n18799 );
nor ( n18801 , n7409 , n11735 );
not ( n18802 , n18801 );
or ( n18803 , n18800 , n18802 );
nand ( n18804 , n18803 , n11618 );
nand ( n18805 , n18798 , n7461 , n18804 );
nor ( n18806 , n18794 , n18805 );
not ( n18807 , n118 );
nor ( n18808 , n18807 , n11689 );
not ( n18809 , n18808 );
nand ( n18810 , n11897 , n15707 );
not ( n18811 , n117 );
nand ( n18812 , n15675 , n7362 , n15637 );
not ( n18813 , n18812 );
or ( n18814 , n18811 , n18813 );
not ( n18815 , n11600 );
not ( n18816 , n112 );
nand ( n18817 , n18816 , n115 );
nand ( n18818 , n18815 , n18817 );
nand ( n18819 , n11597 , n18818 );
nand ( n18820 , n18814 , n18819 );
or ( n18821 , n18810 , n18820 );
nand ( n18822 , n18821 , n118 );
not ( n18823 , n11697 );
not ( n18824 , n11826 );
or ( n18825 , n18823 , n18824 );
not ( n18826 , n117 );
nand ( n18827 , n18825 , n18826 );
nand ( n18828 , n15598 , n7504 , n7364 , n15589 );
nand ( n18829 , n117 , n18828 );
not ( n18830 , n11714 );
not ( n18831 , n113 );
nand ( n18832 , n18831 , n7537 );
not ( n18833 , n18832 );
or ( n18834 , n18830 , n18833 );
nand ( n18835 , n18834 , n117 );
nand ( n18836 , n7375 , n11598 , n18835 );
or ( n18837 , n18836 , n18614 , n18617 );
not ( n18838 , n118 );
nand ( n18839 , n18837 , n18838 );
nand ( n18840 , n18822 , n18827 , n18829 , n18839 );
and ( n18841 , n119 , n18840 );
not ( n18842 , n119 );
or ( n18843 , n116 , n17638 );
or ( n18844 , n117 , n18832 );
nand ( n18845 , n18843 , n18844 );
not ( n18846 , n7336 );
nor ( n18847 , n11765 , n7479 );
nand ( n18848 , n18846 , n18847 , n11697 );
or ( n18849 , n18845 , n18848 );
not ( n18850 , n118 );
nand ( n18851 , n18849 , n18850 );
not ( n18852 , n117 );
and ( n18853 , n7498 , n7452 );
not ( n18854 , n116 );
and ( n18855 , n18854 , n11602 );
nor ( n18856 , n18853 , n18855 );
nand ( n18857 , n115 , n7426 );
nand ( n18858 , n18856 , n7523 , n18857 );
nand ( n18859 , n18852 , n18858 );
not ( n18860 , n118 );
not ( n18861 , n116 );
not ( n18862 , n18861 );
not ( n18863 , n11668 );
or ( n18864 , n18862 , n18863 );
nand ( n18865 , n18864 , n11610 );
nand ( n18866 , n117 , n18865 );
not ( n18867 , n117 );
nand ( n18868 , n18867 , n11902 );
nand ( n18869 , n18866 , n7581 , n18868 );
not ( n18870 , n18869 );
or ( n18871 , n18860 , n18870 );
not ( n18872 , n17590 );
not ( n18873 , n7337 );
or ( n18874 , n18872 , n18873 );
nand ( n18875 , n18874 , n117 );
nand ( n18876 , n18871 , n18875 );
not ( n18877 , n18876 );
nand ( n18878 , n18851 , n18859 , n18877 );
and ( n18879 , n18842 , n18878 );
nor ( n18880 , n18841 , n18879 );
nand ( n18881 , n18806 , n18809 , n18880 );
not ( n18882 , n18881 );
not ( n18883 , n11960 );
and ( n18884 , n144 , n18883 );
not ( n18885 , n144 );
not ( n18886 , n6766 );
nand ( n18887 , n18886 , n141 );
and ( n18888 , n18887 , n11288 , n11330 );
not ( n18889 , n141 );
not ( n18890 , n11956 );
nand ( n18891 , n11258 , n18890 , n11453 );
nand ( n18892 , n18889 , n18891 );
nand ( n18893 , n18888 , n11387 , n18892 );
and ( n18894 , n18885 , n18893 );
nor ( n18895 , n18884 , n18894 );
and ( n18896 , n141 , n11259 );
not ( n18897 , n6795 );
nor ( n18898 , n18897 , n11559 );
nor ( n18899 , n18896 , n18898 , n17541 );
not ( n18900 , n11373 );
not ( n18901 , n142 );
nor ( n18902 , n18901 , n11251 );
or ( n18903 , n18902 , n6778 , n15096 );
nand ( n18904 , n18903 , n11498 );
nand ( n18905 , n18899 , n18900 , n18904 );
not ( n18906 , n18905 );
not ( n18907 , n144 );
not ( n18908 , n141 );
not ( n18909 , n11447 );
nand ( n18910 , n18908 , n18909 );
not ( n18911 , n142 );
not ( n18912 , n18911 );
not ( n18913 , n11362 );
or ( n18914 , n18912 , n18913 );
nand ( n18915 , n18914 , n11318 );
nand ( n18916 , n141 , n18915 );
nand ( n18917 , n6674 , n18910 , n18916 );
not ( n18918 , n18917 );
or ( n18919 , n18907 , n18918 );
not ( n18920 , n141 );
and ( n18921 , n11328 , n6738 );
nor ( n18922 , n142 , n11248 );
nor ( n18923 , n18921 , n18922 );
nand ( n18924 , n140 , n6756 );
nand ( n18925 , n18923 , n6645 , n18924 );
nand ( n18926 , n18920 , n18925 );
nand ( n18927 , n18919 , n18926 );
not ( n18928 , n18927 );
not ( n18929 , n17504 );
not ( n18930 , n6751 );
or ( n18931 , n18929 , n18930 );
nand ( n18932 , n18931 , n141 );
not ( n18933 , n15139 );
nand ( n18934 , n18933 , n6751 );
not ( n18935 , n142 );
and ( n18936 , n18935 , n6613 );
not ( n18937 , n141 );
and ( n18938 , n143 , n140 , n142 );
and ( n18939 , n18937 , n18938 );
nor ( n18940 , n18936 , n18939 );
nand ( n18941 , n142 , n11566 );
nand ( n18942 , n18940 , n18941 , n6725 );
or ( n18943 , n18934 , n18942 );
not ( n18944 , n144 );
nand ( n18945 , n18943 , n18944 );
nand ( n18946 , n6808 , n18928 , n18932 , n18945 );
not ( n18947 , n141 );
not ( n18948 , n15139 );
nand ( n18949 , n18948 , n11526 );
and ( n18950 , n18947 , n18949 );
not ( n18951 , n18947 );
not ( n18952 , n18909 );
not ( n18953 , n11370 );
nand ( n18954 , n6592 , n18952 , n18953 );
and ( n18955 , n18951 , n18954 );
nor ( n18956 , n18950 , n18955 );
not ( n18957 , n144 );
not ( n18958 , n18938 );
nand ( n18959 , n18958 , n11281 );
and ( n18960 , n141 , n18959 );
nand ( n18961 , n140 , n11360 );
nor ( n18962 , n6543 , n18961 );
nor ( n18963 , n18960 , n18962 );
not ( n18964 , n141 );
nand ( n18965 , n18964 , n11265 );
nand ( n18966 , n18963 , n18965 , n11957 , n11928 );
nand ( n18967 , n18957 , n18966 );
nand ( n18968 , n11440 , n15072 );
not ( n18969 , n141 );
not ( n18970 , n15108 );
nand ( n18971 , n18970 , n6716 , n11251 );
not ( n18972 , n18971 );
or ( n18973 , n18969 , n18972 );
not ( n18974 , n140 );
or ( n18975 , n18974 , n138 );
nand ( n18976 , n18975 , n11930 );
nand ( n18977 , n11246 , n18976 );
nand ( n18978 , n18973 , n18977 );
or ( n18979 , n18968 , n18978 );
nand ( n18980 , n18979 , n144 );
nand ( n18981 , n137 , n18956 , n18967 , n18980 );
nand ( n18982 , n18946 , n18981 );
nand ( n18983 , n18895 , n18906 , n18982 );
not ( n18984 , n18983 );
or ( n18985 , n18882 , n18984 );
not ( n18986 , n18881 );
not ( n18987 , n18983 );
nand ( n18988 , n18986 , n18987 );
nand ( n18989 , n18985 , n18988 );
and ( n18990 , n133 , n17928 );
not ( n18991 , n7014 );
nor ( n18992 , n18990 , n17215 , n18991 );
not ( n18993 , n133 );
nand ( n18994 , n7151 , n17229 , n6913 );
nand ( n18995 , n18993 , n18994 );
and ( n18996 , n18992 , n7048 , n18995 );
nor ( n18997 , n18996 , n134 );
not ( n18998 , n133 );
not ( n18999 , n18998 );
not ( n19000 , n6914 );
and ( n19001 , n18999 , n19000 );
nand ( n19002 , n6827 , n15218 );
nand ( n19003 , n19002 , n15219 );
nor ( n19004 , n19001 , n19003 );
not ( n19005 , n132 );
not ( n19006 , n7064 );
or ( n19007 , n19005 , n19006 );
nand ( n19008 , n19007 , n7052 , n17738 );
nand ( n19009 , n7195 , n19008 );
nand ( n19010 , n19004 , n7053 , n19009 );
nor ( n19011 , n18997 , n19010 );
not ( n19012 , n17245 );
nand ( n19013 , n134 , n19012 );
or ( n19014 , n6822 , n129 );
nand ( n19015 , n19014 , n15183 );
nand ( n19016 , n6864 , n19015 );
not ( n19017 , n17750 );
and ( n19018 , n7034 , n6859 );
not ( n19019 , n19018 );
or ( n19020 , n19017 , n19019 );
nand ( n19021 , n19020 , n133 );
nand ( n19022 , n7139 , n15292 , n19016 , n19021 );
and ( n19023 , n134 , n19022 );
nand ( n19024 , n131 , n7027 );
not ( n19025 , n19024 );
nand ( n19026 , n19025 , n7002 );
and ( n19027 , n15196 , n19026 );
not ( n19028 , n133 );
nand ( n19029 , n19028 , n6817 , n6899 );
not ( n19030 , n130 );
nor ( n19031 , n19030 , n6839 );
not ( n19032 , n19031 );
not ( n19033 , n19032 );
not ( n19034 , n6830 );
or ( n19035 , n19033 , n19034 );
nand ( n19036 , n19035 , n133 );
and ( n19037 , n19029 , n17207 , n19036 );
and ( n19038 , n19027 , n19037 );
nor ( n19039 , n19038 , n134 );
nor ( n19040 , n19023 , n19039 );
not ( n19041 , n6982 );
not ( n19042 , n7223 );
or ( n19043 , n19041 , n19042 );
not ( n19044 , n133 );
nand ( n19045 , n19043 , n19044 );
not ( n19046 , n7042 );
not ( n19047 , n7134 );
not ( n19048 , n19047 );
nand ( n19049 , n19046 , n19048 , n7066 );
nand ( n19050 , n133 , n19049 );
nand ( n19051 , n19040 , n19045 , n19050 );
and ( n19052 , n135 , n19051 );
not ( n19053 , n135 );
not ( n19054 , n15186 );
not ( n19055 , n17781 );
or ( n19056 , n19054 , n19055 );
nand ( n19057 , n19056 , n133 );
not ( n19058 , n133 );
not ( n19059 , n19058 );
not ( n19060 , n19047 );
or ( n19061 , n19059 , n19060 );
or ( n19062 , n132 , n7028 );
nand ( n19063 , n19062 , n6953 );
nand ( n19064 , n133 , n19063 );
nand ( n19065 , n19061 , n19064 );
or ( n19066 , n17216 , n19065 );
nand ( n19067 , n19066 , n134 );
not ( n19068 , n133 );
or ( n19069 , n6822 , n15283 );
and ( n19070 , n6873 , n17964 );
not ( n19071 , n132 );
and ( n19072 , n19071 , n6852 );
nor ( n19073 , n19070 , n19072 );
nand ( n19074 , n19069 , n19073 , n6882 );
nand ( n19075 , n19068 , n19074 );
not ( n19076 , n134 );
not ( n19077 , n132 );
and ( n19078 , n19077 , n15264 );
not ( n19079 , n133 );
and ( n19080 , n19079 , n19031 );
nor ( n19081 , n19078 , n19080 );
nand ( n19082 , n132 , n6938 );
and ( n19083 , n19081 , n6982 , n19082 );
nand ( n19084 , n19083 , n17781 , n17969 );
nand ( n19085 , n19076 , n19084 );
nand ( n19086 , n19057 , n19067 , n19075 , n19085 );
and ( n19087 , n19053 , n19086 );
nor ( n19088 , n19052 , n19087 );
nand ( n19089 , n19011 , n19013 , n19088 );
not ( n19090 , n19089 );
and ( n19091 , n19090 , n18538 );
not ( n19092 , n19090 );
and ( n19093 , n19092 , n215 );
nor ( n19094 , n19091 , n19093 );
and ( n19095 , n18989 , n19094 );
not ( n19096 , n18989 );
not ( n19097 , n19094 );
and ( n19098 , n19096 , n19097 );
nor ( n19099 , n19095 , n19098 );
not ( n19100 , n19099 );
nand ( n19101 , n18786 , n19100 );
nand ( n19102 , n18785 , n19099 );
nand ( n19103 , n19101 , n2352 , n19102 );
nand ( n19104 , n18543 , n19103 );
xnor ( n19105 , n217 , n218 );
or ( n19106 , n2352 , n19105 );
not ( n19107 , n218 );
not ( n19108 , n160 );
or ( n19109 , n159 , n10121 );
or ( n19110 , n158 , n9822 );
nand ( n19111 , n19110 , n9884 );
nand ( n19112 , n159 , n19111 );
nand ( n19113 , n19109 , n4259 , n19112 );
not ( n19114 , n19113 );
or ( n19115 , n19108 , n19114 );
not ( n19116 , n16062 );
not ( n19117 , n14766 );
not ( n19118 , n19117 );
or ( n19119 , n19116 , n19118 );
nand ( n19120 , n19119 , n159 );
nand ( n19121 , n19115 , n19120 );
not ( n19122 , n4054 );
and ( n19123 , n9899 , n10063 );
not ( n19124 , n158 );
and ( n19125 , n19124 , n4091 );
not ( n19126 , n159 );
nand ( n19127 , n157 , n4064 );
not ( n19128 , n19127 );
and ( n19129 , n19126 , n19128 );
nor ( n19130 , n19125 , n19129 );
nand ( n19131 , n14767 , n4237 , n19123 , n19130 );
not ( n19132 , n19131 );
or ( n19133 , n19122 , n19132 );
not ( n19134 , n159 );
not ( n19135 , n154 );
or ( n19136 , n19135 , n14803 );
not ( n19137 , n4128 );
not ( n19138 , n4245 );
and ( n19139 , n19137 , n19138 );
not ( n19140 , n158 );
and ( n19141 , n19140 , n10889 );
nor ( n19142 , n19139 , n19141 );
nand ( n19143 , n19136 , n19142 , n4041 );
nand ( n19144 , n19134 , n19143 );
nand ( n19145 , n19133 , n19144 );
nor ( n19146 , n19121 , n19145 );
nor ( n19147 , n161 , n19146 );
not ( n19148 , n19147 );
and ( n19149 , n159 , n4164 );
not ( n19150 , n9919 );
nor ( n19151 , n19149 , n9936 , n19150 );
not ( n19152 , n159 );
nand ( n19153 , n4079 , n10879 , n9811 );
nand ( n19154 , n19152 , n19153 );
nand ( n19155 , n19151 , n9827 , n19154 );
nand ( n19156 , n4054 , n19155 );
nand ( n19157 , n159 , n9814 );
not ( n19158 , n12784 );
and ( n19159 , n19157 , n19158 , n4050 );
not ( n19160 , n158 );
or ( n19161 , n19160 , n9839 );
nand ( n19162 , n19161 , n4085 , n12739 );
and ( n19163 , n10024 , n19162 );
not ( n19164 , n9867 );
nor ( n19165 , n19163 , n19164 );
and ( n19166 , n19156 , n19159 , n19165 );
nand ( n19167 , n160 , n10867 );
not ( n19168 , n159 );
nand ( n19169 , n9899 , n10020 );
and ( n19170 , n19168 , n19169 );
not ( n19171 , n19168 );
not ( n19172 , n9834 );
nand ( n19173 , n10121 , n4138 , n19172 );
and ( n19174 , n19171 , n19173 );
nor ( n19175 , n19170 , n19174 );
not ( n19176 , n19175 );
nor ( n19177 , n4080 , n12772 );
not ( n19178 , n19127 );
not ( n19179 , n9908 );
not ( n19180 , n19179 );
or ( n19181 , n19178 , n19180 );
nand ( n19182 , n19181 , n159 );
nand ( n19183 , n10891 , n19182 );
nor ( n19184 , n12769 , n19183 );
nand ( n19185 , n19177 , n19184 );
and ( n19186 , n4054 , n19185 );
not ( n19187 , n4054 );
and ( n19188 , n10129 , n12704 );
not ( n19189 , n154 );
nor ( n19190 , n19189 , n156 );
or ( n19191 , n19190 , n9956 );
nand ( n19192 , n19191 , n4148 );
not ( n19193 , n4207 );
nand ( n19194 , n14818 , n19193 , n9839 );
nand ( n19195 , n159 , n19194 );
nand ( n19196 , n19188 , n19192 , n19195 );
and ( n19197 , n19187 , n19196 );
nor ( n19198 , n19186 , n19197 );
not ( n19199 , n19198 );
or ( n19200 , n19176 , n19199 );
nand ( n19201 , n19200 , n161 );
nand ( n19202 , n19148 , n19166 , n19167 , n19201 );
not ( n19203 , n19202 );
or ( n19204 , n19107 , n19203 );
not ( n19205 , n218 );
not ( n19206 , n19167 );
not ( n19207 , n19206 );
nand ( n19208 , n19175 , n19198 );
and ( n19209 , n161 , n19208 );
nor ( n19210 , n19209 , n19147 );
nand ( n19211 , n19207 , n19166 , n19210 );
not ( n19212 , n19211 );
nand ( n19213 , n19205 , n19212 );
nand ( n19214 , n19204 , n19213 );
buf ( n19215 , n12823 );
and ( n19216 , n19214 , n19215 );
not ( n19217 , n19214 );
and ( n19218 , n19217 , n18026 );
nor ( n19219 , n19216 , n19218 );
not ( n19220 , n19219 );
not ( n19221 , n17020 );
nand ( n19222 , n172 , n15891 );
and ( n19223 , n19222 , n4718 , n5098 );
nor ( n19224 , n19223 , n4878 );
not ( n19225 , n19224 );
not ( n19226 , n12080 );
nand ( n19227 , n177 , n19226 );
not ( n19228 , n177 );
not ( n19229 , n5017 );
not ( n19230 , n172 );
nand ( n19231 , n19230 , n5129 );
not ( n19232 , n19231 );
or ( n19233 , n19229 , n19232 );
nand ( n19234 , n19233 , n176 );
not ( n19235 , n176 );
nand ( n19236 , n19235 , n12901 );
nand ( n19237 , n19234 , n4579 , n19236 );
not ( n19238 , n19237 );
or ( n19239 , n19228 , n19238 );
not ( n19240 , n172 );
not ( n19241 , n12860 );
nand ( n19242 , n19240 , n19241 );
not ( n19243 , n19242 );
not ( n19244 , n4959 );
or ( n19245 , n19243 , n19244 );
nand ( n19246 , n19245 , n176 );
nand ( n19247 , n19239 , n19246 );
not ( n19248 , n177 );
not ( n19249 , n19248 );
not ( n19250 , n172 );
and ( n19251 , n19250 , n4713 );
not ( n19252 , n176 );
nand ( n19253 , n172 , n171 , n173 );
not ( n19254 , n19253 );
and ( n19255 , n19252 , n19254 );
nor ( n19256 , n19251 , n19255 );
and ( n19257 , n15871 , n4829 );
not ( n19258 , n5011 );
nor ( n19259 , n19258 , n4790 );
nand ( n19260 , n19256 , n19257 , n19259 );
not ( n19261 , n19260 );
or ( n19262 , n19249 , n19261 );
not ( n19263 , n173 );
not ( n19264 , n4809 );
or ( n19265 , n19263 , n19264 );
nand ( n19266 , n19265 , n4748 );
not ( n19267 , n5175 );
not ( n19268 , n4647 );
or ( n19269 , n19267 , n19268 );
or ( n19270 , n172 , n4869 );
nand ( n19271 , n19269 , n19270 );
or ( n19272 , n19266 , n19271 );
not ( n19273 , n176 );
nand ( n19274 , n19272 , n19273 );
nand ( n19275 , n19262 , n19274 );
or ( n19276 , n19247 , n19275 );
nand ( n19277 , n19276 , n4765 );
nand ( n19278 , n19225 , n19227 , n19277 );
not ( n19279 , n19278 );
and ( n19280 , n4660 , n5139 );
not ( n19281 , n5113 );
nand ( n19282 , n19281 , n176 );
not ( n19283 , n176 );
or ( n19284 , n19283 , n4815 );
nand ( n19285 , n19284 , n5070 , n5095 );
not ( n19286 , n176 );
not ( n19287 , n19286 );
nand ( n19288 , n12132 , n4957 , n4706 );
not ( n19289 , n19288 );
or ( n19290 , n19287 , n19289 );
nand ( n19291 , n19290 , n5133 );
or ( n19292 , n19285 , n19291 );
not ( n19293 , n177 );
nand ( n19294 , n19292 , n19293 );
and ( n19295 , n19280 , n12931 , n19282 , n19294 );
not ( n19296 , n15871 );
not ( n19297 , n4915 );
or ( n19298 , n19296 , n19297 );
not ( n19299 , n176 );
nand ( n19300 , n19298 , n19299 );
nand ( n19301 , n4949 , n15884 );
not ( n19302 , n176 );
nand ( n19303 , n4768 , n5150 , n15941 );
not ( n19304 , n19303 );
or ( n19305 , n19302 , n19304 );
not ( n19306 , n173 );
or ( n19307 , n19306 , n175 );
nand ( n19308 , n19307 , n12092 );
nand ( n19309 , n5179 , n19308 );
nand ( n19310 , n19305 , n19309 );
or ( n19311 , n19301 , n19310 );
nand ( n19312 , n19311 , n177 );
nand ( n19313 , n19300 , n19312 );
not ( n19314 , n176 );
not ( n19315 , n5123 );
nand ( n19316 , n12923 , n4760 , n19315 );
not ( n19317 , n19316 );
or ( n19318 , n19314 , n19317 );
and ( n19319 , n4706 , n12919 );
not ( n19320 , n19319 );
not ( n19321 , n19253 );
not ( n19322 , n5071 );
or ( n19323 , n19321 , n19322 );
nand ( n19324 , n19323 , n176 );
and ( n19325 , n12921 , n12085 , n19324 );
not ( n19326 , n19325 );
or ( n19327 , n19320 , n19326 );
not ( n19328 , n177 );
nand ( n19329 , n19327 , n19328 );
nand ( n19330 , n19318 , n19329 );
or ( n19331 , n19313 , n19330 );
nand ( n19332 , n19331 , n178 );
nand ( n19333 , n19279 , n19295 , n19332 );
not ( n19334 , n19333 );
not ( n19335 , n169 );
not ( n19336 , n19335 );
not ( n19337 , n10215 );
and ( n19338 , n167 , n19337 );
not ( n19339 , n5259 );
nor ( n19340 , n19338 , n19339 , n5315 );
not ( n19341 , n167 );
nand ( n19342 , n10704 , n10187 , n5570 );
nand ( n19343 , n19341 , n19342 );
nand ( n19344 , n19340 , n5389 , n19343 );
not ( n19345 , n19344 );
or ( n19346 , n19336 , n19345 );
not ( n19347 , n167 );
nor ( n19348 , n19347 , n5357 );
not ( n19349 , n17101 );
nor ( n19350 , n19348 , n19349 , n15749 );
not ( n19351 , n19350 );
not ( n19352 , n5379 );
not ( n19353 , n166 );
or ( n19354 , n19353 , n5459 );
not ( n19355 , n5427 );
nor ( n19356 , n19355 , n14874 );
nand ( n19357 , n19354 , n19356 );
not ( n19358 , n19357 );
or ( n19359 , n19352 , n19358 );
nand ( n19360 , n19359 , n5414 );
nor ( n19361 , n19351 , n19360 );
nand ( n19362 , n19346 , n19361 );
not ( n19363 , n19362 );
not ( n19364 , n169 );
or ( n19365 , n19364 , n10762 );
not ( n19366 , n15775 );
not ( n19367 , n5573 );
or ( n19368 , n19366 , n19367 );
nand ( n19369 , n19368 , n167 );
not ( n19370 , n5291 );
not ( n19371 , n166 );
not ( n19372 , n5406 );
nand ( n19373 , n19371 , n19372 );
not ( n19374 , n19373 );
or ( n19375 , n19370 , n19374 );
nand ( n19376 , n19375 , n167 );
not ( n19377 , n167 );
not ( n19378 , n5318 );
nand ( n19379 , n19377 , n5248 , n19378 );
nand ( n19380 , n19376 , n5549 , n19379 );
nand ( n19381 , n169 , n19380 );
nand ( n19382 , n19369 , n19381 );
not ( n19383 , n19382 );
not ( n19384 , n167 );
and ( n19385 , n5210 , n10237 );
not ( n19386 , n166 );
and ( n19387 , n19386 , n10683 );
nor ( n19388 , n19385 , n19387 );
nand ( n19389 , n165 , n14891 );
nand ( n19390 , n19388 , n5284 , n19389 );
nand ( n19391 , n19384 , n19390 );
or ( n19392 , n166 , n10268 );
nand ( n19393 , n163 , n5338 );
or ( n19394 , n167 , n19393 );
nand ( n19395 , n19392 , n19394 );
nor ( n19396 , n5658 , n10232 );
nand ( n19397 , n19396 , n14939 , n5573 );
or ( n19398 , n19395 , n19397 );
not ( n19399 , n169 );
nand ( n19400 , n19398 , n19399 );
nand ( n19401 , n19383 , n19391 , n19400 );
and ( n19402 , n5449 , n19401 );
not ( n19403 , n5449 );
not ( n19404 , n19393 );
not ( n19405 , n5245 );
or ( n19406 , n19404 , n19405 );
nand ( n19407 , n19406 , n5478 );
not ( n19408 , n14939 );
not ( n19409 , n5624 );
or ( n19410 , n19408 , n19409 );
not ( n19411 , n167 );
nand ( n19412 , n19410 , n19411 );
nand ( n19413 , n19407 , n19412 );
not ( n19414 , n169 );
not ( n19415 , n19414 );
nor ( n19416 , n17116 , n10679 );
nand ( n19417 , n19416 , n10187 , n17111 );
not ( n19418 , n19417 );
or ( n19419 , n19415 , n19418 );
nand ( n19420 , n19419 , n5343 );
nor ( n19421 , n19413 , n19420 );
not ( n19422 , n5379 );
nand ( n19423 , n5392 , n5459 , n14975 );
not ( n19424 , n19423 );
or ( n19425 , n19422 , n19424 );
nand ( n19426 , n169 , n15838 );
nand ( n19427 , n19425 , n19426 );
not ( n19428 , n19427 );
not ( n19429 , n165 );
nor ( n19430 , n19429 , n164 );
or ( n19431 , n19430 , n10685 );
nand ( n19432 , n19431 , n169 , n5451 );
not ( n19433 , n5504 );
not ( n19434 , n5397 );
or ( n19435 , n19433 , n19434 );
nand ( n19436 , n19435 , n167 );
nand ( n19437 , n19421 , n19428 , n19432 , n19436 );
and ( n19438 , n19403 , n19437 );
nor ( n19439 , n19402 , n19438 );
nand ( n19440 , n19363 , n19365 , n19439 );
not ( n19441 , n19440 );
not ( n19442 , n19441 );
or ( n19443 , n19334 , n19442 );
not ( n19444 , n178 );
not ( n19445 , n19300 );
not ( n19446 , n19445 );
nand ( n19447 , n176 , n19316 );
nand ( n19448 , n19446 , n19447 , n19329 , n19312 );
not ( n19449 , n19448 );
or ( n19450 , n19444 , n19449 );
nand ( n19451 , n19450 , n19295 );
nor ( n19452 , n19278 , n19451 );
nand ( n19453 , n19452 , n19440 );
nand ( n19454 , n19443 , n19453 );
not ( n19455 , n19454 );
and ( n19456 , n19221 , n19455 );
buf ( n19457 , n17020 );
and ( n19458 , n19457 , n19454 );
nor ( n19459 , n19456 , n19458 );
not ( n19460 , n19459 );
nand ( n19461 , n19220 , n19460 );
nand ( n19462 , n19219 , n19459 );
nand ( n19463 , n19461 , n2352 , n19462 );
nand ( n19464 , n19106 , n19463 );
not ( n19465 , n223 );
and ( n19466 , n224 , n19465 );
not ( n19467 , n224 );
and ( n19468 , n19467 , n223 );
nor ( n19469 , n19466 , n19468 );
or ( n19470 , n2352 , n19469 );
not ( n19471 , n194 );
nand ( n19472 , n193 , n12342 );
and ( n19473 , n19472 , n2373 , n2740 );
not ( n19474 , n193 );
nand ( n19475 , n2453 , n2589 , n2797 );
nand ( n19476 , n19474 , n19475 );
nand ( n19477 , n19473 , n16446 , n19476 );
nand ( n19478 , n19471 , n19477 );
and ( n19479 , n193 , n16517 );
nand ( n19480 , n9057 , n2709 );
nor ( n19481 , n19479 , n19480 );
not ( n19482 , n19481 );
not ( n19483 , n2516 );
not ( n19484 , n16464 );
nand ( n19485 , n191 , n19484 );
nand ( n19486 , n19485 , n2531 , n2551 );
not ( n19487 , n19486 );
or ( n19488 , n19483 , n19487 );
nand ( n19489 , n19488 , n16427 );
nor ( n19490 , n19482 , n19489 );
and ( n19491 , n19478 , n19490 );
not ( n19492 , n8963 );
nand ( n19493 , n194 , n19492 );
not ( n19494 , n2689 );
not ( n19495 , n2404 );
or ( n19496 , n19494 , n19495 );
nand ( n19497 , n19496 , n193 );
not ( n19498 , n2887 );
not ( n19499 , n193 );
and ( n19500 , n19499 , n9024 );
not ( n19501 , n19499 );
or ( n19502 , n191 , n9014 );
nand ( n19503 , n19502 , n2720 );
and ( n19504 , n19501 , n19503 );
nor ( n19505 , n19500 , n19504 );
not ( n19506 , n19505 );
or ( n19507 , n19498 , n19506 );
nand ( n19508 , n19507 , n194 );
nand ( n19509 , n19497 , n19508 );
not ( n19510 , n191 );
and ( n19511 , n19510 , n2804 );
not ( n19512 , n193 );
nor ( n19513 , n2376 , n2382 );
and ( n19514 , n19512 , n19513 );
nor ( n19515 , n19511 , n19514 );
and ( n19516 , n2486 , n2404 );
nor ( n19517 , n2861 , n12404 );
and ( n19518 , n19515 , n19516 , n19517 );
or ( n19519 , n194 , n19518 );
not ( n19520 , n193 );
not ( n19521 , n192 );
or ( n19522 , n19521 , n2445 );
not ( n19523 , n191 );
not ( n19524 , n2956 );
and ( n19525 , n19523 , n19524 );
and ( n19526 , n2780 , n12408 );
nor ( n19527 , n19525 , n19526 );
nand ( n19528 , n19522 , n19527 , n12358 );
nand ( n19529 , n19520 , n19528 );
nand ( n19530 , n19519 , n19529 );
or ( n19531 , n19509 , n19530 );
nand ( n19532 , n19531 , n2364 );
not ( n19533 , n193 );
nand ( n19534 , n2486 , n2932 );
and ( n19535 , n19533 , n19534 );
not ( n19536 , n19533 );
nand ( n19537 , n2498 , n12362 , n16443 );
and ( n19538 , n19536 , n19537 );
nor ( n19539 , n19535 , n19538 );
not ( n19540 , n19539 );
not ( n19541 , n194 );
nor ( n19542 , n9025 , n16844 );
or ( n19543 , n19513 , n2528 );
nand ( n19544 , n19543 , n193 );
nand ( n19545 , n2589 , n19542 , n9028 , n19544 );
and ( n19546 , n19541 , n19545 );
not ( n19547 , n19541 );
not ( n19548 , n192 );
or ( n19549 , n19548 , n189 );
not ( n19550 , n2625 );
nand ( n19551 , n19549 , n19550 );
nand ( n19552 , n2585 , n19551 );
not ( n19553 , n2955 );
nand ( n19554 , n19553 , n2576 , n16464 );
nand ( n19555 , n193 , n19554 );
nand ( n19556 , n19552 , n2791 , n19555 );
and ( n19557 , n19547 , n19556 );
nor ( n19558 , n19546 , n19557 );
not ( n19559 , n19558 );
or ( n19560 , n19540 , n19559 );
nand ( n19561 , n19560 , n195 );
nand ( n19562 , n19491 , n19493 , n19532 , n19561 );
not ( n19563 , n19562 );
and ( n19564 , n19563 , n19465 );
not ( n19565 , n19563 );
and ( n19566 , n19565 , n223 );
nor ( n19567 , n19564 , n19566 );
and ( n19568 , n186 , n8903 );
nand ( n19569 , n8822 , n3221 );
nor ( n19570 , n19568 , n19569 );
not ( n19571 , n184 );
or ( n19572 , n19571 , n8850 );
nand ( n19573 , n19572 , n3427 , n8777 );
nand ( n19574 , n3329 , n19573 );
nand ( n19575 , n19570 , n16319 , n19574 );
not ( n19576 , n19575 );
not ( n19577 , n3013 );
not ( n19578 , n11096 );
and ( n19579 , n185 , n19578 );
nand ( n19580 , n9182 , n3251 );
nor ( n19581 , n19579 , n19580 );
not ( n19582 , n185 );
nand ( n19583 , n16881 , n16895 , n3115 );
nand ( n19584 , n19582 , n19583 );
nand ( n19585 , n19581 , n16340 , n19584 );
not ( n19586 , n19585 );
or ( n19587 , n19577 , n19586 );
not ( n19588 , n185 );
or ( n19589 , n19588 , n9138 );
nand ( n19590 , n19587 , n19589 );
not ( n19591 , n19590 );
not ( n19592 , n186 );
nand ( n19593 , n9142 , n3235 , n8850 );
nand ( n19594 , n185 , n19593 );
not ( n19595 , n183 );
not ( n19596 , n3127 );
or ( n19597 , n19595 , n19596 );
nand ( n19598 , n19597 , n16924 );
nand ( n19599 , n3092 , n19598 );
nand ( n19600 , n19594 , n19599 , n3181 , n3184 );
not ( n19601 , n19600 );
or ( n19602 , n19592 , n19601 );
not ( n19603 , n3263 );
not ( n19604 , n3311 );
or ( n19605 , n19603 , n19604 );
not ( n19606 , n185 );
nand ( n19607 , n19605 , n19606 );
nand ( n19608 , n19602 , n19607 );
not ( n19609 , n19608 );
not ( n19610 , n3455 );
not ( n19611 , n16336 );
nand ( n19612 , n19610 , n3222 , n19611 );
nand ( n19613 , n185 , n19612 );
and ( n19614 , n16921 , n3071 , n8799 );
not ( n19615 , n3035 );
nand ( n19616 , n181 , n19615 );
not ( n19617 , n19616 );
not ( n19618 , n3202 );
or ( n19619 , n19617 , n19618 );
nand ( n19620 , n19619 , n185 );
nand ( n19621 , n19614 , n8814 , n19620 );
nand ( n19622 , n3013 , n19621 );
nand ( n19623 , n19609 , n19613 , n19622 );
and ( n19624 , n187 , n19623 );
not ( n19625 , n187 );
not ( n19626 , n3066 );
not ( n19627 , n3341 );
or ( n19628 , n19626 , n19627 );
nand ( n19629 , n19628 , n185 );
nand ( n19630 , n3263 , n3341 );
not ( n19631 , n185 );
not ( n19632 , n19616 );
and ( n19633 , n19631 , n19632 );
not ( n19634 , n184 );
and ( n19635 , n19634 , n3133 );
nor ( n19636 , n19633 , n19635 );
nand ( n19637 , n184 , n16326 );
nand ( n19638 , n19636 , n19637 , n11137 );
or ( n19639 , n19630 , n19638 );
nand ( n19640 , n19639 , n3013 );
not ( n19641 , n183 );
or ( n19642 , n19641 , n3123 );
nand ( n19643 , n19642 , n9135 );
or ( n19644 , n184 , n3276 );
nand ( n19645 , n3130 , n11141 );
nand ( n19646 , n19644 , n19645 );
or ( n19647 , n19643 , n19646 );
not ( n19648 , n185 );
nand ( n19649 , n19647 , n19648 );
not ( n19650 , n3432 );
not ( n19651 , n185 );
and ( n19652 , n19651 , n3455 );
not ( n19653 , n19651 );
not ( n19654 , n184 );
not ( n19655 , n19654 );
not ( n19656 , n8803 );
or ( n19657 , n19655 , n19656 );
nand ( n19658 , n19657 , n3213 );
and ( n19659 , n19653 , n19658 );
nor ( n19660 , n19652 , n19659 );
not ( n19661 , n19660 );
or ( n19662 , n19650 , n19661 );
nand ( n19663 , n19662 , n186 );
nand ( n19664 , n19629 , n19640 , n19649 , n19663 );
and ( n19665 , n19625 , n19664 );
nor ( n19666 , n19624 , n19665 );
nand ( n19667 , n19576 , n19591 , n19666 );
not ( n19668 , n19667 );
not ( n19669 , n19668 );
and ( n19670 , n19567 , n19669 );
not ( n19671 , n19567 );
and ( n19672 , n19671 , n19668 );
nor ( n19673 , n19670 , n19672 );
not ( n19674 , n19673 );
not ( n19675 , n203 );
and ( n19676 , n8312 , n3787 , n3939 );
or ( n19677 , n202 , n19676 );
not ( n19678 , n8381 );
and ( n19679 , n202 , n19678 );
not ( n19680 , n9662 );
nor ( n19681 , n19679 , n3757 , n19680 );
nand ( n19682 , n19677 , n19681 , n12636 );
and ( n19683 , n19675 , n19682 );
not ( n19684 , n19683 );
not ( n19685 , n201 );
or ( n19686 , n19685 , n11030 );
nand ( n19687 , n19686 , n8335 , n3865 );
nand ( n19688 , n3825 , n19687 );
and ( n19689 , n203 , n10967 );
not ( n19690 , n8294 );
nor ( n19691 , n19689 , n19690 );
not ( n19692 , n202 );
or ( n19693 , n19692 , n3948 );
and ( n19694 , n19693 , n11006 , n12632 );
nand ( n19695 , n19688 , n19691 , n19694 );
not ( n19696 , n19695 );
not ( n19697 , n3953 );
nand ( n19698 , n199 , n3759 );
nand ( n19699 , n19697 , n19698 );
nand ( n19700 , n203 , n9760 , n19699 );
and ( n19701 , n9678 , n19700 );
nand ( n19702 , n203 , n9739 );
nand ( n19703 , n3943 , n8346 , n3770 );
nand ( n19704 , n3825 , n19703 );
and ( n19705 , n19701 , n19702 , n19704 );
not ( n19706 , n203 );
nand ( n19707 , n8312 , n11011 , n11002 , n16652 );
and ( n19708 , n19706 , n19707 );
nand ( n19709 , n200 , n3776 );
not ( n19710 , n3938 );
and ( n19711 , n19709 , n19710 );
nor ( n19712 , n19711 , n3853 );
nor ( n19713 , n19708 , n19712 );
not ( n19714 , n9572 );
not ( n19715 , n3881 );
or ( n19716 , n19714 , n19715 );
not ( n19717 , n202 );
nand ( n19718 , n19716 , n19717 );
not ( n19719 , n3894 );
not ( n19720 , n12643 );
not ( n19721 , n19720 );
or ( n19722 , n19719 , n19721 );
nand ( n19723 , n19722 , n202 );
nand ( n19724 , n19705 , n19713 , n19718 , n19723 );
and ( n19725 , n204 , n19724 );
not ( n19726 , n204 );
not ( n19727 , n202 );
and ( n19728 , n19727 , n3893 );
not ( n19729 , n19727 );
not ( n19730 , n201 );
not ( n19731 , n19730 );
not ( n19732 , n11042 );
or ( n19733 , n19731 , n19732 );
nand ( n19734 , n19733 , n9630 );
and ( n19735 , n19729 , n19734 );
nor ( n19736 , n19728 , n19735 );
nand ( n19737 , n8412 , n19736 );
and ( n19738 , n203 , n19737 );
not ( n19739 , n9720 );
not ( n19740 , n3807 );
or ( n19741 , n19739 , n19740 );
nand ( n19742 , n19741 , n202 );
not ( n19743 , n19742 );
nor ( n19744 , n19738 , n19743 );
not ( n19745 , n202 );
or ( n19746 , n3758 , n3791 );
and ( n19747 , n9672 , n8400 );
not ( n19748 , n201 );
and ( n19749 , n19748 , n16655 );
nor ( n19750 , n19747 , n19749 );
nand ( n19751 , n19746 , n19750 , n3995 );
nand ( n19752 , n19745 , n19751 );
not ( n19753 , n203 );
not ( n19754 , n201 );
and ( n19755 , n19754 , n8285 );
not ( n19756 , n202 );
not ( n19757 , n19709 );
and ( n19758 , n19756 , n19757 );
nor ( n19759 , n19755 , n19758 );
nor ( n19760 , n9627 , n8394 );
nand ( n19761 , n19759 , n19760 , n3881 , n3807 );
nand ( n19762 , n19753 , n19761 );
nand ( n19763 , n19744 , n19752 , n19762 );
and ( n19764 , n19726 , n19763 );
nor ( n19765 , n19725 , n19764 );
nand ( n19766 , n19684 , n19696 , n19765 );
not ( n19767 , n19766 );
not ( n19768 , n8766 );
or ( n19769 , n19767 , n19768 );
not ( n19770 , n19766 );
nand ( n19771 , n19770 , n8925 );
nand ( n19772 , n19769 , n19771 );
and ( n19773 , n19772 , n10953 );
not ( n19774 , n19772 );
and ( n19775 , n19774 , n8921 );
nor ( n19776 , n19773 , n19775 );
not ( n19777 , n19776 );
nand ( n19778 , n19674 , n19777 );
nand ( n19779 , n19673 , n19776 );
nand ( n19780 , n19778 , n2352 , n19779 );
nand ( n19781 , n19470 , n19780 );
not ( n19782 , n136 );
and ( n19783 , n145 , n19782 );
not ( n19784 , n145 );
and ( n19785 , n19784 , n136 );
nor ( n19786 , n19783 , n19785 );
or ( n19787 , n2352 , n19786 );
and ( n19788 , n120 , n7812 );
nand ( n19789 , n8171 , n8204 );
nor ( n19790 , n19788 , n19789 );
not ( n19791 , n120 );
nand ( n19792 , n15414 , n8036 , n8106 );
nand ( n19793 , n19791 , n19792 );
and ( n19794 , n19790 , n8117 , n19793 );
not ( n19795 , n126 );
nor ( n19796 , n19794 , n19795 );
nand ( n19797 , n120 , n8226 );
and ( n19798 , n19797 , n18734 , n7671 );
not ( n19799 , n7703 );
nand ( n19800 , n121 , n19799 );
nand ( n19801 , n19800 , n8200 , n7802 );
nand ( n19802 , n8050 , n19801 );
nand ( n19803 , n19798 , n8129 , n19802 );
nor ( n19804 , n19796 , n19803 );
or ( n19805 , n126 , n18704 );
not ( n19806 , n126 );
not ( n19807 , n19806 );
not ( n19808 , n7921 );
not ( n19809 , n121 );
nand ( n19810 , n19809 , n8137 );
not ( n19811 , n19810 );
or ( n19812 , n19808 , n19811 );
nand ( n19813 , n19812 , n120 );
not ( n19814 , n120 );
nand ( n19815 , n19814 , n7994 );
nand ( n19816 , n19813 , n19815 , n7861 );
not ( n19817 , n19816 );
or ( n19818 , n19807 , n19817 );
not ( n19819 , n15334 );
not ( n19820 , n7789 );
or ( n19821 , n19819 , n19820 );
nand ( n19822 , n19821 , n120 );
nand ( n19823 , n19818 , n19822 );
not ( n19824 , n19823 );
not ( n19825 , n120 );
nand ( n19826 , n125 , n15396 );
nand ( n19827 , n8175 , n7845 );
nand ( n19828 , n7664 , n15334 , n19826 , n19827 );
nand ( n19829 , n19825 , n19828 );
not ( n19830 , n121 );
nor ( n19831 , n19830 , n8011 );
not ( n19832 , n19831 );
or ( n19833 , n120 , n19832 );
not ( n19834 , n7717 );
or ( n19835 , n121 , n19834 );
nand ( n19836 , n19833 , n19835 );
nand ( n19837 , n121 , n7756 );
and ( n19838 , n19837 , n7838 );
nand ( n19839 , n19838 , n15556 , n7789 );
or ( n19840 , n19836 , n19839 );
nand ( n19841 , n19840 , n126 );
nand ( n19842 , n19824 , n19829 , n19841 );
and ( n19843 , n7748 , n19842 );
not ( n19844 , n7748 );
not ( n19845 , n126 );
not ( n19846 , n19845 );
not ( n19847 , n8059 );
nand ( n19848 , n125 , n7659 );
nand ( n19849 , n19847 , n19848 );
and ( n19850 , n7813 , n19849 );
not ( n19851 , n19850 );
or ( n19852 , n19846 , n19851 );
or ( n19853 , n15553 , n8119 );
nand ( n19854 , n19853 , n120 );
nand ( n19855 , n19852 , n19854 );
not ( n19856 , n19855 );
not ( n19857 , n120 );
not ( n19858 , n19857 );
not ( n19859 , n8087 );
or ( n19860 , n19858 , n19859 );
or ( n19861 , n19831 , n15357 );
not ( n19862 , n7948 );
nand ( n19863 , n19861 , n19862 );
nand ( n19864 , n19860 , n19863 );
not ( n19865 , n126 );
nor ( n19866 , n8128 , n18756 );
not ( n19867 , n120 );
nand ( n19868 , n19867 , n7880 );
nand ( n19869 , n19866 , n19868 , n18745 );
not ( n19870 , n19869 );
or ( n19871 , n19865 , n19870 );
nand ( n19872 , n19871 , n15428 );
nor ( n19873 , n19864 , n19872 );
not ( n19874 , n8050 );
nand ( n19875 , n7770 , n8106 , n15449 );
not ( n19876 , n19875 );
or ( n19877 , n19874 , n19876 );
not ( n19878 , n126 );
nand ( n19879 , n19878 , n15389 );
nand ( n19880 , n19877 , n19879 );
not ( n19881 , n19880 );
nand ( n19882 , n19856 , n19873 , n19881 );
and ( n19883 , n19844 , n19882 );
nor ( n19884 , n19843 , n19883 );
nand ( n19885 , n19804 , n19805 , n19884 );
not ( n19886 , n19885 );
not ( n19887 , n18808 );
nand ( n19888 , n19887 , n18880 , n18806 );
not ( n19889 , n19888 );
not ( n19890 , n19889 );
or ( n19891 , n19886 , n19890 );
not ( n19892 , n19885 );
nand ( n19893 , n19888 , n19892 );
nand ( n19894 , n19891 , n19893 );
not ( n19895 , n19782 );
not ( n19896 , n7317 );
and ( n19897 , n19895 , n19896 );
and ( n19898 , n19782 , n7317 );
nor ( n19899 , n19897 , n19898 );
not ( n19900 , n11815 );
nand ( n19901 , n19900 , n11867 , n11911 );
not ( n19902 , n19901 );
not ( n19903 , n19902 );
not ( n19904 , n19903 );
not ( n19905 , n11573 );
or ( n19906 , n19904 , n19905 );
or ( n19907 , n11913 , n11573 );
nand ( n19908 , n19906 , n19907 );
and ( n19909 , n19899 , n19908 );
not ( n19910 , n19899 );
not ( n19911 , n19908 );
and ( n19912 , n19910 , n19911 );
nor ( n19913 , n19909 , n19912 );
not ( n19914 , n19913 );
nand ( n19915 , n19894 , n19914 );
not ( n19916 , n19894 );
nand ( n19917 , n19916 , n19913 );
nand ( n19918 , n19915 , n2352 , n19917 );
nand ( n19919 , n19787 , n19918 );
not ( n19920 , n240 );
and ( n19921 , n241 , n19920 );
not ( n19922 , n241 );
and ( n19923 , n19922 , n240 );
nor ( n19924 , n19921 , n19923 );
or ( n19925 , n2352 , n19924 );
not ( n19926 , n19920 );
not ( n19927 , n10926 );
and ( n19928 , n19926 , n19927 );
and ( n19929 , n19920 , n10913 );
nor ( n19930 , n19928 , n19929 );
not ( n19931 , n14864 );
and ( n19932 , n19930 , n19931 );
not ( n19933 , n19930 );
and ( n19934 , n19933 , n14864 );
nor ( n19935 , n19932 , n19934 );
not ( n19936 , n19935 );
not ( n19937 , n16236 );
not ( n19938 , n15022 );
and ( n19939 , n19937 , n19938 );
and ( n19940 , n16236 , n15022 );
nor ( n19941 , n19939 , n19940 );
not ( n19942 , n19941 );
nand ( n19943 , n19936 , n19942 );
nand ( n19944 , n19935 , n19941 );
nand ( n19945 , n19943 , n2352 , n19944 );
nand ( n19946 , n19925 , n19945 );
and ( n19947 , n19090 , n252 );
not ( n19948 , n19090 );
not ( n19949 , n252 );
and ( n19950 , n19948 , n19949 );
nor ( n19951 , n19947 , n19950 );
not ( n19952 , n135 );
not ( n19953 , n134 );
and ( n19954 , n15265 , n6929 );
nand ( n19955 , n19954 , n15292 , n6824 );
not ( n19956 , n19955 );
or ( n19957 , n19953 , n19956 );
not ( n19958 , n133 );
not ( n19959 , n7011 );
nand ( n19960 , n19959 , n7309 , n17237 );
nand ( n19961 , n19958 , n19960 );
nand ( n19962 , n19957 , n19961 );
not ( n19963 , n19962 );
not ( n19964 , n133 );
or ( n19965 , n19964 , n7041 );
nand ( n19966 , n19965 , n6984 );
not ( n19967 , n134 );
not ( n19968 , n19967 );
not ( n19969 , n7230 );
nand ( n19970 , n6840 , n6987 );
not ( n19971 , n19970 );
or ( n19972 , n19969 , n19971 );
nand ( n19973 , n19972 , n133 );
not ( n19974 , n19973 );
not ( n19975 , n133 );
not ( n19976 , n19975 );
not ( n19977 , n6994 );
or ( n19978 , n19976 , n19977 );
not ( n19979 , n7240 );
nand ( n19980 , n19978 , n19979 );
nor ( n19981 , n19974 , n19980 );
nand ( n19982 , n19981 , n7309 , n7041 );
not ( n19983 , n19982 );
or ( n19984 , n19968 , n19983 );
or ( n19985 , n6817 , n6872 );
nand ( n19986 , n19985 , n19024 , n17717 );
nand ( n19987 , n7298 , n19986 );
nand ( n19988 , n19984 , n19987 );
nor ( n19989 , n19966 , n19988 );
and ( n19990 , n17293 , n6834 );
nand ( n19991 , n19963 , n19989 , n19990 );
not ( n19992 , n19991 );
or ( n19993 , n19952 , n19992 );
not ( n19994 , n7007 );
not ( n19995 , n19994 );
not ( n19996 , n7077 );
nand ( n19997 , n19996 , n7195 );
nand ( n19998 , n19995 , n17245 , n19997 , n15250 );
not ( n19999 , n134 );
not ( n20000 , n19999 );
not ( n20001 , n6905 );
not ( n20002 , n7288 );
and ( n20003 , n20001 , n20002 );
nor ( n20004 , n20003 , n6991 );
not ( n20005 , n7041 );
nand ( n20006 , n7208 , n6918 );
not ( n20007 , n20006 );
or ( n20008 , n20005 , n20007 );
nand ( n20009 , n20008 , n133 );
not ( n20010 , n133 );
not ( n20011 , n132 );
nand ( n20012 , n20011 , n7138 );
not ( n20013 , n15270 );
nand ( n20014 , n20012 , n20013 , n7145 );
nand ( n20015 , n20010 , n20014 );
nand ( n20016 , n20004 , n20009 , n20015 );
not ( n20017 , n20016 );
or ( n20018 , n20000 , n20017 );
not ( n20019 , n132 );
not ( n20020 , n19047 );
or ( n20021 , n20019 , n20020 );
not ( n20022 , n133 );
nand ( n20023 , n20022 , n15197 );
nand ( n20024 , n20021 , n20023 );
nand ( n20025 , n134 , n20024 );
nand ( n20026 , n20018 , n20025 );
nor ( n20027 , n19998 , n20026 );
nand ( n20028 , n19993 , n20027 );
not ( n20029 , n20028 );
and ( n20030 , n19026 , n19029 );
not ( n20031 , n134 );
not ( n20032 , n20031 );
not ( n20033 , n132 );
not ( n20034 , n20033 );
not ( n20035 , n7302 );
or ( n20036 , n20034 , n20035 );
not ( n20037 , n17717 );
nand ( n20038 , n6906 , n20037 );
nand ( n20039 , n20036 , n20038 );
not ( n20040 , n20039 );
and ( n20041 , n20040 , n7072 , n19002 );
not ( n20042 , n20041 );
or ( n20043 , n20032 , n20042 );
not ( n20044 , n133 );
not ( n20045 , n20044 );
not ( n20046 , n132 );
nand ( n20047 , n20046 , n6855 );
nand ( n20048 , n20047 , n17807 , n7223 );
not ( n20049 , n20048 );
or ( n20050 , n20045 , n20049 );
nand ( n20051 , n20050 , n17191 );
not ( n20052 , n20051 );
and ( n20053 , n6859 , n7273 );
not ( n20054 , n132 );
or ( n20055 , n20054 , n17728 );
nand ( n20056 , n20053 , n20055 , n7186 );
not ( n20057 , n20056 );
not ( n20058 , n17914 );
not ( n20059 , n7220 );
or ( n20060 , n20058 , n20059 );
nand ( n20061 , n20060 , n133 );
nand ( n20062 , n20052 , n20057 , n20061 , n134 );
nand ( n20063 , n20043 , n20062 );
nand ( n20064 , n20030 , n19048 , n20063 );
not ( n20065 , n132 );
not ( n20066 , n20065 );
not ( n20067 , n7028 );
and ( n20068 , n20066 , n20067 );
nor ( n20069 , n20068 , n15172 );
not ( n20070 , n15224 );
nand ( n20071 , n20069 , n20055 , n20070 );
nand ( n20072 , n133 , n20071 );
nand ( n20073 , n20023 , n20072 );
or ( n20074 , n20064 , n20073 );
nand ( n20075 , n20074 , n7099 );
nand ( n20076 , n20029 , n20075 );
and ( n20077 , n19951 , n20076 );
not ( n20078 , n19951 );
not ( n20079 , n135 );
nor ( n20080 , n20073 , n20064 );
not ( n20081 , n20080 );
and ( n20082 , n20079 , n20081 );
nor ( n20083 , n20082 , n20028 );
and ( n20084 , n20078 , n20083 );
or ( n20085 , n20077 , n20084 );
not ( n20086 , n20085 );
not ( n20087 , n6808 );
nand ( n20088 , n142 , n11362 );
nand ( n20089 , n142 , n11317 );
nand ( n20090 , n6764 , n20088 , n20089 , n17542 );
nand ( n20091 , n141 , n20090 );
nor ( n20092 , n18909 , n18962 );
not ( n20093 , n141 );
nand ( n20094 , n20093 , n11956 );
and ( n20095 , n20091 , n20092 , n20094 , n18965 );
or ( n20096 , n142 , n17481 );
or ( n20097 , n6661 , n15083 );
nand ( n20098 , n20096 , n20097 );
not ( n20099 , n18898 );
nand ( n20100 , n20099 , n6742 );
or ( n20101 , n20098 , n20100 );
not ( n20102 , n144 );
nand ( n20103 , n20101 , n20102 );
nand ( n20104 , n20089 , n6688 , n11561 , n11548 );
not ( n20105 , n141 );
not ( n20106 , n142 );
not ( n20107 , n6623 );
nand ( n20108 , n20106 , n20107 );
nand ( n20109 , n20108 , n11286 , n11526 );
nand ( n20110 , n20105 , n20109 );
not ( n20111 , n6541 );
not ( n20112 , n6672 );
or ( n20113 , n20111 , n20112 );
nand ( n20114 , n20113 , n141 );
nand ( n20115 , n20110 , n11251 , n20114 );
or ( n20116 , n20104 , n20115 );
nand ( n20117 , n20116 , n144 );
nand ( n20118 , n20095 , n20103 , n20117 );
not ( n20119 , n20118 );
or ( n20120 , n20087 , n20119 );
not ( n20121 , n6553 );
or ( n20122 , n142 , n20121 );
nand ( n20123 , n20122 , n11922 , n6674 );
nand ( n20124 , n11268 , n20123 );
nand ( n20125 , n20120 , n20124 );
not ( n20126 , n20125 );
not ( n20127 , n144 );
not ( n20128 , n141 );
not ( n20129 , n6575 );
not ( n20130 , n11282 );
or ( n20131 , n20129 , n20130 );
nand ( n20132 , n20131 , n11369 );
not ( n20133 , n20132 );
or ( n20134 , n20128 , n20133 );
and ( n20135 , n11264 , n11475 );
nor ( n20136 , n20135 , n15096 );
nand ( n20137 , n20134 , n20136 );
nand ( n20138 , n20127 , n20137 );
not ( n20139 , n141 );
nand ( n20140 , n20139 , n11947 );
and ( n20141 , n20140 , n15074 , n11960 );
not ( n20142 , n142 );
not ( n20143 , n18909 );
or ( n20144 , n20142 , n20143 );
nand ( n20145 , n20144 , n20094 );
and ( n20146 , n144 , n20145 );
not ( n20147 , n11398 );
and ( n20148 , n11498 , n20147 );
nor ( n20149 , n20146 , n20148 );
and ( n20150 , n20138 , n20141 , n20149 );
not ( n20151 , n144 );
not ( n20152 , n142 );
not ( n20153 , n6549 );
or ( n20154 , n20152 , n20153 );
nand ( n20155 , n20154 , n6772 );
and ( n20156 , n141 , n20155 );
not ( n20157 , n141 );
and ( n20158 , n20157 , n6591 );
nor ( n20159 , n20156 , n20158 );
nand ( n20160 , n11535 , n11369 , n6702 , n20159 );
and ( n20161 , n20151 , n20160 );
not ( n20162 , n141 );
or ( n20163 , n20162 , n11369 );
not ( n20164 , n12008 );
nand ( n20165 , n20164 , n18961 , n15083 );
not ( n20166 , n141 );
nand ( n20167 , n20165 , n144 , n20166 );
and ( n20168 , n11985 , n20167 );
nand ( n20169 , n11329 , n11274 );
not ( n20170 , n20169 );
nand ( n20171 , n20163 , n20168 , n20170 );
nor ( n20172 , n20161 , n20171 );
not ( n20173 , n11335 );
not ( n20174 , n15076 );
or ( n20175 , n20173 , n20174 );
not ( n20176 , n141 );
nand ( n20177 , n20175 , n20176 );
nand ( n20178 , n17490 , n6611 );
nand ( n20179 , n11294 , n15072 );
or ( n20180 , n20178 , n20179 );
nand ( n20181 , n20180 , n144 );
nand ( n20182 , n20172 , n20177 , n20181 );
nand ( n20183 , n137 , n20182 );
nand ( n20184 , n20126 , n20150 , n20183 );
not ( n20185 , n20184 );
not ( n20186 , n20185 );
and ( n20187 , n19894 , n20186 );
not ( n20188 , n19894 );
not ( n20189 , n20185 );
not ( n20190 , n20189 );
and ( n20191 , n20188 , n20190 );
nor ( n20192 , n20187 , n20191 );
not ( n20193 , n20192 );
or ( n20194 , n20086 , n20193 );
nand ( n20195 , n20194 , n2352 );
nor ( n20196 , n20085 , n20192 );
or ( n20197 , n20195 , n20196 );
and ( n20198 , n253 , n19949 );
not ( n20199 , n253 );
and ( n20200 , n20199 , n252 );
nor ( n20201 , n20198 , n20200 );
or ( n20202 , n2352 , n20201 );
nand ( n20203 , n20197 , n20202 );
not ( n20204 , n260 );
not ( n20205 , n20204 );
not ( n20206 , n19215 );
or ( n20207 , n20205 , n20206 );
or ( n20208 , n20204 , n19215 );
nand ( n20209 , n20207 , n20208 );
and ( n20210 , n20209 , n19457 );
not ( n20211 , n20209 );
not ( n20212 , n19457 );
and ( n20213 , n20211 , n20212 );
nor ( n20214 , n20210 , n20213 );
not ( n20215 , n20214 );
buf ( n20216 , n17151 );
not ( n20217 , n20216 );
not ( n20218 , n20217 );
not ( n20219 , n4852 );
and ( n20220 , n20218 , n20219 );
and ( n20221 , n20217 , n4852 );
nor ( n20222 , n20220 , n20221 );
not ( n20223 , n20222 );
nor ( n20224 , n20215 , n20223 );
or ( n20225 , n20214 , n20222 );
nand ( n20226 , n20225 , n2352 );
or ( n20227 , n20224 , n20226 );
and ( n20228 , n261 , n20204 );
not ( n20229 , n261 );
and ( n20230 , n20229 , n260 );
nor ( n20231 , n20228 , n20230 );
or ( n20232 , n2352 , n20231 );
nand ( n20233 , n20227 , n20232 );
not ( n20234 , n1 );
xor ( n20235 , n265 , n266 );
not ( n20236 , n20235 );
or ( n20237 , n20234 , n20236 );
not ( n20238 , n265 );
not ( n20239 , n2650 );
not ( n20240 , n20239 );
and ( n20241 , n20238 , n20240 );
not ( n20242 , n2654 );
and ( n20243 , n265 , n20242 );
nor ( n20244 , n20241 , n20243 );
not ( n20245 , n16971 );
and ( n20246 , n20244 , n20245 );
not ( n20247 , n20244 );
not ( n20248 , n16985 );
and ( n20249 , n20247 , n20248 );
nor ( n20250 , n20246 , n20249 );
not ( n20251 , n20250 );
not ( n20252 , n4010 );
not ( n20253 , n20252 );
nand ( n20254 , n16551 , n16553 , n16554 , n8660 );
and ( n20255 , n3469 , n20254 );
nor ( n20256 , n20255 , n16621 );
nand ( n20257 , n20256 , n16580 , n16606 );
and ( n20258 , n20257 , n16731 );
not ( n20259 , n20257 );
and ( n20260 , n20259 , n16736 );
nor ( n20261 , n20258 , n20260 );
not ( n20262 , n20261 );
and ( n20263 , n20253 , n20262 );
and ( n20264 , n20252 , n20261 );
nor ( n20265 , n20263 , n20264 );
not ( n20266 , n20265 );
nand ( n20267 , n20251 , n20266 );
nand ( n20268 , n20250 , n20265 );
nand ( n20269 , n20267 , n2352 , n20268 );
nand ( n20270 , n20237 , n20269 );
not ( n20271 , n99 );
and ( n20272 , n269 , n20271 );
not ( n20273 , n269 );
and ( n20274 , n20273 , n99 );
nor ( n20275 , n20272 , n20274 );
or ( n20276 , n2352 , n20275 );
not ( n20277 , n18125 );
not ( n20278 , n16520 );
and ( n20279 , n20277 , n20278 );
and ( n20280 , n16866 , n16748 );
nor ( n20281 , n20279 , n20280 );
and ( n20282 , n12438 , n20271 );
not ( n20283 , n12438 );
and ( n20284 , n20283 , n99 );
nor ( n20285 , n20282 , n20284 );
not ( n20286 , n20285 );
and ( n20287 , n20281 , n20286 );
not ( n20288 , n20281 );
and ( n20289 , n20288 , n20285 );
nor ( n20290 , n20287 , n20289 );
not ( n20291 , n20290 );
not ( n20292 , n8614 );
nand ( n20293 , n16351 , n16373 , n16409 );
not ( n20294 , n20293 );
and ( n20295 , n3462 , n20294 );
not ( n20296 , n3462 );
and ( n20297 , n20296 , n20293 );
or ( n20298 , n20295 , n20297 );
not ( n20299 , n20298 );
or ( n20300 , n20292 , n20299 );
or ( n20301 , n8614 , n20298 );
nand ( n20302 , n20300 , n20301 );
not ( n20303 , n20302 );
nand ( n20304 , n20291 , n20303 );
nand ( n20305 , n20290 , n20302 );
nand ( n20306 , n20304 , n2352 , n20305 );
nand ( n20307 , n20276 , n20306 );
not ( n20308 , n276 );
and ( n20309 , n277 , n20308 );
not ( n20310 , n277 );
and ( n20311 , n20310 , n276 );
nor ( n20312 , n20309 , n20311 );
or ( n20313 , n2352 , n20312 );
not ( n20314 , n17432 );
not ( n20315 , n11409 );
and ( n20316 , n20314 , n20315 );
not ( n20317 , n17430 );
and ( n20318 , n17374 , n17378 , n17381 , n20317 );
and ( n20319 , n11409 , n20318 );
nor ( n20320 , n20316 , n20319 );
and ( n20321 , n7089 , n20308 );
not ( n20322 , n7089 );
and ( n20323 , n20322 , n276 );
nor ( n20324 , n20321 , n20323 );
and ( n20325 , n20320 , n20324 );
not ( n20326 , n20320 );
not ( n20327 , n20324 );
and ( n20328 , n20326 , n20327 );
nor ( n20329 , n20325 , n20328 );
not ( n20330 , n20329 );
not ( n20331 , n126 );
not ( n20332 , n20331 );
or ( n20333 , n7655 , n8057 );
nand ( n20334 , n20333 , n120 );
not ( n20335 , n120 );
nand ( n20336 , n15385 , n15320 , n8136 );
nand ( n20337 , n20335 , n20336 );
nand ( n20338 , n20334 , n8036 , n20337 );
not ( n20339 , n20338 );
or ( n20340 , n20332 , n20339 );
not ( n20341 , n7662 );
and ( n20342 , n120 , n8175 , n20341 );
nor ( n20343 , n20342 , n8128 );
nand ( n20344 , n20340 , n20343 );
not ( n20345 , n20344 );
not ( n20346 , n7928 );
nand ( n20347 , n20346 , n7972 );
nand ( n20348 , n20347 , n7921 );
nand ( n20349 , n126 , n20348 );
nand ( n20350 , n20345 , n18704 , n20349 );
nand ( n20351 , n20350 , n7748 );
not ( n20352 , n20351 );
not ( n20353 , n8050 );
or ( n20354 , n121 , n8011 );
nand ( n20355 , n20354 , n15407 );
not ( n20356 , n20355 );
or ( n20357 , n20353 , n20356 );
nand ( n20358 , n7755 , n7975 );
nand ( n20359 , n20358 , n120 , n7635 );
nand ( n20360 , n20357 , n20359 );
not ( n20361 , n8227 );
and ( n20362 , n20361 , n7736 );
not ( n20363 , n7895 );
nand ( n20364 , n15486 , n7670 );
not ( n20365 , n20364 );
not ( n20366 , n7965 );
or ( n20367 , n20365 , n20366 );
not ( n20368 , n120 );
nand ( n20369 , n20367 , n20368 );
not ( n20370 , n120 );
nand ( n20371 , n20370 , n7897 );
nand ( n20372 , n20363 , n20369 , n20371 );
nor ( n20373 , n20362 , n20372 );
or ( n20374 , n20373 , n126 );
nand ( n20375 , n20374 , n8111 );
nor ( n20376 , n20352 , n20360 , n20375 );
not ( n20377 , n120 );
not ( n20378 , n20377 );
nand ( n20379 , n7961 , n8171 , n7861 );
not ( n20380 , n20379 );
or ( n20381 , n20378 , n20380 );
nand ( n20382 , n20381 , n19868 );
nand ( n20383 , n121 , n15333 );
nand ( n20384 , n121 , n8059 );
nand ( n20385 , n20384 , n7921 , n7898 );
nand ( n20386 , n120 , n20385 );
nand ( n20387 , n20383 , n8228 , n20386 );
or ( n20388 , n20382 , n20387 );
nand ( n20389 , n20388 , n126 );
not ( n20390 , n7923 );
nand ( n20391 , n15414 , n20390 , n15523 );
nand ( n20392 , n8148 , n20391 );
not ( n20393 , n126 );
not ( n20394 , n120 );
not ( n20395 , n123 );
not ( n20396 , n7633 );
not ( n20397 , n20396 );
or ( n20398 , n20395 , n20397 );
nand ( n20399 , n20398 , n8060 );
nand ( n20400 , n20394 , n20399 );
not ( n20401 , n7811 );
nand ( n20402 , n120 , n20401 );
nand ( n20403 , n20400 , n20402 , n15348 );
nand ( n20404 , n20393 , n20403 );
nand ( n20405 , n20392 , n20404 );
and ( n20406 , n7863 , n15352 );
and ( n20407 , n7881 , n7761 );
not ( n20408 , n18675 );
not ( n20409 , n8068 );
and ( n20410 , n120 , n20409 );
not ( n20411 , n120 );
and ( n20412 , n20411 , n8199 );
nor ( n20413 , n20410 , n20412 );
nand ( n20414 , n7718 , n7930 );
nor ( n20415 , n7679 , n20414 );
nand ( n20416 , n20407 , n20408 , n20413 , n20415 );
nand ( n20417 , n126 , n20416 );
nand ( n20418 , n20406 , n15465 , n20417 );
or ( n20419 , n20405 , n20418 );
nand ( n20420 , n20419 , n127 );
nand ( n20421 , n20376 , n20389 , n20420 );
not ( n20422 , n20421 );
not ( n20423 , n8100 );
and ( n20424 , n20422 , n20423 );
not ( n20425 , n20422 );
not ( n20426 , n15439 );
and ( n20427 , n20425 , n20426 );
nor ( n20428 , n20424 , n20427 );
not ( n20429 , n20428 );
and ( n20430 , n11636 , n11657 , n11752 );
not ( n20431 , n20430 );
not ( n20432 , n11913 );
not ( n20433 , n20432 );
and ( n20434 , n20431 , n20433 );
not ( n20435 , n11913 );
and ( n20436 , n20430 , n20435 );
nor ( n20437 , n20434 , n20436 );
not ( n20438 , n20437 );
and ( n20439 , n20429 , n20438 );
and ( n20440 , n20428 , n20437 );
nor ( n20441 , n20439 , n20440 );
not ( n20442 , n20441 );
nand ( n20443 , n20330 , n20442 );
nand ( n20444 , n20329 , n20441 );
nand ( n20445 , n20443 , n2352 , n20444 );
nand ( n20446 , n20313 , n20445 );
not ( n20447 , n18905 );
nand ( n20448 , n20447 , n18895 , n18982 );
xor ( n20449 , n282 , n20448 );
xnor ( n20450 , n20449 , n20083 );
buf ( n20451 , n18774 );
xor ( n20452 , n20451 , n19894 );
nor ( n20453 , n20450 , n20452 );
not ( n20454 , n20450 );
not ( n20455 , n20452 );
or ( n20456 , n20454 , n20455 );
nand ( n20457 , n20456 , n2352 );
or ( n20458 , n20453 , n20457 );
xnor ( n20459 , n282 , n283 );
or ( n20460 , n2352 , n20459 );
nand ( n20461 , n20458 , n20460 );
not ( n20462 , n288 );
and ( n20463 , n289 , n20462 );
not ( n20464 , n289 );
and ( n20465 , n20464 , n288 );
nor ( n20466 , n20463 , n20465 );
or ( n20467 , n2352 , n20466 );
not ( n20468 , n14858 );
not ( n20469 , n20462 );
and ( n20470 , n20468 , n20469 );
and ( n20471 , n20462 , n14864 );
nor ( n20472 , n20470 , n20471 );
not ( n20473 , n20472 );
not ( n20474 , n16105 );
not ( n20475 , n20474 );
not ( n20476 , n10159 );
not ( n20477 , n20476 );
or ( n20478 , n20475 , n20477 );
or ( n20479 , n16106 , n20476 );
nand ( n20480 , n20478 , n20479 );
not ( n20481 , n20480 );
or ( n20482 , n20473 , n20481 );
or ( n20483 , n20472 , n20480 );
nand ( n20484 , n20482 , n20483 );
and ( n20485 , n149 , n10555 );
not ( n20486 , n149 );
nand ( n20487 , n148 , n12237 );
and ( n20488 , n20486 , n20487 );
nor ( n20489 , n20485 , n20488 );
not ( n20490 , n149 );
not ( n20491 , n20490 );
not ( n20492 , n13025 );
not ( n20493 , n150 );
nand ( n20494 , n20492 , n20493 );
nand ( n20495 , n20494 , n10386 , n10378 );
not ( n20496 , n20495 );
or ( n20497 , n20491 , n20496 );
or ( n20498 , n4498 , n12202 );
not ( n20499 , n10332 );
nand ( n20500 , n20498 , n149 , n20499 );
nand ( n20501 , n20497 , n20500 );
not ( n20502 , n4459 );
not ( n20503 , n20502 );
not ( n20504 , n4473 );
not ( n20505 , n20504 );
or ( n20506 , n20503 , n20505 );
nand ( n20507 , n20506 , n20487 );
not ( n20508 , n20507 );
nand ( n20509 , n12200 , n10317 );
nand ( n20510 , n20508 , n20509 , n13057 , n10620 );
nand ( n20511 , n152 , n20510 );
or ( n20512 , n150 , n4305 );
nand ( n20513 , n20512 , n4326 );
nand ( n20514 , n10561 , n20513 );
not ( n20515 , n150 );
not ( n20516 , n20515 );
not ( n20517 , n10633 );
or ( n20518 , n20516 , n20517 );
not ( n20519 , n4313 );
nand ( n20520 , n20518 , n20519 );
nand ( n20521 , n4532 , n20520 );
nand ( n20522 , n20511 , n20514 , n20521 );
nor ( n20523 , n20501 , n20522 );
or ( n20524 , n153 , n20523 );
not ( n20525 , n149 );
not ( n20526 , n150 );
nand ( n20527 , n20526 , n4454 );
nand ( n20528 , n20527 , n4412 , n4509 );
and ( n20529 , n20525 , n20528 );
not ( n20530 , n20525 );
nand ( n20531 , n10437 , n4566 );
and ( n20532 , n20530 , n20531 );
nor ( n20533 , n20529 , n20532 );
nand ( n20534 , n20533 , n12966 , n12265 );
nand ( n20535 , n4532 , n20534 );
nand ( n20536 , n20524 , n20535 );
nor ( n20537 , n20489 , n20536 );
not ( n20538 , n149 );
not ( n20539 , n13059 );
or ( n20540 , n20538 , n20539 );
or ( n20541 , n149 , n12231 );
nand ( n20542 , n20540 , n20541 );
nand ( n20543 , n10430 , n4380 , n4394 , n20542 );
nand ( n20544 , n152 , n20543 );
not ( n20545 , n10448 );
not ( n20546 , n10625 );
or ( n20547 , n20545 , n20546 );
not ( n20548 , n149 );
nand ( n20549 , n20547 , n20548 );
or ( n20550 , n149 , n4464 );
nand ( n20551 , n20550 , n10339 , n10406 );
nand ( n20552 , n152 , n20551 );
and ( n20553 , n10507 , n4422 );
nand ( n20554 , n20553 , n10378 , n12997 );
nand ( n20555 , n149 , n20554 );
nand ( n20556 , n20549 , n20552 , n20555 );
and ( n20557 , n4520 , n4424 );
not ( n20558 , n149 );
not ( n20559 , n150 );
not ( n20560 , n16130 );
or ( n20561 , n20559 , n20560 );
nand ( n20562 , n20561 , n12239 );
nand ( n20563 , n20558 , n20562 );
not ( n20564 , n10317 );
not ( n20565 , n4563 );
or ( n20566 , n20564 , n20565 );
nand ( n20567 , n4350 , n10331 );
and ( n20568 , n20567 , n10515 );
nand ( n20569 , n20566 , n20568 );
not ( n20570 , n149 );
nand ( n20571 , n4442 , n10599 , n16135 );
not ( n20572 , n20571 );
or ( n20573 , n20570 , n20572 );
nand ( n20574 , n20573 , n12995 );
or ( n20575 , n20569 , n20574 );
nand ( n20576 , n20575 , n4532 );
nand ( n20577 , n20557 , n20563 , n20576 );
or ( n20578 , n20556 , n20577 );
nand ( n20579 , n20578 , n153 );
nand ( n20580 , n20537 , n20544 , n20579 );
not ( n20581 , n20580 );
not ( n20582 , n20581 );
not ( n20583 , n10659 );
or ( n20584 , n20582 , n20583 );
nand ( n20585 , n20580 , n10654 );
nand ( n20586 , n20584 , n20585 );
and ( n20587 , n20586 , n15978 );
not ( n20588 , n20586 );
and ( n20589 , n20588 , n15995 );
nor ( n20590 , n20587 , n20589 );
nor ( n20591 , n20484 , n20590 );
not ( n20592 , n20591 );
nand ( n20593 , n20484 , n20590 );
nand ( n20594 , n20592 , n20593 , n2352 );
nand ( n20595 , n20467 , n20594 );
not ( n20596 , n294 );
and ( n20597 , n295 , n20596 );
not ( n20598 , n295 );
and ( n20599 , n20598 , n294 );
nor ( n20600 , n20597 , n20599 );
or ( n20601 , n2352 , n20600 );
xor ( n20602 , n20596 , n2650 );
not ( n20603 , n16987 );
and ( n20604 , n9239 , n20603 );
not ( n20605 , n9239 );
not ( n20606 , n16980 );
and ( n20607 , n20605 , n20606 );
nor ( n20608 , n20604 , n20607 );
and ( n20609 , n20602 , n20608 );
not ( n20610 , n20602 );
not ( n20611 , n20608 );
and ( n20612 , n20610 , n20611 );
nor ( n20613 , n20609 , n20612 );
not ( n20614 , n20613 );
not ( n20615 , n3273 );
not ( n20616 , n9512 );
and ( n20617 , n20615 , n20616 );
and ( n20618 , n3273 , n9509 );
nor ( n20619 , n20617 , n20618 );
not ( n20620 , n20619 );
not ( n20621 , n9369 );
not ( n20622 , n4011 );
or ( n20623 , n20621 , n20622 );
or ( n20624 , n9369 , n20252 );
nand ( n20625 , n20623 , n20624 );
not ( n20626 , n20625 );
and ( n20627 , n20620 , n20626 );
and ( n20628 , n20619 , n20625 );
nor ( n20629 , n20627 , n20628 );
not ( n20630 , n20629 );
nand ( n20631 , n20614 , n20630 );
nand ( n20632 , n20613 , n20629 );
nand ( n20633 , n20631 , n2352 , n20632 );
nand ( n20634 , n20601 , n20633 );
not ( n20635 , n307 );
not ( n20636 , n20635 );
not ( n20637 , n17992 );
or ( n20638 , n20636 , n20637 );
or ( n20639 , n17996 , n20635 );
nand ( n20640 , n20638 , n20639 );
not ( n20641 , n20640 );
not ( n20642 , n6811 );
nor ( n20643 , n7495 , n7621 );
not ( n20644 , n20643 );
and ( n20645 , n20642 , n20644 );
and ( n20646 , n7093 , n20643 );
nor ( n20647 , n20645 , n20646 );
not ( n20648 , n20647 );
not ( n20649 , n20648 );
or ( n20650 , n20641 , n20649 );
not ( n20651 , n20640 );
nand ( n20652 , n20651 , n20647 );
nand ( n20653 , n20650 , n20652 );
not ( n20654 , n8251 );
not ( n20655 , n20318 );
not ( n20656 , n11913 );
not ( n20657 , n20656 );
and ( n20658 , n20655 , n20657 );
and ( n20659 , n20656 , n20318 );
nor ( n20660 , n20658 , n20659 );
not ( n20661 , n20660 );
or ( n20662 , n20654 , n20661 );
or ( n20663 , n8251 , n20660 );
nand ( n20664 , n20662 , n20663 );
or ( n20665 , n20653 , n20664 );
nand ( n20666 , n20665 , n2352 );
not ( n20667 , n20653 );
not ( n20668 , n20664 );
nor ( n20669 , n20667 , n20668 );
or ( n20670 , n20666 , n20669 );
and ( n20671 , n308 , n20635 );
not ( n20672 , n308 );
and ( n20673 , n20672 , n307 );
nor ( n20674 , n20671 , n20673 );
or ( n20675 , n2352 , n20674 );
nand ( n20676 , n20670 , n20675 );
not ( n20677 , n16234 );
and ( n20678 , n313 , n20677 );
not ( n20679 , n313 );
and ( n20680 , n20679 , n16234 );
nor ( n20681 , n20678 , n20680 );
not ( n20682 , n20489 );
not ( n20683 , n20536 );
nand ( n20684 , n20682 , n20683 , n20544 , n20579 );
not ( n20685 , n20684 );
not ( n20686 , n20685 );
not ( n20687 , n176 );
not ( n20688 , n20687 );
not ( n20689 , n172 );
nand ( n20690 , n20689 , n5072 );
nand ( n20691 , n20690 , n4825 , n4588 );
not ( n20692 , n20691 );
or ( n20693 , n20688 , n20692 );
nand ( n20694 , n20693 , n12120 );
or ( n20695 , n12892 , n20694 );
not ( n20696 , n177 );
nand ( n20697 , n20695 , n20696 );
and ( n20698 , n176 , n4995 );
not ( n20699 , n176 );
nor ( n20700 , n4679 , n4699 );
and ( n20701 , n20699 , n20700 );
nor ( n20702 , n20698 , n20701 );
not ( n20703 , n5095 );
not ( n20704 , n4629 );
or ( n20705 , n20703 , n20704 );
nand ( n20706 , n20705 , n5006 );
nand ( n20707 , n4734 , n4660 );
and ( n20708 , n176 , n12913 );
not ( n20709 , n176 );
and ( n20710 , n20709 , n5017 );
or ( n20711 , n20708 , n20710 );
nand ( n20712 , n20711 , n5091 );
or ( n20713 , n20707 , n20712 );
nand ( n20714 , n20713 , n177 );
and ( n20715 , n20697 , n20702 , n20706 , n20714 );
not ( n20716 , n177 );
not ( n20717 , n172 );
not ( n20718 , n20717 );
nand ( n20719 , n4606 , n4841 );
not ( n20720 , n20719 );
or ( n20721 , n20718 , n20720 );
nand ( n20722 , n20721 , n4686 );
nand ( n20723 , n20716 , n20722 );
or ( n20724 , n172 , n4688 );
nand ( n20725 , n20724 , n4782 );
and ( n20726 , n5006 , n20725 );
not ( n20727 , n4593 );
not ( n20728 , n4587 );
not ( n20729 , n20728 );
or ( n20730 , n20727 , n20729 );
not ( n20731 , n176 );
nor ( n20732 , n20731 , n4755 );
nand ( n20733 , n20730 , n20732 );
not ( n20734 , n20733 );
nor ( n20735 , n20726 , n20734 );
nand ( n20736 , n20723 , n20735 );
not ( n20737 , n20736 );
not ( n20738 , n176 );
nand ( n20739 , n19242 , n5085 , n5088 );
nand ( n20740 , n20738 , n20739 );
not ( n20741 , n4889 );
nor ( n20742 , n20741 , n20700 );
not ( n20743 , n4646 );
nand ( n20744 , n20743 , n5179 );
nand ( n20745 , n176 , n4615 );
nand ( n20746 , n20742 , n20744 , n12909 , n20745 );
nand ( n20747 , n177 , n20746 );
nand ( n20748 , n20737 , n20740 , n20747 );
nand ( n20749 , n4765 , n20748 );
not ( n20750 , n177 );
or ( n20751 , n176 , n4833 );
nand ( n20752 , n20751 , n12132 , n5056 );
not ( n20753 , n20752 );
or ( n20754 , n20750 , n20753 );
not ( n20755 , n176 );
nand ( n20756 , n4976 , n4900 );
and ( n20757 , n20755 , n20756 );
not ( n20758 , n20755 );
and ( n20759 , n4949 , n4668 );
nand ( n20760 , n20759 , n5088 , n15884 );
and ( n20761 , n20758 , n20760 );
nor ( n20762 , n20757 , n20761 );
nand ( n20763 , n20754 , n20762 );
nand ( n20764 , n12877 , n4929 );
nor ( n20765 , n175 , n4755 );
not ( n20766 , n20765 );
nand ( n20767 , n5179 , n12928 );
not ( n20768 , n15924 );
nand ( n20769 , n4664 , n4577 );
or ( n20770 , n20768 , n20769 );
nand ( n20771 , n20770 , n176 );
nand ( n20772 , n20766 , n20767 , n20771 );
nor ( n20773 , n20764 , n20772 );
or ( n20774 , n177 , n20773 );
nand ( n20775 , n172 , n15920 );
and ( n20776 , n12066 , n20775 );
or ( n20777 , n176 , n20776 );
not ( n20778 , n15910 );
nor ( n20779 , n20778 , n4670 );
nand ( n20780 , n20774 , n20777 , n20779 );
or ( n20781 , n20763 , n20780 );
nand ( n20782 , n20781 , n178 );
nand ( n20783 , n20715 , n20749 , n20782 );
not ( n20784 , n20783 );
or ( n20785 , n20686 , n20784 );
not ( n20786 , n20783 );
nand ( n20787 , n20580 , n20786 );
nand ( n20788 , n20785 , n20787 );
not ( n20789 , n12161 );
not ( n20790 , n5664 );
or ( n20791 , n20789 , n20790 );
nand ( n20792 , n5040 , n5669 );
nand ( n20793 , n20791 , n20792 );
xor ( n20794 , n20788 , n20793 );
nor ( n20795 , n20681 , n20794 );
not ( n20796 , n20681 );
not ( n20797 , n20794 );
or ( n20798 , n20796 , n20797 );
nand ( n20799 , n20798 , n2352 );
or ( n20800 , n20795 , n20799 );
xnor ( n20801 , n313 , n314 );
or ( n20802 , n2352 , n20801 );
nand ( n20803 , n20800 , n20802 );
not ( n20804 , n316 );
and ( n20805 , n317 , n20804 );
not ( n20806 , n317 );
and ( n20807 , n20806 , n316 );
nor ( n20808 , n20805 , n20807 );
or ( n20809 , n2352 , n20808 );
not ( n20810 , n20804 );
not ( n20811 , n16520 );
or ( n20812 , n20810 , n20811 );
or ( n20813 , n20804 , n16526 );
nand ( n20814 , n20812 , n20813 );
not ( n20815 , n20298 );
and ( n20816 , n20814 , n20815 );
not ( n20817 , n20814 );
and ( n20818 , n20817 , n20298 );
nor ( n20819 , n20816 , n20818 );
not ( n20820 , n20819 );
and ( n20821 , n12674 , n16628 );
not ( n20822 , n12674 );
not ( n20823 , n16628 );
and ( n20824 , n20822 , n20823 );
nor ( n20825 , n20821 , n20824 );
not ( n20826 , n16971 );
not ( n20827 , n9509 );
and ( n20828 , n20826 , n20827 );
and ( n20829 , n16971 , n12449 );
nor ( n20830 , n20828 , n20829 );
and ( n20831 , n20825 , n20830 );
not ( n20832 , n20825 );
not ( n20833 , n20830 );
and ( n20834 , n20832 , n20833 );
nor ( n20835 , n20831 , n20834 );
not ( n20836 , n20835 );
nand ( n20837 , n20820 , n20836 );
nand ( n20838 , n20819 , n20835 );
nand ( n20839 , n20837 , n2352 , n20838 );
nand ( n20840 , n20809 , n20839 );
not ( n20841 , n318 );
not ( n20842 , n20841 );
not ( n20843 , n14858 );
or ( n20844 , n20842 , n20843 );
or ( n20845 , n20841 , n14864 );
nand ( n20846 , n20844 , n20845 );
not ( n20847 , n10654 );
not ( n20848 , n16235 );
or ( n20849 , n20847 , n20848 );
nand ( n20850 , n10659 , n16231 );
nand ( n20851 , n20849 , n20850 );
not ( n20852 , n20851 );
and ( n20853 , n20846 , n20852 );
not ( n20854 , n20846 );
and ( n20855 , n20854 , n20851 );
nor ( n20856 , n20853 , n20855 );
not ( n20857 , n20856 );
not ( n20858 , n20684 );
not ( n20859 , n20858 );
not ( n20860 , n5042 );
or ( n20861 , n20859 , n20860 );
or ( n20862 , n20858 , n5200 );
nand ( n20863 , n20861 , n20862 );
not ( n20864 , n20863 );
not ( n20865 , n20786 );
not ( n20866 , n15974 );
and ( n20867 , n20865 , n20866 );
and ( n20868 , n20786 , n15013 );
nor ( n20869 , n20867 , n20868 );
not ( n20870 , n20869 );
and ( n20871 , n20864 , n20870 );
and ( n20872 , n20863 , n20869 );
nor ( n20873 , n20871 , n20872 );
not ( n20874 , n20873 );
nor ( n20875 , n20857 , n20874 );
or ( n20876 , n20856 , n20873 );
nand ( n20877 , n20876 , n2352 );
or ( n20878 , n20875 , n20877 );
and ( n20879 , n319 , n20841 );
not ( n20880 , n319 );
and ( n20881 , n20880 , n318 );
nor ( n20882 , n20879 , n20881 );
or ( n20883 , n2352 , n20882 );
nand ( n20884 , n20878 , n20883 );
and ( n20885 , n328 , n18080 );
not ( n20886 , n328 );
and ( n20887 , n20886 , n18083 );
nor ( n20888 , n20885 , n20887 );
not ( n20889 , n20888 );
not ( n20890 , n9774 );
not ( n20891 , n9509 );
or ( n20892 , n20890 , n20891 );
or ( n20893 , n18118 , n12449 );
nand ( n20894 , n20892 , n20893 );
and ( n20895 , n3468 , n20894 );
not ( n20896 , n3468 );
not ( n20897 , n20894 );
and ( n20898 , n20896 , n20897 );
nor ( n20899 , n20895 , n20898 );
not ( n20900 , n20899 );
nor ( n20901 , n20889 , n20900 );
or ( n20902 , n20888 , n20899 );
nand ( n20903 , n20902 , n2352 );
or ( n20904 , n20901 , n20903 );
xnor ( n20905 , n328 , n329 );
or ( n20906 , n2352 , n20905 );
nand ( n20907 , n20904 , n20906 );
not ( n20908 , n336 );
and ( n20909 , n337 , n20908 );
not ( n20910 , n337 );
and ( n20911 , n20910 , n336 );
nor ( n20912 , n20909 , n20911 );
or ( n20913 , n2352 , n20912 );
not ( n20914 , n20908 );
not ( n20915 , n14707 );
and ( n20916 , n20914 , n20915 );
and ( n20917 , n20908 , n14707 );
nor ( n20918 , n20916 , n20917 );
not ( n20919 , n20918 );
and ( n20920 , n20788 , n15851 );
not ( n20921 , n20788 );
and ( n20922 , n20921 , n15985 );
nor ( n20923 , n20920 , n20922 );
not ( n20924 , n20923 );
nand ( n20925 , n20919 , n20924 );
nand ( n20926 , n20918 , n20923 );
nand ( n20927 , n20925 , n2352 , n20926 );
nand ( n20928 , n20913 , n20927 );
xor ( n20929 , n363 , n20076 );
xnor ( n20930 , n20929 , n20185 );
and ( n20931 , n20451 , n20647 );
not ( n20932 , n20451 );
and ( n20933 , n20932 , n20648 );
nor ( n20934 , n20931 , n20933 );
nor ( n20935 , n20930 , n20934 );
not ( n20936 , n20930 );
not ( n20937 , n20934 );
or ( n20938 , n20936 , n20937 );
nand ( n20939 , n20938 , n2352 );
or ( n20940 , n20935 , n20939 );
xnor ( n20941 , n363 , n364 );
or ( n20942 , n2352 , n20941 );
nand ( n20943 , n20940 , n20942 );
not ( n20944 , n369 );
and ( n20945 , n12434 , n20944 );
not ( n20946 , n12434 );
and ( n20947 , n20946 , n369 );
nor ( n20948 , n20945 , n20947 );
and ( n20949 , n20948 , n10958 );
not ( n20950 , n20948 );
and ( n20951 , n20950 , n8921 );
nor ( n20952 , n20949 , n20951 );
not ( n20953 , n8436 );
not ( n20954 , n11091 );
not ( n20955 , n20954 );
not ( n20956 , n8766 );
or ( n20957 , n20955 , n20956 );
nand ( n20958 , n11091 , n8925 );
nand ( n20959 , n20957 , n20958 );
and ( n20960 , n20953 , n20959 );
not ( n20961 , n20953 );
not ( n20962 , n20959 );
and ( n20963 , n20961 , n20962 );
nor ( n20964 , n20960 , n20963 );
nor ( n20965 , n20952 , n20964 );
not ( n20966 , n20952 );
not ( n20967 , n20964 );
or ( n20968 , n20966 , n20967 );
nand ( n20969 , n20968 , n2352 );
or ( n20970 , n20965 , n20969 );
and ( n20971 , n370 , n20944 );
not ( n20972 , n370 );
and ( n20973 , n20972 , n369 );
nor ( n20974 , n20971 , n20973 );
or ( n20975 , n2352 , n20974 );
nand ( n20976 , n20970 , n20975 );
not ( n20977 , n380 );
nand ( n20978 , n20977 , n2986 );
not ( n20979 , n20978 );
not ( n20980 , n380 );
nor ( n20981 , n20980 , n18125 );
nor ( n20982 , n20979 , n20981 );
not ( n20983 , n20982 );
not ( n20984 , n16864 );
not ( n20985 , n20984 );
not ( n20986 , n20985 );
not ( n20987 , n16411 );
or ( n20988 , n20986 , n20987 );
not ( n20989 , n20984 );
or ( n20990 , n20989 , n16411 );
nand ( n20991 , n20988 , n20990 );
not ( n20992 , n20991 );
or ( n20993 , n20983 , n20992 );
or ( n20994 , n20982 , n20991 );
nand ( n20995 , n20993 , n20994 );
and ( n20996 , n16738 , n16996 );
not ( n20997 , n16738 );
and ( n20998 , n20997 , n16999 );
nor ( n20999 , n20996 , n20998 );
nor ( n21000 , n20995 , n20999 );
not ( n21001 , n20995 );
not ( n21002 , n20999 );
or ( n21003 , n21001 , n21002 );
nand ( n21004 , n21003 , n2352 );
or ( n21005 , n21000 , n21004 );
xnor ( n21006 , n380 , n381 );
or ( n21007 , n2352 , n21006 );
nand ( n21008 , n21005 , n21007 );
xnor ( n21009 , n63 , n64 );
or ( n21010 , n2352 , n21009 );
not ( n21011 , n13311 );
or ( n21012 , n13228 , n13235 );
nand ( n21013 , n21012 , n793 );
nand ( n21014 , n21013 , n13280 , n13239 , n13276 );
or ( n21015 , n21014 , n13274 );
nand ( n21016 , n21015 , n841 );
nand ( n21017 , n21011 , n13349 , n21016 );
not ( n21018 , n21017 );
not ( n21019 , n21018 );
not ( n21020 , n2336 );
and ( n21021 , n63 , n21020 );
not ( n21022 , n63 );
and ( n21023 , n21022 , n2336 );
nor ( n21024 , n21021 , n21023 );
not ( n21025 , n21024 );
and ( n21026 , n21019 , n21025 );
not ( n21027 , n21017 );
and ( n21028 , n21027 , n21024 );
nor ( n21029 , n21026 , n21028 );
not ( n21030 , n21029 );
not ( n21031 , n1758 );
not ( n21032 , n6308 );
or ( n21033 , n21031 , n21032 );
nand ( n21034 , n1757 , n6480 );
nand ( n21035 , n21033 , n21034 );
and ( n21036 , n21035 , n13617 );
not ( n21037 , n21035 );
and ( n21038 , n21037 , n13616 );
or ( n21039 , n21036 , n21038 );
not ( n21040 , n21039 );
nand ( n21041 , n21030 , n21040 );
nand ( n21042 , n21029 , n21039 );
nand ( n21043 , n21041 , n2352 , n21042 );
nand ( n21044 , n21010 , n21043 );
not ( n21045 , n18 );
and ( n21046 , n35 , n21045 );
not ( n21047 , n35 );
and ( n21048 , n21047 , n18 );
nor ( n21049 , n21046 , n21048 );
and ( n21050 , n1 , n21049 );
not ( n21051 , n1 );
and ( n21052 , n18391 , n21045 );
not ( n21053 , n18391 );
and ( n21054 , n21053 , n18 );
nor ( n21055 , n21052 , n21054 );
not ( n21056 , n3 );
or ( n21057 , n21056 , n1237 );
nor ( n21058 , n1150 , n996 );
nand ( n21059 , n21057 , n21058 );
nand ( n21060 , n1425 , n21059 );
nand ( n21061 , n7 , n1253 );
nand ( n21062 , n1159 , n1290 );
and ( n21063 , n21061 , n21062 , n13664 );
not ( n21064 , n2318 );
nand ( n21065 , n8 , n21064 );
nand ( n21066 , n21060 , n21063 , n1165 , n21065 );
not ( n21067 , n21066 );
not ( n21068 , n13793 );
nand ( n21069 , n21068 , n7 );
and ( n21070 , n21069 , n1066 , n1040 );
not ( n21071 , n7 );
nand ( n21072 , n2283 , n1409 , n1126 );
nand ( n21073 , n21071 , n21072 );
nand ( n21074 , n21070 , n1144 , n21073 );
nand ( n21075 , n992 , n21074 );
not ( n21076 , n1182 );
nand ( n21077 , n21076 , n13203 , n13820 , n1179 );
and ( n21078 , n7 , n21077 );
not ( n21079 , n7 );
nand ( n21080 , n13199 , n1442 );
and ( n21081 , n21079 , n21080 );
nor ( n21082 , n21078 , n21081 );
nand ( n21083 , n4 , n1172 );
not ( n21084 , n21083 );
nand ( n21085 , n21084 , n1164 );
nand ( n21086 , n3 , n2 , n4 );
not ( n21087 , n21086 );
not ( n21088 , n1057 );
or ( n21089 , n21087 , n21088 );
nand ( n21090 , n21089 , n7 );
nand ( n21091 , n21085 , n21090 );
not ( n21092 , n7 );
nand ( n21093 , n21092 , n1271 );
nand ( n21094 , n21093 , n1126 , n2215 );
or ( n21095 , n21091 , n21094 );
nand ( n21096 , n21095 , n992 );
nand ( n21097 , n1359 , n13173 );
not ( n21098 , n7 );
not ( n21099 , n13135 );
not ( n21100 , n1191 );
nand ( n21101 , n21099 , n1177 , n21100 );
not ( n21102 , n21101 );
or ( n21103 , n21098 , n21102 );
or ( n21104 , n1136 , n6 );
nand ( n21105 , n21104 , n2217 );
nand ( n21106 , n1229 , n21105 );
nand ( n21107 , n21103 , n21106 );
or ( n21108 , n21097 , n21107 );
nand ( n21109 , n21108 , n8 );
nand ( n21110 , n21082 , n21096 , n21109 );
and ( n21111 , n9 , n21110 );
not ( n21112 , n9 );
not ( n21113 , n8 );
not ( n21114 , n7 );
nand ( n21115 , n21114 , n1351 );
not ( n21116 , n1122 );
not ( n21117 , n3 );
nand ( n21118 , n21117 , n1174 );
not ( n21119 , n21118 );
or ( n21120 , n21116 , n21119 );
nand ( n21121 , n21120 , n7 );
nand ( n21122 , n1375 , n21115 , n21121 );
not ( n21123 , n21122 );
or ( n21124 , n21113 , n21123 );
not ( n21125 , n4 );
not ( n21126 , n13103 );
or ( n21127 , n21125 , n21126 );
nand ( n21128 , n21127 , n1105 );
or ( n21129 , n3 , n1234 );
nand ( n21130 , n1050 , n13762 );
nand ( n21131 , n21129 , n21130 );
or ( n21132 , n21128 , n21131 );
not ( n21133 , n7 );
nand ( n21134 , n21132 , n21133 );
nand ( n21135 , n21124 , n21134 );
not ( n21136 , n21135 );
not ( n21137 , n13688 );
not ( n21138 , n13211 );
or ( n21139 , n21137 , n21138 );
nand ( n21140 , n21139 , n7 );
nand ( n21141 , n13199 , n13211 );
not ( n21142 , n7 );
not ( n21143 , n21086 );
and ( n21144 , n21142 , n21143 );
not ( n21145 , n3 );
and ( n21146 , n21145 , n13640 );
nor ( n21147 , n21144 , n21146 );
nand ( n21148 , n21147 , n1298 , n13758 );
or ( n21149 , n21141 , n21148 );
nand ( n21150 , n21149 , n992 );
nand ( n21151 , n21136 , n21140 , n21150 );
and ( n21152 , n21112 , n21151 );
nor ( n21153 , n21111 , n21152 );
nand ( n21154 , n21067 , n21075 , n21153 );
and ( n21155 , n21055 , n21154 );
not ( n21156 , n21055 );
not ( n21157 , n21066 );
and ( n21158 , n21157 , n21075 , n21153 );
not ( n21159 , n21158 );
not ( n21160 , n21159 );
and ( n21161 , n21156 , n21160 );
nor ( n21162 , n21155 , n21161 );
or ( n21163 , n1169 , n1324 );
not ( n21164 , n1183 );
nand ( n21165 , n2324 , n1060 );
not ( n21166 , n21165 );
or ( n21167 , n21164 , n21166 );
nand ( n21168 , n21167 , n7 );
nand ( n21169 , n21163 , n997 , n21168 );
and ( n21170 , n992 , n21169 );
not ( n21171 , n1358 );
or ( n21172 , n3 , n21171 );
nand ( n21173 , n21172 , n1293 , n1375 );
and ( n21174 , n1244 , n21173 );
nor ( n21175 , n21170 , n21174 );
not ( n21176 , n3 );
or ( n21177 , n21176 , n1173 );
nand ( n21178 , n21177 , n13701 );
not ( n21179 , n3 );
nor ( n21180 , n21179 , n13150 );
or ( n21181 , n21178 , n21180 , n13665 );
nand ( n21182 , n21181 , n7 );
not ( n21183 , n7 );
nand ( n21184 , n21183 , n1216 );
and ( n21185 , n13203 , n21085 , n21184 , n21093 );
or ( n21186 , n3 , n1042 );
or ( n21187 , n1169 , n13155 );
nand ( n21188 , n21186 , n21187 );
nand ( n21189 , n1201 , n21062 );
or ( n21190 , n21188 , n21189 );
nand ( n21191 , n21190 , n992 );
not ( n21192 , n21180 );
nand ( n21193 , n21192 , n1025 , n1291 , n1278 );
not ( n21194 , n7 );
not ( n21195 , n3 );
nand ( n21196 , n21195 , n1230 );
nand ( n21197 , n21196 , n1064 , n1442 );
nand ( n21198 , n21194 , n21197 );
not ( n21199 , n13828 );
not ( n21200 , n1373 );
or ( n21201 , n21199 , n21200 );
nand ( n21202 , n21201 , n7 );
nand ( n21203 , n21198 , n1237 , n21202 );
or ( n21204 , n21193 , n21203 );
nand ( n21205 , n21204 , n8 );
nand ( n21206 , n21182 , n21185 , n21191 , n21205 );
nand ( n21207 , n1133 , n21206 );
not ( n21208 , n7 );
and ( n21209 , n21208 , n13113 );
not ( n21210 , n13175 );
nor ( n21211 , n21209 , n21210 , n21064 );
not ( n21212 , n3 );
or ( n21213 , n21212 , n13203 );
nand ( n21214 , n21213 , n21184 );
and ( n21215 , n8 , n21214 );
not ( n21216 , n1205 );
and ( n21217 , n1425 , n21216 );
nor ( n21218 , n21215 , n21217 );
and ( n21219 , n21211 , n21218 );
nand ( n21220 , n7 , n1182 );
and ( n21221 , n21220 , n1052 , n1265 );
not ( n21222 , n2252 );
not ( n21223 , n7 );
not ( n21224 , n2269 );
nand ( n21225 , n21224 , n21083 , n13155 );
nand ( n21226 , n8 , n21225 );
nand ( n21227 , n21226 , n1001 , n13149 );
nand ( n21228 , n21223 , n21227 );
nand ( n21229 , n21221 , n21222 , n21228 );
not ( n21230 , n21229 );
and ( n21231 , n13173 , n1262 );
nand ( n21232 , n21231 , n13641 , n1086 );
nand ( n21233 , n8 , n21232 );
and ( n21234 , n1343 , n1183 );
not ( n21235 , n7 );
and ( n21236 , n21235 , n1194 );
not ( n21237 , n21235 );
not ( n21238 , n3 );
not ( n21239 , n1152 );
or ( n21240 , n21238 , n21239 );
not ( n21241 , n1448 );
nand ( n21242 , n21240 , n21241 );
and ( n21243 , n21237 , n21242 );
nor ( n21244 , n21236 , n21243 );
nand ( n21245 , n21234 , n1465 , n21244 );
nand ( n21246 , n992 , n21245 );
nand ( n21247 , n21230 , n21233 , n21246 );
nand ( n21248 , n9 , n21247 );
nand ( n21249 , n21175 , n21207 , n21219 , n21248 );
not ( n21250 , n21249 );
not ( n21251 , n21250 );
not ( n21252 , n21251 );
not ( n21253 , n18498 );
not ( n21254 , n31 );
or ( n21255 , n21254 , n14582 );
nor ( n21256 , n32 , n6002 );
not ( n21257 , n21256 );
nand ( n21258 , n21255 , n21257 );
and ( n21259 , n33 , n21258 );
not ( n21260 , n6136 );
and ( n21261 , n1739 , n21260 );
nor ( n21262 , n21259 , n21261 );
not ( n21263 , n1678 );
not ( n21264 , n21263 );
not ( n21265 , n33 );
not ( n21266 , n2157 );
nand ( n21267 , n21266 , n1515 );
not ( n21268 , n6101 );
nand ( n21269 , n1503 , n6013 );
not ( n21270 , n21269 );
or ( n21271 , n21268 , n21270 );
nand ( n21272 , n21271 , n32 );
nand ( n21273 , n21267 , n14485 , n21272 );
nand ( n21274 , n21265 , n21273 );
and ( n21275 , n21262 , n21264 , n21274 );
not ( n21276 , n14539 );
or ( n21277 , n32 , n21276 );
or ( n21278 , n31 , n2166 );
not ( n21279 , n13506 );
nand ( n21280 , n21279 , n1515 );
nand ( n21281 , n21278 , n21280 );
and ( n21282 , n2074 , n2033 );
nor ( n21283 , n33 , n21281 , n6128 , n21282 );
not ( n21284 , n33 );
and ( n21285 , n6064 , n2192 );
nand ( n21286 , n21285 , n1669 , n2198 );
not ( n21287 , n32 );
not ( n21288 , n31 );
nand ( n21289 , n21288 , n1716 );
nand ( n21290 , n21289 , n14525 , n2146 );
nand ( n21291 , n21287 , n21290 );
not ( n21292 , n31 );
or ( n21293 , n21292 , n14497 );
not ( n21294 , n13966 );
not ( n21295 , n2142 );
or ( n21296 , n21294 , n21295 );
nand ( n21297 , n21296 , n32 );
nand ( n21298 , n21291 , n21293 , n21297 );
nor ( n21299 , n21284 , n21286 , n21298 );
or ( n21300 , n21283 , n21299 );
not ( n21301 , n32 );
nand ( n21302 , n21301 , n6087 );
not ( n21303 , n21302 );
nor ( n21304 , n21256 , n21303 );
nand ( n21305 , n21300 , n21304 , n14582 );
nand ( n21306 , n2155 , n27 , n1704 );
nand ( n21307 , n31 , n1705 );
not ( n21308 , n13548 );
nand ( n21309 , n13524 , n21307 , n21293 , n21308 );
nand ( n21310 , n32 , n21309 );
nand ( n21311 , n21306 , n21310 );
or ( n21312 , n21305 , n21311 );
nand ( n21313 , n21312 , n1673 );
not ( n21314 , n34 );
not ( n21315 , n32 );
not ( n21316 , n21315 );
not ( n21317 , n1573 );
nand ( n21318 , n21317 , n14026 , n1717 );
not ( n21319 , n21318 );
or ( n21320 , n21316 , n21319 );
nand ( n21321 , n21320 , n1586 );
nand ( n21322 , n32 , n6100 );
not ( n21323 , n1494 );
nand ( n21324 , n21322 , n21323 , n6055 );
nor ( n21325 , n21321 , n21324 );
not ( n21326 , n13596 );
not ( n21327 , n6022 );
nor ( n21328 , n21326 , n21327 );
nand ( n21329 , n21328 , n13580 , n6052 );
nand ( n21330 , n33 , n21329 );
nand ( n21331 , n14026 , n6101 );
not ( n21332 , n33 );
nand ( n21333 , n2129 , n13497 );
nand ( n21334 , n32 , n21333 );
not ( n21335 , n32 );
nand ( n21336 , n21335 , n6123 );
nand ( n21337 , n21332 , n21334 , n2105 , n21336 );
or ( n21338 , n21331 , n21337 );
not ( n21339 , n32 );
not ( n21340 , n21339 );
nand ( n21341 , n30 , n6072 );
nand ( n21342 , n27 , n1704 );
nand ( n21343 , n21341 , n21342 , n13506 );
not ( n21344 , n21343 );
or ( n21345 , n21340 , n21344 );
nand ( n21346 , n21345 , n33 );
nand ( n21347 , n21338 , n21346 );
nand ( n21348 , n21325 , n21330 , n21347 );
not ( n21349 , n21348 );
or ( n21350 , n21314 , n21349 );
not ( n21351 , n2055 );
or ( n21352 , n31 , n21351 );
nand ( n21353 , n21352 , n1584 , n1630 );
and ( n21354 , n6091 , n21353 );
not ( n21355 , n13534 );
nor ( n21356 , n21354 , n21355 );
nand ( n21357 , n21350 , n21356 );
not ( n21358 , n21357 );
nand ( n21359 , n21275 , n21277 , n21313 , n21358 );
not ( n21360 , n21359 );
not ( n21361 , n21360 );
and ( n21362 , n21253 , n21361 );
not ( n21363 , n18499 );
nand ( n21364 , n21275 , n21277 , n21313 , n21358 );
not ( n21365 , n21364 );
and ( n21366 , n21363 , n21365 );
nor ( n21367 , n21362 , n21366 );
not ( n21368 , n21367 );
or ( n21369 , n21252 , n21368 );
or ( n21370 , n21251 , n21367 );
nand ( n21371 , n21369 , n21370 );
nor ( n21372 , n21162 , n21371 );
and ( n21373 , n21051 , n21372 );
nor ( n21374 , n21050 , n21373 );
not ( n21375 , n37 );
and ( n21376 , n18391 , n21375 );
not ( n21377 , n18391 );
and ( n21378 , n21377 , n37 );
nor ( n21379 , n21376 , n21378 );
not ( n21380 , n10 );
nand ( n21381 , n15 , n929 );
and ( n21382 , n21381 , n18363 , n13246 );
nor ( n21383 , n21382 , n5854 );
not ( n21384 , n21383 );
and ( n21385 , n16 , n894 );
nor ( n21386 , n21385 , n5777 );
nand ( n21387 , n14274 , n830 );
nand ( n21388 , n926 , n13279 );
or ( n21389 , n21387 , n21388 );
nand ( n21390 , n21389 , n17 );
nand ( n21391 , n21384 , n21386 , n21390 );
not ( n21392 , n21391 );
and ( n21393 , n930 , n836 );
or ( n21394 , n947 , n13243 );
not ( n21395 , n16 );
nand ( n21396 , n21394 , n21395 );
nand ( n21397 , n13329 , n5848 , n5738 );
not ( n21398 , n21397 );
not ( n21399 , n5948 );
not ( n21400 , n14131 );
or ( n21401 , n21399 , n21400 );
nand ( n21402 , n21401 , n16 );
not ( n21403 , n16 );
not ( n21404 , n844 );
nand ( n21405 , n21403 , n21404 );
nand ( n21406 , n21398 , n21402 , n21405 );
nand ( n21407 , n21406 , n793 );
nand ( n21408 , n21392 , n21393 , n21396 , n21407 );
not ( n21409 , n21408 );
or ( n21410 , n21380 , n21409 );
not ( n21411 , n16 );
not ( n21412 , n21411 );
not ( n21413 , n13 );
nand ( n21414 , n21413 , n5896 );
nand ( n21415 , n21414 , n5720 , n5803 );
not ( n21416 , n21415 );
or ( n21417 , n21412 , n21416 );
or ( n21418 , n911 , n5823 );
nand ( n21419 , n21418 , n13329 );
nand ( n21420 , n16 , n21419 );
nand ( n21421 , n21417 , n21420 );
or ( n21422 , n809 , n5858 );
nand ( n21423 , n21422 , n941 );
or ( n21424 , n21421 , n21423 );
nand ( n21425 , n21424 , n793 );
nand ( n21426 , n21410 , n21425 );
not ( n21427 , n21426 );
not ( n21428 , n13 );
or ( n21429 , n21428 , n13316 );
not ( n21430 , n16 );
nand ( n21431 , n21430 , n778 );
nand ( n21432 , n21429 , n21431 );
and ( n21433 , n17 , n21432 );
nor ( n21434 , n21433 , n5719 );
not ( n21435 , n863 );
nand ( n21436 , n21435 , n5839 );
and ( n21437 , n21434 , n21436 , n942 , n13280 );
not ( n21438 , n16 );
and ( n21439 , n13 , n855 );
nor ( n21440 , n21439 , n940 );
nand ( n21441 , n13 , n969 );
not ( n21442 , n14337 );
nand ( n21443 , n21440 , n21441 , n21442 );
not ( n21444 , n21443 );
or ( n21445 , n21438 , n21444 );
not ( n21446 , n13246 );
nand ( n21447 , n21446 , n810 );
not ( n21448 , n13 );
not ( n21449 , n5844 );
nand ( n21450 , n21448 , n21449 );
nand ( n21451 , n21447 , n21450 , n850 , n18300 );
and ( n21452 , n793 , n21451 );
not ( n21453 , n793 );
not ( n21454 , n5887 );
nand ( n21455 , n5814 , n760 );
not ( n21456 , n21455 );
or ( n21457 , n21454 , n21456 );
or ( n21458 , n5887 , n21455 );
nand ( n21459 , n21457 , n21458 );
not ( n21460 , n21459 );
not ( n21461 , n21441 );
not ( n21462 , n5865 );
nor ( n21463 , n21461 , n21462 );
not ( n21464 , n13 );
nand ( n21465 , n21464 , n753 );
nand ( n21466 , n915 , n5956 );
nor ( n21467 , n21465 , n21466 );
not ( n21468 , n21467 );
nand ( n21469 , n21465 , n21466 );
not ( n21470 , n16 );
nand ( n21471 , n21468 , n21469 , n21470 );
not ( n21472 , n14139 );
not ( n21473 , n21472 );
not ( n21474 , n5954 );
or ( n21475 , n21473 , n21474 );
nand ( n21476 , n21475 , n16 );
nand ( n21477 , n21460 , n21463 , n21471 , n21476 );
and ( n21478 , n21453 , n21477 );
nor ( n21479 , n21452 , n21478 );
nand ( n21480 , n21445 , n21479 );
nand ( n21481 , n13316 , n18365 , n21431 , n18372 );
or ( n21482 , n21480 , n21481 );
nand ( n21483 , n21482 , n841 );
nand ( n21484 , n21427 , n21437 , n21483 );
not ( n21485 , n21484 );
buf ( n21486 , n21485 );
not ( n21487 , n21486 );
and ( n21488 , n21379 , n21487 );
not ( n21489 , n21379 );
and ( n21490 , n21489 , n21486 );
nor ( n21491 , n21488 , n21490 );
not ( n21492 , n21249 );
not ( n21493 , n33 );
and ( n21494 , n32 , n13984 );
not ( n21495 , n6043 );
nor ( n21496 , n21494 , n1636 , n21495 );
not ( n21497 , n32 );
nand ( n21498 , n1712 , n1687 , n1534 );
nand ( n21499 , n21497 , n21498 );
nand ( n21500 , n21496 , n6109 , n21499 );
and ( n21501 , n21493 , n21500 );
not ( n21502 , n32 );
or ( n21503 , n21502 , n6083 );
not ( n21504 , n21282 );
and ( n21505 , n21503 , n21504 , n13545 );
not ( n21506 , n31 );
or ( n21507 , n21506 , n6064 );
not ( n21508 , n14484 );
nand ( n21509 , n21507 , n2042 , n21508 );
nand ( n21510 , n1739 , n21509 );
nand ( n21511 , n21505 , n6119 , n21510 );
nor ( n21512 , n21501 , n21511 );
nand ( n21513 , n33 , n21263 );
not ( n21514 , n33 );
not ( n21515 , n2056 );
nor ( n21516 , n21515 , n13579 );
not ( n21517 , n27 );
nor ( n21518 , n21517 , n30 );
or ( n21519 , n21518 , n1611 );
nand ( n21520 , n21519 , n1608 );
nand ( n21521 , n2088 , n6064 , n14472 );
nand ( n21522 , n32 , n21521 );
nand ( n21523 , n21516 , n21520 , n21522 );
not ( n21524 , n21523 );
or ( n21525 , n21514 , n21524 );
not ( n21526 , n2146 );
not ( n21527 , n1493 );
or ( n21528 , n21526 , n21527 );
not ( n21529 , n32 );
nand ( n21530 , n21528 , n21529 );
nand ( n21531 , n21525 , n21530 );
not ( n21532 , n32 );
nand ( n21533 , n14582 , n6124 , n6097 , n6099 );
not ( n21534 , n21533 );
or ( n21535 , n21532 , n21534 );
nand ( n21536 , n21306 , n21302 );
nand ( n21537 , n29 , n1629 );
not ( n21538 , n21537 );
not ( n21539 , n1532 );
or ( n21540 , n21538 , n21539 );
nand ( n21541 , n21540 , n32 );
nand ( n21542 , n21541 , n1609 , n1687 );
or ( n21543 , n21536 , n21542 );
not ( n21544 , n33 );
nand ( n21545 , n21543 , n21544 );
nand ( n21546 , n21535 , n21545 );
nor ( n21547 , n21531 , n21546 );
and ( n21548 , n34 , n21547 );
not ( n21549 , n34 );
not ( n21550 , n33 );
not ( n21551 , n31 );
not ( n21552 , n21551 );
not ( n21553 , n1705 );
or ( n21554 , n21552 , n21553 );
nand ( n21555 , n21554 , n1617 );
nand ( n21556 , n32 , n21555 );
not ( n21557 , n32 );
nand ( n21558 , n21557 , n2039 );
nand ( n21559 , n21556 , n1630 , n21558 );
not ( n21560 , n21559 );
or ( n21561 , n21550 , n21560 );
not ( n21562 , n13508 );
not ( n21563 , n2060 );
or ( n21564 , n21562 , n21563 );
nand ( n21565 , n21564 , n32 );
nand ( n21566 , n21561 , n21565 );
not ( n21567 , n21566 );
not ( n21568 , n27 );
or ( n21569 , n21568 , n1553 );
nand ( n21570 , n21569 , n6076 );
not ( n21571 , n6072 );
not ( n21572 , n14045 );
or ( n21573 , n21571 , n21572 );
or ( n21574 , n31 , n1507 );
nand ( n21575 , n21573 , n21574 );
or ( n21576 , n21570 , n21575 );
not ( n21577 , n32 );
nand ( n21578 , n21576 , n21577 );
nor ( n21579 , n2181 , n14036 );
nand ( n21580 , n21579 , n1493 , n2060 );
not ( n21581 , n1589 );
or ( n21582 , n31 , n21581 );
or ( n21583 , n32 , n21537 );
nand ( n21584 , n21582 , n21583 );
or ( n21585 , n21580 , n21584 );
not ( n21586 , n33 );
nand ( n21587 , n21585 , n21586 );
nand ( n21588 , n21567 , n21578 , n21587 );
not ( n21589 , n21588 );
and ( n21590 , n21549 , n21589 );
or ( n21591 , n21548 , n21590 );
and ( n21592 , n21512 , n21513 , n21591 );
and ( n21593 , n21592 , n18497 );
not ( n21594 , n21592 );
and ( n21595 , n21594 , n18498 );
nor ( n21596 , n21593 , n21595 );
and ( n21597 , n21492 , n21596 );
not ( n21598 , n21492 );
not ( n21599 , n21596 );
and ( n21600 , n21598 , n21599 );
nor ( n21601 , n21597 , n21600 );
nor ( n21602 , n21491 , n21601 );
not ( n21603 , n21491 );
not ( n21604 , n21601 );
or ( n21605 , n21603 , n21604 );
nand ( n21606 , n21605 , n2352 );
or ( n21607 , n21602 , n21606 );
and ( n21608 , n36 , n21375 );
not ( n21609 , n36 );
and ( n21610 , n21609 , n37 );
nor ( n21611 , n21608 , n21610 );
or ( n21612 , n2352 , n21611 );
nand ( n21613 , n21607 , n21612 );
not ( n21614 , n38 );
not ( n21615 , n39 );
and ( n21616 , n21614 , n21615 );
and ( n21617 , n38 , n39 );
nor ( n21618 , n21616 , n21617 );
or ( n21619 , n2352 , n21618 );
not ( n21620 , n21359 );
not ( n21621 , n21620 );
not ( n21622 , n26 );
and ( n21623 , n13424 , n1998 );
nand ( n21624 , n21623 , n14389 , n1956 );
not ( n21625 , n21624 );
or ( n21626 , n21622 , n21625 );
nand ( n21627 , n25 , n1845 );
nand ( n21628 , n21626 , n21627 );
not ( n21629 , n6295 );
nand ( n21630 , n21629 , n13419 );
not ( n21631 , n6444 );
not ( n21632 , n25 );
nand ( n21633 , n21632 , n1833 );
not ( n21634 , n6311 );
not ( n21635 , n13901 );
or ( n21636 , n21634 , n21635 );
nand ( n21637 , n21636 , n25 );
nand ( n21638 , n21631 , n21633 , n21637 );
or ( n21639 , n21630 , n21638 );
not ( n21640 , n26 );
nand ( n21641 , n21639 , n21640 );
and ( n21642 , n1962 , n6265 );
nand ( n21643 , n24 , n1960 );
nand ( n21644 , n21643 , n18486 , n13451 );
nand ( n21645 , n13397 , n21644 );
not ( n21646 , n1927 );
not ( n21647 , n13462 );
or ( n21648 , n21646 , n21647 );
not ( n21649 , n25 );
nand ( n21650 , n21648 , n21649 );
and ( n21651 , n2000 , n21645 , n21650 );
nand ( n21652 , n21641 , n21642 , n21651 );
nor ( n21653 , n21628 , n21652 );
or ( n21654 , n1853 , n21653 );
not ( n21655 , n26 );
not ( n21656 , n23 );
and ( n21657 , n21656 , n6369 );
nor ( n21658 , n21657 , n6188 , n6178 );
or ( n21659 , n25 , n21658 );
not ( n21660 , n1799 );
not ( n21661 , n6434 );
and ( n21662 , n21660 , n21661 );
not ( n21663 , n13418 );
nor ( n21664 , n21662 , n21663 );
not ( n21665 , n1997 );
or ( n21666 , n21665 , n1964 );
nand ( n21667 , n21666 , n13419 );
nand ( n21668 , n25 , n21667 );
nand ( n21669 , n21659 , n21664 , n21668 );
nand ( n21670 , n21655 , n21669 );
nand ( n21671 , n21654 , n21670 );
not ( n21672 , n21671 );
not ( n21673 , n1853 );
not ( n21674 , n25 );
nand ( n21675 , n21674 , n1864 );
not ( n21676 , n26 );
not ( n21677 , n1800 );
not ( n21678 , n14407 );
or ( n21679 , n21677 , n21678 );
nand ( n21680 , n21679 , n18412 );
and ( n21681 , n21676 , n21680 );
nand ( n21682 , n23 , n1899 );
nand ( n21683 , n23 , n1804 );
and ( n21684 , n21682 , n21683 );
not ( n21685 , n25 );
nor ( n21686 , n21684 , n21685 );
nor ( n21687 , n21681 , n21686 );
nand ( n21688 , n18485 , n13402 );
not ( n21689 , n1921 );
not ( n21690 , n14453 );
or ( n21691 , n21689 , n21690 );
nand ( n21692 , n21691 , n25 );
nand ( n21693 , n18488 , n21692 );
nor ( n21694 , n21688 , n21693 );
nand ( n21695 , n21675 , n21687 , n21694 );
not ( n21696 , n21695 );
not ( n21697 , n26 );
not ( n21698 , n6333 );
or ( n21699 , n21665 , n21698 );
nand ( n21700 , n21699 , n1839 );
and ( n21701 , n21697 , n21700 );
not ( n21702 , n21697 );
not ( n21703 , n25 );
not ( n21704 , n21703 );
not ( n21705 , n1968 );
not ( n21706 , n23 );
nand ( n21707 , n21706 , n1857 );
nand ( n21708 , n21705 , n21707 , n6320 );
not ( n21709 , n21708 );
or ( n21710 , n21704 , n21709 );
and ( n21711 , n21682 , n1931 );
nand ( n21712 , n21710 , n21711 );
not ( n21713 , n21712 );
not ( n21714 , n13908 );
not ( n21715 , n6317 );
or ( n21716 , n21714 , n21715 );
nand ( n21717 , n21716 , n25 );
and ( n21718 , n6465 , n6453 );
nand ( n21719 , n21713 , n21717 , n1861 , n21718 );
and ( n21720 , n21702 , n21719 );
nor ( n21721 , n21701 , n21720 );
nand ( n21722 , n21696 , n21721 );
not ( n21723 , n21722 );
or ( n21724 , n21673 , n21723 );
not ( n21725 , n26 );
not ( n21726 , n23 );
not ( n21727 , n21726 );
not ( n21728 , n13402 );
and ( n21729 , n21727 , n21728 );
not ( n21730 , n6317 );
and ( n21731 , n1794 , n21730 );
nor ( n21732 , n21729 , n21731 );
or ( n21733 , n21725 , n21732 );
nand ( n21734 , n21733 , n6193 );
or ( n21735 , n25 , n6253 );
not ( n21736 , n26 );
or ( n21737 , n21736 , n21675 );
nand ( n21738 , n21735 , n21737 , n13433 );
nor ( n21739 , n21734 , n21738 );
nand ( n21740 , n21724 , n21739 );
not ( n21741 , n21740 );
nand ( n21742 , n21672 , n21741 );
not ( n21743 , n21742 );
and ( n21744 , n21621 , n21743 );
and ( n21745 , n21365 , n21742 );
nor ( n21746 , n21744 , n21745 );
not ( n21747 , n21746 );
xor ( n21748 , n39 , n18390 );
not ( n21749 , n21748 );
not ( n21750 , n21592 );
not ( n21751 , n21158 );
or ( n21752 , n21750 , n21751 );
nand ( n21753 , n1673 , n21588 );
or ( n21754 , n21531 , n21546 );
nand ( n21755 , n21754 , n34 );
and ( n21756 , n21512 , n21513 , n21753 , n21755 );
or ( n21757 , n21756 , n21158 );
nand ( n21758 , n21752 , n21757 );
not ( n21759 , n21758 );
or ( n21760 , n21749 , n21759 );
or ( n21761 , n21748 , n21758 );
nand ( n21762 , n21760 , n21761 );
or ( n21763 , n21747 , n21762 );
not ( n21764 , n21620 );
nor ( n21765 , n21671 , n21740 );
not ( n21766 , n21765 );
and ( n21767 , n21764 , n21766 );
and ( n21768 , n21360 , n21765 );
nor ( n21769 , n21767 , n21768 );
buf ( n21770 , n21769 );
nand ( n21771 , n21770 , n21762 );
nand ( n21772 , n21763 , n21771 , n2352 );
nand ( n21773 , n21619 , n21772 );
not ( n21774 , n43 );
not ( n21775 , n5989 );
and ( n21776 , n21774 , n21775 );
and ( n21777 , n43 , n5989 );
nor ( n21778 , n21776 , n21777 );
not ( n21779 , n9104 );
and ( n21780 , n21778 , n21779 );
not ( n21781 , n21778 );
not ( n21782 , n21779 );
and ( n21783 , n21781 , n21782 );
nor ( n21784 , n21780 , n21783 );
not ( n21785 , n21784 );
not ( n21786 , n21756 );
not ( n21787 , n14610 );
and ( n21788 , n21786 , n21787 );
and ( n21789 , n21756 , n14610 );
nor ( n21790 , n21788 , n21789 );
and ( n21791 , n21790 , n21160 );
not ( n21792 , n21790 );
and ( n21793 , n21792 , n21154 );
nor ( n21794 , n21791 , n21793 );
not ( n21795 , n21794 );
nor ( n21796 , n21785 , n21795 );
or ( n21797 , n21784 , n21794 );
nand ( n21798 , n21797 , n2352 );
or ( n21799 , n21796 , n21798 );
xnor ( n21800 , n43 , n44 );
or ( n21801 , n2352 , n21800 );
nand ( n21802 , n21799 , n21801 );
xor ( n21803 , n45 , n5989 );
xor ( n21804 , n21803 , n18392 );
not ( n21805 , n21158 );
not ( n21806 , n18271 );
not ( n21807 , n21806 );
and ( n21808 , n21805 , n21807 );
and ( n21809 , n21160 , n18272 );
nor ( n21810 , n21808 , n21809 );
nor ( n21811 , n21804 , n21810 );
not ( n21812 , n21804 );
not ( n21813 , n21810 );
or ( n21814 , n21812 , n21813 );
nand ( n21815 , n21814 , n2352 );
or ( n21816 , n21811 , n21815 );
xnor ( n21817 , n45 , n46 );
or ( n21818 , n2352 , n21817 );
nand ( n21819 , n21816 , n21818 );
xor ( n21820 , n40 , n21154 );
xnor ( n21821 , n21820 , n21485 );
buf ( n21822 , n21765 );
and ( n21823 , n21822 , n21596 );
not ( n21824 , n21822 );
and ( n21825 , n21824 , n21599 );
nor ( n21826 , n21823 , n21825 );
nor ( n21827 , n21821 , n21826 );
not ( n21828 , n21821 );
not ( n21829 , n21826 );
or ( n21830 , n21828 , n21829 );
nand ( n21831 , n21830 , n2352 );
or ( n21832 , n21827 , n21831 );
xnor ( n21833 , n40 , n47 );
or ( n21834 , n2352 , n21833 );
nand ( n21835 , n21832 , n21834 );
not ( n21836 , n21426 );
nand ( n21837 , n21836 , n21437 , n21483 );
and ( n21838 , n21837 , n51 );
not ( n21839 , n21837 );
not ( n21840 , n51 );
and ( n21841 , n21839 , n21840 );
nor ( n21842 , n21838 , n21841 );
and ( n21843 , n21842 , n21492 );
not ( n21844 , n21842 );
and ( n21845 , n21844 , n21251 );
or ( n21846 , n21843 , n21845 );
xnor ( n21847 , n21822 , n14222 );
nor ( n21848 , n21846 , n21847 );
not ( n21849 , n21846 );
not ( n21850 , n21847 );
or ( n21851 , n21849 , n21850 );
nand ( n21852 , n21851 , n2352 );
or ( n21853 , n21848 , n21852 );
and ( n21854 , n52 , n21840 );
not ( n21855 , n52 );
and ( n21856 , n21855 , n51 );
nor ( n21857 , n21854 , n21856 );
or ( n21858 , n2352 , n21857 );
nand ( n21859 , n21853 , n21858 );
xnor ( n21860 , n55 , n56 );
or ( n21861 , n2352 , n21860 );
not ( n21862 , n2209 );
not ( n21863 , n1472 );
and ( n21864 , n21862 , n21863 );
and ( n21865 , n2209 , n1472 );
nor ( n21866 , n21864 , n21865 );
not ( n21867 , n55 );
not ( n21868 , n5989 );
and ( n21869 , n21867 , n21868 );
and ( n21870 , n55 , n5989 );
nor ( n21871 , n21869 , n21870 );
not ( n21872 , n21871 );
and ( n21873 , n21866 , n21872 );
not ( n21874 , n21866 );
and ( n21875 , n21874 , n21871 );
nor ( n21876 , n21873 , n21875 );
not ( n21877 , n21876 );
nand ( n21878 , n21599 , n21877 );
nand ( n21879 , n21596 , n21876 );
nand ( n21880 , n21878 , n2352 , n21879 );
nand ( n21881 , n21861 , n21880 );
not ( n21882 , n58 );
and ( n21883 , n9084 , n21882 );
not ( n21884 , n9084 );
and ( n21885 , n21884 , n58 );
nor ( n21886 , n21883 , n21885 );
not ( n21887 , n21020 );
not ( n21888 , n1758 );
or ( n21889 , n21887 , n21888 );
or ( n21890 , n2337 , n1758 );
nand ( n21891 , n21889 , n21890 );
not ( n21892 , n21891 );
and ( n21893 , n21886 , n21892 );
not ( n21894 , n21886 );
and ( n21895 , n21894 , n21891 );
nor ( n21896 , n21893 , n21895 );
not ( n21897 , n21896 );
nor ( n21898 , n14596 , n21897 );
or ( n21899 , n14605 , n21896 );
nand ( n21900 , n21899 , n2352 );
or ( n21901 , n21898 , n21900 );
and ( n21902 , n70 , n21882 );
not ( n21903 , n70 );
and ( n21904 , n21903 , n58 );
nor ( n21905 , n21902 , n21904 );
or ( n21906 , n2352 , n21905 );
nand ( n21907 , n21901 , n21906 );
not ( n21908 , n73 );
and ( n21909 , n21908 , n21017 );
not ( n21910 , n21908 );
and ( n21911 , n21910 , n21018 );
nor ( n21912 , n21909 , n21911 );
not ( n21913 , n21912 );
and ( n21914 , n14347 , n14641 );
not ( n21915 , n14347 );
and ( n21916 , n21915 , n5989 );
nor ( n21917 , n21914 , n21916 );
not ( n21918 , n21917 );
and ( n21919 , n21913 , n21918 );
and ( n21920 , n21912 , n21917 );
nor ( n21921 , n21919 , n21920 );
not ( n21922 , n21921 );
not ( n21923 , n14633 );
not ( n21924 , n1472 );
and ( n21925 , n21923 , n21924 );
and ( n21926 , n13718 , n9101 );
nor ( n21927 , n21925 , n21926 );
not ( n21928 , n21927 );
and ( n21929 , n21928 , n14605 );
not ( n21930 , n21928 );
and ( n21931 , n21930 , n14596 );
nor ( n21932 , n21929 , n21931 );
not ( n21933 , n21932 );
nor ( n21934 , n21922 , n21933 );
or ( n21935 , n21921 , n21932 );
nand ( n21936 , n21935 , n2352 );
or ( n21937 , n21934 , n21936 );
and ( n21938 , n74 , n21908 );
not ( n21939 , n74 );
and ( n21940 , n21939 , n73 );
nor ( n21941 , n21938 , n21940 );
or ( n21942 , n2352 , n21941 );
nand ( n21943 , n21937 , n21942 );
and ( n21944 , n14348 , n90 );
not ( n21945 , n14348 );
not ( n21946 , n90 );
and ( n21947 , n21945 , n21946 );
or ( n21948 , n21944 , n21947 );
not ( n21949 , n14467 );
not ( n21950 , n2210 );
and ( n21951 , n21949 , n21950 );
and ( n21952 , n14467 , n2340 );
nor ( n21953 , n21951 , n21952 );
not ( n21954 , n21927 );
and ( n21955 , n21953 , n21954 );
not ( n21956 , n21953 );
and ( n21957 , n21956 , n21927 );
nor ( n21958 , n21955 , n21957 );
nor ( n21959 , n21948 , n21958 );
not ( n21960 , n21948 );
not ( n21961 , n21958 );
or ( n21962 , n21960 , n21961 );
nand ( n21963 , n21962 , n2352 );
or ( n21964 , n21959 , n21963 );
and ( n21965 , n91 , n21946 );
not ( n21966 , n91 );
and ( n21967 , n21966 , n90 );
nor ( n21968 , n21965 , n21967 );
or ( n21969 , n2352 , n21968 );
nand ( n21970 , n21964 , n21969 );
not ( n21971 , n110 );
and ( n21972 , n219 , n21971 );
not ( n21973 , n219 );
and ( n21974 , n21973 , n110 );
nor ( n21975 , n21972 , n21974 );
or ( n21976 , n2352 , n21975 );
not ( n21977 , n21971 );
not ( n21978 , n19211 );
not ( n21979 , n21978 );
and ( n21980 , n21977 , n21979 );
and ( n21981 , n21971 , n19212 );
nor ( n21982 , n21980 , n21981 );
and ( n21983 , n10339 , n4488 , n10539 );
or ( n21984 , n149 , n21983 );
not ( n21985 , n149 );
or ( n21986 , n21985 , n4515 );
and ( n21987 , n21986 , n10372 , n10437 );
not ( n21988 , n10445 );
nand ( n21989 , n21984 , n21987 , n21988 );
and ( n21990 , n4532 , n21989 );
not ( n21991 , n149 );
not ( n21992 , n21991 );
not ( n21993 , n10341 );
and ( n21994 , n21992 , n21993 );
nand ( n21995 , n13036 , n4394 );
nor ( n21996 , n21994 , n21995 );
not ( n21997 , n10470 );
not ( n21998 , n10325 );
nand ( n21999 , n150 , n21998 );
not ( n22000 , n21999 );
and ( n22001 , n4384 , n10426 );
not ( n22002 , n22001 );
or ( n22003 , n22000 , n22002 );
nand ( n22004 , n22003 , n10610 );
nand ( n22005 , n21996 , n21997 , n22004 );
nor ( n22006 , n21990 , n22005 );
not ( n22007 , n12228 );
nand ( n22008 , n152 , n22007 );
nand ( n22009 , n4354 , n12975 , n10485 );
and ( n22010 , n149 , n22009 );
not ( n22011 , n149 );
not ( n22012 , n10554 );
nand ( n22013 , n10603 , n22012 );
and ( n22014 , n22011 , n22013 );
nor ( n22015 , n22010 , n22014 );
not ( n22016 , n10507 );
nor ( n22017 , n22016 , n12963 );
not ( n22018 , n148 );
nor ( n22019 , n22018 , n147 );
or ( n22020 , n22019 , n10319 );
nand ( n22021 , n22020 , n10317 );
nand ( n22022 , n16113 , n4409 , n10323 );
nand ( n22023 , n149 , n22022 );
nand ( n22024 , n22017 , n22021 , n22023 );
and ( n22025 , n152 , n22024 );
not ( n22026 , n152 );
and ( n22027 , n151 , n148 , n150 );
not ( n22028 , n22027 );
nand ( n22029 , n22028 , n4453 );
and ( n22030 , n149 , n22029 );
nor ( n22031 , n22030 , n13065 );
nand ( n22032 , n22031 , n13068 , n4488 , n12288 );
and ( n22033 , n22026 , n22032 );
nor ( n22034 , n22025 , n22033 );
nand ( n22035 , n22015 , n22034 );
and ( n22036 , n153 , n22035 );
not ( n22037 , n153 );
not ( n22038 , n150 );
not ( n22039 , n22038 );
not ( n22040 , n10453 );
not ( n22041 , n22040 );
or ( n22042 , n22039 , n22041 );
nand ( n22043 , n22042 , n10411 );
and ( n22044 , n149 , n22043 );
not ( n22045 , n149 );
and ( n22046 , n22045 , n12974 );
nor ( n22047 , n22044 , n22046 );
nand ( n22048 , n4536 , n22047 );
and ( n22049 , n152 , n22048 );
not ( n22050 , n148 );
not ( n22051 , n4519 );
or ( n22052 , n22050 , n22051 );
nand ( n22053 , n22052 , n4399 );
not ( n22054 , n22053 );
not ( n22055 , n150 );
not ( n22056 , n10320 );
and ( n22057 , n22055 , n22056 );
and ( n22058 , n20499 , n4434 );
nor ( n22059 , n22057 , n22058 );
and ( n22060 , n22054 , n22059 );
nor ( n22061 , n22060 , n149 );
nor ( n22062 , n22049 , n22061 );
not ( n22063 , n20494 );
not ( n22064 , n4525 );
or ( n22065 , n22063 , n22064 );
nand ( n22066 , n22065 , n149 );
nand ( n22067 , n22012 , n4525 );
not ( n22068 , n150 );
and ( n22069 , n22068 , n4369 );
not ( n22070 , n149 );
and ( n22071 , n22070 , n22027 );
nor ( n22072 , n22069 , n22071 );
not ( n22073 , n10570 );
nand ( n22074 , n22072 , n22073 , n4418 );
or ( n22075 , n22067 , n22074 );
nand ( n22076 , n22075 , n4532 );
nand ( n22077 , n22062 , n22066 , n22076 );
and ( n22078 , n22037 , n22077 );
nor ( n22079 , n22036 , n22078 );
and ( n22080 , n22006 , n22008 , n22079 );
not ( n22081 , n22080 );
and ( n22082 , n21982 , n22081 );
not ( n22083 , n21982 );
not ( n22084 , n22081 );
and ( n22085 , n22083 , n22084 );
nor ( n22086 , n22082 , n22085 );
not ( n22087 , n22086 );
not ( n22088 , n19362 );
nand ( n22089 , n22088 , n19365 , n19439 );
not ( n22090 , n12955 );
xor ( n22091 , n22089 , n22090 );
xor ( n22092 , n22091 , n17020 );
not ( n22093 , n22092 );
nand ( n22094 , n22087 , n22093 );
nand ( n22095 , n22086 , n22092 );
nand ( n22096 , n22094 , n2352 , n22095 );
nand ( n22097 , n21976 , n22096 );
and ( n22098 , n19563 , n221 );
not ( n22099 , n19563 );
not ( n22100 , n221 );
and ( n22101 , n22099 , n22100 );
nor ( n22102 , n22098 , n22101 );
not ( n22103 , n19590 );
not ( n22104 , n19575 );
nand ( n22105 , n22103 , n22104 , n19666 );
not ( n22106 , n22105 );
not ( n22107 , n209 );
not ( n22108 , n22107 );
not ( n22109 , n3606 );
and ( n22110 , n22108 , n22109 );
nand ( n22111 , n8690 , n8455 );
nor ( n22112 , n22110 , n22111 );
not ( n22113 , n210 );
or ( n22114 , n22113 , n8703 );
nand ( n22115 , n22114 , n8581 , n3585 );
nand ( n22116 , n3717 , n22115 );
nand ( n22117 , n22112 , n12498 , n22116 );
not ( n22118 , n22117 );
not ( n22119 , n211 );
not ( n22120 , n8660 );
or ( n22121 , n22119 , n22120 );
not ( n22122 , n211 );
nand ( n22123 , n209 , n8595 );
and ( n22124 , n22123 , n3546 , n9328 );
not ( n22125 , n209 );
nand ( n22126 , n3483 , n8569 , n3610 );
nand ( n22127 , n22125 , n22126 );
nand ( n22128 , n22122 , n22124 , n12476 , n22127 );
nand ( n22129 , n22121 , n22128 );
nand ( n22130 , n22118 , n22129 );
not ( n22131 , n22130 );
nand ( n22132 , n9425 , n8522 );
not ( n22133 , n209 );
nand ( n22134 , n206 , n3558 );
not ( n22135 , n22134 );
and ( n22136 , n22133 , n22135 );
not ( n22137 , n210 );
and ( n22138 , n22137 , n8485 );
nor ( n22139 , n22136 , n22138 );
nand ( n22140 , n22139 , n3729 , n3538 );
nor ( n22141 , n22132 , n22140 );
or ( n22142 , n211 , n22141 );
not ( n22143 , n209 );
not ( n22144 , n22143 );
not ( n22145 , n210 );
not ( n22146 , n9448 );
and ( n22147 , n22145 , n22146 );
and ( n22148 , n9271 , n8500 );
nor ( n22149 , n22147 , n22148 );
nand ( n22150 , n208 , n3475 );
nand ( n22151 , n22149 , n8457 , n22150 );
not ( n22152 , n22151 );
or ( n22153 , n22144 , n22152 );
not ( n22154 , n209 );
not ( n22155 , n22154 );
not ( n22156 , n3731 );
or ( n22157 , n22155 , n22156 );
not ( n22158 , n8667 );
not ( n22159 , n210 );
nand ( n22160 , n22158 , n22159 );
nand ( n22161 , n209 , n9428 , n22160 );
nand ( n22162 , n22157 , n22161 );
nand ( n22163 , n8530 , n22162 );
nand ( n22164 , n211 , n22163 );
nand ( n22165 , n22153 , n22164 );
not ( n22166 , n22165 );
not ( n22167 , n9256 );
not ( n22168 , n3538 );
or ( n22169 , n22167 , n22168 );
nand ( n22170 , n22169 , n209 );
nand ( n22171 , n22142 , n22166 , n22170 );
nand ( n22172 , n3469 , n22171 );
not ( n22173 , n209 );
nand ( n22174 , n8699 , n3729 );
and ( n22175 , n22173 , n22174 );
not ( n22176 , n22173 );
nand ( n22177 , n3731 , n8444 , n8556 , n3703 );
and ( n22178 , n22176 , n22177 );
nor ( n22179 , n22175 , n22178 );
not ( n22180 , n22179 );
not ( n22181 , n211 );
not ( n22182 , n22134 );
not ( n22183 , n3487 );
or ( n22184 , n22182 , n22183 );
nand ( n22185 , n22184 , n209 );
and ( n22186 , n8678 , n22185 );
nand ( n22187 , n22186 , n8682 , n16554 , n16612 );
and ( n22188 , n22181 , n22187 );
not ( n22189 , n22181 );
not ( n22190 , n208 );
or ( n22191 , n22190 , n207 );
not ( n22192 , n3622 );
nand ( n22193 , n22191 , n22192 );
nand ( n22194 , n9303 , n22193 );
nand ( n22195 , n8703 , n8517 , n3613 );
nand ( n22196 , n209 , n22195 );
nand ( n22197 , n22194 , n9341 , n22196 );
and ( n22198 , n22189 , n22197 );
nor ( n22199 , n22188 , n22198 );
not ( n22200 , n22199 );
or ( n22201 , n22180 , n22200 );
nand ( n22202 , n22201 , n212 );
and ( n22203 , n22131 , n22172 , n22202 );
and ( n22204 , n22106 , n22203 );
not ( n22205 , n22106 );
not ( n22206 , n22130 );
nand ( n22207 , n22206 , n22172 , n22202 );
and ( n22208 , n22205 , n22207 );
nor ( n22209 , n22204 , n22208 );
xor ( n22210 , n22102 , n22209 );
nor ( n22211 , n20959 , n22210 );
not ( n22212 , n20959 );
not ( n22213 , n22210 );
or ( n22214 , n22212 , n22213 );
nand ( n22215 , n22214 , n2352 );
or ( n22216 , n22211 , n22215 );
and ( n22217 , n220 , n22100 );
not ( n22218 , n220 );
and ( n22219 , n22218 , n221 );
nor ( n22220 , n22217 , n22219 );
or ( n22221 , n2352 , n22220 );
nand ( n22222 , n22216 , n22221 );
not ( n22223 , n225 );
not ( n22224 , n19202 );
or ( n22225 , n22223 , n22224 );
not ( n22226 , n225 );
not ( n22227 , n19202 );
nand ( n22228 , n22226 , n22227 );
nand ( n22229 , n22225 , n22228 );
and ( n22230 , n22006 , n22008 , n22079 );
and ( n22231 , n22230 , n19452 );
not ( n22232 , n22230 );
and ( n22233 , n22232 , n19333 );
nor ( n22234 , n22231 , n22233 );
not ( n22235 , n22234 );
and ( n22236 , n22229 , n22235 );
not ( n22237 , n22229 );
and ( n22238 , n22237 , n22234 );
nor ( n22239 , n22236 , n22238 );
not ( n22240 , n22239 );
nor ( n22241 , n17155 , n22240 );
or ( n22242 , n17156 , n22239 );
nand ( n22243 , n22242 , n2352 );
or ( n22244 , n22241 , n22243 );
xnor ( n22245 , n225 , n226 );
or ( n22246 , n2352 , n22245 );
nand ( n22247 , n22244 , n22246 );
not ( n22248 , n236 );
and ( n22249 , n237 , n22248 );
not ( n22250 , n237 );
and ( n22251 , n22250 , n236 );
nor ( n22252 , n22249 , n22251 );
or ( n22253 , n2352 , n22252 );
not ( n22254 , n22248 );
not ( n22255 , n7317 );
and ( n22256 , n22254 , n22255 );
and ( n22257 , n22248 , n7317 );
nor ( n22258 , n22256 , n22257 );
and ( n22259 , n22258 , n17319 );
not ( n22260 , n22258 );
and ( n22261 , n22260 , n11573 );
nor ( n22262 , n22259 , n22261 );
not ( n22263 , n22262 );
not ( n22264 , n19889 );
not ( n22265 , n8100 );
and ( n22266 , n22264 , n22265 );
and ( n22267 , n18986 , n15440 );
nor ( n22268 , n22266 , n22267 );
buf ( n22269 , n20448 );
and ( n22270 , n22268 , n22269 );
not ( n22271 , n22268 );
not ( n22272 , n22269 );
and ( n22273 , n22271 , n22272 );
nor ( n22274 , n22270 , n22273 );
not ( n22275 , n22274 );
nand ( n22276 , n22263 , n22275 );
nand ( n22277 , n22262 , n22274 );
nand ( n22278 , n22276 , n2352 , n22277 );
nand ( n22279 , n22253 , n22278 );
not ( n22280 , n16279 );
and ( n22281 , n22280 , n17689 );
not ( n22282 , n22280 );
not ( n22283 , n16259 );
and ( n22284 , n22282 , n22283 );
nor ( n22285 , n22281 , n22284 );
not ( n22286 , n22285 );
not ( n22287 , n255 );
not ( n22288 , n22287 );
not ( n22289 , n10164 );
and ( n22290 , n22288 , n22289 );
and ( n22291 , n22287 , n14707 );
nor ( n22292 , n22290 , n22291 );
not ( n22293 , n22292 );
not ( n22294 , n22293 );
not ( n22295 , n19454 );
not ( n22296 , n22295 );
or ( n22297 , n22294 , n22296 );
nand ( n22298 , n22292 , n19454 );
nand ( n22299 , n22297 , n22298 );
not ( n22300 , n22299 );
nor ( n22301 , n22286 , n22300 );
or ( n22302 , n22285 , n22299 );
nand ( n22303 , n22302 , n2352 );
or ( n22304 , n22301 , n22303 );
and ( n22305 , n254 , n22287 );
not ( n22306 , n254 );
and ( n22307 , n22306 , n255 );
nor ( n22308 , n22305 , n22307 );
or ( n22309 , n2352 , n22308 );
nand ( n22310 , n22304 , n22309 );
not ( n22311 , n100 );
xor ( n22312 , n22311 , n9064 );
xor ( n22313 , n22312 , n12439 );
not ( n22314 , n22313 );
not ( n22315 , n18163 );
not ( n22316 , n22315 );
not ( n22317 , n20959 );
and ( n22318 , n22316 , n22317 );
and ( n22319 , n22315 , n20959 );
nor ( n22320 , n22318 , n22319 );
not ( n22321 , n22320 );
nor ( n22322 , n22314 , n22321 );
or ( n22323 , n22313 , n22320 );
nand ( n22324 , n22323 , n2352 );
or ( n22325 , n22322 , n22324 );
and ( n22326 , n268 , n22311 );
not ( n22327 , n268 );
and ( n22328 , n22327 , n100 );
nor ( n22329 , n22326 , n22328 );
or ( n22330 , n2352 , n22329 );
nand ( n22331 , n22325 , n22330 );
not ( n22332 , n17301 );
not ( n22333 , n11409 );
and ( n22334 , n22332 , n22333 );
and ( n22335 , n17307 , n11409 );
nor ( n22336 , n22334 , n22335 );
not ( n22337 , n272 );
xnor ( n22338 , n22337 , n7317 );
xor ( n22339 , n22336 , n22338 );
not ( n22340 , n22339 );
xnor ( n22341 , n20428 , n17436 );
not ( n22342 , n22341 );
or ( n22343 , n22340 , n22342 );
nand ( n22344 , n22343 , n2352 );
nor ( n22345 , n22339 , n22341 );
or ( n22346 , n22344 , n22345 );
and ( n22347 , n273 , n22337 );
not ( n22348 , n273 );
and ( n22349 , n22348 , n272 );
nor ( n22350 , n22347 , n22349 );
or ( n22351 , n2352 , n22350 );
nand ( n22352 , n22346 , n22351 );
not ( n22353 , n278 );
not ( n22354 , n22353 );
not ( n22355 , n17839 );
or ( n22356 , n22354 , n22355 );
or ( n22357 , n22353 , n17839 );
nand ( n22358 , n22356 , n22357 );
not ( n22359 , n22358 );
not ( n22360 , n15298 );
not ( n22361 , n22360 );
not ( n22362 , n7317 );
not ( n22363 , n22362 );
and ( n22364 , n22361 , n22363 );
and ( n22365 , n22360 , n15038 );
nor ( n22366 , n22364 , n22365 );
not ( n22367 , n22366 );
or ( n22368 , n22359 , n22367 );
or ( n22369 , n22358 , n22366 );
nand ( n22370 , n22368 , n22369 );
not ( n22371 , n22370 );
not ( n22372 , n17868 );
not ( n22373 , n11572 );
and ( n22374 , n22372 , n22373 );
and ( n22375 , n17868 , n11573 );
nor ( n22376 , n22374 , n22375 );
and ( n22377 , n22376 , n15737 );
not ( n22378 , n22376 );
and ( n22379 , n22378 , n15717 );
nor ( n22380 , n22377 , n22379 );
nand ( n22381 , n22371 , n2352 , n22380 );
not ( n22382 , n279 );
or ( n22383 , n22353 , n22382 );
or ( n22384 , n278 , n279 );
nand ( n22385 , n22383 , n22384 , n1 );
not ( n22386 , n22380 );
nand ( n22387 , n22386 , n22370 , n2352 );
nand ( n22388 , n22381 , n22385 , n22387 );
not ( n22389 , n284 );
and ( n22390 , n285 , n22389 );
not ( n22391 , n285 );
and ( n22392 , n22391 , n284 );
nor ( n22393 , n22390 , n22392 );
or ( n22394 , n2352 , n22393 );
and ( n22395 , n16234 , n284 );
not ( n22396 , n16234 );
and ( n22397 , n22396 , n22389 );
nor ( n22398 , n22395 , n22397 );
not ( n22399 , n22398 );
not ( n22400 , n15845 );
not ( n22401 , n20786 );
or ( n22402 , n22400 , n22401 );
or ( n22403 , n15849 , n20786 );
nand ( n22404 , n22402 , n22403 );
not ( n22405 , n10654 );
not ( n22406 , n10164 );
or ( n22407 , n22405 , n22406 );
or ( n22408 , n10654 , n10164 );
nand ( n22409 , n22407 , n22408 );
not ( n22410 , n22409 );
and ( n22411 , n22404 , n22410 );
not ( n22412 , n22404 );
and ( n22413 , n22412 , n22409 );
nor ( n22414 , n22411 , n22413 );
not ( n22415 , n22414 );
nand ( n22416 , n22399 , n22415 );
nand ( n22417 , n22398 , n22414 );
nand ( n22418 , n22416 , n2352 , n22417 );
nand ( n22419 , n22394 , n22418 );
and ( n22420 , n297 , n15302 );
not ( n22421 , n297 );
and ( n22422 , n22421 , n15299 );
nor ( n22423 , n22420 , n22422 );
not ( n22424 , n15434 );
not ( n22425 , n19902 );
and ( n22426 , n22424 , n22425 );
not ( n22427 , n15730 );
not ( n22428 , n22427 );
not ( n22429 , n11913 );
and ( n22430 , n22428 , n22429 );
nor ( n22431 , n22426 , n22430 );
not ( n22432 , n22431 );
not ( n22433 , n22376 );
and ( n22434 , n22432 , n22433 );
and ( n22435 , n22431 , n22376 );
nor ( n22436 , n22434 , n22435 );
nor ( n22437 , n22423 , n22436 );
not ( n22438 , n22423 );
not ( n22439 , n22436 );
or ( n22440 , n22438 , n22439 );
nand ( n22441 , n22440 , n2352 );
or ( n22442 , n22437 , n22441 );
xnor ( n22443 , n297 , n298 );
or ( n22444 , n2352 , n22443 );
nand ( n22445 , n22442 , n22444 );
and ( n22446 , n311 , n16234 );
not ( n22447 , n311 );
and ( n22448 , n22447 , n20677 );
nor ( n22449 , n22446 , n22448 );
not ( n22450 , n22449 );
not ( n22451 , n15845 );
not ( n22452 , n5042 );
and ( n22453 , n22451 , n22452 );
and ( n22454 , n15849 , n5200 );
nor ( n22455 , n22453 , n22454 );
not ( n22456 , n22455 );
not ( n22457 , n20586 );
or ( n22458 , n22456 , n22457 );
or ( n22459 , n22455 , n20586 );
nand ( n22460 , n22458 , n22459 );
not ( n22461 , n22460 );
nor ( n22462 , n22450 , n22461 );
or ( n22463 , n22449 , n22460 );
nand ( n22464 , n22463 , n2352 );
or ( n22465 , n22462 , n22464 );
xnor ( n22466 , n311 , n312 );
or ( n22467 , n2352 , n22466 );
nand ( n22468 , n22465 , n22467 );
not ( n22469 , n18163 );
not ( n22470 , n20606 );
and ( n22471 , n22469 , n22470 );
and ( n22472 , n18163 , n16982 );
nor ( n22473 , n22471 , n22472 );
not ( n22474 , n324 );
not ( n22475 , n12435 );
and ( n22476 , n22474 , n22475 );
and ( n22477 , n324 , n12435 );
nor ( n22478 , n22476 , n22477 );
not ( n22479 , n22478 );
and ( n22480 , n22473 , n22479 );
not ( n22481 , n22473 );
and ( n22482 , n22481 , n22478 );
nor ( n22483 , n22480 , n22482 );
not ( n22484 , n22483 );
not ( n22485 , n20953 );
not ( n22486 , n12564 );
and ( n22487 , n22485 , n22486 );
and ( n22488 , n20953 , n12564 );
nor ( n22489 , n22487 , n22488 );
not ( n22490 , n9514 );
not ( n22491 , n16411 );
and ( n22492 , n22490 , n22491 );
and ( n22493 , n12561 , n16411 );
nor ( n22494 , n22492 , n22493 );
and ( n22495 , n22489 , n22494 );
not ( n22496 , n22489 );
not ( n22497 , n22494 );
and ( n22498 , n22496 , n22497 );
nor ( n22499 , n22495 , n22498 );
not ( n22500 , n22499 );
nor ( n22501 , n22484 , n22500 );
or ( n22502 , n22483 , n22499 );
nand ( n22503 , n22502 , n2352 );
or ( n22504 , n22501 , n22503 );
xnor ( n22505 , n324 , n325 );
or ( n22506 , n2352 , n22505 );
nand ( n22507 , n22504 , n22506 );
not ( n22508 , n330 );
not ( n22509 , n2826 );
and ( n22510 , n22508 , n22509 );
and ( n22511 , n330 , n18083 );
nor ( n22512 , n22510 , n22511 );
not ( n22513 , n9507 );
not ( n22514 , n9781 );
or ( n22515 , n22513 , n22514 );
nand ( n22516 , n9508 , n9657 );
nand ( n22517 , n22515 , n22516 );
not ( n22518 , n22517 );
nand ( n22519 , n18194 , n22518 );
not ( n22520 , n22519 );
nor ( n22521 , n18194 , n22518 );
nor ( n22522 , n22520 , n22521 );
nor ( n22523 , n22512 , n22522 );
not ( n22524 , n22512 );
not ( n22525 , n22522 );
or ( n22526 , n22524 , n22525 );
nand ( n22527 , n22526 , n2352 );
or ( n22528 , n22523 , n22527 );
xnor ( n22529 , n330 , n331 );
or ( n22530 , n2352 , n22529 );
nand ( n22531 , n22528 , n22530 );
not ( n22532 , n357 );
and ( n22533 , n358 , n22532 );
not ( n22534 , n358 );
and ( n22535 , n22534 , n357 );
nor ( n22536 , n22533 , n22535 );
or ( n22537 , n2352 , n22536 );
not ( n22538 , n15996 );
not ( n22539 , n22532 );
not ( n22540 , n10926 );
and ( n22541 , n22539 , n22540 );
and ( n22542 , n22532 , n10913 );
nor ( n22543 , n22541 , n22542 );
not ( n22544 , n22543 );
not ( n22545 , n14861 );
not ( n22546 , n15017 );
not ( n22547 , n22546 );
and ( n22548 , n22545 , n22547 );
not ( n22549 , n12300 );
and ( n22550 , n22549 , n22546 );
nor ( n22551 , n22548 , n22550 );
not ( n22552 , n22551 );
or ( n22553 , n22544 , n22552 );
or ( n22554 , n22543 , n22551 );
nand ( n22555 , n22553 , n22554 );
or ( n22556 , n22538 , n22555 );
not ( n22557 , n15978 );
nand ( n22558 , n22557 , n22555 );
nand ( n22559 , n22556 , n22558 , n2352 );
nand ( n22560 , n22537 , n22559 );
not ( n22561 , n353 );
and ( n22562 , n354 , n22561 );
not ( n22563 , n354 );
and ( n22564 , n22563 , n353 );
nor ( n22565 , n22562 , n22564 );
or ( n22566 , n2352 , n22565 );
not ( n22567 , n22561 );
not ( n22568 , n17300 );
not ( n22569 , n22568 );
and ( n22570 , n22567 , n22569 );
and ( n22571 , n22561 , n17301 );
nor ( n22572 , n22570 , n22571 );
not ( n22573 , n12023 );
and ( n22574 , n22572 , n22573 );
not ( n22575 , n22572 );
and ( n22576 , n22575 , n12023 );
nor ( n22577 , n22574 , n22576 );
not ( n22578 , n22577 );
buf ( n22579 , n20421 );
not ( n22580 , n22579 );
and ( n22581 , n15712 , n22580 );
not ( n22582 , n15712 );
and ( n22583 , n22582 , n22579 );
nor ( n22584 , n22581 , n22583 );
and ( n22585 , n22584 , n15158 );
not ( n22586 , n22584 );
and ( n22587 , n22586 , n15157 );
nor ( n22588 , n22585 , n22587 );
not ( n22589 , n22588 );
nand ( n22590 , n22578 , n22589 );
nand ( n22591 , n22577 , n22588 );
nand ( n22592 , n22590 , n2352 , n22591 );
nand ( n22593 , n22566 , n22592 );
not ( n22594 , n6811 );
not ( n22595 , n17316 );
and ( n22596 , n22594 , n22595 );
not ( n22597 , n11580 );
and ( n22598 , n7093 , n22597 );
nor ( n22599 , n22596 , n22598 );
not ( n22600 , n361 );
not ( n22601 , n17991 );
and ( n22602 , n22600 , n22601 );
not ( n22603 , n17992 );
and ( n22604 , n361 , n22603 );
nor ( n22605 , n22602 , n22604 );
and ( n22606 , n22599 , n22605 );
not ( n22607 , n22599 );
not ( n22608 , n22605 );
and ( n22609 , n22607 , n22608 );
nor ( n22610 , n22606 , n22609 );
not ( n22611 , n22610 );
not ( n22612 , n7910 );
not ( n22613 , n17432 );
and ( n22614 , n22612 , n22613 );
and ( n22615 , n7910 , n20318 );
nor ( n22616 , n22614 , n22615 );
and ( n22617 , n11409 , n11913 );
not ( n22618 , n11409 );
and ( n22619 , n22618 , n22429 );
nor ( n22620 , n22617 , n22619 );
not ( n22621 , n22620 );
and ( n22622 , n22616 , n22621 );
not ( n22623 , n22616 );
and ( n22624 , n22623 , n22620 );
nor ( n22625 , n22622 , n22624 );
not ( n22626 , n22625 );
nor ( n22627 , n22611 , n22626 );
or ( n22628 , n22610 , n22625 );
nand ( n22629 , n22628 , n2352 );
or ( n22630 , n22627 , n22629 );
xnor ( n22631 , n361 , n362 );
or ( n22632 , n2352 , n22631 );
nand ( n22633 , n22630 , n22632 );
not ( n22634 , n17690 );
not ( n22635 , n355 );
not ( n22636 , n22635 );
not ( n22637 , n10913 );
and ( n22638 , n22636 , n22637 );
and ( n22639 , n22635 , n10913 );
nor ( n22640 , n22638 , n22639 );
not ( n22641 , n22640 );
or ( n22642 , n22634 , n22641 );
or ( n22643 , n17690 , n22640 );
nand ( n22644 , n22642 , n22643 );
not ( n22645 , n22644 );
not ( n22646 , n10793 );
not ( n22647 , n16231 );
not ( n22648 , n15988 );
or ( n22649 , n22647 , n22648 );
or ( n22650 , n16231 , n15988 );
nand ( n22651 , n22649 , n22650 );
not ( n22652 , n22651 );
not ( n22653 , n22652 );
or ( n22654 , n22646 , n22653 );
nand ( n22655 , n10789 , n22651 );
nand ( n22656 , n22654 , n22655 );
not ( n22657 , n22656 );
nor ( n22658 , n22645 , n22657 );
or ( n22659 , n22644 , n22656 );
nand ( n22660 , n22659 , n2352 );
or ( n22661 , n22658 , n22660 );
and ( n22662 , n356 , n22635 );
not ( n22663 , n356 );
and ( n22664 , n22663 , n355 );
nor ( n22665 , n22662 , n22664 );
or ( n22666 , n2352 , n22665 );
nand ( n22667 , n22661 , n22666 );
xor ( n22668 , n373 , n22080 );
xnor ( n22669 , n22668 , n18026 );
nand ( n22670 , n20216 , n19454 );
not ( n22671 , n22670 );
nor ( n22672 , n20216 , n19454 );
nor ( n22673 , n22671 , n22672 );
nor ( n22674 , n22669 , n22673 );
not ( n22675 , n22669 );
not ( n22676 , n22673 );
or ( n22677 , n22675 , n22676 );
nand ( n22678 , n22677 , n2352 );
or ( n22679 , n22674 , n22678 );
xnor ( n22680 , n373 , n374 );
or ( n22681 , n2352 , n22680 );
nand ( n22682 , n22679 , n22681 );
xnor ( n22683 , n292 , n293 );
or ( n22684 , n2352 , n22683 );
not ( n22685 , n292 );
not ( n22686 , n16981 );
or ( n22687 , n22685 , n22686 );
or ( n22688 , n292 , n20606 );
nand ( n22689 , n22687 , n22688 );
not ( n22690 , n19563 );
and ( n22691 , n22689 , n22690 );
not ( n22692 , n22689 );
not ( n22693 , n22690 );
and ( n22694 , n22692 , n22693 );
nor ( n22695 , n22691 , n22694 );
not ( n22696 , n22695 );
not ( n22697 , n19695 );
not ( n22698 , n19683 );
nand ( n22699 , n22697 , n22698 , n19765 );
not ( n22700 , n22699 );
not ( n22701 , n22700 );
not ( n22702 , n22701 );
not ( n22703 , n22518 );
and ( n22704 , n22702 , n22703 );
and ( n22705 , n22701 , n22518 );
nor ( n22706 , n22704 , n22705 );
not ( n22707 , n22706 );
nand ( n22708 , n22696 , n22707 );
nand ( n22709 , n22695 , n22706 );
nand ( n22710 , n22708 , n2352 , n22709 );
nand ( n22711 , n22684 , n22710 );
not ( n22712 , n246 );
not ( n22713 , n22712 );
not ( n22714 , n17301 );
and ( n22715 , n22713 , n22714 );
not ( n22716 , n17306 );
and ( n22717 , n22716 , n22712 );
nor ( n22718 , n22715 , n22717 );
xor ( n22719 , n17839 , n22718 );
not ( n22720 , n22719 );
and ( n22721 , n20430 , n22579 );
not ( n22722 , n20430 );
not ( n22723 , n22579 );
and ( n22724 , n22722 , n22723 );
nor ( n22725 , n22721 , n22724 );
xnor ( n22726 , n15158 , n22725 );
not ( n22727 , n22726 );
nor ( n22728 , n22720 , n22727 );
or ( n22729 , n22726 , n22719 );
nand ( n22730 , n22729 , n2352 );
or ( n22731 , n22728 , n22730 );
and ( n22732 , n247 , n22712 );
not ( n22733 , n247 );
and ( n22734 , n22733 , n246 );
nor ( n22735 , n22732 , n22734 );
or ( n22736 , n2352 , n22735 );
nand ( n22737 , n22731 , n22736 );
not ( n22738 , n49 );
not ( n22739 , n18207 );
or ( n22740 , n22738 , n22739 );
or ( n22741 , n49 , n18210 );
nand ( n22742 , n22740 , n22741 );
and ( n22743 , n22742 , n21492 );
not ( n22744 , n22742 );
not ( n22745 , n21250 );
and ( n22746 , n22744 , n22745 );
or ( n22747 , n22743 , n22746 );
not ( n22748 , n18228 );
and ( n22749 , n22748 , n21746 );
not ( n22750 , n22748 );
and ( n22751 , n22750 , n21769 );
nor ( n22752 , n22749 , n22751 );
nor ( n22753 , n22747 , n22752 );
not ( n22754 , n22747 );
not ( n22755 , n22752 );
or ( n22756 , n22754 , n22755 );
nand ( n22757 , n22756 , n2352 );
or ( n22758 , n22753 , n22757 );
xnor ( n22759 , n49 , n50 );
or ( n22760 , n2352 , n22759 );
nand ( n22761 , n22758 , n22760 );
not ( n22762 , n21249 );
not ( n22763 , n22762 );
not ( n22764 , n21620 );
and ( n22765 , n22763 , n22764 );
not ( n22766 , n21364 );
and ( n22767 , n21250 , n22766 );
nor ( n22768 , n22765 , n22767 );
and ( n22769 , n21484 , n53 );
not ( n22770 , n21484 );
not ( n22771 , n53 );
and ( n22772 , n22770 , n22771 );
nor ( n22773 , n22769 , n22772 );
and ( n22774 , n22768 , n22773 );
not ( n22775 , n22768 );
not ( n22776 , n22773 );
and ( n22777 , n22775 , n22776 );
nor ( n22778 , n22774 , n22777 );
not ( n22779 , n22778 );
nor ( n22780 , n14077 , n22779 );
buf ( n22781 , n18522 );
or ( n22782 , n22781 , n22778 );
nand ( n22783 , n22782 , n2352 );
or ( n22784 , n22780 , n22783 );
and ( n22785 , n54 , n22771 );
not ( n22786 , n54 );
and ( n22787 , n22786 , n53 );
nor ( n22788 , n22785 , n22787 );
or ( n22789 , n2352 , n22788 );
nand ( n22790 , n22784 , n22789 );
not ( n22791 , n14206 );
not ( n22792 , n48 );
not ( n22793 , n22792 );
not ( n22794 , n21837 );
not ( n22795 , n22794 );
and ( n22796 , n22793 , n22795 );
not ( n22797 , n21484 );
and ( n22798 , n22792 , n22797 );
nor ( n22799 , n22796 , n22798 );
xnor ( n22800 , n22791 , n22799 );
not ( n22801 , n22800 );
buf ( n22802 , n13834 );
not ( n22803 , n22802 );
and ( n22804 , n22803 , n21746 );
not ( n22805 , n22803 );
and ( n22806 , n22805 , n21769 );
nor ( n22807 , n22804 , n22806 );
not ( n22808 , n22807 );
nor ( n22809 , n22801 , n22808 );
or ( n22810 , n22800 , n22807 );
nand ( n22811 , n22810 , n2352 );
or ( n22812 , n22809 , n22811 );
and ( n22813 , n57 , n22792 );
not ( n22814 , n57 );
and ( n22815 , n22814 , n48 );
nor ( n22816 , n22813 , n22815 );
or ( n22817 , n2352 , n22816 );
nand ( n22818 , n22812 , n22817 );
not ( n22819 , n21020 );
xnor ( n22820 , n59 , n9084 );
xor ( n22821 , n22819 , n22820 );
not ( n22822 , n22821 );
not ( n22823 , n14594 );
not ( n22824 , n6480 );
not ( n22825 , n22824 );
not ( n22826 , n22825 );
and ( n22827 , n22823 , n22826 );
and ( n22828 , n22825 , n14594 );
nor ( n22829 , n22827 , n22828 );
buf ( n22830 , n14660 );
and ( n22831 , n22829 , n22830 );
not ( n22832 , n22829 );
not ( n22833 , n22830 );
and ( n22834 , n22832 , n22833 );
nor ( n22835 , n22831 , n22834 );
not ( n22836 , n22835 );
nor ( n22837 , n22822 , n22836 );
or ( n22838 , n22821 , n22835 );
nand ( n22839 , n22838 , n2352 );
or ( n22840 , n22837 , n22839 );
xnor ( n22841 , n59 , n60 );
or ( n22842 , n2352 , n22841 );
nand ( n22843 , n22840 , n22842 );
not ( n22844 , n61 );
and ( n22845 , n62 , n22844 );
not ( n22846 , n62 );
and ( n22847 , n22846 , n61 );
nor ( n22848 , n22845 , n22847 );
or ( n22849 , n2352 , n22848 );
not ( n22850 , n61 );
not ( n22851 , n5835 );
or ( n22852 , n22850 , n22851 );
nand ( n22853 , n22844 , n9084 );
nand ( n22854 , n22852 , n22853 );
and ( n22855 , n22854 , n21027 );
not ( n22856 , n22854 );
not ( n22857 , n21018 );
and ( n22858 , n22856 , n22857 );
nor ( n22859 , n22855 , n22858 );
not ( n22860 , n22859 );
not ( n22861 , n22830 );
not ( n22862 , n21035 );
and ( n22863 , n22861 , n22862 );
and ( n22864 , n22830 , n21035 );
nor ( n22865 , n22863 , n22864 );
not ( n22866 , n22865 );
nand ( n22867 , n22860 , n22866 );
nand ( n22868 , n22859 , n22865 );
nand ( n22869 , n22867 , n2352 , n22868 );
nand ( n22870 , n22849 , n22869 );
and ( n22871 , n80 , n14347 );
not ( n22872 , n80 );
and ( n22873 , n22872 , n14348 );
nor ( n22874 , n22871 , n22873 );
not ( n22875 , n22874 );
not ( n22876 , n14461 );
not ( n22877 , n13613 );
or ( n22878 , n22876 , n22877 );
or ( n22879 , n14467 , n13613 );
nand ( n22880 , n22878 , n22879 );
not ( n22881 , n22880 );
not ( n22882 , n1472 );
not ( n22883 , n5989 );
and ( n22884 , n22882 , n22883 );
and ( n22885 , n9101 , n5989 );
nor ( n22886 , n22884 , n22885 );
not ( n22887 , n22886 );
or ( n22888 , n22881 , n22887 );
or ( n22889 , n22880 , n22886 );
nand ( n22890 , n22888 , n22889 );
not ( n22891 , n22890 );
nor ( n22892 , n22875 , n22891 );
or ( n22893 , n22874 , n22890 );
nand ( n22894 , n22893 , n2352 );
or ( n22895 , n22892 , n22894 );
xnor ( n22896 , n80 , n83 );
or ( n22897 , n2352 , n22896 );
nand ( n22898 , n22895 , n22897 );
xnor ( n22899 , n162 , n179 );
or ( n22900 , n2352 , n22899 );
not ( n22901 , n162 );
not ( n22902 , n10159 );
not ( n22903 , n22902 );
and ( n22904 , n22901 , n22903 );
not ( n22905 , n10159 );
and ( n22906 , n162 , n22905 );
nor ( n22907 , n22904 , n22906 );
and ( n22908 , n22907 , n17689 );
not ( n22909 , n22907 );
and ( n22910 , n22909 , n22283 );
nor ( n22911 , n22908 , n22910 );
not ( n22912 , n22911 );
not ( n22913 , n5665 );
not ( n22914 , n22234 );
and ( n22915 , n22913 , n22914 );
and ( n22916 , n5665 , n22234 );
nor ( n22917 , n22915 , n22916 );
not ( n22918 , n22917 );
nand ( n22919 , n22912 , n22918 );
nand ( n22920 , n22911 , n22917 );
nand ( n22921 , n22919 , n2352 , n22920 );
nand ( n22922 , n22900 , n22921 );
not ( n22923 , n196 );
not ( n22924 , n2985 );
and ( n22925 , n22923 , n22924 );
not ( n22926 , n2990 );
and ( n22927 , n196 , n22926 );
nor ( n22928 , n22925 , n22927 );
not ( n22929 , n16988 );
and ( n22930 , n22928 , n22929 );
not ( n22931 , n22928 );
not ( n22932 , n22929 );
and ( n22933 , n22931 , n22932 );
nor ( n22934 , n22930 , n22933 );
xor ( n22935 , n9782 , n22209 );
nor ( n22936 , n22934 , n22935 );
not ( n22937 , n22934 );
not ( n22938 , n22935 );
or ( n22939 , n22937 , n22938 );
nand ( n22940 , n22939 , n2352 );
or ( n22941 , n22936 , n22940 );
xnor ( n22942 , n196 , n213 );
or ( n22943 , n2352 , n22942 );
nand ( n22944 , n22941 , n22943 );
not ( n22945 , n109 );
and ( n22946 , n214 , n22945 );
not ( n22947 , n214 );
and ( n22948 , n22947 , n109 );
nor ( n22949 , n22946 , n22948 );
or ( n22950 , n2352 , n22949 );
and ( n22951 , n19090 , n22945 );
not ( n22952 , n19090 );
and ( n22953 , n22952 , n109 );
nor ( n22954 , n22951 , n22953 );
and ( n22955 , n22954 , n22269 );
not ( n22956 , n22954 );
not ( n22957 , n22269 );
and ( n22958 , n22956 , n22957 );
nor ( n22959 , n22955 , n22958 );
not ( n22960 , n22959 );
nand ( n22961 , n7748 , n19842 );
not ( n22962 , n19873 );
not ( n22963 , n126 );
nand ( n22964 , n22963 , n7813 , n19849 );
nand ( n22965 , n19881 , n22964 , n19854 );
or ( n22966 , n22962 , n22965 );
nand ( n22967 , n22966 , n127 );
nand ( n22968 , n19804 , n19805 , n22961 , n22967 );
not ( n22969 , n22968 );
not ( n22970 , n18777 );
and ( n22971 , n22969 , n22970 );
not ( n22972 , n22969 );
and ( n22973 , n22972 , n18777 );
nor ( n22974 , n22971 , n22973 );
and ( n22975 , n22974 , n20189 );
not ( n22976 , n22974 );
not ( n22977 , n20186 );
and ( n22978 , n22976 , n22977 );
nor ( n22979 , n22975 , n22978 );
not ( n22980 , n22979 );
nand ( n22981 , n22960 , n22980 );
nand ( n22982 , n22959 , n22979 );
nand ( n22983 , n22981 , n2352 , n22982 );
nand ( n22984 , n22950 , n22983 );
not ( n22985 , n102 );
not ( n22986 , n22926 );
and ( n22987 , n22985 , n22986 );
and ( n22988 , n102 , n22926 );
nor ( n22989 , n22987 , n22988 );
and ( n22990 , n22989 , n22690 );
not ( n22991 , n22989 );
not ( n22992 , n22690 );
and ( n22993 , n22991 , n22992 );
nor ( n22994 , n22990 , n22993 );
and ( n22995 , n19668 , n22517 );
not ( n22996 , n19668 );
and ( n22997 , n22996 , n22518 );
nor ( n22998 , n22995 , n22997 );
nor ( n22999 , n22994 , n22998 );
not ( n23000 , n22994 );
not ( n23001 , n22998 );
or ( n23002 , n23000 , n23001 );
nand ( n23003 , n23002 , n2352 );
or ( n23004 , n22999 , n23003 );
not ( n23005 , n102 );
and ( n23006 , n222 , n23005 );
not ( n23007 , n222 );
and ( n23008 , n23007 , n102 );
nor ( n23009 , n23006 , n23008 );
or ( n23010 , n2352 , n23009 );
nand ( n23011 , n23004 , n23010 );
not ( n23012 , n234 );
not ( n23013 , n23012 );
and ( n23014 , n16863 , n16837 , n16818 );
not ( n23015 , n23014 );
and ( n23016 , n23013 , n23015 );
and ( n23017 , n23012 , n20989 );
nor ( n23018 , n23016 , n23017 );
and ( n23019 , n23018 , n20245 );
not ( n23020 , n23018 );
and ( n23021 , n23020 , n20248 );
nor ( n23022 , n23019 , n23021 );
not ( n23023 , n23022 );
not ( n23024 , n9240 );
xor ( n23025 , n16736 , n23024 );
not ( n23026 , n9239 );
not ( n23027 , n23026 );
xnor ( n23028 , n23025 , n23027 );
not ( n23029 , n23028 );
nor ( n23030 , n23023 , n23029 );
or ( n23031 , n23022 , n23028 );
nand ( n23032 , n23031 , n2352 );
or ( n23033 , n23030 , n23032 );
and ( n23034 , n235 , n23012 );
not ( n23035 , n235 );
and ( n23036 , n23035 , n234 );
nor ( n23037 , n23034 , n23036 );
or ( n23038 , n2352 , n23037 );
nand ( n23039 , n23033 , n23038 );
not ( n23040 , n238 );
not ( n23041 , n23040 );
not ( n23042 , n17306 );
not ( n23043 , n23042 );
and ( n23044 , n23041 , n23043 );
and ( n23045 , n23040 , n22716 );
nor ( n23046 , n23044 , n23045 );
and ( n23047 , n11753 , n12020 );
not ( n23048 , n11753 );
and ( n23049 , n23048 , n12023 );
nor ( n23050 , n23047 , n23049 );
and ( n23051 , n23046 , n23050 );
not ( n23052 , n23046 );
not ( n23053 , n23050 );
and ( n23054 , n23052 , n23053 );
nor ( n23055 , n23051 , n23054 );
not ( n23056 , n23055 );
nor ( n23057 , n15717 , n23056 );
or ( n23058 , n15737 , n23055 );
nand ( n23059 , n23058 , n2352 );
or ( n23060 , n23057 , n23059 );
and ( n23061 , n239 , n23040 );
not ( n23062 , n239 );
and ( n23063 , n23062 , n238 );
nor ( n23064 , n23061 , n23063 );
or ( n23065 , n2352 , n23064 );
nand ( n23066 , n23060 , n23065 );
and ( n23067 , n17838 , n12023 );
not ( n23068 , n17838 );
and ( n23069 , n23068 , n12020 );
nor ( n23070 , n23067 , n23069 );
not ( n23071 , n248 );
and ( n23072 , n23070 , n23071 );
not ( n23073 , n23070 );
and ( n23074 , n23073 , n248 );
nor ( n23075 , n23072 , n23074 );
not ( n23076 , n23075 );
xnor ( n23077 , n15565 , n22725 );
not ( n23078 , n23077 );
nor ( n23079 , n23076 , n23078 );
or ( n23080 , n23077 , n23075 );
nand ( n23081 , n23080 , n2352 );
or ( n23082 , n23079 , n23081 );
and ( n23083 , n249 , n23071 );
not ( n23084 , n249 );
and ( n23085 , n23084 , n248 );
nor ( n23086 , n23083 , n23085 );
or ( n23087 , n2352 , n23086 );
nand ( n23088 , n23082 , n23087 );
xnor ( n23089 , n256 , n257 );
or ( n23090 , n2352 , n23089 );
not ( n23091 , n257 );
not ( n23092 , n10158 );
and ( n23093 , n23091 , n23092 );
and ( n23094 , n257 , n22905 );
nor ( n23095 , n23093 , n23094 );
buf ( n23096 , n19202 );
and ( n23097 , n23095 , n23096 );
not ( n23098 , n23095 );
not ( n23099 , n23096 );
and ( n23100 , n23098 , n23099 );
nor ( n23101 , n23097 , n23100 );
not ( n23102 , n23101 );
not ( n23103 , n22080 );
not ( n23104 , n23103 );
not ( n23105 , n20793 );
and ( n23106 , n23104 , n23105 );
and ( n23107 , n22081 , n20793 );
nor ( n23108 , n23106 , n23107 );
not ( n23109 , n23108 );
nand ( n23110 , n23102 , n23109 );
nand ( n23111 , n23101 , n23108 );
nand ( n23112 , n23110 , n2352 , n23111 );
nand ( n23113 , n23090 , n23112 );
not ( n23114 , n262 );
and ( n23115 , n263 , n23114 );
not ( n23116 , n263 );
and ( n23117 , n23116 , n262 );
nor ( n23118 , n23115 , n23117 );
or ( n23119 , n2352 , n23118 );
and ( n23120 , n22700 , n22203 );
not ( n23121 , n22700 );
and ( n23122 , n23121 , n22207 );
nor ( n23123 , n23120 , n23122 );
not ( n23124 , n23123 );
not ( n23125 , n23114 );
not ( n23126 , n2990 );
or ( n23127 , n23125 , n23126 );
or ( n23128 , n23114 , n2990 );
nand ( n23129 , n23127 , n23128 );
not ( n23130 , n23129 );
not ( n23131 , n9512 );
not ( n23132 , n3466 );
or ( n23133 , n23131 , n23132 );
or ( n23134 , n9509 , n3466 );
nand ( n23135 , n23133 , n23134 );
not ( n23136 , n23135 );
or ( n23137 , n23130 , n23136 );
or ( n23138 , n23129 , n23135 );
nand ( n23139 , n23137 , n23138 );
or ( n23140 , n23124 , n23139 );
not ( n23141 , n22699 );
and ( n23142 , n23141 , n22207 );
not ( n23143 , n23141 );
and ( n23144 , n23143 , n22203 );
nor ( n23145 , n23142 , n23144 );
nand ( n23146 , n23145 , n23139 );
nand ( n23147 , n23140 , n23146 , n2352 );
nand ( n23148 , n23119 , n23147 );
buf ( n23149 , n20242 );
not ( n23150 , n23149 );
not ( n23151 , n23150 );
not ( n23152 , n103 );
not ( n23153 , n23152 );
not ( n23154 , n23014 );
and ( n23155 , n23153 , n23154 );
and ( n23156 , n23152 , n16865 );
nor ( n23157 , n23155 , n23156 );
not ( n23158 , n23157 );
and ( n23159 , n23151 , n23158 );
not ( n23160 , n23149 );
and ( n23161 , n23160 , n23157 );
nor ( n23162 , n23159 , n23161 );
not ( n23163 , n23162 );
not ( n23164 , n23026 );
not ( n23165 , n23164 );
not ( n23166 , n20261 );
or ( n23167 , n23165 , n23166 );
or ( n23168 , n23164 , n20261 );
nand ( n23169 , n23167 , n23168 );
not ( n23170 , n23169 );
nor ( n23171 , n23163 , n23170 );
or ( n23172 , n23162 , n23169 );
nand ( n23173 , n23172 , n2352 );
or ( n23174 , n23171 , n23173 );
and ( n23175 , n264 , n23152 );
not ( n23176 , n264 );
and ( n23177 , n23176 , n103 );
nor ( n23178 , n23175 , n23177 );
or ( n23179 , n2352 , n23178 );
nand ( n23180 , n23174 , n23179 );
and ( n23181 , n274 , n15302 );
not ( n23182 , n274 );
and ( n23183 , n23182 , n15299 );
nor ( n23184 , n23181 , n23183 );
not ( n23185 , n23184 );
not ( n23186 , n22427 );
not ( n23187 , n17862 );
or ( n23188 , n23186 , n23187 );
or ( n23189 , n22427 , n17862 );
nand ( n23190 , n23188 , n23189 );
not ( n23191 , n23190 );
not ( n23192 , n17316 );
not ( n23193 , n7317 );
and ( n23194 , n23192 , n23193 );
and ( n23195 , n22597 , n7317 );
nor ( n23196 , n23194 , n23195 );
not ( n23197 , n23196 );
or ( n23198 , n23191 , n23197 );
or ( n23199 , n23190 , n23196 );
nand ( n23200 , n23198 , n23199 );
not ( n23201 , n23200 );
nor ( n23202 , n23185 , n23201 );
or ( n23203 , n23184 , n23200 );
nand ( n23204 , n23203 , n2352 );
or ( n23205 , n23202 , n23204 );
xnor ( n23206 , n274 , n275 );
or ( n23207 , n2352 , n23206 );
nand ( n23208 , n23205 , n23207 );
not ( n23209 , n7912 );
not ( n23210 , n23209 );
not ( n23211 , n280 );
not ( n23212 , n23211 );
not ( n23213 , n20083 );
or ( n23214 , n23212 , n23213 );
or ( n23215 , n23211 , n20083 );
nand ( n23216 , n23214 , n23215 );
not ( n23217 , n23216 );
not ( n23218 , n18777 );
not ( n23219 , n23218 );
not ( n23220 , n20185 );
and ( n23221 , n23219 , n23220 );
and ( n23222 , n22970 , n20185 );
nor ( n23223 , n23221 , n23222 );
not ( n23224 , n23223 );
or ( n23225 , n23217 , n23224 );
or ( n23226 , n23216 , n23223 );
nand ( n23227 , n23225 , n23226 );
not ( n23228 , n23227 );
nor ( n23229 , n23210 , n23228 );
or ( n23230 , n23209 , n23227 );
nand ( n23231 , n23230 , n2352 );
or ( n23232 , n23229 , n23231 );
and ( n23233 , n281 , n23211 );
not ( n23234 , n281 );
and ( n23235 , n23234 , n280 );
nor ( n23236 , n23233 , n23235 );
or ( n23237 , n2352 , n23236 );
nand ( n23238 , n23232 , n23237 );
not ( n23239 , n101 );
xor ( n23240 , n23239 , n19563 );
xnor ( n23241 , n23240 , n9064 );
and ( n23242 , n10958 , n23123 );
not ( n23243 , n10958 );
and ( n23244 , n23243 , n23145 );
nor ( n23245 , n23242 , n23244 );
nor ( n23246 , n23241 , n23245 );
not ( n23247 , n23241 );
not ( n23248 , n23245 );
or ( n23249 , n23247 , n23248 );
nand ( n23250 , n23249 , n2352 );
or ( n23251 , n23246 , n23250 );
and ( n23252 , n296 , n23239 );
not ( n23253 , n296 );
and ( n23254 , n23253 , n101 );
nor ( n23255 , n23252 , n23254 );
or ( n23256 , n2352 , n23255 );
nand ( n23257 , n23251 , n23256 );
not ( n23258 , n305 );
and ( n23259 , n23258 , n17992 );
not ( n23260 , n23258 );
and ( n23261 , n23260 , n17991 );
or ( n23262 , n23259 , n23261 );
xor ( n23263 , n23262 , n20185 );
xor ( n23264 , n7907 , n18784 );
nor ( n23265 , n23263 , n23264 );
not ( n23266 , n23263 );
not ( n23267 , n23264 );
or ( n23268 , n23266 , n23267 );
nand ( n23269 , n23268 , n2352 );
or ( n23270 , n23265 , n23269 );
and ( n23271 , n306 , n23258 );
not ( n23272 , n306 );
and ( n23273 , n23272 , n305 );
nor ( n23274 , n23271 , n23273 );
or ( n23275 , n2352 , n23274 );
nand ( n23276 , n23270 , n23275 );
not ( n23277 , n346 );
not ( n23278 , n23277 );
not ( n23279 , n14858 );
or ( n23280 , n23278 , n23279 );
or ( n23281 , n23277 , n14864 );
nand ( n23282 , n23280 , n23281 );
xor ( n23283 , n23282 , n22651 );
not ( n23284 , n23283 );
xor ( n23285 , n20786 , n5200 );
and ( n23286 , n23285 , n15851 );
not ( n23287 , n23285 );
and ( n23288 , n23287 , n15985 );
nor ( n23289 , n23286 , n23288 );
not ( n23290 , n23289 );
or ( n23291 , n23284 , n23290 );
nand ( n23292 , n23291 , n2352 );
nor ( n23293 , n23283 , n23289 );
or ( n23294 , n23292 , n23293 );
and ( n23295 , n347 , n23277 );
not ( n23296 , n347 );
and ( n23297 , n23296 , n346 );
nor ( n23298 , n23295 , n23297 );
or ( n23299 , n2352 , n23298 );
nand ( n23300 , n23294 , n23299 );
not ( n23301 , n349 );
and ( n23302 , n350 , n23301 );
not ( n23303 , n350 );
and ( n23304 , n23303 , n349 );
nor ( n23305 , n23302 , n23304 );
or ( n23306 , n2352 , n23305 );
not ( n23307 , n23301 );
not ( n23308 , n7317 );
or ( n23309 , n23307 , n23308 );
or ( n23310 , n23301 , n7317 );
nand ( n23311 , n23309 , n23310 );
buf ( n23312 , n19090 );
and ( n23313 , n23311 , n23312 );
not ( n23314 , n23311 );
not ( n23315 , n23312 );
and ( n23316 , n23314 , n23315 );
nor ( n23317 , n23313 , n23316 );
not ( n23318 , n23317 );
and ( n23319 , n15438 , n19902 );
not ( n23320 , n15438 );
and ( n23321 , n23320 , n19901 );
or ( n23322 , n23319 , n23321 );
and ( n23323 , n23322 , n22269 );
not ( n23324 , n23322 );
and ( n23325 , n23324 , n22957 );
nor ( n23326 , n23323 , n23325 );
not ( n23327 , n23326 );
nand ( n23328 , n23318 , n23327 );
nand ( n23329 , n23317 , n23326 );
nand ( n23330 , n23328 , n2352 , n23329 );
nand ( n23331 , n23306 , n23330 );
not ( n23332 , n365 );
and ( n23333 , n366 , n23332 );
not ( n23334 , n366 );
and ( n23335 , n23334 , n365 );
nor ( n23336 , n23333 , n23335 );
or ( n23337 , n2352 , n23336 );
not ( n23338 , n18097 );
not ( n23339 , n23332 );
not ( n23340 , n23014 );
or ( n23341 , n23339 , n23340 );
or ( n23342 , n23332 , n23014 );
nand ( n23343 , n23341 , n23342 );
not ( n23344 , n23343 );
nand ( n23345 , n16934 , n16970 );
nor ( n23346 , n16919 , n23345 );
not ( n23347 , n23346 );
not ( n23348 , n20257 );
or ( n23349 , n23347 , n23348 );
or ( n23350 , n23346 , n16623 );
nand ( n23351 , n23349 , n23350 );
not ( n23352 , n23351 );
or ( n23353 , n23344 , n23352 );
or ( n23354 , n23343 , n23351 );
nand ( n23355 , n23353 , n23354 );
not ( n23356 , n23355 );
nand ( n23357 , n23338 , n23356 );
nand ( n23358 , n18097 , n23355 );
nand ( n23359 , n23357 , n2352 , n23358 );
nand ( n23360 , n23337 , n23359 );
and ( n23361 , n378 , n15302 );
not ( n23362 , n378 );
and ( n23363 , n23362 , n15299 );
nor ( n23364 , n23361 , n23363 );
not ( n23365 , n17658 );
not ( n23366 , n23322 );
not ( n23367 , n23366 );
and ( n23368 , n23365 , n23367 );
and ( n23369 , n17658 , n23366 );
nor ( n23370 , n23368 , n23369 );
nor ( n23371 , n23364 , n23370 );
not ( n23372 , n23364 );
not ( n23373 , n23370 );
or ( n23374 , n23372 , n23373 );
nand ( n23375 , n23374 , n2352 );
or ( n23376 , n23371 , n23375 );
xnor ( n23377 , n378 , n379 );
or ( n23378 , n2352 , n23377 );
nand ( n23379 , n23376 , n23378 );
not ( n23380 , n23312 );
not ( n23381 , n230 );
not ( n23382 , n23381 );
not ( n23383 , n17316 );
or ( n23384 , n23382 , n23383 );
or ( n23385 , n23381 , n22597 );
nand ( n23386 , n23384 , n23385 );
not ( n23387 , n23386 );
or ( n23388 , n23380 , n23387 );
or ( n23389 , n23312 , n23386 );
nand ( n23390 , n23388 , n23389 );
not ( n23391 , n23390 );
and ( n23392 , n23322 , n22969 );
not ( n23393 , n23322 );
not ( n23394 , n22969 );
and ( n23395 , n23393 , n23394 );
nor ( n23396 , n23392 , n23395 );
not ( n23397 , n23396 );
nor ( n23398 , n23391 , n23397 );
or ( n23399 , n23390 , n23396 );
nand ( n23400 , n23399 , n2352 );
or ( n23401 , n23398 , n23400 );
and ( n23402 , n231 , n23381 );
not ( n23403 , n231 );
and ( n23404 , n23403 , n230 );
nor ( n23405 , n23402 , n23404 );
or ( n23406 , n2352 , n23405 );
nand ( n23407 , n23401 , n23406 );
xor ( n23408 , n244 , n19667 );
xnor ( n23409 , n23408 , n9064 );
and ( n23410 , n11092 , n23145 );
not ( n23411 , n11092 );
and ( n23412 , n23411 , n23123 );
nor ( n23413 , n23410 , n23412 );
nor ( n23414 , n23409 , n23413 );
not ( n23415 , n23409 );
not ( n23416 , n23413 );
or ( n23417 , n23415 , n23416 );
nand ( n23418 , n23417 , n2352 );
or ( n23419 , n23414 , n23418 );
xnor ( n23420 , n244 , n245 );
or ( n23421 , n2352 , n23420 );
nand ( n23422 , n23419 , n23421 );
xor ( n23423 , n299 , n20076 );
not ( n23424 , n17996 );
xnor ( n23425 , n23423 , n23424 );
xor ( n23426 , n7093 , n18784 );
nor ( n23427 , n23425 , n23426 );
not ( n23428 , n23425 );
not ( n23429 , n23426 );
or ( n23430 , n23428 , n23429 );
nand ( n23431 , n23430 , n2352 );
or ( n23432 , n23427 , n23431 );
xnor ( n23433 , n299 , n300 );
or ( n23434 , n2352 , n23433 );
nand ( n23435 , n23432 , n23434 );
not ( n23436 , n351 );
not ( n23437 , n23436 );
not ( n23438 , n10654 );
or ( n23439 , n23437 , n23438 );
or ( n23440 , n23436 , n10654 );
nand ( n23441 , n23439 , n23440 );
and ( n23442 , n23441 , n23096 );
not ( n23443 , n23441 );
not ( n23444 , n23096 );
and ( n23445 , n23443 , n23444 );
nor ( n23446 , n23442 , n23445 );
not ( n23447 , n23446 );
not ( n23448 , n22089 );
not ( n23449 , n20793 );
or ( n23450 , n23448 , n23449 );
or ( n23451 , n22089 , n20793 );
nand ( n23452 , n23450 , n23451 );
not ( n23453 , n23452 );
nor ( n23454 , n23447 , n23453 );
or ( n23455 , n23446 , n23452 );
nand ( n23456 , n23455 , n2352 );
or ( n23457 , n23454 , n23456 );
and ( n23458 , n352 , n23436 );
not ( n23459 , n352 );
and ( n23460 , n23459 , n351 );
nor ( n23461 , n23458 , n23460 );
or ( n23462 , n2352 , n23461 );
nand ( n23463 , n23457 , n23462 );
not ( n23464 , n67 );
not ( n23465 , n2007 );
or ( n23466 , n23464 , n23465 );
or ( n23467 , n67 , n2007 );
nand ( n23468 , n23466 , n23467 );
not ( n23469 , n79 );
not ( n23470 , n14228 );
or ( n23471 , n23469 , n23470 );
or ( n23472 , n79 , n14228 );
nand ( n23473 , n23471 , n23472 );
not ( n23474 , n61 );
not ( n23475 , n2341 );
or ( n23476 , n23474 , n23475 );
not ( n23477 , n22819 );
or ( n23478 , n61 , n23477 );
nand ( n23479 , n23476 , n23478 );
buf ( n23480 , n22833 );
and ( n23481 , n23480 , n21908 );
not ( n23482 , n23480 );
and ( n23483 , n23482 , n73 );
nor ( n23484 , n23481 , n23483 );
not ( n23485 , n40 );
not ( n23486 , n18393 );
or ( n23487 , n23485 , n23486 );
or ( n23488 , n40 , n18393 );
nand ( n23489 , n23487 , n23488 );
and ( n23490 , n39 , n18499 );
not ( n23491 , n39 );
and ( n23492 , n23491 , n18500 );
nor ( n23493 , n23490 , n23492 );
not ( n23494 , n18237 );
and ( n23495 , n95 , n23494 );
not ( n23496 , n95 );
and ( n23497 , n23496 , n18237 );
nor ( n23498 , n23495 , n23497 );
not ( n23499 , n93 );
not ( n23500 , n14348 );
or ( n23501 , n23499 , n23500 );
or ( n23502 , n93 , n14348 );
nand ( n23503 , n23501 , n23502 );
not ( n23504 , n21159 );
and ( n23505 , n23504 , n37 );
not ( n23506 , n23504 );
and ( n23507 , n23506 , n21375 );
nor ( n23508 , n23505 , n23507 );
not ( n23509 , n55 );
not ( n23510 , n14070 );
or ( n23511 , n23509 , n23510 );
or ( n23512 , n55 , n14070 );
nand ( n23513 , n23511 , n23512 );
not ( n23514 , n43 );
not ( n23515 , n14226 );
or ( n23516 , n23514 , n23515 );
or ( n23517 , n43 , n14226 );
nand ( n23518 , n23516 , n23517 );
and ( n23519 , n14631 , n90 );
not ( n23520 , n14631 );
and ( n23521 , n23520 , n21946 );
nor ( n23522 , n23519 , n23521 );
not ( n23523 , n49 );
not ( n23524 , n21486 );
or ( n23525 , n23523 , n23524 );
or ( n23526 , n49 , n21486 );
nand ( n23527 , n23525 , n23526 );
and ( n23528 , n45 , n21779 );
not ( n23529 , n45 );
and ( n23530 , n23529 , n21782 );
nor ( n23531 , n23528 , n23530 );
not ( n23532 , n106 );
not ( n23533 , n111 );
or ( n23534 , n23532 , n23533 );
and ( n23535 , n18 , n21971 );
and ( n23536 , n110 , n21045 );
nor ( n23537 , n23535 , n23536 );
not ( n23538 , n102 );
nor ( n23539 , n23538 , n101 );
nand ( n23540 , n100 , n23539 );
nor ( n23541 , n20271 , n23540 );
nand ( n23542 , n23152 , n23541 );
nor ( n23543 , n23152 , n99 );
nor ( n23544 , n101 , n102 );
and ( n23545 , n23543 , n98 , n23544 );
nor ( n23546 , n98 , n99 );
and ( n23547 , n23546 , n100 , n101 );
nor ( n23548 , n23545 , n23547 );
not ( n23549 , n23539 );
not ( n23550 , n98 );
nor ( n23551 , n23549 , n23550 );
or ( n23552 , n20271 , n23551 );
nand ( n23553 , n101 , n102 );
not ( n23554 , n23553 );
nand ( n23555 , n100 , n23554 );
or ( n23556 , n23152 , n23555 );
nand ( n23557 , n23556 , n20271 );
nand ( n23558 , n23552 , n23557 );
not ( n23559 , n98 );
not ( n23560 , n23540 );
not ( n23561 , n23560 );
or ( n23562 , n23559 , n23561 );
not ( n23563 , n100 );
not ( n23564 , n102 );
nand ( n23565 , n23564 , n101 );
not ( n23566 , n23565 );
nand ( n23567 , n23563 , n23566 );
not ( n23568 , n23567 );
nand ( n23569 , n99 , n23568 );
nand ( n23570 , n23562 , n23569 );
nand ( n23571 , n23152 , n23570 );
nand ( n23572 , n23542 , n23548 , n23558 , n23571 );
and ( n23573 , n2358 , n23572 );
not ( n23574 , n98 );
nand ( n23575 , n20271 , n23560 );
or ( n23576 , n23574 , n23575 );
not ( n23577 , n100 );
nand ( n23578 , n23577 , n23544 );
not ( n23579 , n23578 );
nand ( n23580 , n99 , n23579 );
not ( n23581 , n98 );
nand ( n23582 , n20271 , n23581 , n23544 );
nand ( n23583 , n23576 , n23580 , n23582 );
and ( n23584 , n23583 , n103 , n104 );
nor ( n23585 , n23573 , n23584 );
not ( n23586 , n104 );
nor ( n23587 , n22311 , n23565 );
nand ( n23588 , n99 , n98 , n23587 );
nor ( n23589 , n99 , n23578 );
nand ( n23590 , n23152 , n23589 );
not ( n23591 , n98 );
and ( n23592 , n103 , n23591 , n20271 );
and ( n23593 , n23592 , n22311 , n23005 );
nand ( n23594 , n99 , n103 );
nand ( n23595 , n100 , n102 );
nor ( n23596 , n23594 , n98 , n23595 );
nor ( n23597 , n23593 , n23596 );
nand ( n23598 , n23588 , n23590 , n23597 );
not ( n23599 , n23598 );
or ( n23600 , n23586 , n23599 );
not ( n23601 , n98 );
nor ( n23602 , n100 , n101 );
nand ( n23603 , n20271 , n23601 , n23602 );
not ( n23604 , n23603 );
not ( n23605 , n98 );
nor ( n23606 , n100 , n23553 );
nand ( n23607 , n99 , n23605 , n23606 );
not ( n23608 , n23607 );
or ( n23609 , n23604 , n23608 );
nand ( n23610 , n23609 , n103 );
nand ( n23611 , n23600 , n23610 );
not ( n23612 , n23611 );
or ( n23613 , n23239 , n100 );
not ( n23614 , n100 );
nand ( n23615 , n23614 , n102 );
nand ( n23616 , n23613 , n23615 );
and ( n23617 , n23616 , n98 , n20271 );
not ( n23618 , n98 );
and ( n23619 , n99 , n23618 , n23602 );
nor ( n23620 , n23617 , n23619 );
nand ( n23621 , n98 , n23606 );
not ( n23622 , n98 );
nand ( n23623 , n99 , n23622 , n23587 );
nand ( n23624 , n23620 , n23621 , n23623 );
nand ( n23625 , n23152 , n23624 );
not ( n23626 , n98 );
nor ( n23627 , n99 , n23626 , n23615 );
not ( n23628 , n23152 );
and ( n23629 , n102 , n98 , n99 );
not ( n23630 , n23629 );
or ( n23631 , n23628 , n23630 );
not ( n23632 , n98 );
nand ( n23633 , n20271 , n23632 , n23539 );
nand ( n23634 , n23631 , n23633 );
nor ( n23635 , n23627 , n23634 );
nand ( n23636 , n100 , n23544 );
not ( n23637 , n23636 );
nand ( n23638 , n23637 , n103 , n98 );
nand ( n23639 , n20271 , n23587 );
nand ( n23640 , n23635 , n23638 , n23639 , n23607 );
nand ( n23641 , n2358 , n23640 );
nand ( n23642 , n23612 , n23625 , n23641 );
nand ( n23643 , n18139 , n23642 );
not ( n23644 , n23569 );
and ( n23645 , n103 , n98 , n23644 );
not ( n23646 , n98 );
and ( n23647 , n103 , n23646 , n23579 );
nor ( n23648 , n23645 , n23647 );
not ( n23649 , n98 );
nand ( n23650 , n23649 , n23589 );
not ( n23651 , n23542 );
nand ( n23652 , n23651 , n98 );
not ( n23653 , n98 );
nor ( n23654 , n23653 , n23636 );
nand ( n23655 , n20271 , n23152 , n104 , n23654 );
and ( n23656 , n23648 , n23650 , n23652 , n23655 );
not ( n23657 , n98 );
nand ( n23658 , n99 , n23657 , n100 , n23239 );
nand ( n23659 , n23658 , n23639 );
and ( n23660 , n23152 , n23659 );
not ( n23661 , n23152 );
and ( n23662 , n22311 , n23551 );
nor ( n23663 , n20271 , n23565 );
and ( n23664 , n98 , n23663 );
nor ( n23665 , n23662 , n23664 );
nor ( n23666 , n98 , n23555 );
and ( n23667 , n99 , n23666 );
nor ( n23668 , n23667 , n23589 );
nand ( n23669 , n23665 , n23668 );
and ( n23670 , n23661 , n23669 );
nor ( n23671 , n23660 , n23670 );
not ( n23672 , n23541 );
nand ( n23673 , n20271 , n23606 );
nor ( n23674 , n20271 , n100 );
nand ( n23675 , n23005 , n98 , n23674 );
nand ( n23676 , n23673 , n23675 );
nand ( n23677 , n23152 , n23676 );
or ( n23678 , n98 , n23636 );
nand ( n23679 , n23678 , n23152 );
not ( n23680 , n23629 );
nand ( n23681 , n103 , n23680 , n23567 );
nand ( n23682 , n23679 , n23681 );
nand ( n23683 , n23672 , n23677 , n2358 , n23682 );
not ( n23684 , n103 );
or ( n23685 , n98 , n23673 );
not ( n23686 , n23663 );
nand ( n23687 , n23685 , n23686 , n23575 );
not ( n23688 , n23687 );
or ( n23689 , n23684 , n23688 );
not ( n23690 , n98 );
or ( n23691 , n20271 , n23690 , n23636 );
not ( n23692 , n98 );
or ( n23693 , n99 , n23692 , n23595 );
nand ( n23694 , n23691 , n23693 );
not ( n23695 , n23674 );
not ( n23696 , n23602 );
and ( n23697 , n23695 , n23696 );
not ( n23698 , n98 );
nand ( n23699 , n23698 , n23152 );
nor ( n23700 , n23697 , n23699 );
nor ( n23701 , n23694 , n2358 , n23700 );
nand ( n23702 , n23689 , n23701 );
nand ( n23703 , n23683 , n23702 );
nand ( n23704 , n23671 , n23703 );
nand ( n23705 , n105 , n23704 );
nand ( n23706 , n23585 , n23643 , n23656 , n23705 );
and ( n23707 , n23706 , n22945 );
not ( n23708 , n23706 );
and ( n23709 , n23708 , n109 );
nor ( n23710 , n23707 , n23709 );
nor ( n23711 , n23537 , n23710 );
not ( n23712 , n23711 );
not ( n23713 , n106 );
nand ( n23714 , n23537 , n23710 );
nand ( n23715 , n23712 , n23713 , n23714 );
nand ( n23716 , n23534 , n23715 );
not ( n23717 , n51 );
not ( n23718 , n22766 );
or ( n23719 , n23717 , n23718 );
or ( n23720 , n51 , n22766 );
nand ( n23721 , n23719 , n23720 );
or ( n23722 , n22771 , n21742 );
or ( n23723 , n53 , n21765 );
nand ( n23724 , n23722 , n23723 );
or ( n23725 , n21882 , n6308 );
not ( n23726 , n22824 );
or ( n23727 , n58 , n23726 );
nand ( n23728 , n23725 , n23727 );
not ( n23729 , n69 );
not ( n23730 , n13617 );
or ( n23731 , n23729 , n23730 );
or ( n23732 , n69 , n13617 );
nand ( n23733 , n23731 , n23732 );
not ( n23734 , n77 );
not ( n23735 , n14467 );
or ( n23736 , n23734 , n23735 );
or ( n23737 , n77 , n14467 );
nand ( n23738 , n23736 , n23737 );
buf ( n23739 , n22802 );
and ( n23740 , n23739 , n81 );
not ( n23741 , n23739 );
and ( n23742 , n23741 , n18511 );
nor ( n23743 , n23740 , n23742 );
not ( n23744 , n65 );
not ( n23745 , n987 );
or ( n23746 , n23744 , n23745 );
or ( n23747 , n65 , n987 );
nand ( n23748 , n23746 , n23747 );
not ( n23749 , n86 );
not ( n23750 , n14210 );
or ( n23751 , n23749 , n23750 );
or ( n23752 , n86 , n22791 );
nand ( n23753 , n23751 , n23752 );
not ( n23754 , n106 );
not ( n23755 , n108 );
or ( n23756 , n23754 , n23755 );
and ( n23757 , n18 , n22945 );
and ( n23758 , n109 , n21045 );
nor ( n23759 , n23757 , n23758 );
not ( n23760 , n23706 );
or ( n23761 , n23759 , n23760 );
not ( n23762 , n23759 );
not ( n23763 , n23760 );
or ( n23764 , n23762 , n23763 );
nand ( n23765 , n23764 , n23713 );
not ( n23766 , n23765 );
nand ( n23767 , n23761 , n23766 );
nand ( n23768 , n23756 , n23767 );
not ( n23769 , n106 );
not ( n23770 , n227 );
or ( n23771 , n23769 , n23770 );
and ( n23772 , n109 , n21971 );
and ( n23773 , n110 , n22945 );
nor ( n23774 , n23772 , n23773 );
and ( n23775 , n18 , n19465 );
and ( n23776 , n223 , n21045 );
nor ( n23777 , n23775 , n23776 );
xnor ( n23778 , n23774 , n23777 );
or ( n23779 , n23778 , n23760 );
not ( n23780 , n23778 );
not ( n23781 , n23760 );
or ( n23782 , n23780 , n23781 );
nand ( n23783 , n23782 , n23713 );
not ( n23784 , n23783 );
nand ( n23785 , n23779 , n23784 );
nand ( n23786 , n23771 , n23785 );
not ( n23787 , n75 );
buf ( n23788 , n14594 );
not ( n23789 , n23788 );
or ( n23790 , n23787 , n23789 );
or ( n23791 , n75 , n23788 );
nand ( n23792 , n23790 , n23791 );
not ( n23793 , n59 );
not ( n23794 , n1758 );
or ( n23795 , n23793 , n23794 );
or ( n23796 , n59 , n1758 );
nand ( n23797 , n23795 , n23796 );
not ( n23798 , n41 );
buf ( n23799 , n13730 );
not ( n23800 , n23799 );
or ( n23801 , n23798 , n23800 );
or ( n23802 , n41 , n23799 );
nand ( n23803 , n23801 , n23802 );
and ( n23804 , n22748 , n14091 );
not ( n23805 , n22748 );
and ( n23806 , n23805 , n78 );
nor ( n23807 , n23804 , n23806 );
not ( n23808 , n106 );
not ( n23809 , n107 );
or ( n23810 , n23808 , n23809 );
or ( n23811 , n21045 , n23760 );
or ( n23812 , n18 , n23706 );
nand ( n23813 , n23811 , n23812 , n23713 );
nand ( n23814 , n23810 , n23813 );
not ( n23815 , n71 );
not ( n23816 , n21027 );
or ( n23817 , n23815 , n23816 );
or ( n23818 , n71 , n21027 );
nand ( n23819 , n23817 , n23818 );
not ( n23820 , n48 );
not ( n23821 , n21250 );
or ( n23822 , n23820 , n23821 );
or ( n23823 , n48 , n21492 );
nand ( n23824 , n23822 , n23823 );
not ( n23825 , n80 );
not ( n23826 , n13718 );
or ( n23827 , n23825 , n23826 );
or ( n23828 , n80 , n13718 );
nand ( n23829 , n23827 , n23828 );
not ( n23830 , n63 );
not ( n23831 , n9084 );
or ( n23832 , n23830 , n23831 );
or ( n23833 , n63 , n9084 );
nand ( n23834 , n23832 , n23833 );
not ( n23835 , n18 );
not ( n23836 , n21756 );
or ( n23837 , n23835 , n23836 );
or ( n23838 , n18 , n21756 );
nand ( n23839 , n23837 , n23838 );
not ( n23840 , n84 );
not ( n23841 , n14057 );
or ( n23842 , n23840 , n23841 );
or ( n23843 , n84 , n14057 );
nand ( n23844 , n23842 , n23843 );
nand ( n23845 , n401 , n434 );
xor ( n23846 , n439 , n23845 );
nor ( n23847 , n106 , n23846 );
xnor ( n23848 , n401 , n434 );
nor ( n23849 , n106 , n23848 );
not ( n23850 , n106 );
not ( n23851 , n423 );
or ( n23852 , n23850 , n23851 );
or ( n23853 , n22382 , n106 );
nand ( n23854 , n23852 , n23853 );
and ( n23855 , n106 , n428 );
not ( n23856 , n106 );
and ( n23857 , n23856 , n62 );
or ( n23858 , n23855 , n23857 );
and ( n23859 , n106 , n404 );
not ( n23860 , n106 );
and ( n23861 , n23860 , n341 );
or ( n23862 , n23859 , n23861 );
and ( n23863 , n106 , n394 );
not ( n23864 , n106 );
and ( n23865 , n23864 , n345 );
or ( n23866 , n23863 , n23865 );
and ( n23867 , n106 , n413 );
not ( n23868 , n106 );
and ( n23869 , n23868 , n263 );
or ( n23870 , n23867 , n23869 );
and ( n23871 , n106 , n431 );
not ( n23872 , n106 );
and ( n23873 , n23872 , n391 );
or ( n23874 , n23871 , n23873 );
and ( n23875 , n106 , n450 );
not ( n23876 , n106 );
and ( n23877 , n23876 , n268 );
or ( n23878 , n23875 , n23877 );
and ( n23879 , n106 , n440 );
not ( n23880 , n106 );
and ( n23881 , n23880 , n325 );
or ( n23882 , n23879 , n23881 );
and ( n23883 , n106 , n406 );
not ( n23884 , n106 );
and ( n23885 , n23884 , n226 );
or ( n23886 , n23883 , n23885 );
and ( n23887 , n106 , n444 );
not ( n23888 , n106 );
and ( n23889 , n23888 , n222 );
or ( n23890 , n23887 , n23889 );
and ( n23891 , n106 , n407 );
not ( n23892 , n106 );
and ( n23893 , n23892 , n216 );
or ( n23894 , n23891 , n23893 );
and ( n23895 , n106 , n429 );
not ( n23896 , n106 );
and ( n23897 , n23896 , n50 );
or ( n23898 , n23895 , n23897 );
and ( n23899 , n106 , n418 );
not ( n23900 , n106 );
and ( n23901 , n23900 , n347 );
or ( n23902 , n23899 , n23901 );
and ( n23903 , n106 , n445 );
not ( n23904 , n106 );
and ( n23905 , n23904 , n285 );
or ( n23906 , n23903 , n23905 );
and ( n23907 , n106 , n415 );
not ( n23908 , n106 );
and ( n23909 , n23908 , n89 );
or ( n23910 , n23907 , n23909 );
and ( n23911 , n106 , n416 );
not ( n23912 , n106 );
and ( n23913 , n23912 , n92 );
or ( n23914 , n23911 , n23913 );
and ( n23915 , n106 , n446 );
not ( n23916 , n106 );
and ( n23917 , n23916 , n329 );
or ( n23918 , n23915 , n23917 );
and ( n23919 , n106 , n396 );
not ( n23920 , n106 );
and ( n23921 , n23920 , n374 );
or ( n23922 , n23919 , n23921 );
and ( n23923 , n106 , n402 );
not ( n23924 , n106 );
and ( n23925 , n23924 , n52 );
or ( n23926 , n23923 , n23925 );
and ( n23927 , n106 , n405 );
not ( n23928 , n106 );
and ( n23929 , n23928 , n312 );
or ( n23930 , n23927 , n23929 );
and ( n23931 , n106 , n399 );
not ( n23932 , n106 );
and ( n23933 , n23932 , n370 );
or ( n23934 , n23931 , n23933 );
and ( n23935 , n106 , n397 );
not ( n23936 , n106 );
and ( n23937 , n23936 , n372 );
or ( n23938 , n23935 , n23937 );
and ( n23939 , n106 , n398 );
not ( n23940 , n106 );
and ( n23941 , n23940 , n224 );
or ( n23942 , n23939 , n23941 );
and ( n23943 , n106 , n427 );
not ( n23944 , n106 );
and ( n23945 , n23944 , n377 );
or ( n23946 , n23943 , n23945 );
and ( n23947 , n106 , n412 );
not ( n23948 , n106 );
and ( n23949 , n23948 , n70 );
or ( n23950 , n23947 , n23949 );
and ( n23951 , n106 , n424 );
not ( n23952 , n106 );
and ( n23953 , n23952 , n281 );
or ( n23954 , n23951 , n23953 );
and ( n23955 , n106 , n432 );
not ( n23956 , n106 );
and ( n23957 , n23956 , n266 );
or ( n23958 , n23955 , n23957 );
and ( n23959 , n106 , n414 );
not ( n23960 , n106 );
and ( n23961 , n23960 , n64 );
or ( n23962 , n23959 , n23961 );
and ( n23963 , n106 , n435 );
not ( n23964 , n106 );
and ( n23965 , n23964 , n259 );
or ( n23966 , n23963 , n23965 );
and ( n23967 , n106 , n437 );
not ( n23968 , n106 );
and ( n23969 , n23968 , n302 );
or ( n23970 , n23967 , n23969 );
and ( n23971 , n106 , n443 );
not ( n23972 , n106 );
and ( n23973 , n23972 , n97 );
or ( n23974 , n23971 , n23973 );
and ( n23975 , n106 , n426 );
not ( n23976 , n106 );
and ( n23977 , n23976 , n335 );
or ( n23978 , n23975 , n23977 );
and ( n23979 , n106 , n425 );
not ( n23980 , n106 );
and ( n23981 , n23980 , n91 );
or ( n23982 , n23979 , n23981 );
and ( n23983 , n106 , n442 );
not ( n23984 , n106 );
and ( n23985 , n23984 , n289 );
or ( n23986 , n23983 , n23985 );
and ( n23987 , n106 , n400 );
not ( n23988 , n106 );
and ( n23989 , n23988 , n360 );
or ( n23990 , n23987 , n23989 );
and ( n23991 , n106 , n436 );
not ( n23992 , n106 );
and ( n23993 , n23992 , n379 );
or ( n23994 , n23991 , n23993 );
and ( n23995 , n106 , n403 );
not ( n23996 , n106 );
and ( n23997 , n23996 , n57 );
or ( n23998 , n23995 , n23997 );
and ( n23999 , n106 , n419 );
not ( n24000 , n106 );
and ( n24001 , n24000 , n323 );
or ( n24002 , n23999 , n24001 );
and ( n24003 , n106 , n348 );
not ( n24004 , n106 );
and ( n24005 , n24004 , n35 );
or ( n24006 , n24003 , n24005 );
and ( n24007 , n106 , n408 );
not ( n24008 , n106 );
and ( n24009 , n24008 , n76 );
or ( n24010 , n24007 , n24009 );
and ( n24011 , n106 , n410 );
not ( n24012 , n106 );
and ( n24013 , n24012 , n47 );
or ( n24014 , n24011 , n24013 );
and ( n24015 , n106 , n409 );
not ( n24016 , n106 );
and ( n24017 , n24016 , n310 );
or ( n24018 , n24015 , n24017 );
and ( n24019 , n106 , n411 );
not ( n24020 , n106 );
and ( n24021 , n24020 , n44 );
or ( n24022 , n24019 , n24021 );
and ( n24023 , n106 , n393 );
not ( n24024 , n106 );
and ( n24025 , n24024 , n237 );
or ( n24026 , n24023 , n24025 );
and ( n24027 , n106 , n441 );
not ( n24028 , n106 );
and ( n24029 , n24028 , n233 );
or ( n24030 , n24027 , n24029 );
and ( n24031 , n106 , n433 );
not ( n24032 , n106 );
and ( n24033 , n24032 , n54 );
or ( n24034 , n24031 , n24033 );
and ( n24035 , n106 , n448 );
not ( n24036 , n106 );
and ( n24037 , n24036 , n362 );
or ( n24038 , n24035 , n24037 );
and ( n24039 , n106 , n417 );
not ( n24040 , n106 );
and ( n24041 , n24040 , n145 );
or ( n24042 , n24039 , n24041 );
and ( n24043 , n106 , n438 );
not ( n24044 , n106 );
and ( n24045 , n24044 , n337 );
or ( n24046 , n24043 , n24045 );
and ( n24047 , n106 , n420 );
not ( n24048 , n106 );
and ( n24049 , n24048 , n60 );
or ( n24050 , n24047 , n24049 );
and ( n24051 , n106 , n430 );
not ( n24052 , n106 );
and ( n24053 , n24052 , n275 );
or ( n24054 , n24051 , n24053 );
and ( n24055 , n106 , n395 );
not ( n24056 , n106 );
and ( n24057 , n24056 , n231 );
or ( n24058 , n24055 , n24057 );
and ( n24059 , n106 , n422 );
not ( n24060 , n106 );
and ( n24061 , n24060 , n356 );
or ( n24062 , n24059 , n24061 );
and ( n24063 , n106 , n421 );
not ( n24064 , n106 );
and ( n24065 , n24064 , n87 );
or ( n24066 , n24063 , n24065 );
and ( n24067 , n106 , n447 );
not ( n24068 , n106 );
and ( n24069 , n24068 , n247 );
or ( n24070 , n24067 , n24069 );
and ( n24071 , n106 , n449 );
not ( n24072 , n106 );
and ( n24073 , n24072 , n88 );
or ( n24074 , n24071 , n24073 );
nor ( n24075 , n106 , n401 );
endmodule
