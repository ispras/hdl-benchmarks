//NOTE: no-implementation module stub

module DEC (
    input T_RST,
    input DSPCLK,
    input [23:0] CM_rd,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input PPclr_h,
    input GO_D,
    input GO_Ex,
    input GO_Cx,
    input Prderr_Eg,
    input ICE_ST,
    input redoSTI_h,
    input [7:0] ASTAT,
    input Ctrue,
    input Upd_IR,
    input [23:0] SPC,
    input SBP_EN,
    input enTYP3,
    input [23:0] IR,
    input [19:0] IRE,
    input EX_en,
    input EX_enc,
    input Dummy_E,
    input Dummy_R,
    input DU_R,
    input dBR_R,
    input idBR_R,
    input RET_R,
    input RTS_R,
    input EXIT_E,
    input DU_Eg,
    input Call_Ed,
    input RTI_Ed,
    input RTS_Ed,
    input BR_Ed,
    input RET_Ed,
    input Nseq_Ed,
    input IDLE_Eg,
    input MACdep_Eg,
    input MTCNTR_Eg,
    input MTOWRCNTR_Eg,
    input MTtoppcs_Eg,
    input MTIMASK_Eg,
    input MTICNTL_Eg,
    input MTIFC_Eg,
    input MTMSTAT_Eg,
    input MFPSQ_E,
    input MFtoppcs_E,
    input MFIMASK_E,
    input MFICNTL_E,
    input MFSSTAT_E,
    input MFMSTAT_E,
    input MFCNTR_E,
    input Stkctl_Eg,
    input Modctl_Eg,
    input MpopLP_Eg,
    input imm16_E,
    input imm14_E,
    input Long_Eg,
    input Nrti_Ed,
    input [3:0] ALUop_E,
    input cdAM_E,
    input [7:0] MTAX0_E,
    input [7:0] MTAX1_E,
    input [7:0] MTAY0_E,
    input [7:0] MTAY1_E,
    input [7:0] MTAR_E,
    input [7:0] MTASTAT_E,
    input [7:0] MFAX0_E,
    input [7:0] MFAX1_E,
    input [7:0] MFAY0_E,
    input [7:0] MFAY1_E,
    input [7:0] MFAR_E,
    input [7:0] MFASTAT_E,
    input [7:0] MFALU_E,
    input pMFALU_E,
    input [7:0] DIVQ_E,
    input [7:0] DIVS_E,
    input updAR_E,
    input updAF_E,
    input [3:0] ALUop_R,
    input type9,
    input [7:0] DIVQ_R,
    input [7:0] DIVS_R,
    input MACop_E,
    input satMR_Eg,
    input Rbyp_Rg,
    input Xbyp_Rg,
    input Ybyp_Rg,
    input [7:0] MTMX0_Eg,
    input [7:0] MTMX1_Eg,
    input [7:0] MTMY0_Eg,
    input [7:0] MTMY1_Eg,
    input [7:0] MTMR0_Eg,
    input [7:0] MTMR1_Eg,
    input [7:0] MTMR2_Eg,
    input [7:0] MFMX0_E,
    input [7:0] MFMX1_E,
    input [7:0] MFMY0_E,
    input [7:0] MFMY1_E,
    input [7:0] MFMR0_E,
    input [7:0] MFMR1_E,
    input [7:0] MFMR2_E,
    input MFMAC_E,
    input pMFMAC_E,
    input updMR_E,
    input updMF_E,
    input Squ_Rx,
    input MACop_R,
    input [7:0] SHTop_E,
    input imSHT_E,
    input MTSI_E,
    input MTSE_E,
    input MTSR0_E,
    input MTSR1_E,
    input MTSB_E,
    input MFSI_E,
    input MFSE_E,
    input MFSR0_E,
    input MFSR1_E,
    input MFSB_E,
    input MFSHT_E,
    input pMFSHT_E,
    input updSR0_Eg,
    input updSR1_Eg,
    input updSR_E,
    input [7:0] MTIreg_E,
    input [7:0] MTLreg_E,
    input [7:0] MTMreg_E,
    input [7:0] MFIreg_E,
    input [7:0] MFLreg_E,
    input [7:0] MFMreg_E,
    input MFDAG1_E,
    input MFDAG2_E,
    input accPM_E,
    input Double_R,
    input Double_E,
    input Post1_E,
    input Post2_E,
    input DAG1D_R,
    input DAG2D_R,
    input imAddr_R,
    input DAG1_EN,
    input DAG2_EN,
    input DAG2P_R,
    input DMAen_R,
    input Pread_R,
    input Pwrite_R,
    input Dread_R,
    input Dwrite_R,
    input IOcmd_R,
    input IOread_R,
    input IOwrite_R,
    input IDLE_R,
    input MTPMOVL_E,
    input MTDMOVL_E,
    input MFPMOVL_E,
    input MFDMOVL_E,
    input MFSPT_E,
    input MFRX0_E,
    input MFTX0_E,
    input MFRX1_E,
    input MFTX1_E,
    input MTRX0_E,
    input MTTX0_E,
    input MTRX1_E,
    input MTTX1_E,
    input SBP_R,
    input MFIDR_E,
    input MTIDR_Eg,
    input nNOP_Eg,
    input accCM_R,
    input accCM_E,
    input wrCM_R,
    input rdCM_E
);

endmodule
