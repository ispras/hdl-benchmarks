module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 ;
wire n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n320434 , n320435 , n320436 , n320437 , n320438 , n320439 , n320440 , n320441 , n320442 , 
 n320443 , n320444 , n320445 , n320446 , n320447 , n320448 , n320449 , n320450 , n320451 , n320452 , 
 n320453 , n320454 , n320455 , n320456 , n320457 , n320458 , n320459 , n320460 , n320461 , n320462 , 
 n320463 , n320464 , n320465 , n320466 , n320467 , n320468 , n320469 , n320470 , n320471 , n320472 , 
 n320473 , n320474 , n320475 , n320476 , n320477 , n320478 , n320479 , n320480 , n320481 , n320482 , 
 n320483 , n320484 , n320485 , n320486 , n320487 , n320488 , n320489 , n320490 , n320491 , n320492 , 
 n320493 , n320494 , n320495 , n320496 , n320497 , n320498 , n320499 , n320500 , n320501 , n320502 , 
 n320503 , n320504 , n320505 , n320506 , n320507 , n320508 , n320509 , n320510 , n320511 , n320512 , 
 n320513 , n320514 , n320515 , n320516 , n320517 , n320518 , n320519 , n320520 , n320521 , n320522 , 
 n320523 , n320524 , n320525 , n320526 , n320527 , n320528 , n320529 , n320530 , n320531 , n320532 , 
 n320533 , n320534 , n320535 , n320536 , n320537 , n320538 , n320539 , n320540 , n320541 , n320542 , 
 n320543 , n320544 , n320545 , n320546 , n320547 , n320548 , n320549 , n320550 , n320551 , n320552 , 
 n320553 , n320554 , n320555 , n320556 , n320557 , n320558 , n320559 , n320560 , n320561 , n823 , 
 n320563 , n825 , n320565 , n320566 , n320567 , n829 , n320569 , n320570 , n832 , n833 , 
 n320573 , n835 , n320575 , n320576 , n838 , n320578 , n320579 , n841 , n320581 , n843 , 
 n320583 , n320584 , n320585 , n320586 , n320587 , n320588 , n320589 , n320590 , n320591 , n320592 , 
 n320593 , n855 , n320595 , n320596 , n858 , n320598 , n860 , n320600 , n320601 , n863 , 
 n320603 , n320604 , n320605 , n320606 , n320607 , n320608 , n320609 , n320610 , n320611 , n873 , 
 n320613 , n875 , n876 , n320616 , n320617 , n879 , n320619 , n320620 , n320621 , n883 , 
 n320623 , n320624 , n886 , n320626 , n320627 , n320628 , n890 , n891 , n892 , n893 , 
 n320633 , n895 , n320635 , n320636 , n898 , n320638 , n900 , n320640 , n902 , n320642 , 
 n320643 , n320644 , n320645 , n320646 , n320647 , n320648 , n320649 , n320650 , n320651 , n320652 , 
 n320653 , n320654 , n320655 , n320656 , n320657 , n320658 , n320659 , n921 , n320661 , n923 , 
 n320663 , n320664 , n926 , n320666 , n928 , n929 , n320669 , n320670 , n320671 , n933 , 
 n320673 , n320674 , n320675 , n320676 , n320677 , n320678 , n320679 , n320680 , n320681 , n320682 , 
 n944 , n320684 , n320685 , n947 , n320687 , n320688 , n320689 , n320690 , n320691 , n320692 , 
 n320693 , n320694 , n320695 , n320696 , n320697 , n959 , n320699 , n320700 , n320701 , n320702 , 
 n320703 , n320704 , n320705 , n320706 , n320707 , n320708 , n970 , n971 , n320711 , n973 , 
 n320713 , n320714 , n976 , n320716 , n320717 , n320718 , n320719 , n320720 , n320721 , n983 , 
 n320723 , n320724 , n320725 , n987 , n320727 , n320728 , n320729 , n991 , n992 , n320732 , 
 n320733 , n995 , n320735 , n320736 , n998 , n320738 , n320739 , n320740 , n320741 , n1003 , 
 n320743 , n320744 , n320745 , n320746 , n320747 , n320748 , n320749 , n320750 , n320751 , n320752 , 
 n320753 , n320754 , n320755 , n1017 , n320757 , n1019 , n1020 , n320760 , n320761 , n1023 , 
 n1024 , n1025 , n1026 , n320766 , n320767 , n1029 , n320769 , n1031 , n320771 , n1033 , 
 n1034 , n320774 , n1036 , n320776 , n320777 , n320778 , n320779 , n1041 , n320781 , n320782 , 
 n320783 , n320784 , n1046 , n320786 , n320787 , n320788 , n320789 , n320790 , n320791 , n1053 , 
 n320793 , n320794 , n320795 , n320796 , n320797 , n320798 , n320799 , n320800 , n1062 , n320802 , 
 n320803 , n320804 , n320805 , n320806 , n320807 , n320808 , n1070 , n1071 , n1072 , n320812 , 
 n320813 , n320814 , n320815 , n1077 , n1078 , n1079 , n320819 , n1081 , n1082 , n320822 , 
 n1084 , n320824 , n1086 , n320826 , n1088 , n1089 , n1090 , n320830 , n320831 , n1093 , 
 n1094 , n1095 , n1096 , n1097 , n320837 , n320838 , n320839 , n1101 , n320841 , n320842 , 
 n1104 , n1105 , n320845 , n1107 , n320847 , n320848 , n320849 , n320850 , n1112 , n320852 , 
 n320853 , n320854 , n320855 , n320856 , n320857 , n320858 , n320859 , n320860 , n320861 , n320862 , 
 n320863 , n320864 , n320865 , n320866 , n320867 , n320868 , n1130 , n320870 , n320871 , n320872 , 
 n1134 , n320874 , n320875 , n1137 , n320877 , n320878 , n320879 , n1141 , n320881 , n320882 , 
 n320883 , n1145 , n320885 , n320886 , n320887 , n1149 , n320889 , n1151 , n320891 , n320892 , 
 n1154 , n320894 , n320895 , n1157 , n320897 , n320898 , n1160 , n1161 , n320901 , n320902 , 
 n320903 , n320904 , n320905 , n320906 , n1168 , n320908 , n1170 , n320910 , n320911 , n320912 , 
 n320913 , n1175 , n320915 , n320916 , n320917 , n1179 , n320919 , n1181 , n320921 , n320922 , 
 n320923 , n320924 , n320925 , n320926 , n320927 , n320928 , n320929 , n320930 , n320931 , n320932 , 
 n320933 , n1195 , n320935 , n1197 , n1198 , n1199 , n1200 , n320940 , n320941 , n320942 , 
 n1204 , n320944 , n320945 , n320946 , n320947 , n320948 , n320949 , n1211 , n320951 , n320952 , 
 n1214 , n1215 , n1216 , n320956 , n320957 , n1219 , n1220 , n1221 , n320961 , n320962 , 
 n320963 , n320964 , n1226 , n320966 , n320967 , n1229 , n320969 , n320970 , n1232 , n320972 , 
 n1234 , n320974 , n320975 , n320976 , n320977 , n320978 , n320979 , n320980 , n1242 , n1243 , 
 n320983 , n320984 , n1246 , n320986 , n320987 , n1249 , n320989 , n320990 , n1252 , n320992 , 
 n320993 , n320994 , n320995 , n1257 , n320997 , n320998 , n1260 , n321000 , n1262 , n1263 , 
 n321003 , n321004 , n321005 , n321006 , n321007 , n1269 , n321009 , n321010 , n321011 , n321012 , 
 n321013 , n321014 , n321015 , n321016 , n321017 , n1279 , n321019 , n1281 , n321021 , n321022 , 
 n1284 , n321024 , n1286 , n321026 , n321027 , n321028 , n1290 , n1291 , n321031 , n321032 , 
 n1294 , n321034 , n321035 , n321036 , n321037 , n321038 , n321039 , n1301 , n1302 , n1303 , 
 n321043 , n1305 , n321045 , n1307 , n321047 , n321048 , n321049 , n321050 , n1312 , n321052 , 
 n1314 , n1315 , n1316 , n321056 , n1318 , n321058 , n321059 , n321060 , n321061 , n321062 , 
 n321063 , n321064 , n1326 , n321066 , n1328 , n321068 , n321069 , n321070 , n1332 , n321072 , 
 n321073 , n1335 , n321075 , n1337 , n1338 , n1339 , n321079 , n321080 , n321081 , n321082 , 
 n321083 , n321084 , n1346 , n321086 , n321087 , n1349 , n321089 , n321090 , n1352 , n321092 , 
 n1354 , n321094 , n321095 , n321096 , n321097 , n321098 , n1360 , n321100 , n321101 , n1363 , 
 n1364 , n321104 , n321105 , n1367 , n321107 , n321108 , n1370 , n321110 , n321111 , n1373 , 
 n1374 , n321114 , n1376 , n321116 , n1378 , n1379 , n321119 , n321120 , n321121 , n321122 , 
 n321123 , n321124 , n1386 , n321126 , n321127 , n321128 , n1390 , n321130 , n321131 , n321132 , 
 n321133 , n321134 , n1396 , n321136 , n1398 , n1399 , n321139 , n321140 , n321141 , n321142 , 
 n321143 , n321144 , n321145 , n1407 , n321147 , n321148 , n321149 , n1411 , n321151 , n321152 , 
 n321153 , n321154 , n321155 , n1417 , n321157 , n321158 , n1420 , n1421 , n321161 , n321162 , 
 n321163 , n321164 , n321165 , n321166 , n321167 , n321168 , n1430 , n321170 , n321171 , n1433 , 
 n321173 , n321174 , n1436 , n321176 , n321177 , n321178 , n1440 , n1441 , n321181 , n1443 , 
 n321183 , n321184 , n321185 , n321186 , n1448 , n321188 , n321189 , n1451 , n321191 , n321192 , 
 n1454 , n321194 , n321195 , n1457 , n321197 , n321198 , n321199 , n321200 , n1462 , n321202 , 
 n321203 , n321204 , n1466 , n321206 , n321207 , n1469 , n321209 , n1471 , n1472 , n1473 , 
 n1474 , n1475 , n321215 , n321216 , n321217 , n321218 , n321219 , n321220 , n321221 , n321222 , 
 n1484 , n321224 , n321225 , n1487 , n321227 , n1489 , n321229 , n321230 , n321231 , n321232 , 
 n1494 , n1495 , n321235 , n321236 , n321237 , n321238 , n321239 , n1501 , n1502 , n321242 , 
 n1504 , n321244 , n321245 , n321246 , n321247 , n321248 , n321249 , n321250 , n321251 , n321252 , 
 n321253 , n321254 , n1516 , n321256 , n1518 , n321258 , n321259 , n321260 , n321261 , n321262 , 
 n321263 , n321264 , n321265 , n321266 , n321267 , n321268 , n1530 , n1531 , n321271 , n1533 , 
 n321273 , n321274 , n321275 , n321276 , n321277 , n321278 , n321279 , n1541 , n1542 , n1543 , 
 n1544 , n1545 , n321285 , n321286 , n1548 , n321288 , n321289 , n321290 , n321291 , n321292 , 
 n1554 , n321294 , n321295 , n1557 , n1558 , n321298 , n1560 , n321300 , n321301 , n321302 , 
 n321303 , n321304 , n321305 , n1567 , n1568 , n1569 , n321309 , n321310 , n321311 , n321312 , 
 n1574 , n321314 , n1576 , n1577 , n321317 , n321318 , n1580 , n321320 , n321321 , n321322 , 
 n321323 , n321324 , n321325 , n321326 , n1588 , n321328 , n321329 , n321330 , n321331 , n321332 , 
 n321333 , n1595 , n321335 , n321336 , n321337 , n321338 , n1600 , n321340 , n321341 , n1603 , 
 n321343 , n321344 , n1606 , n321346 , n321347 , n1609 , n321349 , n1611 , n321351 , n321352 , 
 n321353 , n1615 , n1616 , n321356 , n1618 , n321358 , n321359 , n1621 , n1622 , n321362 , 
 n321363 , n321364 , n1626 , n1627 , n321367 , n1629 , n321369 , n321370 , n1632 , n1633 , 
 n321373 , n321374 , n1636 , n321376 , n321377 , n1639 , n1640 , n321380 , n1642 , n321382 , 
 n1644 , n321384 , n321385 , n1647 , n321387 , n1649 , n1650 , n1651 , n321391 , n321392 , 
 n1654 , n321394 , n1656 , n1657 , n1658 , n321398 , n1660 , n321400 , n321401 , n1663 , 
 n321403 , n1665 , n321405 , n321406 , n1668 , n1669 , n321409 , n321410 , n1672 , n321412 , 
 n321413 , n1675 , n321415 , n321416 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , 
 n321423 , n1685 , n1686 , n321426 , n321427 , n1689 , n321429 , n321430 , n1692 , n321432 , 
 n1694 , n321434 , n321435 , n1697 , n321437 , n1699 , n1700 , n1701 , n1702 , n1703 , 
 n1704 , n1705 , n1706 , n1707 , n321447 , n1709 , n321449 , n1711 , n321451 , n321452 , 
 n1714 , n321454 , n321455 , n321456 , n1718 , n321458 , n321459 , n321460 , n321461 , n1723 , 
 n321463 , n321464 , n321465 , n1727 , n321467 , n321468 , n1730 , n321470 , n1732 , n1733 , 
 n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n321480 , n321481 , n1743 , 
 n321483 , n1745 , n1746 , n1747 , n1748 , n321488 , n1750 , n321490 , n321491 , n321492 , 
 n1754 , n321494 , n321495 , n321496 , n321497 , n1759 , n321499 , n321500 , n1762 , n321502 , 
 n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , 
 n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n321520 , n1782 , n321522 , 
 n321523 , n1785 , n321525 , n321526 , n1788 , n321528 , n1790 , n321530 , n1792 , n321532 , 
 n321533 , n1795 , n321535 , n1797 , n1798 , n1799 , n321539 , n1801 , n321541 , n321542 , 
 n321543 , n1805 , n321545 , n1807 , n321547 , n1809 , n321549 , n321550 , n321551 , n1813 , 
 n321553 , n321554 , n1816 , n321556 , n1818 , n1819 , n1820 , n1821 , n321561 , n1823 , 
 n321563 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , 
 n1834 , n1835 , n321575 , n321576 , n1838 , n321578 , n321579 , n1841 , n1842 , n1843 , 
 n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n321590 , n1852 , n321592 , 
 n321593 , n1855 , n1856 , n1857 , n321597 , n321598 , n321599 , n1861 , n321601 , n321602 , 
 n1864 , n321604 , n321605 , n1867 , n321607 , n321608 , n321609 , n321610 , n1872 , n321612 , 
 n321613 , n1875 , n321615 , n1877 , n1878 , n321618 , n321619 , n321620 , n1882 , n321622 , 
 n321623 , n1885 , n321625 , n321626 , n1888 , n321628 , n321629 , n1891 , n321631 , n321632 , 
 n1894 , n321634 , n321635 , n321636 , n321637 , n321638 , n321639 , n321640 , n321641 , n321642 , 
 n321643 , n321644 , n321645 , n321646 , n321647 , n321648 , n321649 , n321650 , n321651 , n321652 , 
 n321653 , n321654 , n321655 , n321656 , n321657 , n321658 , n321659 , n321660 , n321661 , n321662 , 
 n321663 , n321664 , n321665 , n321666 , n321667 , n321668 , n321669 , n321670 , n321671 , n321672 , 
 n321673 , n321674 , n321675 , n321676 , n1900 , n321678 , n321679 , n321680 , n321681 , n321682 , 
 n321683 , n321684 , n321685 , n321686 , n1910 , n321688 , n1912 , n1913 , n321691 , n1914 , 
 n321693 , n321694 , n321695 , n321696 , n321697 , n321698 , n321699 , n321700 , n321701 , n321702 , 
 n321703 , n321704 , n321705 , n321706 , n321707 , n321708 , n321709 , n321710 , n1929 , n1930 , 
 n1931 , n1932 , n321715 , n1934 , n1935 , n321718 , n1937 , n321720 , n321721 , n1940 , 
 n1941 , n321724 , n1943 , n321726 , n1945 , n321728 , n1947 , n1948 , n321731 , n321732 , 
 n321733 , n1952 , n321735 , n321736 , n1955 , n321738 , n321739 , n1958 , n321741 , n1960 , 
 n1961 , n1962 , n321745 , n321746 , n1965 , n321748 , n1967 , n321750 , n321751 , n1970 , 
 n321753 , n1972 , n321755 , n321756 , n1975 , n1976 , n321759 , n321760 , n321761 , n321762 , 
 n321763 , n321764 , n1983 , n321766 , n321767 , n321768 , n321769 , n321770 , n321771 , n321772 , 
 n321773 , n321774 , n321775 , n321776 , n321777 , n1996 , n1997 , n321780 , n1999 , n2000 , 
 n321783 , n2002 , n321785 , n2004 , n321787 , n2006 , n2007 , n321790 , n2009 , n2010 , 
 n2011 , n2012 , n321795 , n321796 , n321797 , n321798 , n2017 , n321800 , n321801 , n2020 , 
 n321803 , n2022 , n321805 , n321806 , n321807 , n321808 , n321809 , n321810 , n321811 , n321812 , 
 n321813 , n321814 , n321815 , n321816 , n321817 , n2036 , n2037 , n321820 , n2039 , n321822 , 
 n321823 , n2042 , n2043 , n321826 , n2045 , n321828 , n321829 , n321830 , n321831 , n321832 , 
 n321833 , n321834 , n321835 , n321836 , n321837 , n2056 , n321839 , n321840 , n2059 , n321842 , 
 n321843 , n321844 , n2063 , n321846 , n321847 , n2066 , n321849 , n321850 , n321851 , n321852 , 
 n321853 , n321854 , n2073 , n321856 , n321857 , n321858 , n321859 , n321860 , n321861 , n321862 , 
 n321863 , n321864 , n321865 , n321866 , n2085 , n2086 , n321869 , n321870 , n2089 , n321872 , 
 n321873 , n321874 , n2093 , n321876 , n2095 , n321878 , n321879 , n321880 , n2099 , n321882 , 
 n321883 , n2102 , n321885 , n2104 , n2105 , n2106 , n321889 , n321890 , n321891 , n321892 , 
 n2111 , n321894 , n2113 , n321896 , n321897 , n2116 , n321899 , n321900 , n2119 , n2120 , 
 n321903 , n2122 , n2123 , n321906 , n321907 , n321908 , n321909 , n321910 , n321911 , n321912 , 
 n321913 , n321914 , n321915 , n321916 , n321917 , n321918 , n321919 , n321920 , n321921 , n321922 , 
 n321923 , n2142 , n321925 , n321926 , n321927 , n321928 , n2147 , n321930 , n321931 , n2150 , 
 n321933 , n321934 , n321935 , n321936 , n321937 , n321938 , n2157 , n321940 , n321941 , n2160 , 
 n321943 , n321944 , n321945 , n321946 , n321947 , n321948 , n321949 , n321950 , n2169 , n321952 , 
 n321953 , n321954 , n321955 , n321956 , n321957 , n2176 , n321959 , n2178 , n321961 , n2180 , 
 n321963 , n2182 , n2183 , n321966 , n321967 , n321968 , n321969 , n321970 , n321971 , n321972 , 
 n321973 , n321974 , n2193 , n321976 , n2195 , n321978 , n321979 , n2198 , n321981 , n321982 , 
 n321983 , n321984 , n321985 , n321986 , n321987 , n321988 , n321989 , n321990 , n2209 , n321992 , 
 n321993 , n321994 , n321995 , n2214 , n321997 , n2216 , n321999 , n322000 , n2219 , n2220 , 
 n322003 , n322004 , n2223 , n2224 , n322007 , n2226 , n322009 , n2228 , n322011 , n2230 , 
 n322013 , n2232 , n2233 , n322016 , n322017 , n2236 , n322019 , n322020 , n2239 , n322022 , 
 n322023 , n2242 , n322025 , n322026 , n2245 , n2246 , n322029 , n2248 , n2249 , n2250 , 
 n2251 , n2252 , n2253 , n2254 , n322037 , n2256 , n2257 , n322040 , n2259 , n322042 , 
 n2261 , n2262 , n322045 , n322046 , n2265 , n322048 , n322049 , n2268 , n322051 , n322052 , 
 n2271 , n322054 , n322055 , n322056 , n2275 , n322058 , n2277 , n322060 , n322061 , n2280 , 
 n322063 , n322064 , n2283 , n322066 , n322067 , n2286 , n2287 , n2288 , n322071 , n322072 , 
 n322073 , n2292 , n322075 , n2294 , n2295 , n322078 , n322079 , n322080 , n2299 , n322082 , 
 n322083 , n2302 , n322085 , n322086 , n2305 , n322088 , n322089 , n322090 , n2309 , n322092 , 
 n2311 , n2312 , n322095 , n322096 , n322097 , n2316 , n322099 , n322100 , n2319 , n322102 , 
 n322103 , n322104 , n322105 , n322106 , n322107 , n322108 , n322109 , n322110 , n322111 , n322112 , 
 n322113 , n322114 , n322115 , n322116 , n322117 , n322118 , n322119 , n322120 , n322121 , n2320 , 
 n322123 , n322124 , n322125 , n322126 , n322127 , n322128 , n322129 , n2324 , n322131 , n322132 , 
 n322133 , n322134 , n322135 , n322136 , n322137 , n322138 , n322139 , n322140 , n322141 , n322142 , 
 n322143 , n322144 , n322145 , n2327 , n322147 , n2329 , n322149 , n2330 , n2331 , n322152 , 
 n322153 , n322154 , n2335 , n322156 , n322157 , n2338 , n322159 , n322160 , n322161 , n322162 , 
 n322163 , n2342 , n322165 , n322166 , n2345 , n322168 , n322169 , n2347 , n322171 , n2349 , 
 n322173 , n322174 , n2352 , n322176 , n322177 , n2355 , n2356 , n322180 , n322181 , n322182 , 
 n2360 , n2361 , n322185 , n2363 , n2364 , n322188 , n2366 , n322190 , n322191 , n322192 , 
 n322193 , n322194 , n322195 , n322196 , n322197 , n322198 , n2376 , n322200 , n322201 , n322202 , 
 n322203 , n322204 , n322205 , n322206 , n2381 , n322208 , n322209 , n2384 , n322211 , n322212 , 
 n322213 , n322214 , n2389 , n322216 , n2391 , n322218 , n322219 , n322220 , n322221 , n322222 , 
 n322223 , n2398 , n322225 , n322226 , n2401 , n322228 , n322229 , n322230 , n322231 , n322232 , 
 n322233 , n322234 , n322235 , n322236 , n322237 , n2412 , n322239 , n322240 , n322241 , n322242 , 
 n322243 , n2418 , n322245 , n322246 , n322247 , n322248 , n322249 , n322250 , n2425 , n322252 , 
 n322253 , n322254 , n322255 , n2430 , n322257 , n322258 , n2433 , n322260 , n322261 , n2436 , 
 n2437 , n322264 , n2439 , n2440 , n322267 , n322268 , n2443 , n322270 , n322271 , n322272 , 
 n322273 , n322274 , n322275 , n322276 , n2451 , n322278 , n322279 , n322280 , n322281 , n322282 , 
 n322283 , n322284 , n2459 , n2460 , n322287 , n322288 , n322289 , n322290 , n322291 , n322292 , 
 n322293 , n322294 , n322295 , n2470 , n2471 , n322298 , n322299 , n322300 , n322301 , n2476 , 
 n322303 , n2478 , n2479 , n322306 , n322307 , n322308 , n322309 , n2484 , n322311 , n322312 , 
 n2487 , n322314 , n322315 , n322316 , n322317 , n322318 , n2493 , n322320 , n2495 , n2496 , 
 n2497 , n322324 , n322325 , n322326 , n322327 , n322328 , n322329 , n322330 , n322331 , n322332 , 
 n2504 , n322334 , n322335 , n2505 , n2506 , n322338 , n2508 , n322340 , n322341 , n322342 , 
 n322343 , n2513 , n322345 , n322346 , n322347 , n322348 , n2518 , n2519 , n322351 , n322352 , 
 n322353 , n322354 , n322355 , n322356 , n322357 , n322358 , n322359 , n322360 , n322361 , n322362 , 
 n322363 , n322364 , n2534 , n322366 , n322367 , n322368 , n322369 , n2539 , n322371 , n322372 , 
 n322373 , n322374 , n322375 , n2544 , n322377 , n2546 , n322379 , n2548 , n322381 , n322382 , 
 n322383 , n322384 , n2549 , n322386 , n322387 , n322388 , n322389 , n322390 , n322391 , n322392 , 
 n322393 , n322394 , n322395 , n322396 , n2561 , n2562 , n322399 , n2564 , n2565 , n322402 , 
 n322403 , n2568 , n322405 , n322406 , n322407 , n322408 , n322409 , n322410 , n2570 , n322412 , 
 n322413 , n322414 , n322415 , n2575 , n322417 , n322418 , n2578 , n2579 , n322421 , n322422 , 
 n322423 , n322424 , n322425 , n2585 , n322427 , n322428 , n322429 , n2589 , n2590 , n2591 , 
 n322433 , n322434 , n2594 , n322436 , n322437 , n322438 , n322439 , n322440 , n2600 , n322442 , 
 n322443 , n322444 , n322445 , n322446 , n322447 , n2607 , n322449 , n322450 , n322451 , n322452 , 
 n322453 , n322454 , n322455 , n322456 , n322457 , n322458 , n322459 , n322460 , n322461 , n2621 , 
 n322463 , n322464 , n322465 , n2625 , n322467 , n322468 , n322469 , n322470 , n322471 , n322472 , 
 n322473 , n322474 , n322475 , n322476 , n322477 , n322478 , n322479 , n322480 , n2640 , n322482 , 
 n2642 , n2643 , n322485 , n322486 , n2646 , n322488 , n322489 , n322490 , n322491 , n322492 , 
 n322493 , n2653 , n322495 , n322496 , n322497 , n322498 , n2658 , n322500 , n322501 , n322502 , 
 n322503 , n322504 , n322505 , n322506 , n322507 , n322508 , n2668 , n322510 , n322511 , n2671 , 
 n2672 , n322514 , n322515 , n2675 , n322517 , n322518 , n322519 , n322520 , n322521 , n322522 , 
 n322523 , n322524 , n322525 , n322526 , n322527 , n322528 , n322529 , n322530 , n2690 , n2691 , 
 n2692 , n2693 , n2694 , n322536 , n2696 , n322538 , n2698 , n322540 , n322541 , n322542 , 
 n322543 , n322544 , n2704 , n322546 , n322547 , n322548 , n322549 , n322550 , n322551 , n322552 , 
 n2711 , n322554 , n322555 , n2714 , n2715 , n322558 , n322559 , n322560 , n2719 , n322562 , 
 n322563 , n2722 , n322565 , n322566 , n322567 , n2726 , n322569 , n322570 , n2729 , n322572 , 
 n2731 , n2732 , n322575 , n322576 , n322577 , n322578 , n322579 , n322580 , n322581 , n2740 , 
 n322583 , n322584 , n322585 , n322586 , n322587 , n322588 , n322589 , n322590 , n2749 , n322592 , 
 n322593 , n2752 , n322595 , n322596 , n322597 , n322598 , n322599 , n322600 , n322601 , n2760 , 
 n322603 , n322604 , n2763 , n322606 , n2765 , n322608 , n322609 , n2768 , n322611 , n322612 , 
 n322613 , n2772 , n2773 , n322616 , n322617 , n322618 , n322619 , n322620 , n2779 , n322622 , 
 n322623 , n322624 , n322625 , n322626 , n2785 , n2786 , n2787 , n322630 , n2789 , n322632 , 
 n322633 , n322634 , n2793 , n2794 , n322637 , n322638 , n322639 , n2798 , n322641 , n322642 , 
 n322643 , n322644 , n322645 , n2804 , n2805 , n322648 , n322649 , n322650 , n2809 , n2810 , 
 n322653 , n322654 , n2813 , n322656 , n322657 , n322658 , n322659 , n322660 , n322661 , n2820 , 
 n322663 , n322664 , n2823 , n322666 , n322667 , n322668 , n322669 , n322670 , n322671 , n322672 , 
 n322673 , n2832 , n322675 , n322676 , n2835 , n322678 , n322679 , n322680 , n322681 , n2840 , 
 n2841 , n2842 , n2843 , n322686 , n2845 , n322688 , n2847 , n322690 , n322691 , n322692 , 
 n322693 , n322694 , n2853 , n322696 , n2855 , n322698 , n322699 , n322700 , n322701 , n322702 , 
 n322703 , n322704 , n322705 , n322706 , n322707 , n322708 , n2867 , n322710 , n322711 , n322712 , 
 n322713 , n2872 , n322715 , n322716 , n322717 , n322718 , n322719 , n2878 , n322721 , n322722 , 
 n2881 , n2882 , n322725 , n2884 , n322727 , n322728 , n322729 , n322730 , n322731 , n322732 , 
 n322733 , n322734 , n322735 , n2893 , n322737 , n2895 , n322739 , n322740 , n322741 , n322742 , 
 n2900 , n322744 , n322745 , n2903 , n2904 , n2905 , n322749 , n322750 , n2908 , n2909 , 
 n322753 , n322754 , n322755 , n2913 , n2914 , n2915 , n322759 , n322760 , n322761 , n322762 , 
 n322763 , n2921 , n2922 , n322766 , n322767 , n2925 , n2926 , n2927 , n2928 , n2929 , 
 n2930 , n322774 , n2932 , n322776 , n322777 , n2935 , n322779 , n322780 , n2938 , n322782 , 
 n2940 , n2941 , n2942 , n322786 , n322787 , n2945 , n322789 , n2947 , n322791 , n322792 , 
 n2950 , n322794 , n2952 , n2953 , n2954 , n2955 , n322799 , n2957 , n322801 , n2959 , 
 n322803 , n322804 , n2962 , n322806 , n2964 , n2965 , n2966 , n2967 , n322811 , n2969 , 
 n322813 , n2971 , n2972 , n322816 , n322817 , n2975 , n322819 , n322820 , n2978 , n322822 , 
 n2980 , n2981 , n322825 , n2983 , n322827 , n2985 , n322829 , n322830 , n2988 , n322832 , 
 n322833 , n322834 , n2992 , n322836 , n322837 , n2995 , n2996 , n2997 , n2998 , n2999 , 
 n3000 , n3001 , n322845 , n322846 , n3004 , n322848 , n3006 , n322850 , n3008 , n3009 , 
 n3010 , n322854 , n322855 , n322856 , n3014 , n322858 , n322859 , n3017 , n322861 , n322862 , 
 n3020 , n322864 , n322865 , n3023 , n322867 , n3025 , n3026 , n322870 , n3028 , n322872 , 
 n3030 , n3031 , n322875 , n322876 , n322877 , n3035 , n322879 , n322880 , n3038 , n322882 , 
 n322883 , n3041 , n322885 , n3043 , n322887 , n3045 , n3046 , n3047 , n3048 , n322892 , 
 n322893 , n322894 , n3052 , n322896 , n322897 , n3055 , n322899 , n3057 , n3058 , n3059 , 
 n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n322910 , n3068 , n322912 , 
 n3070 , n3071 , n322915 , n322916 , n3074 , n322918 , n3076 , n3077 , n3078 , n322922 , 
 n3080 , n322924 , n3082 , n322926 , n3084 , n3085 , n3086 , n322930 , n3088 , n3089 , 
 n3090 , n3091 , n3092 , n322936 , n322937 , n3095 , n322939 , n3097 , n3098 , n322942 , 
 n322943 , n322944 , n3102 , n322946 , n322947 , n3105 , n322949 , n3107 , n322951 , n3109 , 
 n3110 , n3111 , n3112 , n322956 , n3114 , n322958 , n3116 , n322960 , n3118 , n322962 , 
 n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n322971 , n3129 , 
 n322973 , n322974 , n3132 , n322976 , n3134 , n3135 , n322979 , n3137 , n322981 , n322982 , 
 n3140 , n322984 , n322985 , n322986 , n322987 , n3145 , n322989 , n3147 , n322991 , n322992 , 
 n3150 , n322994 , n322995 , n322996 , n3154 , n322998 , n3156 , n3157 , n3158 , n3159 , 
 n323003 , n323004 , n3162 , n323006 , n323007 , n3165 , n323009 , n323010 , n323011 , n323012 , 
 n3170 , n323014 , n323015 , n3173 , n323017 , n3175 , n323019 , n323020 , n323021 , n3179 , 
 n323023 , n323024 , n3182 , n323026 , n3184 , n3185 , n3186 , n323030 , n323031 , n3189 , 
 n323033 , n323034 , n3192 , n323036 , n323037 , n3195 , n323039 , n323040 , n3198 , n323042 , 
 n3200 , n323044 , n323045 , n323046 , n323047 , n3205 , n323049 , n323050 , n323051 , n3209 , 
 n323053 , n323054 , n323055 , n323056 , n3214 , n323058 , n323059 , n3217 , n323061 , n3219 , 
 n3220 , n323064 , n323065 , n3223 , n323067 , n323068 , n323069 , n3227 , n323071 , n323072 , 
 n3230 , n323074 , n323075 , n3233 , n323077 , n323078 , n3236 , n323080 , n323081 , n3239 , 
 n3240 , n323084 , n3242 , n3243 , n323087 , n323088 , n323089 , n3247 , n323091 , n3249 , 
 n3250 , n323094 , n323095 , n3253 , n323097 , n323098 , n3256 , n323100 , n323101 , n323102 , 
 n3260 , n323104 , n3262 , n3263 , n323107 , n323108 , n323109 , n3267 , n323111 , n323112 , 
 n3270 , n323114 , n323115 , n3273 , n323117 , n323118 , n3276 , n323120 , n323121 , n3279 , 
 n323123 , n323124 , n323125 , n3283 , n323127 , n323128 , n3286 , n323130 , n323131 , n3289 , 
 n323133 , n323134 , n3292 , n3293 , n3294 , n323138 , n323139 , n3297 , n3298 , n3299 , 
 n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n323149 , n323150 , n3308 , n323152 , 
 n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n323161 , n323162 , 
 n323163 , n3321 , n323165 , n323166 , n3324 , n323168 , n3326 , n3327 , n3328 , n3329 , 
 n3330 , n323174 , n3332 , n3333 , n3334 , n323178 , n323179 , n3337 , n3338 , n3339 , 
 n323183 , n323184 , n3342 , n3343 , n3344 , n3345 , n3346 , n323190 , n323191 , n3349 , 
 n3350 , n3351 , n323195 , n3353 , n323197 , n3355 , n323199 , n3357 , n323201 , n323202 , 
 n3360 , n323204 , n3362 , n323206 , n323207 , n323208 , n323209 , n3367 , n323211 , n323212 , 
 n323213 , n3371 , n323215 , n323216 , n323217 , n3375 , n323219 , n3377 , n3378 , n323222 , 
 n323223 , n323224 , n323225 , n323226 , n323227 , n3385 , n323229 , n323230 , n323231 , n323232 , 
 n323233 , n323234 , n323235 , n3393 , n323237 , n3395 , n323239 , n3397 , n323241 , n323242 , 
 n323243 , n323244 , n323245 , n323246 , n3404 , n323248 , n323249 , n323250 , n3408 , n323252 , 
 n323253 , n323254 , n323255 , n323256 , n323257 , n323258 , n323259 , n323260 , n323261 , n323262 , 
 n323263 , n323264 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n323272 , 
 n323273 , n323274 , n323275 , n3433 , n323277 , n323278 , n3436 , n3437 , n323281 , n323282 , 
 n323283 , n323284 , n323285 , n3443 , n323287 , n3445 , n3446 , n3447 , n3448 , n3449 , 
 n3450 , n323294 , n323295 , n323296 , n323297 , n323298 , n3456 , n323300 , n323301 , n323302 , 
 n323303 , n323304 , n323305 , n323306 , n3464 , n323308 , n323309 , n323310 , n323311 , n323312 , 
 n323313 , n323314 , n323315 , n323316 , n3474 , n323318 , n3476 , n323320 , n323321 , n323322 , 
 n323323 , n323324 , n323325 , n3483 , n323327 , n323328 , n323329 , n3487 , n323331 , n3489 , 
 n3490 , n323334 , n323335 , n323336 , n3494 , n323338 , n323339 , n323340 , n323341 , n323342 , 
 n3500 , n323344 , n323345 , n323346 , n3504 , n323348 , n323349 , n323350 , n323351 , n323352 , 
 n323353 , n323354 , n3512 , n323356 , n323357 , n3515 , n323359 , n323360 , n3518 , n323362 , 
 n323363 , n3521 , n323365 , n323366 , n3524 , n323368 , n3526 , n323370 , n323371 , n3529 , 
 n323373 , n323374 , n3532 , n323376 , n323377 , n323378 , n323379 , n323380 , n3538 , n323382 , 
 n3540 , n323384 , n323385 , n3543 , n323387 , n323388 , n3546 , n323390 , n323391 , n323392 , 
 n323393 , n323394 , n323395 , n323396 , n323397 , n3555 , n323399 , n323400 , n323401 , n323402 , 
 n323403 , n323404 , n3562 , n323406 , n323407 , n323408 , n3566 , n323410 , n323411 , n323412 , 
 n323413 , n3571 , n323415 , n3573 , n323417 , n323418 , n323419 , n3577 , n323421 , n323422 , 
 n323423 , n3581 , n323425 , n323426 , n3584 , n323428 , n323429 , n3587 , n3588 , n323432 , 
 n323433 , n3591 , n323435 , n323436 , n323437 , n323438 , n3596 , n323440 , n323441 , n3599 , 
 n323443 , n323444 , n3602 , n323446 , n323447 , n323448 , n323449 , n3607 , n3608 , n323452 , 
 n323453 , n323454 , n323455 , n323456 , n323457 , n3615 , n323459 , n323460 , n3618 , n3619 , 
 n323463 , n323464 , n323465 , n3623 , n3624 , n323468 , n323469 , n323470 , n323471 , n3629 , 
 n3630 , n323474 , n323475 , n323476 , n323477 , n3635 , n323479 , n323480 , n3638 , n323482 , 
 n323483 , n323484 , n323485 , n323486 , n323487 , n323488 , n323489 , n323490 , n323491 , n323492 , 
 n323493 , n323494 , n3652 , n3653 , n3654 , n323498 , n323499 , n323500 , n323501 , n323502 , 
 n323503 , n323504 , n3662 , n323506 , n3664 , n323508 , n3666 , n3667 , n323511 , n323512 , 
 n323513 , n323514 , n323515 , n323516 , n3674 , n323518 , n323519 , n3677 , n323521 , n323522 , 
 n3680 , n323524 , n323525 , n3683 , n323527 , n323528 , n323529 , n323530 , n323531 , n3689 , 
 n323533 , n323534 , n323535 , n3693 , n3694 , n323538 , n3696 , n323540 , n3698 , n323542 , 
 n323543 , n3701 , n3702 , n3703 , n3704 , n323548 , n323549 , n323550 , n323551 , n323552 , 
 n3710 , n323554 , n323555 , n323556 , n3714 , n323558 , n323559 , n323560 , n323561 , n323562 , 
 n323563 , n3721 , n323565 , n3723 , n323567 , n323568 , n3726 , n3727 , n323571 , n3729 , 
 n323573 , n323574 , n323575 , n323576 , n323577 , n3735 , n323579 , n323580 , n3738 , n323582 , 
 n323583 , n3741 , n323585 , n323586 , n323587 , n323588 , n323589 , n323590 , n323591 , n323592 , 
 n3750 , n323594 , n3752 , n323596 , n3754 , n3755 , n3756 , n3757 , n323601 , n323602 , 
 n323603 , n323604 , n323605 , n323606 , n323607 , n323608 , n323609 , n323610 , n323611 , n323612 , 
 n3770 , n323614 , n323615 , n323616 , n323617 , n323618 , n323619 , n323620 , n323621 , n323622 , 
 n323623 , n323624 , n323625 , n323626 , n323627 , n3785 , n323629 , n323630 , n3788 , n323632 , 
 n323633 , n3791 , n3792 , n323636 , n323637 , n3795 , n323639 , n323640 , n323641 , n3799 , 
 n323643 , n3801 , n3802 , n323646 , n323647 , n323648 , n3806 , n323650 , n323651 , n323652 , 
 n323653 , n323654 , n3812 , n323656 , n323657 , n323658 , n323659 , n323660 , n323661 , n3819 , 
 n323663 , n3821 , n323665 , n323666 , n323667 , n323668 , n323669 , n323670 , n323671 , n323672 , 
 n323673 , n323674 , n323675 , n3833 , n3834 , n3835 , n3836 , n323680 , n3838 , n323682 , 
 n323683 , n3841 , n323685 , n3843 , n323687 , n3845 , n323689 , n323690 , n323691 , n323692 , 
 n323693 , n3851 , n323695 , n323696 , n3854 , n323698 , n323699 , n3857 , n3858 , n3859 , 
 n323703 , n323704 , n323705 , n323706 , n323707 , n3865 , n323709 , n3867 , n3868 , n3869 , 
 n323713 , n323714 , n323715 , n323716 , n3874 , n3875 , n3876 , n323720 , n323721 , n3879 , 
 n3880 , n323724 , n3882 , n3883 , n323727 , n323728 , n323729 , n323730 , n323731 , n323732 , 
 n323733 , n323734 , n3892 , n323736 , n3894 , n3895 , n3896 , n3897 , n323741 , n323742 , 
 n323743 , n323744 , n323745 , n323746 , n323747 , n323748 , n3906 , n323750 , n3908 , n323752 , 
 n323753 , n3911 , n323755 , n3913 , n323757 , n323758 , n323759 , n323760 , n323761 , n323762 , 
 n323763 , n323764 , n323765 , n323766 , n323767 , n323768 , n323769 , n3927 , n323771 , n3929 , 
 n3930 , n323774 , n323775 , n323776 , n323777 , n323778 , n323779 , n3937 , n323781 , n323782 , 
 n323783 , n323784 , n323785 , n323786 , n323787 , n323788 , n323789 , n323790 , n3948 , n323792 , 
 n323793 , n3951 , n323795 , n323796 , n3954 , n323798 , n323799 , n323800 , n323801 , n323802 , 
 n323803 , n323804 , n323805 , n3963 , n323807 , n323808 , n3966 , n323810 , n323811 , n3969 , 
 n323813 , n323814 , n323815 , n3973 , n323817 , n323818 , n323819 , n3977 , n3978 , n323822 , 
 n323823 , n323824 , n323825 , n323826 , n3984 , n323828 , n323829 , n323830 , n323831 , n323832 , 
 n323833 , n323834 , n323835 , n323836 , n3994 , n323838 , n323839 , n323840 , n323841 , n323842 , 
 n323843 , n323844 , n323845 , n323846 , n323847 , n4005 , n323849 , n323850 , n4008 , n323852 , 
 n4010 , n323854 , n4012 , n4013 , n323857 , n323858 , n323859 , n4017 , n323861 , n323862 , 
 n4020 , n323864 , n323865 , n4023 , n323867 , n323868 , n4026 , n323870 , n323871 , n4029 , 
 n323873 , n4031 , n323875 , n323876 , n323877 , n323878 , n323879 , n323880 , n4038 , n323882 , 
 n323883 , n323884 , n4042 , n323886 , n323887 , n323888 , n4046 , n323890 , n323891 , n323892 , 
 n323893 , n323894 , n323895 , n323896 , n323897 , n323898 , n323899 , n323900 , n323901 , n4059 , 
 n323903 , n323904 , n323905 , n4063 , n323907 , n323908 , n323909 , n323910 , n323911 , n323912 , 
 n323913 , n323914 , n323915 , n323916 , n323917 , n323918 , n4076 , n323920 , n323921 , n4079 , 
 n4080 , n323924 , n323925 , n323926 , n323927 , n323928 , n323929 , n323930 , n323931 , n4089 , 
 n323933 , n4091 , n323935 , n323936 , n323937 , n323938 , n323939 , n323940 , n323941 , n323942 , 
 n323943 , n323944 , n323945 , n4103 , n4104 , n323948 , n323949 , n323950 , n4108 , n323952 , 
 n323953 , n323954 , n323955 , n4113 , n4114 , n323958 , n323959 , n323960 , n323961 , n323962 , 
 n4120 , n323964 , n323965 , n4123 , n323967 , n323968 , n323969 , n323970 , n4128 , n323972 , 
 n4130 , n323974 , n323975 , n323976 , n323977 , n323978 , n323979 , n4137 , n323981 , n323982 , 
 n4140 , n323984 , n4142 , n323986 , n323987 , n323988 , n4146 , n4147 , n4148 , n323992 , 
 n323993 , n323994 , n323995 , n323996 , n4154 , n4155 , n4156 , n324000 , n324001 , n324002 , 
 n324003 , n4161 , n324005 , n324006 , n4164 , n324008 , n4166 , n324010 , n324011 , n324012 , 
 n324013 , n4171 , n324015 , n324016 , n324017 , n324018 , n324019 , n324020 , n4178 , n324022 , 
 n4180 , n4181 , n324025 , n324026 , n4184 , n324028 , n324029 , n324030 , n4188 , n324032 , 
 n324033 , n4191 , n4192 , n324036 , n324037 , n324038 , n324039 , n324040 , n324041 , n4199 , 
 n4200 , n324044 , n324045 , n324046 , n324047 , n324048 , n324049 , n324050 , n324051 , n324052 , 
 n4210 , n324054 , n324055 , n324056 , n4214 , n4215 , n324059 , n324060 , n4218 , n324062 , 
 n324063 , n4221 , n4222 , n324066 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
 n4230 , n4231 , n324075 , n324076 , n324077 , n324078 , n4236 , n4237 , n324081 , n324082 , 
 n324083 , n324084 , n4242 , n324086 , n324087 , n324088 , n324089 , n324090 , n324091 , n324092 , 
 n4250 , n324094 , n324095 , n4253 , n324097 , n4255 , n4256 , n4257 , n324101 , n4259 , 
 n324103 , n4261 , n324105 , n324106 , n324107 , n324108 , n324109 , n324110 , n324111 , n4269 , 
 n324113 , n324114 , n324115 , n324116 , n4274 , n4275 , n4276 , n4277 , n324121 , n324122 , 
 n324123 , n324124 , n324125 , n324126 , n324127 , n324128 , n4286 , n324130 , n324131 , n4289 , 
 n324133 , n4291 , n324135 , n324136 , n324137 , n324138 , n324139 , n324140 , n324141 , n324142 , 
 n324143 , n324144 , n324145 , n324146 , n4304 , n324148 , n4306 , n4307 , n324151 , n324152 , 
 n324153 , n324154 , n324155 , n324156 , n324157 , n324158 , n324159 , n324160 , n324161 , n4319 , 
 n324163 , n324164 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n324171 , n4329 , 
 n324173 , n4331 , n4332 , n4333 , n324177 , n324178 , n4336 , n324180 , n324181 , n324182 , 
 n4340 , n324184 , n324185 , n4343 , n324187 , n324188 , n4346 , n324190 , n324191 , n4349 , 
 n324193 , n324194 , n324195 , n324196 , n4354 , n324198 , n324199 , n4357 , n324201 , n324202 , 
 n324203 , n4361 , n324205 , n324206 , n4364 , n324208 , n324209 , n4367 , n324211 , n324212 , 
 n324213 , n324214 , n324215 , n324216 , n324217 , n324218 , n324219 , n324220 , n324221 , n4379 , 
 n4380 , n324224 , n324225 , n4383 , n324227 , n324228 , n324229 , n324230 , n324231 , n324232 , 
 n4390 , n324234 , n324235 , n324236 , n324237 , n324238 , n324239 , n324240 , n324241 , n324242 , 
 n324243 , n324244 , n324245 , n324246 , n324247 , n324248 , n324249 , n4407 , n324251 , n4409 , 
 n4410 , n324254 , n324255 , n324256 , n324257 , n324258 , n4416 , n4417 , n4418 , n4419 , 
 n324263 , n324264 , n324265 , n324266 , n324267 , n324268 , n4426 , n324270 , n324271 , n324272 , 
 n324273 , n324274 , n324275 , n324276 , n324277 , n4435 , n4436 , n324280 , n324281 , n324282 , 
 n4440 , n324284 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n324291 , n324292 , 
 n324293 , n324294 , n324295 , n324296 , n4454 , n324298 , n4456 , n4457 , n324301 , n4459 , 
 n324303 , n4461 , n324305 , n324306 , n324307 , n324308 , n324309 , n4467 , n324311 , n4469 , 
 n324313 , n324314 , n4472 , n4473 , n4474 , n4475 , n4476 , n324320 , n324321 , n324322 , 
 n324323 , n4481 , n324325 , n324326 , n324327 , n324328 , n324329 , n4487 , n4488 , n4489 , 
 n4490 , n324334 , n324335 , n4493 , n4494 , n4495 , n324339 , n324340 , n4498 , n324342 , 
 n324343 , n324344 , n324345 , n4503 , n4504 , n324348 , n4506 , n4507 , n324351 , n324352 , 
 n324353 , n4511 , n324355 , n324356 , n324357 , n324358 , n4516 , n4517 , n324361 , n324362 , 
 n4520 , n324364 , n324365 , n4523 , n4524 , n324368 , n324369 , n4527 , n4528 , n324372 , 
 n324373 , n324374 , n4532 , n324376 , n324377 , n324378 , n324379 , n324380 , n4538 , n324382 , 
 n324383 , n324384 , n324385 , n4543 , n324387 , n324388 , n324389 , n4547 , n324391 , n324392 , 
 n324393 , n324394 , n4552 , n4553 , n4554 , n4555 , n4556 , n324400 , n324401 , n324402 , 
 n324403 , n4561 , n324405 , n4563 , n324407 , n324408 , n324409 , n324410 , n324411 , n4569 , 
 n4570 , n324414 , n324415 , n324416 , n4574 , n324418 , n324419 , n4577 , n324421 , n324422 , 
 n324423 , n324424 , n4582 , n324426 , n324427 , n324428 , n4586 , n4587 , n4588 , n4589 , 
 n324433 , n4591 , n324435 , n324436 , n4594 , n324438 , n324439 , n4597 , n324441 , n324442 , 
 n324443 , n324444 , n324445 , n324446 , n324447 , n4605 , n324449 , n324450 , n324451 , n324452 , 
 n324453 , n324454 , n4612 , n324456 , n324457 , n4615 , n324459 , n4617 , n4618 , n4619 , 
 n324463 , n4621 , n324465 , n324466 , n324467 , n324468 , n324469 , n4627 , n324471 , n324472 , 
 n324473 , n324474 , n324475 , n324476 , n324477 , n324478 , n324479 , n4637 , n4638 , n4639 , 
 n324483 , n324484 , n4642 , n324486 , n4644 , n4645 , n4646 , n4647 , n324491 , n4649 , 
 n324493 , n4651 , n4652 , n4653 , n4654 , n324498 , n4656 , n4657 , n4658 , n4659 , 
 n4660 , n324504 , n324505 , n4663 , n324507 , n4665 , n324509 , n4667 , n324511 , n324512 , 
 n324513 , n324514 , n4672 , n324516 , n324517 , n324518 , n324519 , n4677 , n324521 , n324522 , 
 n4680 , n4681 , n4682 , n324526 , n4684 , n324528 , n324529 , n4687 , n324531 , n324532 , 
 n324533 , n324534 , n324535 , n324536 , n324537 , n4695 , n324539 , n324540 , n4698 , n4699 , 
 n324543 , n4701 , n324545 , n4703 , n4704 , n324548 , n324549 , n324550 , n324551 , n324552 , 
 n324553 , n324554 , n324555 , n324556 , n324557 , n324558 , n324559 , n4717 , n4718 , n4719 , 
 n324563 , n324564 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
 n4730 , n4731 , n4732 , n4733 , n324577 , n324578 , n4736 , n324580 , n324581 , n4739 , 
 n324583 , n324584 , n324585 , n324586 , n324587 , n4742 , n324589 , n324590 , n324591 , n4746 , 
 n324593 , n324594 , n4749 , n324596 , n4751 , n4752 , n4753 , n324600 , n4755 , n324602 , 
 n324603 , n324604 , n4759 , n324606 , n324607 , n4762 , n324609 , n324610 , n4765 , n324612 , 
 n4767 , n4768 , n324615 , n324616 , n4771 , n324618 , n4773 , n324620 , n4775 , n324622 , 
 n324623 , n4778 , n324625 , n4780 , n324627 , n4782 , n324629 , n4784 , n324631 , n4786 , 
 n4787 , n4788 , n324635 , n324636 , n4791 , n324638 , n4793 , n324640 , n4795 , n4796 , 
 n324643 , n324644 , n324645 , n4800 , n324647 , n4802 , n4803 , n4804 , n324651 , n324652 , 
 n324653 , n324654 , n324655 , n324656 , n324657 , n324658 , n324659 , n4814 , n4815 , n324662 , 
 n324663 , n4818 , n324665 , n324666 , n324667 , n324668 , n324669 , n324670 , n4825 , n324672 , 
 n324673 , n324674 , n324675 , n4830 , n324677 , n4832 , n324679 , n324680 , n4835 , n4836 , 
 n324683 , n324684 , n4839 , n324686 , n324687 , n324688 , n324689 , n324690 , n324691 , n324692 , 
 n4847 , n324694 , n324695 , n4850 , n324697 , n324698 , n324699 , n324700 , n324701 , n324702 , 
 n4857 , n324704 , n4859 , n324706 , n324707 , n324708 , n324709 , n324710 , n324711 , n324712 , 
 n324713 , n324714 , n324715 , n324716 , n324717 , n324718 , n324719 , n324720 , n324721 , n324722 , 
 n324723 , n324724 , n324725 , n4880 , n324727 , n324728 , n324729 , n4884 , n324731 , n4886 , 
 n324733 , n324734 , n324735 , n324736 , n324737 , n324738 , n324739 , n324740 , n4895 , n4896 , 
 n324743 , n4898 , n4899 , n324746 , n4901 , n324748 , n324749 , n324750 , n324751 , n324752 , 
 n324753 , n4908 , n324755 , n4910 , n4911 , n324758 , n324759 , n4914 , n324761 , n324762 , 
 n4917 , n324764 , n324765 , n324766 , n324767 , n324768 , n324769 , n324770 , n4925 , n324772 , 
 n324773 , n324774 , n324775 , n324776 , n324777 , n324778 , n324779 , n324780 , n324781 , n324782 , 
 n324783 , n4938 , n4939 , n324786 , n324787 , n324788 , n324789 , n324790 , n324791 , n324792 , 
 n324793 , n324794 , n324795 , n324796 , n4951 , n4952 , n4953 , n324800 , n324801 , n324802 , 
 n4957 , n324804 , n324805 , n4960 , n324807 , n324808 , n324809 , n4964 , n324811 , n324812 , 
 n324813 , n324814 , n4969 , n324816 , n324817 , n324818 , n324819 , n324820 , n4975 , n4976 , 
 n324823 , n4978 , n324825 , n324826 , n324827 , n324828 , n324829 , n324830 , n324831 , n324832 , 
 n324833 , n324834 , n324835 , n324836 , n324837 , n324838 , n324839 , n324840 , n4995 , n324842 , 
 n324843 , n4998 , n324845 , n5000 , n5001 , n324848 , n5003 , n324850 , n5005 , n324852 , 
 n5007 , n5008 , n324855 , n324856 , n324857 , n324858 , n324859 , n324860 , n324861 , n324862 , 
 n324863 , n5018 , n5019 , n5020 , n324867 , n324868 , n324869 , n324870 , n324871 , n324872 , 
 n324873 , n5028 , n324875 , n324876 , n5031 , n324878 , n5033 , n5034 , n324881 , n5036 , 
 n324883 , n5038 , n324885 , n324886 , n5041 , n324888 , n324889 , n324890 , n324891 , n324892 , 
 n324893 , n324894 , n324895 , n324896 , n324897 , n324898 , n324899 , n5054 , n324901 , n5056 , 
 n5057 , n324904 , n324905 , n5060 , n324907 , n324908 , n324909 , n5064 , n5065 , n324912 , 
 n324913 , n324914 , n5069 , n324916 , n324917 , n5072 , n324919 , n324920 , n5075 , n324922 , 
 n5077 , n324924 , n324925 , n5080 , n5081 , n324928 , n324929 , n5084 , n324931 , n5086 , 
 n324933 , n5088 , n324935 , n5090 , n324937 , n5092 , n5093 , n324940 , n324941 , n324942 , 
 n5097 , n324944 , n324945 , n5100 , n324947 , n324948 , n5103 , n324950 , n5105 , n5106 , 
 n324953 , n5108 , n324955 , n5110 , n5111 , n324958 , n324959 , n324960 , n5115 , n324962 , 
 n324963 , n5118 , n324965 , n324966 , n5121 , n324968 , n5123 , n324970 , n324971 , n324972 , 
 n5127 , n324974 , n324975 , n324976 , n324977 , n5132 , n324979 , n5134 , n5135 , n5136 , 
 n324983 , n5138 , n5139 , n5140 , n324987 , n5142 , n324989 , n324990 , n5145 , n324992 , 
 n324993 , n5148 , n324995 , n324996 , n5151 , n324998 , n324999 , n5154 , n325001 , n325002 , 
 n325003 , n5158 , n325005 , n325006 , n325007 , n5162 , n325009 , n5164 , n5165 , n5166 , 
 n5167 , n325014 , n5169 , n325016 , n5171 , n325018 , n325019 , n325020 , n5175 , n325022 , 
 n325023 , n5178 , n325025 , n325026 , n5181 , n325028 , n325029 , n5184 , n325031 , n325032 , 
 n5187 , n325034 , n325035 , n5190 , n325037 , n5192 , n5193 , n325040 , n325041 , n5196 , 
 n325043 , n325044 , n5199 , n325046 , n325047 , n5202 , n325049 , n325050 , n5205 , n5206 , 
 n5207 , n325054 , n5209 , n325056 , n325057 , n325058 , n325059 , n5214 , n325061 , n325062 , 
 n5217 , n325064 , n325065 , n5220 , n5221 , n325068 , n325069 , n5224 , n325071 , n5226 , 
 n325073 , n5228 , n5229 , n325076 , n325077 , n5232 , n325079 , n325080 , n5235 , n325082 , 
 n325083 , n325084 , n5239 , n5240 , n325087 , n5242 , n5243 , n325090 , n325091 , n5246 , 
 n5247 , n5248 , n325095 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
 n5257 , n5258 , n5259 , n5260 , n325107 , n325108 , n5263 , n325110 , n325111 , n325112 , 
 n5267 , n325114 , n325115 , n5270 , n5271 , n325118 , n5273 , n325120 , n5275 , n5276 , 
 n325123 , n325124 , n5279 , n325126 , n325127 , n5282 , n325129 , n325130 , n5285 , n5286 , 
 n5287 , n325134 , n5289 , n5290 , n325137 , n5292 , n325139 , n5294 , n5295 , n5296 , 
 n325143 , n325144 , n5299 , n325146 , n5301 , n5302 , n5303 , n325150 , n325151 , n5306 , 
 n325153 , n5308 , n325155 , n5310 , n5311 , n325158 , n5313 , n325160 , n5315 , n5316 , 
 n325163 , n325164 , n5319 , n325166 , n325167 , n5322 , n325169 , n325170 , n5325 , n5326 , 
 n325173 , n325174 , n5329 , n5330 , n325177 , n5332 , n325179 , n5334 , n5335 , n325182 , 
 n325183 , n5338 , n325185 , n325186 , n5341 , n325188 , n325189 , n5344 , n325191 , n325192 , 
 n5347 , n325194 , n5349 , n5350 , n325197 , n5352 , n5353 , n325200 , n325201 , n5356 , 
 n325203 , n325204 , n5359 , n325206 , n325207 , n325208 , n5363 , n325210 , n5365 , n5366 , 
 n325213 , n325214 , n5369 , n325216 , n325217 , n5372 , n325219 , n325220 , n5375 , n325222 , 
 n325223 , n325224 , n325225 , n325226 , n325227 , n325228 , n5383 , n325230 , n325231 , n325232 , 
 n325233 , n325234 , n325235 , n325236 , n5391 , n325238 , n325239 , n5394 , n5395 , n5396 , 
 n325243 , n325244 , n5399 , n325246 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
 n5407 , n325254 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n325262 , 
 n5417 , n325264 , n325265 , n325266 , n325267 , n5422 , n325269 , n325270 , n325271 , n325272 , 
 n325273 , n325274 , n5429 , n5430 , n325277 , n5432 , n5433 , n325280 , n325281 , n325282 , 
 n325283 , n5438 , n325285 , n325286 , n325287 , n325288 , n5443 , n325290 , n325291 , n5445 , 
 n325293 , n5447 , n5448 , n5449 , n5450 , n5451 , n325299 , n325300 , n5454 , n325302 , 
 n325303 , n325304 , n325305 , n325306 , n325307 , n325308 , n325309 , n325310 , n325311 , n325312 , 
 n325313 , n5467 , n325315 , n325316 , n325317 , n325318 , n325319 , n5473 , n325321 , n325322 , 
 n325323 , n325324 , n325325 , n325326 , n325327 , n325328 , n325329 , n325330 , n325331 , n325332 , 
 n5486 , n325334 , n325335 , n5489 , n325337 , n325338 , n325339 , n325340 , n325341 , n325342 , 
 n325343 , n325344 , n325345 , n5499 , n5500 , n325348 , n325349 , n5503 , n325351 , n325352 , 
 n5506 , n325354 , n325355 , n5509 , n325357 , n325358 , n325359 , n325360 , n325361 , n5515 , 
 n325363 , n5516 , n325365 , n325366 , n5519 , n325368 , n325369 , n325370 , n5523 , n325372 , 
 n325373 , n5526 , n325375 , n325376 , n325377 , n325378 , n325379 , n5532 , n325381 , n5534 , 
 n5535 , n325384 , n325385 , n5538 , n325387 , n325388 , n325389 , n325390 , n325391 , n325392 , 
 n5545 , n325394 , n5547 , n325396 , n325397 , n5550 , n325399 , n325400 , n325401 , n325402 , 
 n5555 , n325404 , n325405 , n5558 , n325407 , n325408 , n5561 , n325410 , n325411 , n5564 , 
 n5565 , n5566 , n325415 , n325416 , n325417 , n5570 , n325419 , n325420 , n325421 , n325422 , 
 n325423 , n5576 , n325425 , n325426 , n5579 , n5580 , n325429 , n325430 , n325431 , n325432 , 
 n325433 , n325434 , n325435 , n325436 , n325437 , n5590 , n325439 , n325440 , n325441 , n325442 , 
 n5595 , n325444 , n325445 , n5598 , n325447 , n5600 , n325449 , n325450 , n325451 , n325452 , 
 n325453 , n325454 , n325455 , n325456 , n325457 , n325458 , n325459 , n325460 , n325461 , n325462 , 
 n325463 , n325464 , n325465 , n325466 , n325467 , n325468 , n325469 , n325470 , n5623 , n325472 , 
 n325473 , n5626 , n5627 , n325476 , n5629 , n5630 , n325479 , n325480 , n325481 , n325482 , 
 n325483 , n325484 , n325485 , n325486 , n325487 , n325488 , n325489 , n325490 , n325491 , n325492 , 
 n325493 , n325494 , n325495 , n325496 , n325497 , n5650 , n325499 , n5652 , n325501 , n325502 , 
 n325503 , n325504 , n5657 , n325506 , n325507 , n5660 , n325509 , n325510 , n5663 , n325512 , 
 n325513 , n325514 , n325515 , n325516 , n325517 , n325518 , n325519 , n5672 , n325521 , n5674 , 
 n5675 , n325524 , n325525 , n325526 , n5679 , n325528 , n325529 , n325530 , n325531 , n325532 , 
 n325533 , n325534 , n325535 , n325536 , n325537 , n325538 , n5691 , n325540 , n325541 , n325542 , 
 n5695 , n5696 , n5697 , n5698 , n325547 , n5700 , n325549 , n5702 , n5703 , n5704 , 
 n325553 , n325554 , n5707 , n325556 , n325557 , n5710 , n325559 , n5712 , n325561 , n325562 , 
 n325563 , n5716 , n325565 , n5718 , n5719 , n325568 , n5721 , n325570 , n5723 , n325572 , 
 n325573 , n325574 , n325575 , n325576 , n325577 , n325578 , n5731 , n325580 , n325581 , n5734 , 
 n325583 , n325584 , n325585 , n325586 , n325587 , n325588 , n5741 , n325590 , n325591 , n5744 , 
 n325593 , n5746 , n5747 , n325596 , n325597 , n5750 , n325599 , n5752 , n5753 , n5754 , 
 n325603 , n325604 , n325605 , n325606 , n5759 , n325608 , n5761 , n5762 , n5763 , n5764 , 
 n325613 , n325614 , n325615 , n325616 , n325617 , n325618 , n325619 , n325620 , n5773 , n325622 , 
 n325623 , n5776 , n325625 , n325626 , n325627 , n325628 , n325629 , n325630 , n325631 , n325632 , 
 n5785 , n5786 , n5787 , n325636 , n325637 , n5790 , n325639 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n325647 , n325648 , n325649 , n325650 , n325651 , n325652 , 
 n325653 , n325654 , n325655 , n5808 , n325657 , n325658 , n5811 , n325660 , n325661 , n5814 , 
 n325663 , n325664 , n5817 , n325666 , n5819 , n5820 , n5821 , n5822 , n325671 , n325672 , 
 n325673 , n5826 , n325675 , n325676 , n5829 , n325678 , n325679 , n5832 , n325681 , n325682 , 
 n325683 , n5836 , n325685 , n325686 , n5839 , n325688 , n325689 , n5842 , n325691 , n325692 , 
 n5845 , n325694 , n5847 , n325696 , n325697 , n5850 , n325699 , n325700 , n325701 , n325702 , 
 n325703 , n325704 , n325705 , n325706 , n325707 , n325708 , n325709 , n325710 , n325711 , n325712 , 
 n325713 , n325714 , n325715 , n5868 , n325717 , n325718 , n5871 , n325720 , n325721 , n5874 , 
 n325723 , n5876 , n325725 , n5878 , n325727 , n5880 , n325729 , n325730 , n325731 , n325732 , 
 n5885 , n325734 , n325735 , n5888 , n325737 , n325738 , n325739 , n5892 , n325741 , n325742 , 
 n5895 , n325744 , n325745 , n325746 , n325747 , n325748 , n325749 , n325750 , n325751 , n325752 , 
 n325753 , n325754 , n325755 , n5908 , n5909 , n325758 , n325759 , n5912 , n325761 , n325762 , 
 n325763 , n325764 , n325765 , n325766 , n5919 , n325768 , n5921 , n325770 , n325771 , n5924 , 
 n5925 , n325774 , n325775 , n325776 , n325777 , n5930 , n325779 , n325780 , n5933 , n325782 , 
 n325783 , n5936 , n325785 , n5938 , n5939 , n5940 , n325789 , n5942 , n325791 , n325792 , 
 n325793 , n325794 , n5947 , n5948 , n5949 , n5950 , n325799 , n325800 , n5953 , n325802 , 
 n5955 , n325804 , n325805 , n325806 , n325807 , n325808 , n325809 , n5962 , n325811 , n325812 , 
 n5965 , n325814 , n325815 , n325816 , n325817 , n325818 , n325819 , n325820 , n5973 , n325822 , 
 n325823 , n325824 , n5977 , n325826 , n325827 , n5980 , n325829 , n325830 , n325831 , n325832 , 
 n325833 , n325834 , n325835 , n325836 , n325837 , n5990 , n325839 , n325840 , n5993 , n325842 , 
 n5995 , n5996 , n325845 , n325846 , n325847 , n6000 , n325849 , n325850 , n325851 , n325852 , 
 n325853 , n325854 , n6007 , n325856 , n325857 , n325858 , n325859 , n325860 , n6013 , n325862 , 
 n6015 , n325864 , n325865 , n6018 , n325867 , n325868 , n6021 , n6022 , n325871 , n325872 , 
 n6025 , n6026 , n325875 , n325876 , n325877 , n325878 , n325879 , n325880 , n325881 , n325882 , 
 n325883 , n325884 , n325885 , n6038 , n325887 , n325888 , n6041 , n325890 , n325891 , n325892 , 
 n6045 , n6046 , n6047 , n325896 , n325897 , n325898 , n325899 , n6052 , n325901 , n325902 , 
 n325903 , n325904 , n325905 , n325906 , n325907 , n325908 , n6061 , n6062 , n325911 , n6064 , 
 n325913 , n325914 , n6067 , n325916 , n325917 , n6070 , n325919 , n325920 , n325921 , n6074 , 
 n325923 , n325924 , n6077 , n325926 , n6079 , n325928 , n6081 , n325930 , n325931 , n6084 , 
 n325933 , n325934 , n325935 , n325936 , n325937 , n325938 , n325939 , n325940 , n325941 , n325942 , 
 n325943 , n325944 , n325945 , n325946 , n325947 , n325948 , n6101 , n325950 , n325951 , n325952 , 
 n325953 , n6106 , n325955 , n325956 , n325957 , n325958 , n325959 , n325960 , n325961 , n325962 , 
 n6115 , n325964 , n6117 , n6118 , n325967 , n6120 , n6121 , n325970 , n6123 , n325972 , 
 n6125 , n6126 , n325975 , n325976 , n325977 , n325978 , n6131 , n325980 , n6133 , n6134 , 
 n6135 , n325984 , n6137 , n325986 , n325987 , n325988 , n6141 , n325990 , n325991 , n325992 , 
 n325993 , n325994 , n325995 , n6148 , n325997 , n325998 , n325999 , n326000 , n326001 , n6154 , 
 n326003 , n6156 , n6157 , n326006 , n326007 , n6160 , n326009 , n326010 , n6163 , n326012 , 
 n326013 , n6166 , n6167 , n6168 , n326017 , n326018 , n6171 , n326020 , n6173 , n326022 , 
 n6175 , n6176 , n326025 , n326026 , n6179 , n326028 , n326029 , n6182 , n326031 , n6184 , 
 n326033 , n326034 , n326035 , n326036 , n326037 , n6190 , n326039 , n6192 , n6193 , n326042 , 
 n326043 , n326044 , n326045 , n326046 , n6199 , n326048 , n6201 , n326050 , n6203 , n6204 , 
 n6205 , n326054 , n326055 , n6208 , n326057 , n6210 , n326059 , n326060 , n6213 , n6214 , 
 n326063 , n326064 , n6217 , n326066 , n6219 , n326068 , n326069 , n6222 , n326071 , n326072 , 
 n326073 , n6226 , n326075 , n326076 , n326077 , n326078 , n326079 , n326080 , n326081 , n6234 , 
 n326083 , n6236 , n326085 , n6238 , n6239 , n326088 , n326089 , n6242 , n326091 , n326092 , 
 n326093 , n326094 , n326095 , n326096 , n6249 , n6250 , n326099 , n6252 , n326101 , n6254 , 
 n6255 , n6256 , n326105 , n6258 , n326107 , n326108 , n6261 , n326110 , n6263 , n326112 , 
 n6265 , n326114 , n6267 , n326116 , n6269 , n6270 , n326119 , n326120 , n326121 , n6274 , 
 n326123 , n326124 , n326125 , n326126 , n326127 , n6280 , n326129 , n6282 , n326131 , n326132 , 
 n326133 , n326134 , n6287 , n326136 , n326137 , n6290 , n326139 , n6292 , n326141 , n6294 , 
 n6295 , n6296 , n326145 , n326146 , n326147 , n326148 , n326149 , n326150 , n326151 , n6304 , 
 n326153 , n326154 , n6307 , n6308 , n326157 , n6310 , n326159 , n6312 , n6313 , n326162 , 
 n326163 , n326164 , n326165 , n326166 , n326167 , n326168 , n326169 , n326170 , n326171 , n326172 , 
 n326173 , n326174 , n6327 , n6328 , n6329 , n326178 , n6331 , n6332 , n6333 , n6334 , 
 n326183 , n326184 , n326185 , n326186 , n326187 , n326188 , n326189 , n6342 , n326191 , n326192 , 
 n6345 , n326194 , n6347 , n326196 , n6349 , n326198 , n326199 , n6352 , n326201 , n326202 , 
 n326203 , n326204 , n326205 , n326206 , n326207 , n6360 , n326209 , n326210 , n326211 , n326212 , 
 n326213 , n326214 , n326215 , n326216 , n326217 , n6370 , n6371 , n326220 , n326221 , n326222 , 
 n326223 , n6376 , n326225 , n326226 , n326227 , n326228 , n6381 , n326230 , n326231 , n6384 , 
 n326233 , n6386 , n326235 , n326236 , n6389 , n326238 , n6391 , n326240 , n326241 , n326242 , 
 n326243 , n6396 , n326245 , n6398 , n6399 , n326248 , n6401 , n326250 , n326251 , n6404 , 
 n326253 , n6406 , n6407 , n6408 , n326257 , n326258 , n326259 , n6412 , n326261 , n326262 , 
 n326263 , n326264 , n326265 , n6418 , n326267 , n326268 , n6421 , n326270 , n326271 , n326272 , 
 n6425 , n326274 , n6427 , n326276 , n326277 , n326278 , n6431 , n326280 , n326281 , n6434 , 
 n326283 , n326284 , n6437 , n326286 , n6439 , n6440 , n6441 , n326290 , n326291 , n6444 , 
 n6445 , n6446 , n6447 , n6448 , n6449 , n326298 , n6451 , n326300 , n326301 , n6454 , 
 n326303 , n6456 , n326305 , n326306 , n6459 , n6460 , n6461 , n6462 , n326311 , n6464 , 
 n326313 , n6466 , n326315 , n6468 , n6469 , n6470 , n6471 , n6472 , n326321 , n6474 , 
 n326323 , n326324 , n326325 , n6478 , n6479 , n326328 , n6481 , n6482 , n326331 , n326332 , 
 n326333 , n6486 , n326335 , n326336 , n6489 , n326338 , n326339 , n6492 , n326341 , n326342 , 
 n326343 , n6496 , n326345 , n6498 , n6499 , n6500 , n326349 , n326350 , n6503 , n326352 , 
 n326353 , n326354 , n326355 , n326356 , n326357 , n326358 , n326359 , n6512 , n326361 , n326362 , 
 n6515 , n326364 , n326365 , n326366 , n326367 , n6520 , n6521 , n326370 , n326371 , n6524 , 
 n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n326379 , n326380 , n326381 , n326382 , 
 n326383 , n326384 , n326385 , n326386 , n6539 , n326388 , n326389 , n6542 , n326391 , n326392 , 
 n326393 , n326394 , n326395 , n326396 , n326397 , n326398 , n326399 , n6552 , n326401 , n326402 , 
 n6555 , n326404 , n326405 , n6558 , n326407 , n326408 , n6561 , n326410 , n326411 , n326412 , 
 n326413 , n326414 , n6567 , n326416 , n326417 , n326418 , n6571 , n6572 , n326421 , n326422 , 
 n326423 , n6576 , n6577 , n326426 , n326427 , n326428 , n326429 , n6582 , n326431 , n326432 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n326439 , n6592 , n6593 , n326442 , 
 n326443 , n326444 , n326445 , n6598 , n326447 , n326448 , n326449 , n6602 , n326451 , n6604 , 
 n6605 , n326454 , n326455 , n326456 , n6609 , n326458 , n326459 , n6612 , n326461 , n326462 , 
 n326463 , n326464 , n6617 , n326466 , n6619 , n326468 , n326469 , n6622 , n326471 , n326472 , 
 n326473 , n326474 , n326475 , n326476 , n6629 , n326478 , n326479 , n6632 , n326481 , n326482 , 
 n326483 , n6636 , n326485 , n6638 , n326487 , n6640 , n6641 , n6642 , n326491 , n326492 , 
 n6645 , n6646 , n326495 , n6648 , n326497 , n326498 , n326499 , n6652 , n326501 , n326502 , 
 n326503 , n6656 , n6657 , n326506 , n326507 , n326508 , n326509 , n6662 , n6663 , n6664 , 
 n326513 , n326514 , n6667 , n326516 , n6669 , n326518 , n6671 , n6672 , n6673 , n326522 , 
 n6675 , n6676 , n6677 , n6678 , n326527 , n6680 , n326529 , n326530 , n326531 , n6684 , 
 n326533 , n326534 , n326535 , n326536 , n326537 , n6690 , n6691 , n326540 , n6693 , n326542 , 
 n326543 , n326544 , n326545 , n326546 , n326547 , n326548 , n326549 , n326550 , n326551 , n326552 , 
 n6705 , n326554 , n6707 , n6708 , n6709 , n6710 , n6711 , n326560 , n326561 , n326562 , 
 n326563 , n326564 , n6717 , n326566 , n6719 , n326568 , n326569 , n326570 , n326571 , n326572 , 
 n6725 , n326574 , n326575 , n326576 , n326577 , n326578 , n326579 , n326580 , n326581 , n6734 , 
 n326583 , n6736 , n326585 , n6738 , n326587 , n6740 , n326589 , n6742 , n326591 , n326592 , 
 n6745 , n326594 , n326595 , n6748 , n6749 , n6750 , n326599 , n6752 , n326601 , n6754 , 
 n326603 , n326604 , n6757 , n6758 , n326607 , n326608 , n6761 , n326610 , n326611 , n326612 , 
 n6765 , n326614 , n326615 , n326616 , n326617 , n326618 , n6771 , n326620 , n326621 , n6774 , 
 n326623 , n6776 , n6777 , n326626 , n326627 , n326628 , n6781 , n326630 , n326631 , n6784 , 
 n326633 , n326634 , n6787 , n326636 , n326637 , n326638 , n326639 , n6792 , n6793 , n6794 , 
 n326643 , n326644 , n326645 , n326646 , n6799 , n326648 , n326649 , n6802 , n6803 , n6804 , 
 n326653 , n326654 , n6807 , n326656 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n326664 , n326665 , n326666 , n326667 , n326668 , n326669 , n326670 , n326671 , n326672 , 
 n326673 , n326674 , n326675 , n6828 , n326677 , n326678 , n326679 , n6832 , n326681 , n326682 , 
 n326683 , n326684 , n326685 , n6838 , n326687 , n326688 , n6841 , n326690 , n6843 , n6844 , 
 n326693 , n326694 , n326695 , n6848 , n6849 , n326698 , n6851 , n326700 , n326701 , n6854 , 
 n326703 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n326712 , 
 n6865 , n326714 , n6867 , n326716 , n6869 , n326718 , n326719 , n6872 , n6873 , n6874 , 
 n6875 , n326724 , n326725 , n6878 , n326727 , n326728 , n6881 , n326730 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n326739 , n6892 , n326741 , n326742 , 
 n326743 , n326744 , n326745 , n326746 , n326747 , n326748 , n6901 , n326750 , n326751 , n6904 , 
 n326753 , n326754 , n6907 , n326756 , n326757 , n6910 , n326759 , n326760 , n6913 , n6914 , 
 n326763 , n6916 , n326765 , n6918 , n6919 , n326768 , n6921 , n326770 , n6923 , n6924 , 
 n326773 , n326774 , n326775 , n6928 , n326777 , n326778 , n6931 , n326780 , n326781 , n6934 , 
 n326783 , n326784 , n6937 , n326786 , n326787 , n6940 , n326789 , n326790 , n326791 , n6944 , 
 n326793 , n6946 , n6947 , n326796 , n326797 , n326798 , n6951 , n326800 , n326801 , n6954 , 
 n326803 , n326804 , n6957 , n326806 , n326807 , n326808 , n326809 , n6962 , n326811 , n6964 , 
 n326813 , n326814 , n6967 , n326816 , n6969 , n326818 , n6971 , n6972 , n326821 , n326822 , 
 n326823 , n6976 , n326825 , n326826 , n6979 , n326828 , n326829 , n6982 , n326831 , n326832 , 
 n6985 , n326834 , n326835 , n6988 , n326837 , n326838 , n6991 , n326840 , n6993 , n6994 , 
 n326843 , n326844 , n6997 , n326846 , n6999 , n326848 , n326849 , n7002 , n326851 , n326852 , 
 n7005 , n326854 , n326855 , n7008 , n326857 , n326858 , n326859 , n7012 , n326861 , n7014 , 
 n7015 , n326864 , n326865 , n326866 , n7019 , n326868 , n326869 , n7022 , n326871 , n326872 , 
 n7025 , n326874 , n326875 , n7028 , n326877 , n7030 , n7031 , n326880 , n7033 , n7034 , 
 n326883 , n326884 , n326885 , n7038 , n326887 , n326888 , n7041 , n326890 , n326891 , n7044 , 
 n326893 , n326894 , n7047 , n326896 , n326897 , n7050 , n326899 , n326900 , n7053 , n326902 , 
 n326903 , n7056 , n7057 , n7058 , n7059 , n7060 , n326909 , n326910 , n7063 , n326912 , 
 n326913 , n7066 , n326915 , n326916 , n7069 , n7070 , n326919 , n7072 , n7073 , n326922 , 
 n326923 , n7076 , n326925 , n326926 , n7079 , n7080 , n7081 , n7082 , n7083 , n326932 , 
 n326933 , n7086 , n7087 , n326936 , n326937 , n7090 , n326939 , n326940 , n7093 , n326942 , 
 n326943 , n7096 , n326945 , n326946 , n7099 , n326948 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n326959 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n326965 , n326966 , n326967 , n7120 , n326969 , n7122 , n7123 , n326972 , 
 n326973 , n326974 , n7127 , n326976 , n326977 , n7130 , n326979 , n326980 , n7133 , n326982 , 
 n7135 , n7136 , n7137 , n326986 , n326987 , n7140 , n326989 , n7142 , n7143 , n326992 , 
 n7145 , n326994 , n7147 , n7148 , n326997 , n326998 , n326999 , n7152 , n327001 , n327002 , 
 n7155 , n327004 , n327005 , n7158 , n327007 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n327013 , n7166 , n7167 , n7168 , n7169 , n7170 , n327019 , n327020 , n7173 , n327022 , 
 n327023 , n7176 , n7177 , n7178 , n7179 , n327028 , n327029 , n7182 , n327031 , n327032 , 
 n7185 , n327034 , n327035 , n327036 , n7189 , n327038 , n7191 , n7192 , n327041 , n327042 , 
 n327043 , n7196 , n327045 , n327046 , n7199 , n327048 , n327049 , n7202 , n327051 , n327052 , 
 n7205 , n327054 , n7207 , n327056 , n7209 , n7210 , n327059 , n327060 , n327061 , n7214 , 
 n327063 , n327064 , n7217 , n327066 , n327067 , n7220 , n327069 , n327070 , n7223 , n327072 , 
 n327073 , n7226 , n327075 , n327076 , n7229 , n7230 , n7231 , n7232 , n327081 , n327082 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n327088 , n327089 , n7242 , n327091 , n327092 , 
 n7245 , n327094 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n327103 , n327104 , n7257 , n7258 , n7259 , n7260 , n327109 , n327110 , n327111 , n7264 , 
 n327113 , n7266 , n7267 , n327116 , n327117 , n327118 , n7271 , n327120 , n327121 , n7274 , 
 n327123 , n327124 , n7277 , n327126 , n327127 , n327128 , n7281 , n327130 , n7283 , n7284 , 
 n327133 , n327134 , n327135 , n7288 , n327137 , n327138 , n7291 , n327140 , n327141 , n7294 , 
 n327143 , n327144 , n7297 , n327146 , n327147 , n7300 , n327149 , n7302 , n327151 , n327152 , 
 n7305 , n327154 , n327155 , n7308 , n327157 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n327164 , n7317 , n327166 , n327167 , n7320 , n327169 , n327170 , n327171 , n7324 , 
 n327173 , n7326 , n7327 , n327176 , n327177 , n327178 , n7331 , n327180 , n327181 , n7334 , 
 n327183 , n327184 , n7337 , n327186 , n327187 , n7340 , n327189 , n7342 , n327191 , n7344 , 
 n7345 , n327194 , n327195 , n327196 , n7349 , n327198 , n327199 , n7352 , n327201 , n327202 , 
 n7355 , n327204 , n327205 , n7358 , n327207 , n327208 , n7361 , n327210 , n327211 , n7364 , 
 n327213 , n327214 , n7367 , n7368 , n7369 , n7370 , n7371 , n327220 , n327221 , n7374 , 
 n327223 , n327224 , n7377 , n7378 , n7379 , n7380 , n327229 , n327230 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n327244 , n7397 , n7398 , n7399 , n7400 , n327249 , n327250 , n7403 , n327252 , 
 n327253 , n7406 , n7407 , n327256 , n7409 , n7410 , n327259 , n327260 , n327261 , n327262 , 
 n7415 , n327264 , n327265 , n327266 , n7419 , n327268 , n7421 , n7422 , n7423 , n327272 , 
 n7425 , n7426 , n7427 , n7428 , n327277 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n327287 , n327288 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n327296 , n327297 , n7450 , n327299 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n327329 , n7482 , n327331 , n327332 , 
 n327333 , n7486 , n327335 , n327336 , n7489 , n327338 , n327339 , n7492 , n7493 , n327342 , 
 n327343 , n7496 , n7497 , n327346 , n7499 , n7500 , n7501 , n7502 , n7503 , n327352 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n327366 , n7519 , n7520 , n7521 , n327370 , n7523 , n7524 , 
 n7525 , n327374 , n327375 , n7528 , n7529 , n7530 , n327379 , n7532 , n7533 , n7534 , 
 n327383 , n327384 , n7537 , n7538 , n7539 , n327388 , n327389 , n7542 , n7543 , n7544 , 
 n327393 , n327394 , n7547 , n7548 , n327397 , n327398 , n7551 , n327400 , n7553 , n7554 , 
 n7555 , n7556 , n327405 , n7558 , n327407 , n327408 , n327409 , n327410 , n327411 , n7564 , 
 n7565 , n327414 , n327415 , n7568 , n327417 , n327418 , n327419 , n327420 , n327421 , n7574 , 
 n327423 , n327424 , n327425 , n327426 , n7579 , n327428 , n327429 , n7582 , n7583 , n327432 , 
 n7585 , n7586 , n327435 , n327436 , n7589 , n7590 , n7591 , n7592 , n7593 , n327442 , 
 n7595 , n7596 , n327445 , n327446 , n327447 , n327448 , n7601 , n7602 , n7603 , n327452 , 
 n7605 , n327454 , n327455 , n327456 , n327457 , n7610 , n7611 , n7612 , n327461 , n7614 , 
 n7615 , n327464 , n327465 , n327466 , n327467 , n327468 , n327469 , n327470 , n327471 , n7624 , 
 n327473 , n327474 , n327475 , n7628 , n327477 , n7630 , n327479 , n327480 , n327481 , n327482 , 
 n327483 , n7636 , n327485 , n7638 , n7639 , n327488 , n7641 , n7642 , n327491 , n327492 , 
 n7645 , n7646 , n327495 , n327496 , n7649 , n7650 , n7651 , n7652 , n327501 , n327502 , 
 n327503 , n7656 , n7657 , n327506 , n7659 , n327508 , n327509 , n327510 , n327511 , n327512 , 
 n327513 , n7666 , n327515 , n327516 , n7669 , n327518 , n327519 , n7672 , n327521 , n327522 , 
 n7675 , n327524 , n327525 , n7678 , n7679 , n327528 , n327529 , n7682 , n327531 , n327532 , 
 n327533 , n327534 , n327535 , n7688 , n327537 , n7690 , n7691 , n7692 , n7693 , n327542 , 
 n327543 , n7696 , n7697 , n327546 , n327547 , n327548 , n327549 , n327550 , n7703 , n327552 , 
 n327553 , n327554 , n327555 , n327556 , n327557 , n327558 , n7711 , n327560 , n327561 , n327562 , 
 n7715 , n327564 , n327565 , n7718 , n327567 , n327568 , n327569 , n7722 , n327571 , n327572 , 
 n7725 , n7726 , n327575 , n7728 , n7729 , n327578 , n327579 , n327580 , n327581 , n327582 , 
 n7735 , n327584 , n327585 , n327586 , n327587 , n7740 , n327589 , n327590 , n327591 , n327592 , 
 n7745 , n327594 , n327595 , n327596 , n7749 , n327598 , n327599 , n327600 , n7753 , n327602 , 
 n327603 , n327604 , n327605 , n327606 , n327607 , n7760 , n7761 , n327610 , n7763 , n327612 , 
 n327613 , n327614 , n7767 , n327616 , n327617 , n7770 , n327619 , n327620 , n7773 , n7774 , 
 n327623 , n7776 , n327625 , n327626 , n7779 , n327628 , n327629 , n7782 , n327631 , n327632 , 
 n7785 , n327634 , n327635 , n327636 , n7789 , n7790 , n327639 , n327640 , n327641 , n7794 , 
 n327643 , n327644 , n7797 , n327646 , n7799 , n7800 , n7801 , n327650 , n7803 , n327652 , 
 n7805 , n327654 , n327655 , n7808 , n327657 , n7810 , n327659 , n7812 , n327661 , n7814 , 
 n7815 , n327664 , n7817 , n327666 , n7819 , n327668 , n327669 , n327670 , n327671 , n7824 , 
 n327673 , n7826 , n7827 , n7828 , n7829 , n327678 , n327679 , n7832 , n327681 , n7834 , 
 n7835 , n7836 , n7837 , n327686 , n7839 , n327688 , n327689 , n327690 , n327691 , n327692 , 
 n7845 , n327694 , n7847 , n327696 , n327697 , n327698 , n327699 , n327700 , n327701 , n7854 , 
 n327703 , n327704 , n327705 , n327706 , n327707 , n7860 , n327709 , n7862 , n327711 , n327712 , 
 n327713 , n327714 , n327715 , n7868 , n327717 , n327718 , n7871 , n7872 , n327721 , n327722 , 
 n7875 , n327724 , n327725 , n327726 , n7879 , n327728 , n327729 , n7882 , n327731 , n327732 , 
 n7885 , n7886 , n327735 , n7888 , n327737 , n327738 , n327739 , n7892 , n327741 , n327742 , 
 n327743 , n7896 , n327745 , n327746 , n327747 , n327748 , n7901 , n327750 , n327751 , n327752 , 
 n327753 , n327754 , n327755 , n327756 , n327757 , n327758 , n7911 , n327760 , n7913 , n7914 , 
 n327763 , n327764 , n327765 , n7918 , n327767 , n327768 , n7921 , n327770 , n327771 , n7924 , 
 n327773 , n327774 , n327775 , n327776 , n327777 , n327778 , n7931 , n327780 , n327781 , n7934 , 
 n327783 , n327784 , n7937 , n327786 , n327787 , n327788 , n327789 , n327790 , n327791 , n7944 , 
 n327793 , n327794 , n7947 , n327796 , n327797 , n327798 , n327799 , n7952 , n327801 , n7954 , 
 n327803 , n7956 , n327805 , n327806 , n327807 , n327808 , n7961 , n327810 , n327811 , n327812 , 
 n7965 , n327814 , n7967 , n327816 , n327817 , n327818 , n327819 , n7972 , n327821 , n327822 , 
 n7975 , n327824 , n327825 , n327826 , n327827 , n327828 , n327829 , n327830 , n7983 , n327832 , 
 n327833 , n7986 , n327835 , n327836 , n327837 , n327838 , n327839 , n327840 , n327841 , n327842 , 
 n327843 , n327844 , n327845 , n327846 , n327847 , n327848 , n327849 , n327850 , n327851 , n8004 , 
 n327853 , n327854 , n327855 , n327856 , n8009 , n327858 , n327859 , n327860 , n8013 , n8014 , 
 n327863 , n8016 , n327865 , n327866 , n327867 , n327868 , n327869 , n327870 , n327871 , n327872 , 
 n327873 , n327874 , n327875 , n327876 , n327877 , n327878 , n327879 , n327880 , n327881 , n327882 , 
 n327883 , n327884 , n327885 , n327886 , n8039 , n8040 , n8041 , n8042 , n327891 , n8044 , 
 n327893 , n8046 , n327895 , n327896 , n8049 , n327898 , n327899 , n8052 , n327901 , n327902 , 
 n327903 , n8056 , n327905 , n8058 , n327907 , n327908 , n327909 , n327910 , n327911 , n8064 , 
 n327913 , n327914 , n8067 , n327916 , n8069 , n327918 , n8071 , n8072 , n327921 , n327922 , 
 n327923 , n327924 , n327925 , n327926 , n8079 , n327928 , n327929 , n327930 , n327931 , n327932 , 
 n327933 , n327934 , n8087 , n327936 , n8089 , n8090 , n327939 , n8092 , n8093 , n8094 , 
 n327943 , n327944 , n327945 , n327946 , n8099 , n327948 , n327949 , n8102 , n327951 , n8104 , 
 n327953 , n327954 , n8107 , n327956 , n327957 , n8110 , n8111 , n8112 , n8113 , n327962 , 
 n327963 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n327974 , n8127 , n327976 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n327984 , n8137 , n327986 , n8139 , n327988 , n8141 , n327990 , n8143 , n8144 , 
 n327993 , n327994 , n327995 , n8148 , n327997 , n327998 , n8151 , n328000 , n328001 , n8154 , 
 n328003 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n328019 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n328026 , n328027 , n8180 , n328029 , n8182 , n8183 , n328032 , 
 n328033 , n8186 , n328035 , n8188 , n328037 , n328038 , n328039 , n8192 , n328041 , n328042 , 
 n8195 , n328044 , n8197 , n8198 , n328047 , n328048 , n328049 , n8202 , n328051 , n328052 , 
 n8205 , n328054 , n8207 , n8208 , n8209 , n8210 , n8211 , n328060 , n328061 , n328062 , 
 n8215 , n328064 , n328065 , n8218 , n328067 , n8220 , n8221 , n328070 , n8223 , n328072 , 
 n328073 , n8226 , n328075 , n328076 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n328088 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n328098 , n328099 , n328100 , n8253 , n328102 , 
 n8255 , n328104 , n328105 , n328106 , n328107 , n8260 , n328109 , n328110 , n328111 , n8264 , 
 n328113 , n328114 , n328115 , n8268 , n328117 , n8270 , n8271 , n328120 , n328121 , n8274 , 
 n328123 , n328124 , n328125 , n8278 , n328127 , n328128 , n8281 , n328130 , n328131 , n8284 , 
 n328133 , n328134 , n328135 , n8288 , n328137 , n8290 , n8291 , n328140 , n8293 , n328142 , 
 n328143 , n8296 , n328145 , n8298 , n328147 , n328148 , n8301 , n328150 , n328151 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n328157 , n328158 , n8311 , n328160 , n328161 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n328167 , n328168 , n8321 , n328170 , n328171 , n8324 , 
 n328173 , n328174 , n8327 , n328176 , n328177 , n8330 , n328179 , n328180 , n8333 , n8334 , 
 n8335 , n8336 , n328185 , n328186 , n8339 , n328188 , n8341 , n328190 , n8343 , n328192 , 
 n328193 , n328194 , n8347 , n328196 , n328197 , n8350 , n328199 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8559 , n328408 , n8561 , n8562 , n8563 , n8564 , 
 n8565 , n8566 , n328415 , n328416 , n328417 , n8570 , n328419 , n328420 , n328421 , n8574 , 
 n328423 , n328424 , n8577 , n328426 , n328427 , n8580 , n328429 , n328430 , n8583 , n328432 , 
 n328433 , n8586 , n328435 , n328436 , n328437 , n8590 , n328439 , n8592 , n328441 , n8594 , 
 n328443 , n328444 , n8597 , n8598 , n328447 , n8600 , n328449 , n8602 , n328451 , n328452 , 
 n8605 , n328454 , n328455 , n8608 , n8609 , n328458 , n8611 , n328460 , n8613 , n8614 , 
 n328463 , n328464 , n8617 , n328466 , n328467 , n8620 , n328469 , n328470 , n328471 , n8624 , 
 n328473 , n328474 , n8627 , n328476 , n328477 , n8630 , n8631 , n328480 , n328481 , n8634 , 
 n328483 , n8636 , n328485 , n8638 , n8639 , n328488 , n8641 , n8642 , n328491 , n328492 , 
 n8645 , n328494 , n328495 , n8648 , n328497 , n328498 , n8651 , n8652 , n328501 , n8654 , 
 n328503 , n8656 , n8657 , n328506 , n328507 , n8660 , n328509 , n328510 , n8663 , n328512 , 
 n328513 , n328514 , n8667 , n328516 , n328517 , n8670 , n328519 , n328520 , n8673 , n8674 , 
 n8675 , n328524 , n328525 , n328526 , n8679 , n328528 , n8681 , n328530 , n8683 , n328532 , 
 n328533 , n8686 , n8687 , n328536 , n328537 , n8690 , n328539 , n328540 , n8693 , n328542 , 
 n328543 , n8696 , n8697 , n328546 , n8699 , n328548 , n8701 , n8702 , n328551 , n328552 , 
 n8705 , n328554 , n328555 , n8708 , n328557 , n328558 , n328559 , n8712 , n328561 , n328562 , 
 n8715 , n328564 , n328565 , n8718 , n328567 , n8720 , n328569 , n8722 , n8723 , n328572 , 
 n328573 , n8726 , n328575 , n328576 , n8729 , n328578 , n328579 , n328580 , n8733 , n328582 , 
 n8735 , n8736 , n328585 , n328586 , n8739 , n328588 , n328589 , n8742 , n328591 , n328592 , 
 n8745 , n8746 , n8747 , n328596 , n328597 , n8750 , n328599 , n328600 , n8753 , n8754 , 
 n8755 , n328604 , n328605 , n8758 , n8759 , n8760 , n8761 , n8762 , n328611 , n328612 , 
 n8765 , n8766 , n328615 , n328616 , n8769 , n328618 , n8771 , n328620 , n8773 , n8774 , 
 n328623 , n328624 , n8777 , n328626 , n328627 , n8780 , n328629 , n328630 , n8783 , n328632 , 
 n328633 , n8786 , n8787 , n8788 , n328637 , n328638 , n8791 , n8792 , n8793 , n8794 , 
 n8795 , n328644 , n328645 , n328646 , n8799 , n8800 , n8801 , n8802 , n8803 , n328652 , 
 n328653 , n328654 , n8807 , n328656 , n8809 , n328658 , n328659 , n8812 , n328661 , n8814 , 
 n8815 , n328664 , n328665 , n8818 , n328667 , n8820 , n328669 , n328670 , n8823 , n328672 , 
 n8825 , n8826 , n328675 , n8828 , n328677 , n8830 , n8831 , n328680 , n8833 , n328682 , 
 n8835 , n8836 , n328685 , n328686 , n8839 , n328688 , n8841 , n8842 , n8843 , n328692 , 
 n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n328702 , 
 n8855 , n328704 , n8857 , n8858 , n8859 , n8860 , n328709 , n8862 , n328711 , n328712 , 
 n8865 , n328714 , n328715 , n8868 , n8869 , n328718 , n328719 , n8872 , n328721 , n328722 , 
 n328723 , n8876 , n328725 , n8878 , n8879 , n328728 , n8881 , n328730 , n8883 , n8884 , 
 n328733 , n8886 , n328735 , n8888 , n8889 , n328738 , n328739 , n328740 , n8893 , n328742 , 
 n328743 , n8896 , n328745 , n328746 , n8899 , n328748 , n8901 , n8902 , n8903 , n8904 , 
 n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n328759 , n328760 , n328761 , n8914 , 
 n328763 , n328764 , n8917 , n328766 , n8919 , n328768 , n8921 , n328770 , n8923 , n8924 , 
 n328773 , n328774 , n328775 , n8928 , n328777 , n328778 , n8931 , n328780 , n328781 , n8934 , 
 n328783 , n8936 , n328785 , n8938 , n328787 , n8940 , n8941 , n328790 , n328791 , n328792 , 
 n8945 , n328794 , n328795 , n8948 , n328797 , n328798 , n8951 , n328800 , n8953 , n328802 , 
 n8955 , n328804 , n8957 , n8958 , n328807 , n328808 , n8961 , n328810 , n8963 , n328812 , 
 n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n328822 , 
 n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n328832 , 
 n8985 , n328834 , n8987 , n328836 , n8989 , n8990 , n328839 , n328840 , n328841 , n8994 , 
 n328843 , n328844 , n8997 , n328846 , n328847 , n9000 , n328849 , n328850 , n9003 , n328852 , 
 n328853 , n9006 , n328855 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , 
 n328863 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , 
 n328873 , n328874 , n9027 , n328876 , n328877 , n9030 , n328879 , n9032 , n9033 , n328882 , 
 n328883 , n9036 , n328885 , n9038 , n328887 , n328888 , n9041 , n328890 , n9043 , n328892 , 
 n9045 , n328894 , n328895 , n9048 , n328897 , n328898 , n9051 , n9052 , n328901 , n9054 , 
 n328903 , n9056 , n328905 , n328906 , n9059 , n328908 , n9061 , n9062 , n9063 , n328912 , 
 n328913 , n328914 , n9067 , n328916 , n328917 , n9070 , n328919 , n9072 , n9073 , n9074 , 
 n9075 , n9076 , n328925 , n9078 , n328927 , n9080 , n328929 , n9082 , n9083 , n328932 , 
 n9085 , n328934 , n9087 , n9088 , n328937 , n328938 , n9091 , n328940 , n328941 , n9094 , 
 n328943 , n328944 , n328945 , n9098 , n328947 , n9100 , n328949 , n9102 , n328951 , n9104 , 
 n9105 , n328954 , n328955 , n9108 , n328957 , n328958 , n328959 , n9112 , n328961 , n328962 , 
 n9115 , n328964 , n9117 , n9118 , n9119 , n328968 , n9121 , n328970 , n9123 , n9124 , 
 n328973 , n328974 , n328975 , n9128 , n328977 , n328978 , n9131 , n328980 , n328981 , n9134 , 
 n328983 , n328984 , n328985 , n9138 , n328987 , n9140 , n9141 , n328990 , n328991 , n328992 , 
 n9145 , n328994 , n328995 , n9148 , n328997 , n328998 , n9151 , n329000 , n329001 , n9154 , 
 n329003 , n9156 , n329005 , n9158 , n9159 , n329008 , n329009 , n329010 , n9163 , n329012 , 
 n329013 , n9166 , n329015 , n329016 , n9169 , n329018 , n329019 , n9172 , n329021 , n329022 , 
 n9175 , n329024 , n9177 , n329026 , n9179 , n9180 , n9181 , n9182 , n329031 , n329032 , 
 n9185 , n9186 , n9187 , n9188 , n9189 , n329038 , n329039 , n329040 , n9193 , n329042 , 
 n9195 , n9196 , n329045 , n9198 , n329047 , n329048 , n329049 , n9202 , n329051 , n9204 , 
 n329053 , n329054 , n9207 , n329056 , n329057 , n9210 , n9211 , n329060 , n329061 , n9214 , 
 n9215 , n9216 , n9217 , n329066 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , 
 n9225 , n329074 , n9227 , n329076 , n329077 , n9230 , n329079 , n329080 , n9233 , n329082 , 
 n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , 
 n329093 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n329100 , n9253 , n329102 , 
 n329103 , n9256 , n329105 , n329106 , n329107 , n9260 , n329109 , n329110 , n9263 , n9264 , 
 n329113 , n329114 , n9267 , n329116 , n329117 , n9270 , n329119 , n9272 , n329121 , n329122 , 
 n9275 , n329124 , n329125 , n9278 , n329127 , n329128 , n329129 , n329130 , n9283 , n329132 , 
 n9285 , n329134 , n329135 , n329136 , n329137 , n329138 , n9291 , n329140 , n329141 , n9294 , 
 n329143 , n329144 , n9297 , n329146 , n329147 , n9300 , n329149 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n329378 , n9531 , n9532 , n329381 , n329382 , 
 n9535 , n329384 , n329385 , n9538 , n329387 , n329388 , n9541 , n329390 , n9543 , n329392 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n329537 , n329538 , n329539 , n329540 , n9693 , n329542 , 
 n329543 , n9696 , n9697 , n329546 , n329547 , n9700 , n329549 , n9702 , n9703 , n9704 , 
 n9705 , n329554 , n9707 , n329556 , n329557 , n9710 , n329559 , n329560 , n9713 , n329562 , 
 n9715 , n329564 , n9717 , n9718 , n329567 , n329568 , n329569 , n9722 , n329571 , n329572 , 
 n9725 , n329574 , n329575 , n9728 , n329577 , n329578 , n9731 , n329580 , n9733 , n9734 , 
 n329583 , n329584 , n329585 , n9738 , n329587 , n329588 , n9741 , n329590 , n329591 , n9744 , 
 n329593 , n9746 , n329595 , n9748 , n329597 , n9750 , n9751 , n329600 , n9753 , n329602 , 
 n9755 , n329604 , n329605 , n9758 , n329607 , n9760 , n9761 , n9762 , n9763 , n9764 , 
 n329613 , n9766 , n9767 , n9768 , n9769 , n329618 , n9771 , n329620 , n329621 , n9774 , 
 n9775 , n9776 , n9777 , n329626 , n9779 , n329628 , n329629 , n9782 , n9783 , n329632 , 
 n9785 , n9786 , n329635 , n9788 , n9789 , n329638 , n9791 , n329640 , n9793 , n9794 , 
 n329643 , n9796 , n9797 , n9798 , n329647 , n9800 , n9801 , n329650 , n329651 , n329652 , 
 n9805 , n329654 , n329655 , n9808 , n329657 , n329658 , n9811 , n329660 , n329661 , n9814 , 
 n329663 , n9816 , n9817 , n329666 , n329667 , n329668 , n9821 , n329670 , n329671 , n9824 , 
 n329673 , n329674 , n9827 , n329676 , n9829 , n329678 , n9831 , n329680 , n9833 , n9834 , 
 n329683 , n329684 , n329685 , n9838 , n329687 , n329688 , n9841 , n329690 , n329691 , n9844 , 
 n329693 , n9846 , n329695 , n9848 , n329697 , n329698 , n9851 , n329700 , n329701 , n9854 , 
 n9855 , n329704 , n329705 , n9858 , n329707 , n329708 , n9861 , n329710 , n329711 , n9864 , 
 n9865 , n329714 , n9867 , n329716 , n9869 , n329718 , n329719 , n9872 , n9873 , n9874 , 
 n9875 , n9876 , n329725 , n329726 , n9879 , n329728 , n9881 , n9882 , n9883 , n9884 , 
 n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n329739 , n9892 , n329741 , n9894 , 
 n329743 , n329744 , n9897 , n329746 , n9899 , n9900 , n329749 , n329750 , n9903 , n329752 , 
 n9905 , n329754 , n329755 , n9908 , n329757 , n329758 , n9911 , n329760 , n9913 , n329762 , 
 n9915 , n9916 , n329765 , n329766 , n9919 , n329768 , n9921 , n329770 , n329771 , n9924 , 
 n329773 , n329774 , n9927 , n9928 , n9929 , n9930 , n329779 , n329780 , n9933 , n329782 , 
 n329783 , n9936 , n329785 , n329786 , n329787 , n9940 , n329789 , n9942 , n329791 , n329792 , 
 n9945 , n329794 , n329795 , n9948 , n9949 , n329798 , n9951 , n329800 , n329801 , n9954 , 
 n329803 , n9956 , n329805 , n329806 , n9959 , n329808 , n329809 , n9962 , n329811 , n329812 , 
 n329813 , n9966 , n329815 , n9968 , n9969 , n329818 , n9971 , n329820 , n9973 , n329822 , 
 n329823 , n9976 , n329825 , n329826 , n9979 , n329828 , n329829 , n9982 , n329831 , n9984 , 
 n9985 , n329834 , n329835 , n329836 , n9989 , n329838 , n329839 , n9992 , n329841 , n329842 , 
 n9995 , n329844 , n9997 , n9998 , n9999 , n10000 , n329849 , n329850 , n10003 , n329852 , 
 n329853 , n329854 , n10007 , n329856 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , 
 n10015 , n329864 , n10017 , n10018 , n10019 , n10020 , n10021 , n329870 , n329871 , n10024 , 
 n329873 , n329874 , n10027 , n10028 , n10029 , n10030 , n329879 , n329880 , n10033 , n329882 , 
 n10035 , n329884 , n10037 , n10038 , n329887 , n10040 , n329889 , n10042 , n329891 , n329892 , 
 n10045 , n329894 , n329895 , n329896 , n10049 , n329898 , n10051 , n10052 , n329901 , n10054 , 
 n329903 , n10056 , n329905 , n329906 , n10059 , n329908 , n329909 , n10062 , n329911 , n10064 , 
 n329913 , n10066 , n10067 , n329916 , n10069 , n329918 , n10071 , n329920 , n329921 , n10074 , 
 n329923 , n329924 , n10077 , n329926 , n329927 , n10080 , n329929 , n329930 , n329931 , n10084 , 
 n329933 , n10086 , n329935 , n329936 , n10089 , n10090 , n10091 , n10092 , n329941 , n10094 , 
 n329943 , n329944 , n10097 , n329946 , n10099 , n329948 , n10101 , n329950 , n10103 , n329952 , 
 n329953 , n10106 , n10107 , n329956 , n10109 , n329958 , n10111 , n329960 , n329961 , n10114 , 
 n329963 , n329964 , n329965 , n329966 , n10119 , n329968 , n10121 , n329970 , n329971 , n329972 , 
 n329973 , n10126 , n329975 , n329976 , n10129 , n329978 , n329979 , n10132 , n10133 , n10134 , 
 n10135 , n329984 , n329985 , n10138 , n329987 , n329988 , n10141 , n329990 , n10143 , n10144 , 
 n329993 , n10146 , n329995 , n329996 , n10149 , n329998 , n329999 , n10152 , n330001 , n330002 , 
 n10155 , n330004 , n330005 , n10158 , n330007 , n10160 , n10161 , n10162 , n10163 , n10164 , 
 n10165 , n10166 , n10167 , n10168 , n330017 , n330018 , n10171 , n330020 , n10173 , n10174 , 
 n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , 
 n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , 
 n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , 
 n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , 
 n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , 
 n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , 
 n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , 
 n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , 
 n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , 
 n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , 
 n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , 
 n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , 
 n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , 
 n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , 
 n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , 
 n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n330182 , 
 n10335 , n330184 , n10337 , n330186 , n330187 , n10340 , n330189 , n330190 , n330191 , n10344 , 
 n330193 , n10346 , n10347 , n330196 , n10349 , n330198 , n10351 , n330200 , n330201 , n10354 , 
 n330203 , n330204 , n10357 , n330206 , n10359 , n330208 , n10361 , n10362 , n330211 , n330212 , 
 n330213 , n10366 , n330215 , n330216 , n10369 , n330218 , n330219 , n10372 , n330221 , n330222 , 
 n10375 , n330224 , n330225 , n330226 , n10379 , n10380 , n330229 , n10382 , n10383 , n330232 , 
 n330233 , n330234 , n10387 , n330236 , n330237 , n10390 , n330239 , n330240 , n10393 , n330242 , 
 n330243 , n330244 , n10397 , n330246 , n10399 , n330248 , n10401 , n10402 , n330251 , n330252 , 
 n10405 , n330254 , n330255 , n10408 , n330257 , n330258 , n10411 , n330260 , n330261 , n10414 , 
 n330263 , n330264 , n10417 , n10418 , n10419 , n10420 , n10421 , n330270 , n330271 , n10424 , 
 n330273 , n330274 , n330275 , n10428 , n330277 , n10430 , n330279 , n330280 , n10433 , n10434 , 
 n330283 , n10436 , n330285 , n330286 , n330287 , n10440 , n330289 , n10442 , n330291 , n330292 , 
 n10445 , n330294 , n330295 , n10448 , n330297 , n330298 , n10451 , n330300 , n330301 , n330302 , 
 n10455 , n330304 , n330305 , n10458 , n330307 , n330308 , n10461 , n330310 , n330311 , n330312 , 
 n330313 , n10466 , n330315 , n10468 , n10469 , n10470 , n10471 , n10472 , n330321 , n330322 , 
 n10475 , n330324 , n10477 , n10478 , n10479 , n10480 , n330329 , n10482 , n330331 , n330332 , 
 n10485 , n330334 , n10487 , n330336 , n10489 , n10490 , n10491 , n10492 , n330341 , n10494 , 
 n330343 , n330344 , n330345 , n10498 , n330347 , n10500 , n10501 , n330350 , n330351 , n330352 , 
 n10505 , n330354 , n330355 , n10508 , n330357 , n330358 , n10511 , n330360 , n330361 , n10514 , 
 n330363 , n10516 , n330365 , n10518 , n10519 , n330368 , n330369 , n330370 , n10523 , n330372 , 
 n330373 , n10526 , n330375 , n330376 , n10529 , n330378 , n330379 , n10532 , n330381 , n330382 , 
 n10535 , n330384 , n330385 , n10538 , n10539 , n10540 , n330389 , n330390 , n330391 , n10544 , 
 n330393 , n330394 , n10547 , n330396 , n330397 , n10550 , n330399 , n330400 , n10553 , n330402 , 
 n330403 , n10556 , n10557 , n10558 , n10559 , n330408 , n330409 , n10562 , n10563 , n330412 , 
 n10565 , n330414 , n10567 , n10568 , n10569 , n10570 , n10571 , n330420 , n10573 , n10574 , 
 n10575 , n10576 , n330425 , n330426 , n10579 , n330428 , n10581 , n330430 , n10583 , n10584 , 
 n330433 , n330434 , n330435 , n10588 , n330437 , n330438 , n10591 , n330440 , n330441 , n10594 , 
 n330443 , n330444 , n330445 , n330446 , n10599 , n330448 , n330449 , n10602 , n330451 , n330452 , 
 n10605 , n10606 , n330455 , n10608 , n10609 , n330458 , n330459 , n10612 , n330461 , n10614 , 
 n10615 , n330464 , n10617 , n330466 , n10619 , n330468 , n330469 , n10622 , n330471 , n10624 , 
 n330473 , n330474 , n10627 , n330476 , n10629 , n10630 , n330479 , n330480 , n330481 , n10634 , 
 n330483 , n330484 , n10637 , n330486 , n330487 , n10640 , n330489 , n330490 , n330491 , n10644 , 
 n330493 , n10646 , n10647 , n330496 , n330497 , n10650 , n330499 , n330500 , n10653 , n330502 , 
 n330503 , n10656 , n330505 , n330506 , n10659 , n330508 , n10661 , n330510 , n330511 , n10664 , 
 n10665 , n10666 , n10667 , n10668 , n330517 , n330518 , n10671 , n330520 , n330521 , n10674 , 
 n10675 , n10676 , n10677 , n330526 , n330527 , n10680 , n10681 , n10682 , n10683 , n10684 , 
 n330533 , n330534 , n10687 , n10688 , n10689 , n10690 , n330539 , n330540 , n330541 , n10694 , 
 n330543 , n10696 , n10697 , n330546 , n10699 , n330548 , n10701 , n10702 , n330551 , n10704 , 
 n330553 , n330554 , n10707 , n330556 , n330557 , n10710 , n330559 , n330560 , n10713 , n330562 , 
 n10715 , n10716 , n10717 , n10718 , n10719 , n330568 , n330569 , n10722 , n330571 , n10724 , 
 n10725 , n330574 , n330575 , n330576 , n10729 , n330578 , n330579 , n10732 , n330581 , n330582 , 
 n10735 , n330584 , n330585 , n10738 , n330587 , n10740 , n330589 , n10742 , n10743 , n330592 , 
 n10745 , n330594 , n10747 , n330596 , n330597 , n10750 , n330599 , n330600 , n10753 , n330602 , 
 n330603 , n10756 , n330605 , n330606 , n10759 , n10760 , n10761 , n10762 , n10763 , n330612 , 
 n330613 , n10766 , n330615 , n330616 , n10769 , n330618 , n330619 , n10772 , n330621 , n330622 , 
 n10775 , n330624 , n10777 , n10778 , n10779 , n10780 , n330629 , n10782 , n330631 , n330632 , 
 n10785 , n330634 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , 
 n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , 
 n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , 
 n10815 , n10816 , n10817 , n10818 , n10819 , n330668 , n10821 , n330670 , n10823 , n10824 , 
 n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n330680 , n10833 , n10834 , 
 n330683 , n10836 , n330685 , n10838 , n330687 , n330688 , n10841 , n330690 , n330691 , n10844 , 
 n10845 , n330694 , n10847 , n10848 , n10849 , n10850 , n10851 , n330700 , n10853 , n330702 , 
 n10855 , n10856 , n10857 , n10858 , n330707 , n10860 , n330709 , n330710 , n10863 , n10864 , 
 n330713 , n330714 , n10867 , n330716 , n330717 , n10870 , n330719 , n330720 , n330721 , n330722 , 
 n10875 , n330724 , n330725 , n10878 , n330727 , n330728 , n10881 , n330730 , n330731 , n10884 , 
 n330733 , n330734 , n10887 , n330736 , n330737 , n10890 , n330739 , n330740 , n10893 , n330742 , 
 n330743 , n10896 , n330745 , n10898 , n330747 , n10900 , n10901 , n10902 , n10903 , n10904 , 
 n10905 , n10906 , n330755 , n330756 , n10909 , n330758 , n330759 , n10912 , n330761 , n330762 , 
 n330763 , n10916 , n330765 , n10918 , n10919 , n330768 , n330769 , n10922 , n330771 , n10924 , 
 n10925 , n330774 , n330775 , n10928 , n330777 , n330778 , n10931 , n330780 , n330781 , n10934 , 
 n330783 , n330784 , n10937 , n330786 , n330787 , n10940 , n10941 , n330790 , n330791 , n10944 , 
 n10945 , n330794 , n10947 , n330796 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , 
 n330803 , n330804 , n10957 , n330806 , n330807 , n10960 , n330809 , n330810 , n10963 , n10964 , 
 n10965 , n330814 , n330815 , n10968 , n10969 , n10970 , n330819 , n10972 , n330821 , n10974 , 
 n10975 , n330824 , n330825 , n10978 , n330827 , n330828 , n10981 , n330830 , n330831 , n330832 , 
 n10985 , n330834 , n10987 , n330836 , n10989 , n10990 , n10991 , n330840 , n330841 , n10994 , 
 n10995 , n10996 , n330845 , n330846 , n330847 , n11000 , n330849 , n11002 , n11003 , n11004 , 
 n11005 , n11006 , n11007 , n11008 , n330857 , n11010 , n330859 , n11012 , n11013 , n11014 , 
 n11015 , n330864 , n330865 , n11018 , n330867 , n330868 , n11021 , n330870 , n330871 , n11024 , 
 n11025 , n11026 , n330875 , n330876 , n11029 , n11030 , n11031 , n330880 , n330881 , n11034 , 
 n11035 , n11036 , n330885 , n330886 , n11039 , n11040 , n11041 , n330890 , n330891 , n11044 , 
 n330893 , n330894 , n11047 , n330896 , n11049 , n330898 , n11051 , n330900 , n11053 , n330902 , 
 n11055 , n11056 , n330905 , n330906 , n11059 , n330908 , n330909 , n11062 , n330911 , n330912 , 
 n11065 , n11066 , n330915 , n11068 , n330917 , n11070 , n11071 , n330920 , n330921 , n11074 , 
 n330923 , n330924 , n11077 , n330926 , n330927 , n330928 , n11081 , n330930 , n330931 , n11084 , 
 n330933 , n330934 , n330935 , n11088 , n330937 , n11090 , n11091 , n330940 , n11093 , n330942 , 
 n11095 , n330944 , n330945 , n11098 , n11099 , n330948 , n11101 , n330950 , n330951 , n330952 , 
 n11105 , n330954 , n330955 , n11108 , n330957 , n330958 , n330959 , n11112 , n330961 , n330962 , 
 n11115 , n330964 , n330965 , n330966 , n11119 , n330968 , n11121 , n11122 , n330971 , n11124 , 
 n330973 , n11126 , n11127 , n330976 , n330977 , n11130 , n330979 , n330980 , n11133 , n330982 , 
 n330983 , n330984 , n11137 , n330986 , n330987 , n11140 , n330989 , n330990 , n11143 , n11144 , 
 n330993 , n330994 , n11147 , n11148 , n11149 , n330998 , n330999 , n331000 , n11153 , n331002 , 
 n11155 , n11156 , n331005 , n11158 , n331007 , n11160 , n11161 , n331010 , n331011 , n11164 , 
 n331013 , n331014 , n11167 , n331016 , n331017 , n331018 , n11171 , n331020 , n331021 , n11174 , 
 n331023 , n331024 , n11177 , n331026 , n11179 , n331028 , n11181 , n11182 , n331031 , n331032 , 
 n11185 , n11186 , n331035 , n331036 , n331037 , n11190 , n331039 , n11192 , n11193 , n331042 , 
 n11195 , n331044 , n11197 , n11198 , n331047 , n331048 , n11201 , n331050 , n331051 , n11204 , 
 n331053 , n331054 , n331055 , n11208 , n331057 , n331058 , n11211 , n331060 , n331061 , n11214 , 
 n331063 , n331064 , n11217 , n331066 , n331067 , n11220 , n331069 , n331070 , n11223 , n11224 , 
 n11225 , n11226 , n331075 , n331076 , n11229 , n331078 , n11231 , n11232 , n11233 , n331082 , 
 n331083 , n11236 , n331085 , n331086 , n11239 , n331088 , n11241 , n11242 , n331091 , n331092 , 
 n331093 , n11246 , n11247 , n331096 , n331097 , n11250 , n11251 , n331100 , n11253 , n331102 , 
 n331103 , n331104 , n11257 , n331106 , n11259 , n331108 , n331109 , n331110 , n331111 , n11264 , 
 n331113 , n11266 , n331115 , n331116 , n11269 , n331118 , n331119 , n11272 , n11273 , n331122 , 
 n331123 , n11276 , n331125 , n11278 , n331127 , n11280 , n11281 , n11282 , n331131 , n11284 , 
 n331133 , n331134 , n11287 , n331136 , n11288 , n331138 , n331139 , n11291 , n11292 , n11293 , 
 n331143 , n331144 , n11296 , n11297 , n11298 , n331148 , n331149 , n11301 , n331151 , n331152 , 
 n11304 , n331154 , n11306 , n331156 , n11308 , n331158 , n11310 , n11311 , n331161 , n331162 , 
 n11314 , n331164 , n331165 , n11317 , n331167 , n331168 , n11320 , n11321 , n331171 , n11323 , 
 n331173 , n11325 , n11326 , n331176 , n331177 , n11329 , n331179 , n331180 , n11332 , n331182 , 
 n331183 , n331184 , n11336 , n331186 , n331187 , n11339 , n331189 , n331190 , n11342 , n11343 , 
 n11344 , n331194 , n331195 , n331196 , n11348 , n331198 , n331199 , n11351 , n11352 , n331202 , 
 n11354 , n11355 , n331205 , n331206 , n11358 , n11359 , n11360 , n11361 , n331211 , n11363 , 
 n331213 , n11365 , n11366 , n331216 , n331217 , n11369 , n331219 , n331220 , n11372 , n331222 , 
 n331223 , n11375 , n11376 , n11377 , n11378 , n11379 , n331229 , n331230 , n331231 , n11383 , 
 n331233 , n11385 , n11386 , n331236 , n331237 , n11389 , n331239 , n331240 , n11392 , n331242 , 
 n331243 , n11395 , n11396 , n11397 , n331247 , n331248 , n11400 , n331250 , n331251 , n11403 , 
 n11404 , n11405 , n331255 , n331256 , n11408 , n11409 , n11410 , n11411 , n11412 , n331262 , 
 n331263 , n11415 , n11416 , n331266 , n331267 , n11419 , n331269 , n11421 , n331271 , n11423 , 
 n11424 , n331274 , n331275 , n11427 , n331277 , n331278 , n11430 , n331280 , n331281 , n11433 , 
 n331283 , n331284 , n11436 , n331286 , n331287 , n331288 , n11440 , n331290 , n11442 , n11443 , 
 n331293 , n11445 , n331295 , n11447 , n11448 , n331298 , n331299 , n11451 , n331301 , n331302 , 
 n11454 , n331304 , n331305 , n331306 , n331307 , n331308 , n331309 , n331310 , n331311 , n331312 , 
 n11464 , n11465 , n331315 , n331316 , n11468 , n331318 , n331319 , n331320 , n331321 , n11473 , 
 n331323 , n11475 , n331325 , n331326 , n11478 , n331328 , n331329 , n11481 , n11482 , n331332 , 
 n11484 , n331334 , n331335 , n331336 , n331337 , n331338 , n331339 , n11491 , n331341 , n331342 , 
 n11494 , n11495 , n331345 , n331346 , n11498 , n331348 , n331349 , n331350 , n331351 , n331352 , 
 n11504 , n331354 , n11506 , n11507 , n331357 , n11509 , n331359 , n11511 , n331361 , n11513 , 
 n331363 , n331364 , n331365 , n331366 , n331367 , n331368 , n331369 , n331370 , n11522 , n331372 , 
 n331373 , n331374 , n331375 , n331376 , n331377 , n331378 , n11530 , n331380 , n331381 , n11533 , 
 n331383 , n331384 , n11536 , n331386 , n331387 , n331388 , n11540 , n331390 , n11542 , n331392 , 
 n331393 , n331394 , n331395 , n331396 , n331397 , n11549 , n331399 , n11551 , n11552 , n331402 , 
 n331403 , n331404 , n331405 , n331406 , n331407 , n11559 , n331409 , n331410 , n331411 , n331412 , 
 n331413 , n331414 , n331415 , n331416 , n331417 , n331418 , n331419 , n331420 , n331421 , n11573 , 
 n331423 , n331424 , n11576 , n331426 , n331427 , n331428 , n331429 , n331430 , n331431 , n331432 , 
 n331433 , n11585 , n331435 , n331436 , n331437 , n331438 , n11590 , n331440 , n331441 , n331442 , 
 n331443 , n331444 , n331445 , n11597 , n331447 , n331448 , n11600 , n331450 , n331451 , n331452 , 
 n331453 , n331454 , n11603 , n11604 , n11605 , n11606 , n331459 , n331460 , n11608 , n11609 , 
 n331463 , n331464 , n331465 , n331466 , n331467 , n331468 , n331469 , n11614 , n331471 , n331472 , 
 n11617 , n331474 , n331475 , n331476 , n331477 , n331478 , n331479 , n331480 , n331481 , n331482 , 
 n11626 , n331484 , n331485 , n331486 , n331487 , n331488 , n331489 , n331490 , n331491 , n11635 , 
 n331493 , n11637 , n331495 , n331496 , n11640 , n331498 , n331499 , n331500 , n331501 , n331502 , 
 n331503 , n11647 , n331505 , n331506 , n11650 , n331508 , n331509 , n331510 , n331511 , n331512 , 
 n11656 , n331514 , n11658 , n331516 , n331517 , n11661 , n331519 , n331520 , n331521 , n331522 , 
 n331523 , n331524 , n331525 , n331526 , n331527 , n331528 , n331529 , n331530 , n331531 , n331532 , 
 n331533 , n11677 , n11678 , n331536 , n331537 , n331538 , n331539 , n331540 , n331541 , n11685 , 
 n331543 , n331544 , n11688 , n331546 , n331547 , n11691 , n11692 , n331550 , n331551 , n331552 , 
 n331553 , n331554 , n331555 , n331556 , n331557 , n11701 , n11702 , n331560 , n11704 , n331562 , 
 n331563 , n11707 , n331565 , n331566 , n331567 , n331568 , n11712 , n11713 , n11714 , n11715 , 
 n331573 , n11717 , n331575 , n331576 , n11720 , n331578 , n11722 , n11723 , n11724 , n331582 , 
 n331583 , n331584 , n11728 , n331586 , n11730 , n11731 , n331589 , n11733 , n331591 , n11735 , 
 n11736 , n331594 , n331595 , n11739 , n331597 , n331598 , n11742 , n331600 , n331601 , n331602 , 
 n11746 , n331604 , n331605 , n11749 , n331607 , n331608 , n331609 , n11753 , n331611 , n11755 , 
 n11756 , n331614 , n11758 , n11759 , n331617 , n11761 , n11762 , n331620 , n11764 , n331622 , 
 n11766 , n331624 , n331625 , n11769 , n331627 , n331628 , n331629 , n11773 , n331631 , n331632 , 
 n11776 , n331634 , n331635 , n11779 , n11780 , n11781 , n331639 , n331640 , n11784 , n11785 , 
 n11786 , n331644 , n331645 , n11789 , n11790 , n331648 , n331649 , n11793 , n331651 , n11795 , 
 n331653 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n331662 , 
 n331663 , n11807 , n331665 , n331666 , n11810 , n331668 , n331669 , n11813 , n11814 , n11815 , 
 n331673 , n331674 , n11818 , n331676 , n11820 , n11821 , n331679 , n11823 , n331681 , n11825 , 
 n331683 , n11827 , n11828 , n331686 , n331687 , n11831 , n331689 , n331690 , n11834 , n331692 , 
 n331693 , n11837 , n11838 , n331696 , n11840 , n331698 , n11842 , n11843 , n331701 , n331702 , 
 n11846 , n331704 , n331705 , n11849 , n331707 , n331708 , n331709 , n331710 , n331711 , n331712 , 
 n331713 , n331714 , n331715 , n331716 , n331717 , n331718 , n331719 , n331720 , n11864 , n11865 , 
 n331723 , n331724 , n331725 , n331726 , n331727 , n11871 , n11872 , n331730 , n331731 , n331732 , 
 n11876 , n11877 , n11878 , n11879 , n331737 , n11881 , n331739 , n331740 , n331741 , n11885 , 
 n331743 , n331744 , n331745 , n331746 , n331747 , n11891 , n331749 , n331750 , n331751 , n11895 , 
 n331753 , n11897 , n331755 , n331756 , n331757 , n331758 , n331759 , n11903 , n331761 , n331762 , 
 n331763 , n331764 , n331765 , n331766 , n11910 , n11911 , n11912 , n331770 , n331771 , n331772 , 
 n331773 , n331774 , n11918 , n331776 , n331777 , n11921 , n11922 , n331780 , n331781 , n331782 , 
 n331783 , n331784 , n331785 , n331786 , n331787 , n331788 , n331789 , n331790 , n331791 , n331792 , 
 n331793 , n331794 , n331795 , n331796 , n331797 , n331798 , n331799 , n331800 , n11944 , n331802 , 
 n331803 , n331804 , n331805 , n331806 , n331807 , n331808 , n331809 , n331810 , n331811 , n11955 , 
 n11956 , n11957 , n331815 , n331816 , n11960 , n331818 , n331819 , n11963 , n331821 , n11965 , 
 n331823 , n331824 , n331825 , n331826 , n11969 , n331828 , n11971 , n331830 , n331831 , n331832 , 
 n11975 , n11976 , n331835 , n11978 , n331837 , n331838 , n11981 , n331840 , n11983 , n331842 , 
 n331843 , n11986 , n331845 , n331846 , n331847 , n331848 , n331849 , n11992 , n331851 , n331852 , 
 n331853 , n331854 , n331855 , n331856 , n11999 , n12000 , n331859 , n12002 , n331861 , n12004 , 
 n331863 , n331864 , n12007 , n331866 , n331867 , n331868 , n331869 , n331870 , n331871 , n331872 , 
 n331873 , n331874 , n331875 , n331876 , n331877 , n331878 , n331879 , n331880 , n331881 , n331882 , 
 n331883 , n331884 , n331885 , n12028 , n12029 , n331888 , n331889 , n331890 , n331891 , n331892 , 
 n12035 , n331894 , n331895 , n331896 , n331897 , n331898 , n331899 , n12042 , n331901 , n331902 , 
 n12045 , n331904 , n331905 , n331906 , n331907 , n331908 , n331909 , n331910 , n331911 , n331912 , 
 n331913 , n12056 , n331915 , n331916 , n331917 , n331918 , n12061 , n331920 , n331921 , n331922 , 
 n331923 , n12066 , n331925 , n12068 , n331927 , n12070 , n331929 , n331930 , n331931 , n331932 , 
 n331933 , n331934 , n12077 , n331936 , n12079 , n331938 , n331939 , n331940 , n331941 , n331942 , 
 n331943 , n331944 , n331945 , n331946 , n12089 , n331948 , n331949 , n12092 , n12093 , n331952 , 
 n12095 , n331954 , n331955 , n331956 , n331957 , n331958 , n12101 , n12102 , n12103 , n12104 , 
 n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n331969 , n331970 , n331971 , n331972 , 
 n331973 , n331974 , n331975 , n331976 , n331977 , n331978 , n331979 , n331980 , n12123 , n331982 , 
 n331983 , n331984 , n331985 , n331986 , n331987 , n331988 , n12131 , n331990 , n331991 , n331992 , 
 n331993 , n331994 , n331995 , n12138 , n331997 , n331998 , n331999 , n332000 , n332001 , n332002 , 
 n332003 , n332004 , n332005 , n12148 , n12149 , n12150 , n12151 , n12152 , n332011 , n332012 , 
 n332013 , n12156 , n332015 , n332016 , n332017 , n332018 , n332019 , n332020 , n332021 , n332022 , 
 n332023 , n12166 , n12167 , n332026 , n332027 , n332028 , n332029 , n12172 , n332031 , n332032 , 
 n12175 , n332034 , n332035 , n12178 , n332037 , n332038 , n332039 , n12182 , n332041 , n332042 , 
 n332043 , n332044 , n332045 , n332046 , n332047 , n332048 , n332049 , n12192 , n332051 , n332052 , 
 n332053 , n332054 , n12197 , n332056 , n12199 , n332058 , n332059 , n12202 , n332061 , n332062 , 
 n332063 , n332064 , n332065 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n332072 , 
 n332073 , n332074 , n332075 , n332076 , n332077 , n332078 , n332079 , n12222 , n12223 , n332082 , 
 n332083 , n332084 , n12227 , n332086 , n332087 , n332088 , n332089 , n332090 , n332091 , n332092 , 
 n332093 , n12236 , n12237 , n12238 , n12239 , n12240 , n332099 , n332100 , n12243 , n332102 , 
 n332103 , n12246 , n332105 , n332106 , n12249 , n332108 , n332109 , n332110 , n12253 , n332112 , 
 n332113 , n332114 , n12257 , n12258 , n332117 , n332118 , n332119 , n332120 , n332121 , n332122 , 
 n12265 , n12266 , n12267 , n12268 , n12269 , n332128 , n332129 , n332130 , n332131 , n332132 , 
 n332133 , n332134 , n332135 , n332136 , n332137 , n332138 , n332139 , n332140 , n332141 , n332142 , 
 n12285 , n332144 , n12287 , n332146 , n12289 , n12290 , n332149 , n12292 , n332151 , n12294 , 
 n332153 , n332154 , n12297 , n332156 , n332157 , n12300 , n12301 , n332160 , n332161 , n12304 , 
 n12305 , n332164 , n12307 , n12308 , n332167 , n332168 , n332169 , n12312 , n332171 , n332172 , 
 n12315 , n332174 , n332175 , n12318 , n332177 , n332178 , n12321 , n332180 , n12323 , n332182 , 
 n332183 , n332184 , n332185 , n12328 , n12329 , n332188 , n12331 , n332190 , n332191 , n12334 , 
 n332193 , n332194 , n12337 , n332196 , n332197 , n12340 , n332199 , n12342 , n332201 , n12344 , 
 n12345 , n332204 , n332205 , n12348 , n332207 , n332208 , n12351 , n332210 , n332211 , n12354 , 
 n332213 , n12355 , n332215 , n332216 , n12358 , n12359 , n12360 , n332220 , n332221 , n12363 , 
 n12364 , n12365 , n332225 , n332226 , n12368 , n12369 , n12370 , n332230 , n12372 , n12373 , 
 n332233 , n12375 , n12376 , n12377 , n332237 , n12379 , n332239 , n12381 , n332241 , n332242 , 
 n12384 , n12385 , n332245 , n12387 , n12388 , n332248 , n332249 , n12391 , n12392 , n12393 , 
 n12394 , n12395 , n332255 , n332256 , n12398 , n332258 , n12400 , n332260 , n332261 , n12403 , 
 n332263 , n332264 , n12406 , n332266 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , 
 n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n332282 , 
 n12424 , n332284 , n332285 , n332286 , n12428 , n332288 , n12430 , n332290 , n332291 , n332292 , 
 n332293 , n332294 , n12436 , n12437 , n332297 , n332298 , n332299 , n332300 , n12442 , n332302 , 
 n332303 , n12445 , n332305 , n332306 , n332307 , n12449 , n332309 , n12451 , n12452 , n332312 , 
 n332313 , n12455 , n332315 , n332316 , n12458 , n332318 , n332319 , n332320 , n12462 , n332322 , 
 n12464 , n332324 , n12466 , n332326 , n332327 , n12469 , n332329 , n332330 , n332331 , n332332 , 
 n12474 , n332334 , n332335 , n12477 , n332337 , n332338 , n12480 , n332340 , n332341 , n332342 , 
 n12484 , n332344 , n332345 , n12487 , n332347 , n332348 , n12490 , n12491 , n332351 , n332352 , 
 n332353 , n332354 , n332355 , n332356 , n332357 , n332358 , n12500 , n332360 , n332361 , n12503 , 
 n332363 , n332364 , n332365 , n332366 , n332367 , n332368 , n12509 , n332370 , n332371 , n12512 , 
 n332373 , n332374 , n12515 , n332376 , n12517 , n332378 , n12519 , n332380 , n332381 , n332382 , 
 n332383 , n332384 , n332385 , n12526 , n332387 , n332388 , n12529 , n332390 , n332391 , n332392 , 
 n332393 , n332394 , n332395 , n12536 , n332397 , n12538 , n332399 , n332400 , n12541 , n332402 , 
 n12543 , n12544 , n332405 , n332406 , n332407 , n12548 , n332409 , n332410 , n12551 , n12552 , 
 n12553 , n332414 , n332415 , n332416 , n12557 , n332418 , n332419 , n332420 , n332421 , n332422 , 
 n12563 , n12564 , n332425 , n12566 , n332427 , n332428 , n332429 , n332430 , n332431 , n332432 , 
 n332433 , n332434 , n332435 , n332436 , n332437 , n332438 , n332439 , n332440 , n332441 , n332442 , 
 n332443 , n12584 , n332445 , n332446 , n12587 , n12588 , n332449 , n12590 , n12591 , n332452 , 
 n332453 , n332454 , n12595 , n332456 , n332457 , n12598 , n332459 , n332460 , n12601 , n332462 , 
 n332463 , n332464 , n12605 , n12606 , n12607 , n12608 , n332469 , n332470 , n12611 , n332472 , 
 n332473 , n332474 , n12615 , n332476 , n332477 , n12618 , n332479 , n332480 , n12621 , n332482 , 
 n12623 , n332484 , n332485 , n332486 , n332487 , n332488 , n12629 , n332490 , n12631 , n332492 , 
 n12633 , n332494 , n12635 , n12636 , n332497 , n12638 , n332499 , n332500 , n12641 , n332502 , 
 n332503 , n332504 , n12645 , n332506 , n332507 , n332508 , n12649 , n332510 , n332511 , n12652 , 
 n332513 , n332514 , n332515 , n332516 , n332517 , n332518 , n12659 , n332520 , n332521 , n12662 , 
 n332523 , n332524 , n332525 , n332526 , n332527 , n332528 , n332529 , n332530 , n332531 , n12672 , 
 n332533 , n332534 , n12675 , n332536 , n332537 , n332538 , n332539 , n332540 , n332541 , n332542 , 
 n332543 , n332544 , n332545 , n12686 , n332547 , n332548 , n332549 , n332550 , n332551 , n332552 , 
 n332553 , n332554 , n332555 , n332556 , n332557 , n332558 , n332559 , n332560 , n332561 , n332562 , 
 n332563 , n332564 , n332565 , n332566 , n332567 , n12708 , n332569 , n332570 , n12711 , n332572 , 
 n332573 , n12714 , n332575 , n332576 , n12717 , n332578 , n332579 , n332580 , n332581 , n332582 , 
 n332583 , n12724 , n332585 , n332586 , n12727 , n332588 , n332589 , n332590 , n332591 , n332592 , 
 n332593 , n12734 , n332595 , n332596 , n12737 , n12738 , n332599 , n332600 , n12741 , n332602 , 
 n12743 , n12744 , n12745 , n332606 , n12747 , n332608 , n12749 , n12750 , n332611 , n332612 , 
 n332613 , n332614 , n12755 , n12756 , n12757 , n12758 , n332619 , n332620 , n12761 , n332622 , 
 n332623 , n12764 , n332625 , n332626 , n12767 , n332628 , n332629 , n332630 , n332631 , n332632 , 
 n12773 , n332634 , n332635 , n12776 , n332637 , n332638 , n12779 , n332640 , n332641 , n12782 , 
 n332643 , n332644 , n332645 , n332646 , n12787 , n332648 , n332649 , n332650 , n332651 , n12792 , 
 n332653 , n332654 , n332655 , n332656 , n332657 , n332658 , n12799 , n332660 , n12801 , n12802 , 
 n332663 , n332664 , n12805 , n332666 , n332667 , n332668 , n332669 , n332670 , n12811 , n332672 , 
 n332673 , n332674 , n332675 , n332676 , n332677 , n332678 , n12819 , n332680 , n12821 , n12822 , 
 n332683 , n332684 , n12825 , n332686 , n332687 , n12828 , n12829 , n12830 , n12831 , n12832 , 
 n332693 , n332694 , n12835 , n332696 , n332697 , n332698 , n332699 , n12840 , n332701 , n12842 , 
 n332703 , n332704 , n12845 , n332706 , n12847 , n12848 , n12849 , n332710 , n12851 , n12852 , 
 n332713 , n12854 , n332715 , n332716 , n332717 , n12858 , n12859 , n332720 , n12861 , n332722 , 
 n332723 , n332724 , n332725 , n12866 , n332727 , n332728 , n332729 , n332730 , n332731 , n332732 , 
 n332733 , n12874 , n332735 , n332736 , n12877 , n332738 , n332739 , n332740 , n332741 , n332742 , 
 n12883 , n12884 , n332745 , n12886 , n332747 , n332748 , n332749 , n332750 , n332751 , n332752 , 
 n332753 , n12894 , n332755 , n332756 , n12897 , n332758 , n12899 , n12900 , n332761 , n332762 , 
 n12903 , n332764 , n332765 , n12906 , n332767 , n12908 , n332769 , n332770 , n332771 , n12912 , 
 n332773 , n332774 , n12915 , n332776 , n12917 , n332778 , n332779 , n12920 , n332781 , n332782 , 
 n12923 , n12924 , n12925 , n12926 , n12927 , n332788 , n332789 , n332790 , n332791 , n332792 , 
 n332793 , n332794 , n332795 , n332796 , n12937 , n332798 , n12939 , n332800 , n332801 , n332802 , 
 n12943 , n332804 , n332805 , n12946 , n332807 , n332808 , n12949 , n332810 , n332811 , n12952 , 
 n12953 , n12954 , n12955 , n332816 , n332817 , n332818 , n332819 , n332820 , n332821 , n332822 , 
 n12963 , n12964 , n332825 , n12966 , n332827 , n12968 , n332829 , n332830 , n332831 , n12972 , 
 n332833 , n332834 , n12975 , n332836 , n332837 , n12978 , n12979 , n332840 , n332841 , n12982 , 
 n332843 , n332844 , n12985 , n332846 , n332847 , n12988 , n332849 , n332850 , n12991 , n332852 , 
 n332853 , n12994 , n332855 , n332856 , n12997 , n332858 , n332859 , n13000 , n13001 , n13002 , 
 n13003 , n332864 , n332865 , n13006 , n13007 , n13008 , n13009 , n13010 , n332871 , n332872 , 
 n332873 , n13014 , n13015 , n13016 , n13017 , n13018 , n332879 , n13020 , n13021 , n332882 , 
 n332883 , n13024 , n332885 , n332886 , n13027 , n332888 , n332889 , n13030 , n332891 , n13032 , 
 n332893 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , 
 n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n332911 , n332912 , 
 n332913 , n332914 , n13055 , n332916 , n332917 , n332918 , n13059 , n332920 , n13061 , n13062 , 
 n332923 , n332924 , n332925 , n13066 , n332927 , n332928 , n13069 , n332930 , n332931 , n13072 , 
 n332933 , n332934 , n13075 , n332936 , n13077 , n332938 , n13079 , n13080 , n332941 , n13082 , 
 n332943 , n13084 , n332945 , n332946 , n13087 , n332948 , n332949 , n13090 , n332951 , n332952 , 
 n13093 , n13094 , n13095 , n13096 , n332957 , n332958 , n332959 , n13100 , n332961 , n332962 , 
 n13103 , n332964 , n13105 , n13106 , n332967 , n13108 , n332969 , n13110 , n13111 , n332972 , 
 n332973 , n332974 , n13115 , n332976 , n332977 , n13118 , n332979 , n332980 , n13121 , n332982 , 
 n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n332992 , 
 n13133 , n332994 , n332995 , n13136 , n13137 , n13138 , n13139 , n333000 , n333001 , n13142 , 
 n13143 , n13144 , n13145 , n13146 , n333007 , n333008 , n13149 , n13150 , n13151 , n13152 , 
 n333013 , n13154 , n13155 , n333016 , n333017 , n13158 , n333019 , n333020 , n13161 , n333022 , 
 n333023 , n333024 , n333025 , n13166 , n333027 , n333028 , n333029 , n333030 , n333031 , n333032 , 
 n333033 , n333034 , n333035 , n333036 , n333037 , n333038 , n13179 , n13180 , n333041 , n13182 , 
 n333043 , n13184 , n333045 , n13186 , n13187 , n333048 , n333049 , n333050 , n13191 , n333052 , 
 n333053 , n13194 , n333055 , n333056 , n13197 , n333058 , n333059 , n13200 , n333061 , n333062 , 
 n13203 , n333064 , n333065 , n13206 , n13207 , n13208 , n333069 , n333070 , n333071 , n333072 , 
 n333073 , n333074 , n333075 , n333076 , n333077 , n333078 , n333079 , n13220 , n333081 , n333082 , 
 n333083 , n333084 , n13225 , n13226 , n13227 , n13228 , n13229 , n333090 , n333091 , n13232 , 
 n13233 , n13234 , n13235 , n333096 , n333097 , n13238 , n13239 , n13240 , n13241 , n333102 , 
 n333103 , n333104 , n333105 , n333106 , n13247 , n333108 , n333109 , n13250 , n13251 , n13252 , 
 n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n333121 , n13262 , 
 n333123 , n13264 , n333125 , n13266 , n13267 , n333128 , n13269 , n333130 , n13271 , n333132 , 
 n333133 , n13274 , n333135 , n333136 , n13277 , n333138 , n333139 , n13280 , n333141 , n13282 , 
 n333143 , n13284 , n13285 , n333146 , n333147 , n333148 , n13289 , n333150 , n333151 , n13292 , 
 n333153 , n333154 , n333155 , n333156 , n333157 , n333158 , n13299 , n333160 , n13301 , n13302 , 
 n333163 , n13304 , n333165 , n333166 , n333167 , n333168 , n13309 , n13310 , n333171 , n13312 , 
 n333173 , n333174 , n333175 , n13316 , n333177 , n333178 , n13319 , n333180 , n333181 , n13322 , 
 n13323 , n13324 , n13325 , n333186 , n333187 , n13328 , n13329 , n13330 , n13331 , n13332 , 
 n333193 , n333194 , n333195 , n333196 , n13337 , n333198 , n13339 , n333200 , n333201 , n333202 , 
 n333203 , n13344 , n333205 , n333206 , n13347 , n333208 , n333209 , n13350 , n333211 , n13352 , 
 n13353 , n333214 , n333215 , n13356 , n333217 , n333218 , n333219 , n13360 , n13361 , n333222 , 
 n333223 , n333224 , n13365 , n333226 , n333227 , n13368 , n333229 , n333230 , n13371 , n333232 , 
 n333233 , n13374 , n333235 , n13376 , n13377 , n333238 , n333239 , n333240 , n13381 , n333242 , 
 n333243 , n13384 , n333245 , n333246 , n13387 , n333248 , n13389 , n13390 , n333251 , n13392 , 
 n333253 , n13394 , n333255 , n333256 , n333257 , n333258 , n333259 , n333260 , n13401 , n333262 , 
 n333263 , n13404 , n13405 , n13406 , n13407 , n13408 , n333269 , n333270 , n13411 , n333272 , 
 n333273 , n13414 , n333275 , n333276 , n13417 , n333278 , n333279 , n13420 , n333281 , n13422 , 
 n13423 , n13424 , n13425 , n333286 , n13427 , n13428 , n333289 , n333290 , n13431 , n333292 , 
 n13433 , n13434 , n13435 , n333296 , n333297 , n333298 , n333299 , n13440 , n333301 , n333302 , 
 n333303 , n333304 , n13445 , n333306 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , 
 n333313 , n333314 , n13455 , n333316 , n13457 , n333318 , n13459 , n333320 , n13461 , n333322 , 
 n333323 , n13464 , n333325 , n333326 , n13467 , n333328 , n13469 , n13470 , n13471 , n13472 , 
 n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , 
 n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , 
 n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n333360 , n333361 , n13502 , 
 n333363 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , 
 n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , 
 n333383 , n333384 , n13525 , n333386 , n13527 , n333388 , n333389 , n333390 , n13531 , n333392 , 
 n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , 
 n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , 
 n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n333421 , n13562 , 
 n333423 , n13564 , n13565 , n13566 , n13567 , n13568 , n333429 , n13570 , n333431 , n13572 , 
 n333433 , n333434 , n13575 , n333436 , n333437 , n333438 , n13579 , n333440 , n13581 , n13582 , 
 n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n333450 , n13591 , n333452 , 
 n333453 , n333454 , n13595 , n333456 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , 
 n333463 , n13604 , n333465 , n333466 , n13607 , n13608 , n333469 , n13610 , n333471 , n333472 , 
 n333473 , n13614 , n333475 , n333476 , n13617 , n333478 , n333479 , n13620 , n13621 , n333482 , 
 n333483 , n13624 , n333485 , n333486 , n13627 , n333488 , n333489 , n13630 , n333491 , n333492 , 
 n13633 , n333494 , n13635 , n13636 , n13637 , n13638 , n333499 , n13640 , n333501 , n333502 , 
 n333503 , n333504 , n333505 , n333506 , n13647 , n13648 , n333509 , n13650 , n333511 , n13652 , 
 n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , 
 n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , 
 n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , 
 n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n333549 , n13690 , n333551 , n333552 , 
 n13693 , n333554 , n13695 , n333556 , n13697 , n333558 , n333559 , n333560 , n13701 , n333562 , 
 n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , 
 n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , 
 n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n333591 , n333592 , 
 n13733 , n333594 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n333601 , n333602 , 
 n333603 , n13744 , n333605 , n333606 , n13747 , n333608 , n333609 , n333610 , n333611 , n13752 , 
 n333613 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , 
 n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , 
 n13773 , n13774 , n13775 , n13776 , n13777 , n333638 , n333639 , n13780 , n333641 , n13782 , 
 n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , 
 n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , 
 n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , 
 n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , 
 n13823 , n333684 , n13825 , n333686 , n13827 , n333688 , n13829 , n13830 , n13831 , n13832 , 
 n13833 , n333694 , n333695 , n13836 , n13837 , n13838 , n13839 , n333700 , n333701 , n13842 , 
 n13843 , n13844 , n13845 , n13846 , n333707 , n333708 , n333709 , n13850 , n333711 , n13852 , 
 n13853 , n333714 , n333715 , n13856 , n333717 , n333718 , n13859 , n333720 , n333721 , n13862 , 
 n333723 , n333724 , n13865 , n13866 , n13867 , n13868 , n333729 , n333730 , n13871 , n13872 , 
 n13873 , n13874 , n13875 , n333736 , n333737 , n13878 , n333739 , n333740 , n333741 , n333742 , 
 n13883 , n333744 , n333745 , n13886 , n333747 , n333748 , n333749 , n333750 , n333751 , n333752 , 
 n13893 , n333754 , n333755 , n13896 , n333757 , n333758 , n333759 , n333760 , n13901 , n333762 , 
 n333763 , n333764 , n13905 , n333766 , n13907 , n13908 , n333769 , n333770 , n333771 , n333772 , 
 n333773 , n333774 , n13915 , n333776 , n333777 , n13918 , n13919 , n333780 , n13921 , n333782 , 
 n333783 , n333784 , n13925 , n13926 , n333787 , n13928 , n13929 , n333790 , n333791 , n333792 , 
 n13933 , n333794 , n333795 , n13936 , n333797 , n333798 , n13939 , n333800 , n333801 , n13942 , 
 n333803 , n333804 , n13945 , n333806 , n13947 , n333808 , n13949 , n13950 , n333811 , n333812 , 
 n333813 , n13954 , n333815 , n333816 , n13957 , n333818 , n333819 , n13960 , n333821 , n333822 , 
 n333823 , n13964 , n333825 , n13966 , n13967 , n333828 , n333829 , n333830 , n13971 , n333832 , 
 n333833 , n13974 , n333835 , n333836 , n13977 , n333838 , n333839 , n333840 , n333841 , n333842 , 
 n333843 , n13984 , n13985 , n333846 , n333847 , n333848 , n13989 , n333850 , n333851 , n13992 , 
 n333853 , n333854 , n13995 , n333856 , n333857 , n13998 , n333859 , n333860 , n14001 , n333862 , 
 n333863 , n14004 , n333865 , n333866 , n14007 , n333868 , n333869 , n14010 , n14011 , n14012 , 
 n14013 , n333874 , n333875 , n14016 , n14017 , n14018 , n14019 , n14020 , n333881 , n333882 , 
 n14023 , n14024 , n14025 , n14026 , n333887 , n333888 , n14029 , n14030 , n14031 , n14032 , 
 n14033 , n333894 , n333895 , n333896 , n14037 , n333898 , n14039 , n14040 , n333901 , n333902 , 
 n14043 , n333904 , n333905 , n14046 , n333907 , n333908 , n14049 , n333910 , n333911 , n14052 , 
 n14053 , n14054 , n14055 , n333916 , n333917 , n14058 , n333919 , n333920 , n14061 , n333922 , 
 n14063 , n333924 , n333925 , n333926 , n333927 , n14068 , n333929 , n333930 , n14071 , n333932 , 
 n333933 , n14074 , n333935 , n333936 , n14077 , n14078 , n14079 , n14080 , n333941 , n333942 , 
 n14083 , n333944 , n14085 , n333946 , n14087 , n14088 , n333949 , n333950 , n14091 , n333952 , 
 n14093 , n333954 , n333955 , n14096 , n333957 , n333958 , n14099 , n14100 , n14101 , n14102 , 
 n333963 , n333964 , n333965 , n14106 , n333967 , n333968 , n14109 , n333970 , n14111 , n14112 , 
 n14113 , n14114 , n14115 , n333976 , n333977 , n333978 , n14119 , n333980 , n333981 , n14122 , 
 n333983 , n14124 , n14125 , n333986 , n14127 , n14128 , n14129 , n14130 , n333991 , n333992 , 
 n333993 , n14134 , n333995 , n333996 , n14137 , n333998 , n14139 , n334000 , n14141 , n334002 , 
 n14143 , n14144 , n334005 , n14146 , n334007 , n14148 , n334009 , n334010 , n14151 , n334012 , 
 n14153 , n334014 , n334015 , n14156 , n334017 , n14158 , n14159 , n14160 , n14161 , n14162 , 
 n14163 , n334024 , n14165 , n334026 , n334027 , n14168 , n334029 , n334030 , n14171 , n14172 , 
 n14173 , n14174 , n14175 , n334036 , n334037 , n14178 , n334039 , n334040 , n14181 , n334042 , 
 n334043 , n14184 , n334045 , n334046 , n14187 , n334048 , n334049 , n14190 , n14191 , n14192 , 
 n14193 , n334054 , n334055 , n14196 , n334057 , n334058 , n14199 , n334060 , n334061 , n14202 , 
 n334063 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n334070 , n14211 , n334072 , 
 n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , 
 n334083 , n14224 , n334085 , n14226 , n14227 , n334088 , n14229 , n334090 , n14231 , n334092 , 
 n14233 , n334094 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , 
 n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , 
 n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , 
 n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , 
 n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , 
 n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , 
 n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , 
 n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , 
 n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , 
 n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , 
 n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , 
 n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , 
 n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , 
 n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n334232 , 
 n14373 , n334234 , n14375 , n334236 , n14377 , n334238 , n334239 , n14380 , n14381 , n14382 , 
 n14383 , n14384 , n14385 , n334246 , n14387 , n334248 , n334249 , n14390 , n334251 , n14392 , 
 n14393 , n14394 , n14395 , n334256 , n334257 , n334258 , n14399 , n334260 , n14401 , n14402 , 
 n334263 , n334264 , n334265 , n14406 , n334267 , n334268 , n14409 , n334270 , n334271 , n14412 , 
 n334273 , n334274 , n334275 , n14416 , n334277 , n14418 , n334279 , n334280 , n14421 , n14422 , 
 n334283 , n334284 , n334285 , n14426 , n334287 , n334288 , n14429 , n334290 , n334291 , n14432 , 
 n334293 , n334294 , n14435 , n334296 , n334297 , n14438 , n334299 , n14440 , n334301 , n334302 , 
 n14443 , n334304 , n334305 , n14446 , n334307 , n14448 , n334309 , n14450 , n14451 , n334312 , 
 n334313 , n334314 , n14455 , n334316 , n334317 , n14458 , n334319 , n334320 , n14461 , n334322 , 
 n334323 , n334324 , n14465 , n334326 , n14467 , n14468 , n334329 , n334330 , n334331 , n14472 , 
 n334333 , n334334 , n14475 , n334336 , n334337 , n14478 , n334339 , n334340 , n14481 , n334342 , 
 n14483 , n334344 , n14485 , n14486 , n334347 , n334348 , n334349 , n14490 , n334351 , n334352 , 
 n14493 , n334354 , n334355 , n14496 , n334357 , n334358 , n14499 , n334360 , n334361 , n14502 , 
 n334363 , n334364 , n14505 , n14506 , n14507 , n14508 , n334369 , n334370 , n14511 , n334372 , 
 n334373 , n14514 , n334375 , n334376 , n334377 , n14518 , n14519 , n14520 , n14521 , n14522 , 
 n334383 , n334384 , n14525 , n334386 , n334387 , n14528 , n14529 , n14530 , n14531 , n334392 , 
 n334393 , n14534 , n14535 , n14536 , n14537 , n14538 , n334399 , n334400 , n14541 , n334402 , 
 n334403 , n14544 , n334405 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , 
 n14553 , n334414 , n334415 , n334416 , n14557 , n334418 , n14559 , n334420 , n334421 , n334422 , 
 n14563 , n334424 , n14565 , n14566 , n14567 , n14568 , n334429 , n14570 , n334431 , n334432 , 
 n14573 , n334434 , n14575 , n334436 , n14577 , n14578 , n334439 , n334440 , n334441 , n14582 , 
 n334443 , n334444 , n14585 , n334446 , n334447 , n14588 , n334449 , n334450 , n14591 , n334452 , 
 n334453 , n14594 , n334455 , n14596 , n334457 , n14598 , n14599 , n334460 , n334461 , n334462 , 
 n14603 , n334464 , n334465 , n14606 , n334467 , n334468 , n14609 , n334470 , n334471 , n334472 , 
 n14613 , n334474 , n14615 , n334476 , n334477 , n14618 , n14619 , n334480 , n334481 , n334482 , 
 n14623 , n334484 , n334485 , n14626 , n334487 , n334488 , n14629 , n334490 , n334491 , n14632 , 
 n334493 , n14634 , n334495 , n14636 , n334497 , n334498 , n14639 , n14640 , n334501 , n334502 , 
 n334503 , n14644 , n334505 , n334506 , n14647 , n334508 , n334509 , n14650 , n334511 , n334512 , 
 n14653 , n334514 , n334515 , n14656 , n334517 , n334518 , n334519 , n334520 , n14661 , n334522 , 
 n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n334531 , n14672 , 
 n14673 , n14674 , n14675 , n334536 , n334537 , n14678 , n14679 , n14680 , n14681 , n14682 , 
 n334543 , n334544 , n14685 , n334546 , n334547 , n14688 , n14689 , n14690 , n14691 , n14692 , 
 n334553 , n334554 , n14695 , n334556 , n14697 , n14698 , n14699 , n14700 , n334561 , n334562 , 
 n14703 , n334564 , n14705 , n14706 , n334567 , n14708 , n14709 , n14710 , n14711 , n14712 , 
 n14713 , n334574 , n14715 , n334576 , n14717 , n334578 , n334579 , n14720 , n14721 , n14722 , 
 n14723 , n334584 , n334585 , n14726 , n334587 , n334588 , n14729 , n334590 , n334591 , n14732 , 
 n334593 , n14734 , n14735 , n334596 , n14737 , n334598 , n14739 , n14740 , n14741 , n14742 , 
 n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n334610 , n14751 , n334612 , 
 n14753 , n334614 , n334615 , n14756 , n334617 , n334618 , n14759 , n334620 , n14761 , n14762 , 
 n334623 , n14764 , n334625 , n14766 , n14767 , n14768 , n334629 , n334630 , n14771 , n334632 , 
 n334633 , n14774 , n334635 , n14776 , n334637 , n334638 , n14779 , n14780 , n14781 , n14782 , 
 n334643 , n334644 , n14785 , n334646 , n334647 , n334648 , n14789 , n334650 , n14791 , n14792 , 
 n334653 , n334654 , n334655 , n14796 , n334657 , n334658 , n14799 , n334660 , n334661 , n334662 , 
 n334663 , n334664 , n14805 , n334666 , n334667 , n14808 , n334669 , n334670 , n334671 , n334672 , 
 n334673 , n334674 , n334675 , n14816 , n14817 , n334678 , n14819 , n334680 , n334681 , n14822 , 
 n334683 , n14824 , n334685 , n334686 , n334687 , n334688 , n334689 , n334690 , n334691 , n14832 , 
 n334693 , n334694 , n334695 , n334696 , n14837 , n14838 , n14839 , n334700 , n334701 , n334702 , 
 n334703 , n14844 , n14845 , n14846 , n14847 , n334708 , n334709 , n334710 , n334711 , n334712 , 
 n334713 , n334714 , n334715 , n334716 , n334717 , n14858 , n334719 , n14860 , n14861 , n334722 , 
 n334723 , n334724 , n334725 , n14866 , n334727 , n334728 , n334729 , n334730 , n334731 , n14872 , 
 n334733 , n334734 , n334735 , n334736 , n14877 , n334738 , n334739 , n334740 , n334741 , n334742 , 
 n334743 , n334744 , n14885 , n334746 , n14887 , n334748 , n14889 , n14890 , n14891 , n334752 , 
 n334753 , n334754 , n334755 , n14896 , n14897 , n14898 , n334759 , n14900 , n334761 , n334762 , 
 n334763 , n14904 , n334765 , n334766 , n14907 , n334768 , n334769 , n14910 , n14911 , n334772 , 
 n14913 , n334774 , n14915 , n334776 , n334777 , n334778 , n334779 , n334780 , n14921 , n334782 , 
 n14923 , n14924 , n334785 , n334786 , n334787 , n14928 , n334789 , n334790 , n334791 , n334792 , 
 n334793 , n14934 , n334795 , n334796 , n14937 , n14938 , n14939 , n334800 , n14941 , n334802 , 
 n334803 , n334804 , n334805 , n334806 , n334807 , n14948 , n14949 , n334810 , n14951 , n334812 , 
 n334813 , n14954 , n334815 , n14956 , n14957 , n14958 , n334819 , n14960 , n334821 , n334822 , 
 n14963 , n334824 , n334825 , n334826 , n334827 , n334828 , n334829 , n14970 , n14971 , n334832 , 
 n14973 , n334834 , n334835 , n14976 , n334837 , n334838 , n14979 , n14980 , n334841 , n334842 , 
 n334843 , n334844 , n334845 , n334846 , n334847 , n334848 , n14989 , n334850 , n334851 , n334852 , 
 n334853 , n334854 , n14995 , n334856 , n334857 , n334858 , n334859 , n334860 , n334861 , n334862 , 
 n334863 , n334864 , n334865 , n15006 , n334867 , n334868 , n15009 , n334870 , n15011 , n15012 , 
 n334873 , n334874 , n334875 , n15016 , n334877 , n334878 , n334879 , n334880 , n334881 , n334882 , 
 n334883 , n334884 , n334885 , n334886 , n334887 , n15028 , n334889 , n334890 , n334891 , n334892 , 
 n334893 , n334894 , n334895 , n334896 , n334897 , n334898 , n15039 , n334900 , n334901 , n334902 , 
 n334903 , n334904 , n334905 , n334906 , n334907 , n334908 , n334909 , n15050 , n334911 , n334912 , 
 n334913 , n334914 , n334915 , n334916 , n334917 , n15058 , n15059 , n334920 , n15061 , n334922 , 
 n334923 , n334924 , n334925 , n15066 , n334927 , n334928 , n15069 , n334930 , n334931 , n15072 , 
 n334933 , n15074 , n334935 , n334936 , n334937 , n15078 , n334939 , n15080 , n15081 , n15082 , 
 n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n334949 , n334950 , n15091 , n334952 , 
 n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , 
 n15103 , n15104 , n15105 , n334966 , n15107 , n15108 , n15109 , n334970 , n15111 , n334972 , 
 n15113 , n15114 , n15115 , n334976 , n15117 , n334978 , n15119 , n334980 , n15121 , n334982 , 
 n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n334990 , n15131 , n334992 , 
 n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n334999 , n15140 , n335001 , n15142 , 
 n335003 , n335004 , n15145 , n15146 , n335007 , n335008 , n15149 , n335010 , n335011 , n15152 , 
 n335013 , n335014 , n15155 , n15156 , n335017 , n335018 , n15159 , n335020 , n15161 , n15162 , 
 n15163 , n15164 , n335025 , n15166 , n335027 , n15168 , n335029 , n15170 , n15171 , n15172 , 
 n335033 , n335034 , n15175 , n335036 , n335037 , n15178 , n15179 , n15180 , n15181 , n15182 , 
 n15183 , n15184 , n15185 , n15186 , n335047 , n335048 , n15189 , n335050 , n15191 , n335052 , 
 n15193 , n15194 , n335055 , n335056 , n15197 , n335058 , n335059 , n15200 , n335061 , n335062 , 
 n15203 , n15204 , n335065 , n335066 , n15207 , n335068 , n335069 , n15210 , n335071 , n335072 , 
 n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , 
 n15223 , n335084 , n15225 , n335086 , n335087 , n15228 , n335089 , n335090 , n15231 , n335092 , 
 n15233 , n15234 , n335095 , n15236 , n335097 , n15238 , n15239 , n335100 , n335101 , n335102 , 
 n15243 , n15244 , n335105 , n15246 , n15247 , n335108 , n335109 , n15250 , n335111 , n335112 , 
 n15253 , n335114 , n335115 , n15256 , n15257 , n15258 , n335119 , n15260 , n335121 , n15262 , 
 n15263 , n15264 , n335125 , n335126 , n15267 , n335128 , n15269 , n335130 , n15271 , n15272 , 
 n15273 , n335134 , n15275 , n335136 , n15277 , n335138 , n335139 , n15280 , n335141 , n335142 , 
 n15283 , n335144 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , 
 n15293 , n15294 , n335155 , n15296 , n15297 , n335158 , n15299 , n15300 , n335161 , n15302 , 
 n335163 , n335164 , n15305 , n15306 , n335167 , n335168 , n15309 , n335170 , n335171 , n15312 , 
 n335173 , n335174 , n335175 , n15316 , n335177 , n335178 , n335179 , n15320 , n335181 , n15322 , 
 n15323 , n15324 , n335185 , n15326 , n335187 , n335188 , n15329 , n15330 , n335191 , n335192 , 
 n15333 , n335194 , n15335 , n335196 , n15337 , n335198 , n335199 , n15340 , n15341 , n15342 , 
 n335203 , n335204 , n335205 , n335206 , n335207 , n335208 , n335209 , n15350 , n335211 , n335212 , 
 n15353 , n335214 , n335215 , n15356 , n335217 , n335218 , n335219 , n335220 , n15361 , n335222 , 
 n335223 , n15364 , n15365 , n15366 , n15367 , n15368 , n335229 , n335230 , n335231 , n15372 , 
 n15373 , n15374 , n335235 , n335236 , n335237 , n335238 , n335239 , n335240 , n15381 , n335242 , 
 n335243 , n15384 , n15385 , n335246 , n15387 , n335248 , n335249 , n335250 , n15391 , n335252 , 
 n335253 , n335254 , n335255 , n335256 , n335257 , n335258 , n335259 , n335260 , n335261 , n335262 , 
 n335263 , n335264 , n335265 , n335266 , n335267 , n335268 , n335269 , n335270 , n335271 , n15412 , 
 n15413 , n15414 , n335275 , n335276 , n335277 , n15418 , n335279 , n335280 , n15421 , n335282 , 
 n335283 , n335284 , n335285 , n335286 , n335287 , n335288 , n335289 , n15430 , n335291 , n335292 , 
 n335293 , n335294 , n335295 , n335296 , n335297 , n15438 , n15439 , n335300 , n335301 , n15442 , 
 n15443 , n335304 , n335305 , n335306 , n335307 , n335308 , n335309 , n335310 , n335311 , n15452 , 
 n335313 , n335314 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n335321 , n15462 , 
 n15463 , n335324 , n335325 , n335326 , n335327 , n15468 , n335329 , n15470 , n15471 , n335332 , 
 n335333 , n15474 , n335335 , n335336 , n15477 , n335338 , n15479 , n15480 , n15481 , n335342 , 
 n335343 , n335344 , n335345 , n335346 , n335347 , n335348 , n15489 , n15490 , n335351 , n15492 , 
 n335353 , n15494 , n335355 , n335356 , n15497 , n15498 , n335359 , n335360 , n335361 , n335362 , 
 n335363 , n15504 , n335365 , n335366 , n15507 , n335368 , n335369 , n335370 , n335371 , n335372 , 
 n15513 , n15514 , n15515 , n335376 , n15517 , n335378 , n335379 , n335380 , n335381 , n335382 , 
 n15523 , n335384 , n335385 , n335386 , n335387 , n15528 , n335389 , n335390 , n15531 , n335392 , 
 n335393 , n15534 , n335395 , n15536 , n335397 , n15538 , n335399 , n335400 , n335401 , n335402 , 
 n335403 , n335404 , n335405 , n335406 , n15547 , n335408 , n335409 , n335410 , n335411 , n335412 , 
 n335413 , n15554 , n335415 , n335416 , n335417 , n335418 , n335419 , n335420 , n335421 , n335422 , 
 n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n335431 , n335432 , 
 n15573 , n335434 , n335435 , n15576 , n335437 , n15578 , n335439 , n335440 , n335441 , n335442 , 
 n15583 , n335444 , n335445 , n15586 , n335447 , n335448 , n335449 , n335450 , n335451 , n335452 , 
 n15593 , n335454 , n335455 , n15596 , n335457 , n335458 , n335459 , n335460 , n335461 , n15602 , 
 n15603 , n15604 , n335465 , n15606 , n335467 , n15608 , n15609 , n335470 , n335471 , n335472 , 
 n335473 , n335474 , n335475 , n335476 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , 
 n15623 , n335484 , n335485 , n335486 , n335487 , n335488 , n335489 , n335490 , n15631 , n335492 , 
 n335493 , n15634 , n335495 , n335496 , n335497 , n15638 , n15639 , n15640 , n335501 , n15642 , 
 n335503 , n335504 , n335505 , n15646 , n335507 , n15648 , n335509 , n15650 , n15651 , n335512 , 
 n15653 , n335514 , n335515 , n15656 , n335517 , n15658 , n335519 , n335520 , n15661 , n335522 , 
 n335523 , n15664 , n15665 , n335526 , n335527 , n15668 , n335529 , n335530 , n15671 , n335532 , 
 n335533 , n15674 , n335535 , n15676 , n15677 , n15678 , n15679 , n15680 , n335541 , n15682 , 
 n15683 , n335544 , n335545 , n15686 , n335547 , n335548 , n15689 , n335550 , n335551 , n15692 , 
 n335553 , n335554 , n15695 , n335556 , n15697 , n15698 , n15699 , n15700 , n15701 , n335562 , 
 n335563 , n15704 , n335565 , n335566 , n15707 , n335568 , n335569 , n15710 , n15711 , n335572 , 
 n15713 , n15714 , n335575 , n335576 , n15717 , n15718 , n335579 , n15720 , n335581 , n15722 , 
 n335583 , n335584 , n15725 , n335586 , n15727 , n15728 , n335589 , n15730 , n335591 , n15732 , 
 n15733 , n335594 , n335595 , n15736 , n15737 , n335598 , n335599 , n335600 , n15741 , n15742 , 
 n335603 , n15744 , n335605 , n335606 , n15747 , n335608 , n15749 , n15750 , n335611 , n335612 , 
 n15753 , n335614 , n335615 , n15756 , n335617 , n335618 , n15759 , n15760 , n15761 , n15762 , 
 n15763 , n15764 , n15765 , n15766 , n15767 , n335628 , n335629 , n15770 , n335631 , n15772 , 
 n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , 
 n15783 , n15784 , n15785 , n335646 , n15787 , n335648 , n15789 , n335650 , n335651 , n15792 , 
 n335653 , n15794 , n15795 , n15796 , n335657 , n15798 , n335659 , n15800 , n335661 , n15802 , 
 n15803 , n335664 , n335665 , n15806 , n335667 , n335668 , n15809 , n335670 , n335671 , n15812 , 
 n15813 , n335674 , n335675 , n335676 , n335677 , n335678 , n15819 , n335680 , n15821 , n335682 , 
 n335683 , n335684 , n335685 , n15826 , n335687 , n15828 , n335689 , n335690 , n335691 , n335692 , 
 n335693 , n15834 , n335695 , n335696 , n335697 , n335698 , n335699 , n335700 , n335701 , n15842 , 
 n15843 , n335704 , n335705 , n15846 , n335707 , n335708 , n335709 , n335710 , n15851 , n335712 , 
 n15853 , n15854 , n335715 , n335716 , n335717 , n335718 , n335719 , n335720 , n335721 , n335722 , 
 n335723 , n15864 , n335725 , n335726 , n335727 , n335728 , n335729 , n335730 , n335731 , n335732 , 
 n335733 , n335734 , n335735 , n335736 , n335737 , n335738 , n335739 , n335740 , n335741 , n335742 , 
 n335743 , n15884 , n335745 , n335746 , n335747 , n15888 , n335749 , n335750 , n15891 , n15892 , 
 n335753 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n335762 , 
 n15903 , n15904 , n335765 , n15906 , n335767 , n15908 , n335769 , n335770 , n15911 , n335772 , 
 n335773 , n15914 , n335775 , n15916 , n335777 , n15918 , n335779 , n335780 , n15921 , n335782 , 
 n335783 , n15924 , n15925 , n335786 , n335787 , n335788 , n335789 , n335790 , n15931 , n15932 , 
 n335793 , n335794 , n335795 , n15936 , n335797 , n335798 , n15939 , n335800 , n335801 , n335802 , 
 n15943 , n335804 , n15945 , n335806 , n15947 , n335808 , n335809 , n15950 , n15951 , n335812 , 
 n335813 , n335814 , n335815 , n335816 , n335817 , n335818 , n335819 , n335820 , n335821 , n335822 , 
 n335823 , n15964 , n335825 , n335826 , n335827 , n335828 , n335829 , n335830 , n335831 , n15972 , 
 n335833 , n335834 , n15975 , n335836 , n335837 , n15978 , n335839 , n335840 , n335841 , n335842 , 
 n335843 , n335844 , n335845 , n335846 , n335847 , n335848 , n335849 , n335850 , n335851 , n15992 , 
 n335853 , n335854 , n335855 , n335856 , n335857 , n15998 , n335859 , n16000 , n16001 , n16002 , 
 n16003 , n335864 , n335865 , n335866 , n335867 , n335868 , n335869 , n335870 , n335871 , n335872 , 
 n335873 , n16014 , n335875 , n16016 , n335877 , n335878 , n335879 , n335880 , n335881 , n335882 , 
 n335883 , n335884 , n335885 , n335886 , n335887 , n335888 , n335889 , n335890 , n335891 , n16032 , 
 n16033 , n16034 , n335895 , n335896 , n335897 , n16038 , n335899 , n335900 , n16041 , n335902 , 
 n16043 , n16044 , n16045 , n335906 , n16047 , n16048 , n335909 , n16050 , n335911 , n335912 , 
 n16053 , n335914 , n335915 , n335916 , n16057 , n335918 , n335919 , n16060 , n335921 , n335922 , 
 n16063 , n335924 , n335925 , n335926 , n335927 , n335928 , n335929 , n335930 , n335931 , n335932 , 
 n335933 , n335934 , n16075 , n335936 , n335937 , n335938 , n335939 , n335940 , n335941 , n335942 , 
 n335943 , n16084 , n335945 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , 
 n16093 , n16094 , n16095 , n335956 , n16097 , n335958 , n16099 , n335960 , n335961 , n16102 , 
 n335963 , n335964 , n16105 , n335966 , n16107 , n335968 , n335969 , n335970 , n335971 , n335972 , 
 n335973 , n335974 , n16115 , n335976 , n16117 , n16118 , n335979 , n335980 , n335981 , n335982 , 
 n16123 , n335984 , n335985 , n335986 , n335987 , n16128 , n16129 , n335990 , n16131 , n335992 , 
 n16133 , n16134 , n335995 , n16136 , n335997 , n16138 , n335999 , n336000 , n336001 , n336002 , 
 n16143 , n336004 , n336005 , n16146 , n336007 , n336008 , n336009 , n16150 , n16151 , n336012 , 
 n16153 , n336014 , n336015 , n16156 , n16157 , n336018 , n336019 , n336020 , n336021 , n336022 , 
 n16163 , n336024 , n336025 , n16166 , n16167 , n336028 , n16169 , n336030 , n336031 , n336032 , 
 n16173 , n336034 , n336035 , n336036 , n336037 , n336038 , n336039 , n336040 , n336041 , n336042 , 
 n336043 , n16184 , n336045 , n16186 , n336047 , n336048 , n16189 , n336050 , n336051 , n336052 , 
 n336053 , n336054 , n16195 , n336056 , n336057 , n16198 , n16199 , n16200 , n16201 , n336062 , 
 n336063 , n336064 , n336065 , n16206 , n336067 , n336068 , n336069 , n16210 , n336071 , n336072 , 
 n16213 , n336074 , n336075 , n336076 , n336077 , n336078 , n336079 , n336080 , n16221 , n16222 , 
 n16223 , n16224 , n16225 , n16226 , n16227 , n336088 , n336089 , n336090 , n336091 , n336092 , 
 n336093 , n336094 , n336095 , n16236 , n16237 , n336098 , n16239 , n336100 , n336101 , n16242 , 
 n16243 , n336104 , n16245 , n336106 , n336107 , n336108 , n336109 , n336110 , n336111 , n336112 , 
 n16253 , n16254 , n336115 , n16256 , n336117 , n336118 , n16259 , n336120 , n336121 , n16262 , 
 n336123 , n336124 , n336125 , n16266 , n336127 , n336128 , n16269 , n336130 , n336131 , n16272 , 
 n336133 , n16274 , n336135 , n336136 , n16277 , n16278 , n336139 , n336140 , n16281 , n336142 , 
 n336143 , n16284 , n336145 , n336146 , n336147 , n336148 , n336149 , n336150 , n336151 , n336152 , 
 n336153 , n336154 , n336155 , n336156 , n336157 , n336158 , n16299 , n336160 , n16301 , n16302 , 
 n336163 , n336164 , n336165 , n16306 , n336167 , n336168 , n16309 , n336170 , n336171 , n336172 , 
 n336173 , n336174 , n336175 , n16316 , n336177 , n336178 , n336179 , n336180 , n336181 , n336182 , 
 n16323 , n336184 , n336185 , n336186 , n16327 , n336188 , n16329 , n336190 , n16331 , n336192 , 
 n336193 , n336194 , n336195 , n16336 , n336197 , n336198 , n336199 , n16340 , n336201 , n16342 , 
 n336203 , n336204 , n16345 , n336206 , n336207 , n336208 , n336209 , n336210 , n16351 , n16352 , 
 n16353 , n16354 , n16355 , n16356 , n336217 , n16358 , n336219 , n336220 , n16361 , n336222 , 
 n16363 , n336224 , n336225 , n16366 , n336227 , n336228 , n336229 , n336230 , n336231 , n336232 , 
 n16373 , n336234 , n336235 , n336236 , n336237 , n336238 , n336239 , n16380 , n336241 , n16382 , 
 n336243 , n336244 , n16385 , n336246 , n16387 , n336248 , n336249 , n336250 , n336251 , n336252 , 
 n336253 , n336254 , n336255 , n336256 , n336257 , n336258 , n336259 , n336260 , n16401 , n336262 , 
 n336263 , n336264 , n336265 , n336266 , n16407 , n16408 , n336269 , n16410 , n16411 , n336272 , 
 n336273 , n16414 , n336275 , n336276 , n336277 , n336278 , n336279 , n336280 , n336281 , n336282 , 
 n336283 , n336284 , n16425 , n336286 , n336287 , n336288 , n336289 , n16430 , n336291 , n336292 , 
 n336293 , n336294 , n336295 , n336296 , n336297 , n336298 , n336299 , n336300 , n336301 , n336302 , 
 n336303 , n16444 , n336305 , n16446 , n16447 , n16448 , n16449 , n16450 , n336311 , n16452 , 
 n16453 , n336314 , n16455 , n16456 , n336317 , n16458 , n336319 , n336320 , n16461 , n16462 , 
 n336323 , n336324 , n16465 , n336326 , n336327 , n16468 , n336329 , n336330 , n336331 , n16472 , 
 n336333 , n336334 , n16475 , n336336 , n336337 , n336338 , n336339 , n16480 , n336341 , n336342 , 
 n16483 , n16484 , n336345 , n16486 , n16487 , n336348 , n336349 , n16490 , n336351 , n336352 , 
 n16493 , n336354 , n336355 , n16496 , n336357 , n336358 , n336359 , n16500 , n336361 , n336362 , 
 n16503 , n16504 , n16505 , n16506 , n16507 , n336368 , n16509 , n16510 , n336371 , n336372 , 
 n16513 , n336374 , n336375 , n16516 , n336377 , n336378 , n16519 , n336380 , n16521 , n336382 , 
 n16523 , n16524 , n16525 , n16526 , n16527 , n336388 , n16529 , n16530 , n336391 , n336392 , 
 n16533 , n336394 , n336395 , n16536 , n336397 , n16538 , n16539 , n16540 , n336401 , n16542 , 
 n336403 , n336404 , n16545 , n16546 , n16547 , n16548 , n336409 , n336410 , n16551 , n16552 , 
 n16553 , n16554 , n16555 , n336416 , n336417 , n336418 , n336419 , n336420 , n336421 , n16562 , 
 n336423 , n336424 , n336425 , n336426 , n336427 , n16568 , n336429 , n336430 , n336431 , n336432 , 
 n336433 , n336434 , n16575 , n16576 , n336437 , n336438 , n336439 , n336440 , n336441 , n336442 , 
 n336443 , n336444 , n336445 , n336446 , n16587 , n336448 , n16589 , n16590 , n336451 , n16592 , 
 n336453 , n336454 , n336455 , n336456 , n336457 , n336458 , n336459 , n336460 , n16601 , n16602 , 
 n336463 , n336464 , n336465 , n336466 , n336467 , n336468 , n16609 , n336470 , n336471 , n336472 , 
 n336473 , n336474 , n336475 , n336476 , n336477 , n16618 , n336479 , n336480 , n16621 , n336482 , 
 n336483 , n16624 , n16625 , n336486 , n336487 , n16628 , n336489 , n336490 , n16631 , n336492 , 
 n336493 , n16634 , n336495 , n336496 , n16637 , n336498 , n336499 , n16640 , n336501 , n336502 , 
 n16643 , n336504 , n16645 , n336506 , n16647 , n336508 , n16649 , n336510 , n336511 , n336512 , 
 n336513 , n336514 , n336515 , n16656 , n336517 , n336518 , n16659 , n16660 , n336521 , n336522 , 
 n16663 , n336524 , n336525 , n16666 , n16667 , n336528 , n16669 , n336530 , n336531 , n16672 , 
 n336533 , n336534 , n336535 , n16676 , n16677 , n336538 , n336539 , n336540 , n336541 , n16682 , 
 n336543 , n16684 , n336545 , n16686 , n336547 , n16688 , n336549 , n336550 , n336551 , n336552 , 
 n16693 , n336554 , n336555 , n16696 , n336557 , n336558 , n16699 , n336560 , n336561 , n16702 , 
 n16703 , n336564 , n336565 , n336566 , n16707 , n336568 , n336569 , n336570 , n336571 , n336572 , 
 n336573 , n336574 , n16715 , n336576 , n336577 , n16718 , n16719 , n16720 , n16721 , n336582 , 
 n336583 , n16724 , n336585 , n336586 , n16727 , n336588 , n336589 , n16730 , n16731 , n16732 , 
 n336593 , n16734 , n16735 , n336596 , n336597 , n16738 , n336599 , n336600 , n336601 , n336602 , 
 n336603 , n16744 , n336605 , n16746 , n336607 , n336608 , n336609 , n16750 , n336611 , n336612 , 
 n336613 , n16754 , n336615 , n336616 , n16757 , n336618 , n336619 , n336620 , n16761 , n336622 , 
 n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n336629 , n336630 , n16771 , n336632 , 
 n16773 , n16774 , n16775 , n336636 , n16777 , n336638 , n16779 , n16780 , n336641 , n336642 , 
 n16783 , n336644 , n336645 , n16786 , n336647 , n16788 , n16789 , n16790 , n16791 , n16792 , 
 n336653 , n16794 , n16795 , n336656 , n16797 , n16798 , n16799 , n336660 , n16801 , n336662 , 
 n336663 , n16804 , n336665 , n336666 , n16807 , n336668 , n16809 , n336670 , n336671 , n16812 , 
 n336673 , n16814 , n336675 , n336676 , n336677 , n16818 , n336679 , n16820 , n336681 , n16822 , 
 n16823 , n16824 , n16825 , n336686 , n336687 , n16828 , n336689 , n336690 , n16831 , n336692 , 
 n336693 , n16834 , n336695 , n336696 , n16837 , n16838 , n16839 , n16840 , n336701 , n16842 , 
 n16843 , n336704 , n16845 , n16846 , n336707 , n336708 , n16849 , n336710 , n336711 , n16852 , 
 n336713 , n336714 , n336715 , n16856 , n336717 , n16858 , n336719 , n16860 , n16861 , n336722 , 
 n16863 , n336724 , n16865 , n336726 , n336727 , n16868 , n336729 , n336730 , n16871 , n16872 , 
 n16873 , n16874 , n336735 , n16876 , n336737 , n16878 , n16879 , n336740 , n336741 , n16882 , 
 n336743 , n336744 , n16885 , n336746 , n336747 , n336748 , n16889 , n336750 , n16891 , n16892 , 
 n336753 , n16894 , n336755 , n336756 , n336757 , n336758 , n16899 , n336760 , n336761 , n16902 , 
 n336763 , n16904 , n336765 , n336766 , n16907 , n336768 , n16909 , n16910 , n336771 , n336772 , 
 n336773 , n16914 , n336775 , n16916 , n336777 , n336778 , n16919 , n336780 , n336781 , n336782 , 
 n336783 , n336784 , n16925 , n336786 , n336787 , n16928 , n336789 , n336790 , n336791 , n16932 , 
 n16933 , n336794 , n16935 , n336796 , n336797 , n336798 , n336799 , n336800 , n16941 , n336802 , 
 n336803 , n16944 , n336805 , n16946 , n336807 , n336808 , n16949 , n336810 , n16951 , n336812 , 
 n336813 , n16954 , n336815 , n16956 , n16957 , n336818 , n336819 , n336820 , n16961 , n336822 , 
 n336823 , n16964 , n336825 , n336826 , n336827 , n336828 , n336829 , n336830 , n16971 , n336832 , 
 n16973 , n16974 , n336835 , n336836 , n336837 , n336838 , n336839 , n336840 , n16981 , n16982 , 
 n16983 , n16984 , n336845 , n336846 , n16987 , n336848 , n336849 , n16990 , n336851 , n16992 , 
 n16993 , n336854 , n16995 , n336856 , n16997 , n16998 , n336859 , n336860 , n336861 , n17002 , 
 n336863 , n336864 , n336865 , n336866 , n336867 , n336868 , n336869 , n17010 , n17011 , n336872 , 
 n336873 , n17014 , n336875 , n336876 , n17017 , n336878 , n336879 , n336880 , n336881 , n336882 , 
 n17023 , n336884 , n336885 , n336886 , n336887 , n336888 , n17029 , n336890 , n336891 , n336892 , 
 n336893 , n336894 , n336895 , n336896 , n336897 , n336898 , n336899 , n17040 , n17041 , n336902 , 
 n17043 , n336904 , n336905 , n17046 , n336907 , n336908 , n336909 , n336910 , n17051 , n336912 , 
 n336913 , n336914 , n17055 , n336916 , n17057 , n17058 , n17059 , n336920 , n336921 , n336922 , 
 n336923 , n17064 , n17065 , n17066 , n17067 , n17068 , n336929 , n336930 , n336931 , n336932 , 
 n336933 , n17074 , n336935 , n336936 , n336937 , n336938 , n336939 , n336940 , n336941 , n17082 , 
 n336943 , n17084 , n336945 , n336946 , n336947 , n336948 , n17089 , n336950 , n336951 , n336952 , 
 n336953 , n336954 , n336955 , n17096 , n336957 , n336958 , n336959 , n336960 , n17101 , n336962 , 
 n336963 , n17104 , n336965 , n336966 , n17107 , n336968 , n336969 , n17110 , n17111 , n336972 , 
 n336973 , n17114 , n336975 , n336976 , n17117 , n336978 , n336979 , n17120 , n336981 , n17122 , 
 n336983 , n17124 , n17125 , n336986 , n17127 , n336988 , n17129 , n336990 , n17131 , n17132 , 
 n336993 , n17134 , n336995 , n17136 , n17137 , n336998 , n336999 , n17140 , n337001 , n337002 , 
 n17143 , n337004 , n337005 , n17146 , n337007 , n17148 , n337009 , n17150 , n337011 , n17152 , 
 n17153 , n17154 , n17155 , n337016 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , 
 n17163 , n17164 , n17165 , n17166 , n17167 , n337028 , n337029 , n17170 , n337031 , n337032 , 
 n17173 , n337034 , n17175 , n17176 , n337037 , n337038 , n17179 , n337040 , n17181 , n337042 , 
 n337043 , n17184 , n337045 , n17186 , n337047 , n337048 , n17189 , n337050 , n337051 , n337052 , 
 n337053 , n337054 , n337055 , n337056 , n337057 , n337058 , n337059 , n337060 , n337061 , n17202 , 
 n337063 , n17204 , n337065 , n337066 , n337067 , n17208 , n337069 , n17210 , n17211 , n337072 , 
 n337073 , n337074 , n17215 , n337076 , n337077 , n337078 , n337079 , n17220 , n337081 , n337082 , 
 n337083 , n17224 , n337085 , n337086 , n17227 , n337088 , n337089 , n337090 , n17231 , n337092 , 
 n337093 , n17234 , n337095 , n337096 , n337097 , n337098 , n337099 , n17240 , n337101 , n337102 , 
 n337103 , n337104 , n337105 , n337106 , n337107 , n337108 , n337109 , n337110 , n337111 , n337112 , 
 n17253 , n17254 , n337115 , n337116 , n17257 , n337118 , n337119 , n17260 , n337121 , n17262 , 
 n17263 , n337124 , n337125 , n17266 , n337127 , n337128 , n337129 , n337130 , n337131 , n17272 , 
 n337133 , n17274 , n337135 , n337136 , n337137 , n337138 , n17279 , n337140 , n17281 , n337142 , 
 n17283 , n337144 , n337145 , n337146 , n337147 , n17288 , n337149 , n337150 , n17291 , n337152 , 
 n337153 , n17294 , n337155 , n337156 , n17297 , n17298 , n17299 , n17300 , n337161 , n17302 , 
 n337163 , n17304 , n337165 , n337166 , n337167 , n17308 , n337169 , n337170 , n337171 , n337172 , 
 n337173 , n337174 , n337175 , n17316 , n337177 , n17318 , n17319 , n337180 , n337181 , n17322 , 
 n337183 , n337184 , n337185 , n17326 , n337187 , n337188 , n17329 , n337190 , n337191 , n17332 , 
 n337193 , n17334 , n337195 , n337196 , n337197 , n337198 , n337199 , n337200 , n337201 , n337202 , 
 n337203 , n337204 , n17345 , n337206 , n337207 , n17348 , n337209 , n17350 , n337211 , n17352 , 
 n17353 , n17354 , n337215 , n17356 , n337217 , n17358 , n17359 , n337220 , n17361 , n337222 , 
 n17363 , n17364 , n337225 , n337226 , n17367 , n337228 , n337229 , n17370 , n337231 , n17372 , 
 n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , 
 n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n337250 , n17391 , n337252 , 
 n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n337261 , n337262 , 
 n17403 , n337264 , n17405 , n337266 , n17407 , n337268 , n17409 , n17410 , n17411 , n17412 , 
 n17413 , n17414 , n17415 , n17416 , n337277 , n337278 , n337279 , n337280 , n17421 , n337282 , 
 n337283 , n337284 , n337285 , n337286 , n17427 , n17428 , n337289 , n17430 , n337291 , n17432 , 
 n17433 , n337294 , n17435 , n337296 , n337297 , n337298 , n337299 , n17440 , n337301 , n337302 , 
 n337303 , n17444 , n337305 , n337306 , n17447 , n337308 , n17449 , n17450 , n337311 , n337312 , 
 n337313 , n337314 , n17455 , n17456 , n337317 , n337318 , n337319 , n337320 , n337321 , n337322 , 
 n337323 , n337324 , n337325 , n337326 , n337327 , n17468 , n17469 , n337330 , n17471 , n337332 , 
 n337333 , n17474 , n337335 , n337336 , n337337 , n337338 , n17479 , n337340 , n17481 , n337342 , 
 n337343 , n337344 , n337345 , n337346 , n337347 , n337348 , n337349 , n337350 , n337351 , n337352 , 
 n17493 , n337354 , n337355 , n337356 , n337357 , n337358 , n337359 , n337360 , n337361 , n337362 , 
 n337363 , n337364 , n337365 , n337366 , n17507 , n337368 , n337369 , n337370 , n337371 , n17512 , 
 n337373 , n337374 , n337375 , n337376 , n337377 , n337378 , n337379 , n17520 , n17521 , n337382 , 
 n17523 , n337384 , n337385 , n337386 , n337387 , n337388 , n337389 , n337390 , n337391 , n337392 , 
 n17533 , n337394 , n337395 , n337396 , n17537 , n337398 , n17539 , n17540 , n337401 , n337402 , 
 n337403 , n17544 , n337405 , n17546 , n337407 , n337408 , n337409 , n337410 , n337411 , n337412 , 
 n337413 , n337414 , n17555 , n337416 , n337417 , n337418 , n337419 , n17560 , n337421 , n337422 , 
 n17563 , n337424 , n337425 , n17566 , n17567 , n337428 , n17569 , n337430 , n337431 , n337432 , 
 n337433 , n337434 , n337435 , n337436 , n337437 , n337438 , n337439 , n337440 , n337441 , n17582 , 
 n337443 , n337444 , n337445 , n337446 , n337447 , n337448 , n337449 , n337450 , n337451 , n337452 , 
 n337453 , n17594 , n17595 , n337456 , n337457 , n337458 , n17599 , n337460 , n17601 , n17602 , 
 n337463 , n337464 , n337465 , n337466 , n17607 , n337468 , n337469 , n337470 , n337471 , n337472 , 
 n337473 , n337474 , n17615 , n17616 , n337477 , n337478 , n337479 , n337480 , n17621 , n337482 , 
 n337483 , n17624 , n17625 , n337486 , n337487 , n17628 , n337489 , n337490 , n337491 , n17632 , 
 n337493 , n337494 , n337495 , n337496 , n17637 , n337498 , n337499 , n337500 , n17641 , n337502 , 
 n337503 , n337504 , n337505 , n337506 , n17647 , n337508 , n337509 , n337510 , n337511 , n337512 , 
 n337513 , n337514 , n337515 , n337516 , n17657 , n337518 , n337519 , n337520 , n337521 , n17662 , 
 n337523 , n337524 , n17665 , n17666 , n17667 , n17668 , n17669 , n337530 , n337531 , n17672 , 
 n337533 , n337534 , n17675 , n17676 , n17677 , n337538 , n17679 , n337540 , n337541 , n17682 , 
 n337543 , n337544 , n337545 , n337546 , n337547 , n337548 , n337549 , n17690 , n337551 , n337552 , 
 n337553 , n337554 , n17695 , n337556 , n17697 , n17698 , n337559 , n337560 , n337561 , n17702 , 
 n337563 , n337564 , n17705 , n337566 , n337567 , n17708 , n337569 , n17710 , n337571 , n17712 , 
 n17713 , n337574 , n17715 , n337576 , n17717 , n17718 , n337579 , n337580 , n17721 , n337582 , 
 n337583 , n17724 , n337585 , n337586 , n337587 , n17728 , n337589 , n337590 , n17731 , n337592 , 
 n337593 , n17734 , n17735 , n337596 , n337597 , n17738 , n17739 , n17740 , n17741 , n17742 , 
 n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , 
 n337613 , n337614 , n17755 , n337616 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , 
 n17763 , n337624 , n17765 , n337626 , n17767 , n17768 , n17769 , n17770 , n17771 , n337632 , 
 n337633 , n17774 , n337635 , n337636 , n17777 , n337638 , n337639 , n17780 , n17781 , n337642 , 
 n337643 , n17784 , n337645 , n17786 , n337647 , n17788 , n17789 , n17790 , n17791 , n17792 , 
 n337653 , n17794 , n337655 , n17796 , n337657 , n17798 , n337659 , n337660 , n17801 , n337662 , 
 n337663 , n17804 , n337665 , n337666 , n17807 , n17808 , n17809 , n337670 , n337671 , n337672 , 
 n17813 , n337674 , n17815 , n17816 , n337677 , n337678 , n17819 , n337680 , n17821 , n17822 , 
 n17823 , n17824 , n337685 , n17826 , n337687 , n337688 , n17829 , n337690 , n337691 , n17832 , 
 n337693 , n17834 , n337695 , n337696 , n337697 , n337698 , n17839 , n337700 , n337701 , n17842 , 
 n337703 , n337704 , n337705 , n337706 , n17847 , n337708 , n337709 , n337710 , n337711 , n17852 , 
 n17853 , n337714 , n337715 , n337716 , n337717 , n337718 , n17859 , n17860 , n337721 , n17862 , 
 n17863 , n337724 , n337725 , n337726 , n337727 , n17868 , n337729 , n337730 , n337731 , n337732 , 
 n337733 , n337734 , n337735 , n337736 , n337737 , n337738 , n337739 , n337740 , n17881 , n337742 , 
 n17883 , n337744 , n337745 , n17886 , n337747 , n337748 , n337749 , n337750 , n17891 , n337752 , 
 n337753 , n337754 , n17895 , n337756 , n337757 , n337758 , n337759 , n17900 , n337761 , n337762 , 
 n337763 , n337764 , n337765 , n337766 , n337767 , n337768 , n337769 , n337770 , n337771 , n337772 , 
 n17913 , n337774 , n337775 , n337776 , n337777 , n337778 , n337779 , n337780 , n337781 , n337782 , 
 n17923 , n337784 , n17925 , n17926 , n17927 , n17928 , n337789 , n17930 , n17931 , n337792 , 
 n17933 , n17934 , n337795 , n337796 , n17937 , n17938 , n337799 , n337800 , n17941 , n337802 , 
 n337803 , n17944 , n337805 , n337806 , n17947 , n17948 , n337809 , n17950 , n337811 , n337812 , 
 n17953 , n337814 , n337815 , n17956 , n337817 , n337818 , n337819 , n17960 , n337821 , n337822 , 
 n17963 , n337824 , n337825 , n17966 , n337827 , n17968 , n337829 , n337830 , n17971 , n337832 , 
 n337833 , n17974 , n337835 , n337836 , n17977 , n337838 , n17979 , n17980 , n337841 , n17982 , 
 n337843 , n337844 , n337845 , n17986 , n337847 , n17988 , n17989 , n17990 , n17991 , n17992 , 
 n17993 , n337854 , n17995 , n17996 , n17997 , n17998 , n337859 , n337860 , n337861 , n18002 , 
 n337863 , n18004 , n18005 , n337866 , n337867 , n18008 , n337869 , n337870 , n18011 , n337872 , 
 n337873 , n18014 , n337875 , n18016 , n337877 , n18018 , n18019 , n337880 , n337881 , n18022 , 
 n337883 , n337884 , n18025 , n337886 , n337887 , n18028 , n337889 , n337890 , n18031 , n337892 , 
 n18033 , n337894 , n337895 , n18036 , n337897 , n18038 , n18039 , n337900 , n18041 , n337902 , 
 n337903 , n337904 , n18045 , n18046 , n337907 , n337908 , n18049 , n337910 , n18051 , n18052 , 
 n337913 , n337914 , n18055 , n18056 , n337917 , n337918 , n18059 , n337920 , n18061 , n18062 , 
 n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , 
 n18073 , n18074 , n18075 , n18076 , n18077 , n337938 , n18079 , n18080 , n18081 , n18082 , 
 n18083 , n337944 , n18085 , n18086 , n337947 , n18088 , n337949 , n18090 , n18091 , n337952 , 
 n337953 , n18094 , n337955 , n337956 , n18097 , n337958 , n337959 , n337960 , n18101 , n337962 , 
 n337963 , n18104 , n337965 , n337966 , n18107 , n18108 , n337969 , n337970 , n337971 , n18112 , 
 n337973 , n18114 , n337975 , n18116 , n18117 , n337978 , n337979 , n18120 , n337981 , n337982 , 
 n18123 , n337984 , n337985 , n18126 , n18127 , n337988 , n18129 , n337990 , n18131 , n18132 , 
 n18133 , n18134 , n337995 , n18136 , n337997 , n337998 , n18139 , n18140 , n338001 , n338002 , 
 n18143 , n18144 , n18145 , n18146 , n18147 , n338008 , n18149 , n18150 , n338011 , n18152 , 
 n338013 , n18154 , n338015 , n338016 , n18157 , n18158 , n338019 , n338020 , n18161 , n338022 , 
 n338023 , n18164 , n338025 , n338026 , n338027 , n338028 , n338029 , n338030 , n18171 , n338032 , 
 n338033 , n338034 , n338035 , n18176 , n338037 , n18178 , n338039 , n338040 , n338041 , n338042 , 
 n18183 , n338044 , n18185 , n338046 , n338047 , n18188 , n338049 , n338050 , n18191 , n338052 , 
 n338053 , n18194 , n338055 , n18196 , n338057 , n18198 , n18199 , n338060 , n338061 , n18202 , 
 n338063 , n338064 , n18205 , n18206 , n338067 , n338068 , n338069 , n18210 , n338071 , n338072 , 
 n18213 , n338074 , n338075 , n18216 , n18217 , n338078 , n338079 , n338080 , n338081 , n338082 , 
 n18223 , n338084 , n338085 , n338086 , n338087 , n338088 , n18229 , n338090 , n338091 , n338092 , 
 n338093 , n338094 , n338095 , n338096 , n338097 , n338098 , n338099 , n338100 , n338101 , n18242 , 
 n338103 , n338104 , n338105 , n18246 , n18247 , n338108 , n338109 , n18250 , n338111 , n338112 , 
 n18253 , n338114 , n338115 , n338116 , n338117 , n338118 , n338119 , n18260 , n338121 , n338122 , 
 n18263 , n338124 , n338125 , n18266 , n18267 , n338128 , n18269 , n338130 , n338131 , n338132 , 
 n338133 , n18274 , n18275 , n338136 , n338137 , n338138 , n338139 , n18280 , n338141 , n338142 , 
 n338143 , n18284 , n338145 , n338146 , n338147 , n338148 , n338149 , n338150 , n18291 , n338152 , 
 n18293 , n338154 , n338155 , n338156 , n338157 , n338158 , n338159 , n338160 , n338161 , n338162 , 
 n338163 , n338164 , n338165 , n338166 , n338167 , n18308 , n18309 , n338170 , n18311 , n18312 , 
 n338173 , n338174 , n18315 , n338176 , n338177 , n18318 , n18319 , n338180 , n338181 , n338182 , 
 n338183 , n338184 , n338185 , n338186 , n338187 , n18328 , n338189 , n338190 , n18331 , n338192 , 
 n338193 , n338194 , n338195 , n338196 , n338197 , n338198 , n338199 , n338200 , n338201 , n18342 , 
 n18343 , n18344 , n338205 , n338206 , n338207 , n338208 , n338209 , n338210 , n338211 , n18352 , 
 n18353 , n18354 , n338215 , n338216 , n18357 , n338218 , n18359 , n338220 , n338221 , n338222 , 
 n338223 , n18364 , n18365 , n338226 , n338227 , n338228 , n338229 , n338230 , n338231 , n338232 , 
 n18373 , n338234 , n338235 , n338236 , n18377 , n338238 , n338239 , n18380 , n338241 , n338242 , 
 n338243 , n338244 , n338245 , n338246 , n338247 , n338248 , n338249 , n18390 , n338251 , n338252 , 
 n338253 , n18394 , n338255 , n338256 , n338257 , n338258 , n338259 , n338260 , n18401 , n338262 , 
 n338263 , n18404 , n338265 , n18406 , n338267 , n18408 , n338269 , n338270 , n338271 , n338272 , 
 n338273 , n338274 , n338275 , n18416 , n338277 , n18418 , n338279 , n18420 , n338281 , n338282 , 
 n338283 , n338284 , n338285 , n338286 , n338287 , n338288 , n338289 , n338290 , n338291 , n338292 , 
 n338293 , n338294 , n338295 , n338296 , n18437 , n338298 , n18439 , n338300 , n18441 , n338302 , 
 n338303 , n18444 , n338305 , n18446 , n338307 , n338308 , n338309 , n338310 , n338311 , n338312 , 
 n338313 , n338314 , n18455 , n338316 , n338317 , n338318 , n338319 , n18460 , n338321 , n338322 , 
 n18463 , n338324 , n338325 , n338326 , n338327 , n338328 , n338329 , n338330 , n18471 , n338332 , 
 n338333 , n338334 , n338335 , n338336 , n338337 , n338338 , n338339 , n338340 , n338341 , n338342 , 
 n338343 , n338344 , n338345 , n338346 , n338347 , n338348 , n338349 , n338350 , n338351 , n338352 , 
 n18493 , n338354 , n18495 , n338356 , n338357 , n338358 , n18499 , n338360 , n338361 , n338362 , 
 n18503 , n338364 , n338365 , n338366 , n18507 , n338368 , n338369 , n338370 , n338371 , n338372 , 
 n18513 , n338374 , n338375 , n18516 , n338377 , n338378 , n18519 , n338380 , n338381 , n18522 , 
 n338383 , n338384 , n338385 , n338386 , n18527 , n338388 , n338389 , n338390 , n338391 , n338392 , 
 n338393 , n338394 , n338395 , n18536 , n338397 , n338398 , n338399 , n338400 , n338401 , n338402 , 
 n338403 , n18544 , n18545 , n338406 , n338407 , n338408 , n338409 , n18550 , n338411 , n338412 , 
 n338413 , n338414 , n338415 , n18556 , n338417 , n338418 , n18559 , n18560 , n338421 , n18562 , 
 n338423 , n18564 , n18565 , n338426 , n338427 , n18568 , n338429 , n338430 , n338431 , n18572 , 
 n338433 , n338434 , n338435 , n338436 , n338437 , n338438 , n338439 , n338440 , n338441 , n338442 , 
 n338443 , n338444 , n338445 , n338446 , n338447 , n18588 , n338449 , n18590 , n18591 , n338452 , 
 n338453 , n18594 , n338455 , n18596 , n338457 , n338458 , n338459 , n338460 , n18601 , n18602 , 
 n338463 , n18604 , n338465 , n338466 , n338467 , n18608 , n18609 , n338470 , n18611 , n338472 , 
 n18613 , n338474 , n338475 , n338476 , n338477 , n338478 , n338479 , n338480 , n338481 , n18622 , 
 n338483 , n338484 , n338485 , n338486 , n18627 , n338488 , n338489 , n18630 , n338491 , n18632 , 
 n338493 , n338494 , n338495 , n338496 , n338497 , n338498 , n338499 , n338500 , n338501 , n338502 , 
 n338503 , n338504 , n338505 , n338506 , n338507 , n338508 , n338509 , n338510 , n18651 , n338512 , 
 n338513 , n338514 , n338515 , n338516 , n338517 , n338518 , n338519 , n338520 , n338521 , n338522 , 
 n18663 , n338524 , n338525 , n18666 , n18667 , n338528 , n338529 , n338530 , n338531 , n338532 , 
 n18673 , n18674 , n338535 , n18676 , n338537 , n338538 , n18679 , n338540 , n18681 , n338542 , 
 n338543 , n18684 , n338545 , n338546 , n338547 , n18688 , n18689 , n18690 , n338551 , n18692 , 
 n338553 , n338554 , n338555 , n338556 , n338557 , n338558 , n338559 , n18700 , n338561 , n338562 , 
 n18703 , n338564 , n338565 , n338566 , n338567 , n18708 , n18709 , n18710 , n18711 , n338572 , 
 n338573 , n338574 , n338575 , n338576 , n338577 , n338578 , n338579 , n338580 , n338581 , n18722 , 
 n338583 , n18724 , n338585 , n338586 , n338587 , n338588 , n18729 , n338590 , n338591 , n338592 , 
 n338593 , n338594 , n338595 , n338596 , n338597 , n338598 , n18739 , n338600 , n338601 , n18742 , 
 n338603 , n338604 , n18745 , n338606 , n338607 , n18748 , n338609 , n338610 , n338611 , n338612 , 
 n18753 , n338614 , n338615 , n338616 , n338617 , n338618 , n18759 , n338620 , n338621 , n338622 , 
 n338623 , n338624 , n338625 , n338626 , n338627 , n18768 , n18769 , n18770 , n338631 , n18772 , 
 n338633 , n338634 , n338635 , n18776 , n338637 , n338638 , n338639 , n338640 , n338641 , n338642 , 
 n338643 , n338644 , n338645 , n338646 , n338647 , n18788 , n338649 , n338650 , n18791 , n338652 , 
 n338653 , n338654 , n18795 , n338656 , n338657 , n18798 , n338659 , n338660 , n338661 , n338662 , 
 n338663 , n338664 , n338665 , n338666 , n18807 , n338668 , n338669 , n338670 , n18811 , n338672 , 
 n338673 , n338674 , n338675 , n338676 , n338677 , n18818 , n18819 , n338680 , n18821 , n338682 , 
 n18823 , n338684 , n338685 , n18826 , n18827 , n18828 , n338689 , n338690 , n18831 , n18832 , 
 n338693 , n18834 , n338695 , n338696 , n338697 , n338698 , n18839 , n338700 , n338701 , n338702 , 
 n338703 , n338704 , n18845 , n18846 , n18847 , n18848 , n338709 , n18850 , n338711 , n338712 , 
 n18853 , n338714 , n338715 , n338716 , n338717 , n338718 , n338719 , n338720 , n338721 , n338722 , 
 n338723 , n338724 , n338725 , n338726 , n18867 , n18868 , n18869 , n338730 , n338731 , n338732 , 
 n18873 , n338734 , n338735 , n338736 , n338737 , n338738 , n338739 , n338740 , n338741 , n338742 , 
 n18883 , n18884 , n18885 , n338746 , n18887 , n338748 , n338749 , n18890 , n338751 , n338752 , 
 n18893 , n338754 , n338755 , n338756 , n338757 , n338758 , n338759 , n338760 , n338761 , n338762 , 
 n338763 , n338764 , n338765 , n338766 , n338767 , n18908 , n338769 , n338770 , n18911 , n338772 , 
 n338773 , n338774 , n338775 , n338776 , n18917 , n338778 , n338779 , n338780 , n338781 , n338782 , 
 n18923 , n18924 , n338785 , n338786 , n338787 , n338788 , n338789 , n18930 , n338791 , n18932 , 
 n338793 , n338794 , n18935 , n338796 , n18937 , n338798 , n338799 , n18940 , n338801 , n18942 , 
 n338803 , n338804 , n338805 , n18946 , n338807 , n338808 , n18949 , n18950 , n338811 , n338812 , 
 n338813 , n338814 , n338815 , n338816 , n18957 , n338818 , n338819 , n338820 , n338821 , n338822 , 
 n18963 , n338824 , n18965 , n18966 , n18967 , n338828 , n18969 , n18970 , n338831 , n338832 , 
 n338833 , n338834 , n338835 , n338836 , n338837 , n338838 , n338839 , n338840 , n338841 , n338842 , 
 n338843 , n18984 , n338845 , n338846 , n338847 , n18988 , n338849 , n18990 , n338851 , n338852 , 
 n338853 , n338854 , n338855 , n338856 , n18997 , n338858 , n338859 , n338860 , n338861 , n338862 , 
 n338863 , n338864 , n19005 , n338866 , n338867 , n338868 , n19009 , n19010 , n338871 , n338872 , 
 n338873 , n338874 , n338875 , n338876 , n338877 , n338878 , n19019 , n338880 , n338881 , n338882 , 
 n338883 , n19024 , n338885 , n338886 , n19027 , n338888 , n338889 , n338890 , n338891 , n19032 , 
 n338893 , n338894 , n338895 , n19036 , n338897 , n338898 , n338899 , n338900 , n338901 , n338902 , 
 n338903 , n338904 , n338905 , n338906 , n338907 , n338908 , n338909 , n338910 , n19051 , n338912 , 
 n338913 , n19054 , n338915 , n338916 , n338917 , n338918 , n19059 , n338920 , n338921 , n19062 , 
 n338923 , n338924 , n338925 , n338926 , n19067 , n338928 , n338929 , n19070 , n338931 , n338932 , 
 n19073 , n338934 , n338935 , n19076 , n19077 , n338938 , n19079 , n338940 , n19081 , n338942 , 
 n19083 , n19084 , n338945 , n338946 , n19087 , n338948 , n338949 , n338950 , n338951 , n338952 , 
 n338953 , n338954 , n338955 , n338956 , n338957 , n19098 , n338959 , n338960 , n19101 , n338962 , 
 n19103 , n338964 , n338965 , n19106 , n338967 , n338968 , n338969 , n338970 , n19111 , n338972 , 
 n19113 , n338974 , n338975 , n19116 , n338977 , n19118 , n19119 , n338980 , n338981 , n338982 , 
 n338983 , n338984 , n338985 , n338986 , n338987 , n338988 , n338989 , n338990 , n338991 , n19132 , 
 n19133 , n338994 , n19135 , n19136 , n338997 , n338998 , n19139 , n19140 , n19141 , n339002 , 
 n339003 , n19144 , n339005 , n339006 , n339007 , n339008 , n339009 , n339010 , n19151 , n19152 , 
 n339013 , n19154 , n339015 , n19156 , n339017 , n339018 , n339019 , n339020 , n19161 , n339022 , 
 n339023 , n19164 , n339025 , n339026 , n339027 , n339028 , n19169 , n339030 , n339031 , n19172 , 
 n339033 , n339034 , n339035 , n19176 , n339037 , n19178 , n19179 , n19180 , n339041 , n339042 , 
 n19183 , n339044 , n19185 , n339046 , n339047 , n339048 , n339049 , n339050 , n19191 , n339052 , 
 n339053 , n19194 , n339055 , n19196 , n339057 , n339058 , n19199 , n339060 , n19201 , n19202 , 
 n339063 , n339064 , n19205 , n339066 , n339067 , n339068 , n19209 , n339070 , n339071 , n19212 , 
 n339073 , n339074 , n19215 , n339076 , n339077 , n339078 , n339079 , n19220 , n19221 , n339082 , 
 n19223 , n339084 , n339085 , n339086 , n339087 , n339088 , n339089 , n339090 , n339091 , n19232 , 
 n339093 , n339094 , n339095 , n339096 , n339097 , n339098 , n339099 , n339100 , n339101 , n339102 , 
 n339103 , n339104 , n339105 , n339106 , n339107 , n339108 , n19249 , n339110 , n339111 , n19252 , 
 n19253 , n339114 , n19255 , n19256 , n339117 , n339118 , n339119 , n339120 , n339121 , n339122 , 
 n339123 , n19264 , n339125 , n339126 , n19267 , n339128 , n339129 , n19270 , n339131 , n19272 , 
 n339133 , n339134 , n339135 , n19276 , n339137 , n339138 , n19279 , n339140 , n339141 , n339142 , 
 n339143 , n339144 , n19285 , n339146 , n339147 , n339148 , n339149 , n339150 , n19291 , n339152 , 
 n339153 , n339154 , n19295 , n339156 , n339157 , n339158 , n339159 , n339160 , n339161 , n339162 , 
 n339163 , n339164 , n19305 , n339166 , n339167 , n339168 , n339169 , n339170 , n339171 , n339172 , 
 n339173 , n339174 , n339175 , n19316 , n339177 , n339178 , n339179 , n339180 , n339181 , n339182 , 
 n339183 , n339184 , n339185 , n339186 , n339187 , n19328 , n339189 , n19330 , n339191 , n339192 , 
 n19333 , n339194 , n339195 , n19336 , n339197 , n339198 , n339199 , n339200 , n339201 , n19342 , 
 n339203 , n339204 , n339205 , n339206 , n339207 , n19348 , n339209 , n339210 , n339211 , n339212 , 
 n339213 , n19354 , n339215 , n19356 , n19357 , n19358 , n339219 , n339220 , n19361 , n339222 , 
 n339223 , n339224 , n19365 , n19366 , n339227 , n339228 , n19369 , n339230 , n339231 , n339232 , 
 n339233 , n339234 , n339235 , n339236 , n339237 , n339238 , n339239 , n339240 , n339241 , n339242 , 
 n19383 , n339244 , n339245 , n19386 , n339247 , n339248 , n19389 , n19390 , n339251 , n339252 , 
 n19393 , n339254 , n339255 , n339256 , n339257 , n339258 , n19399 , n339260 , n339261 , n19402 , 
 n339263 , n19404 , n19405 , n19406 , n19407 , n339268 , n339269 , n339270 , n339271 , n339272 , 
 n19413 , n339274 , n339275 , n339276 , n339277 , n339278 , n339279 , n19420 , n339281 , n339282 , 
 n339283 , n339284 , n339285 , n339286 , n339287 , n339288 , n19429 , n339290 , n339291 , n19432 , 
 n339293 , n339294 , n339295 , n19436 , n339297 , n339298 , n339299 , n19440 , n339301 , n19442 , 
 n339303 , n339304 , n19445 , n339306 , n339307 , n339308 , n339309 , n339310 , n19451 , n339312 , 
 n339313 , n339314 , n19455 , n339316 , n339317 , n19458 , n339319 , n19460 , n339321 , n339322 , 
 n19463 , n339324 , n339325 , n339326 , n339327 , n339328 , n19469 , n19470 , n339331 , n19472 , 
 n339333 , n19474 , n19475 , n339336 , n339337 , n339338 , n19479 , n339340 , n339341 , n339342 , 
 n339343 , n339344 , n339345 , n339346 , n339347 , n339348 , n19489 , n339350 , n19491 , n339352 , 
 n19493 , n339354 , n339355 , n19496 , n339357 , n339358 , n19499 , n19500 , n339361 , n339362 , 
 n19503 , n339364 , n339365 , n339366 , n339367 , n339368 , n19509 , n339370 , n19511 , n339372 , 
 n19513 , n339374 , n339375 , n19516 , n339377 , n339378 , n19519 , n339380 , n339381 , n19522 , 
 n19523 , n339384 , n339385 , n339386 , n339387 , n339388 , n339389 , n339390 , n339391 , n339392 , 
 n339393 , n339394 , n339395 , n339396 , n339397 , n339398 , n339399 , n339400 , n339401 , n339402 , 
 n19543 , n339404 , n339405 , n339406 , n339407 , n19548 , n339409 , n339410 , n19551 , n339412 , 
 n339413 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , 
 n339423 , n339424 , n19565 , n339426 , n339427 , n339428 , n339429 , n339430 , n339431 , n339432 , 
 n19573 , n339434 , n19575 , n19576 , n339437 , n19578 , n339439 , n19580 , n19581 , n339442 , 
 n339443 , n19584 , n339445 , n339446 , n339447 , n339448 , n339449 , n339450 , n339451 , n339452 , 
 n339453 , n339454 , n339455 , n339456 , n19597 , n339458 , n19599 , n339460 , n339461 , n339462 , 
 n339463 , n339464 , n19605 , n19606 , n339467 , n19608 , n339469 , n19610 , n339471 , n339472 , 
 n339473 , n19614 , n339475 , n339476 , n19617 , n339478 , n339479 , n339480 , n19621 , n339482 , 
 n339483 , n19624 , n339485 , n339486 , n339487 , n339488 , n339489 , n339490 , n339491 , n339492 , 
 n339493 , n339494 , n19635 , n339496 , n339497 , n339498 , n339499 , n339500 , n339501 , n339502 , 
 n19643 , n339504 , n339505 , n19646 , n339507 , n339508 , n339509 , n339510 , n339511 , n339512 , 
 n19653 , n19654 , n339515 , n339516 , n19657 , n339518 , n339519 , n339520 , n339521 , n339522 , 
 n339523 , n19664 , n339525 , n339526 , n19667 , n19668 , n339529 , n19670 , n339531 , n19672 , 
 n339533 , n19674 , n19675 , n339536 , n339537 , n339538 , n339539 , n19680 , n339541 , n339542 , 
 n19683 , n339544 , n339545 , n19686 , n339547 , n339548 , n339549 , n339550 , n339551 , n339552 , 
 n339553 , n339554 , n339555 , n339556 , n19697 , n339558 , n339559 , n339560 , n339561 , n339562 , 
 n339563 , n19704 , n19705 , n339566 , n19707 , n339568 , n339569 , n19710 , n339571 , n339572 , 
 n19713 , n339574 , n339575 , n19716 , n19717 , n339578 , n339579 , n339580 , n339581 , n339582 , 
 n19723 , n339584 , n339585 , n339586 , n339587 , n19728 , n339589 , n339590 , n19731 , n339592 , 
 n19733 , n339594 , n339595 , n19736 , n339597 , n19738 , n339599 , n339600 , n19741 , n339602 , 
 n19743 , n339604 , n339605 , n339606 , n339607 , n19748 , n339609 , n339610 , n19751 , n339612 , 
 n339613 , n339614 , n19755 , n339616 , n19757 , n339618 , n339619 , n339620 , n19761 , n19762 , 
 n339623 , n19764 , n339625 , n339626 , n339627 , n339628 , n339629 , n339630 , n339631 , n339632 , 
 n339633 , n339634 , n339635 , n339636 , n339637 , n339638 , n339639 , n19780 , n339641 , n19782 , 
 n339643 , n339644 , n339645 , n339646 , n19787 , n339648 , n339649 , n339650 , n339651 , n339652 , 
 n339653 , n339654 , n339655 , n19796 , n339657 , n339658 , n339659 , n339660 , n339661 , n19802 , 
 n19803 , n339664 , n339665 , n339666 , n19807 , n339668 , n339669 , n339670 , n19811 , n19812 , 
 n19813 , n339674 , n339675 , n19816 , n339677 , n339678 , n19819 , n19820 , n339681 , n19822 , 
 n19823 , n339684 , n19825 , n339686 , n339687 , n339688 , n339689 , n339690 , n339691 , n19832 , 
 n339693 , n339694 , n339695 , n339696 , n19837 , n19838 , n339699 , n339700 , n339701 , n339702 , 
 n339703 , n339704 , n339705 , n339706 , n339707 , n339708 , n339709 , n339710 , n339711 , n19852 , 
 n339713 , n339714 , n339715 , n339716 , n339717 , n339718 , n339719 , n339720 , n19861 , n339722 , 
 n19863 , n339724 , n339725 , n19866 , n339727 , n339728 , n19869 , n339730 , n339731 , n19872 , 
 n19873 , n339734 , n339735 , n339736 , n339737 , n339738 , n19879 , n19880 , n339741 , n19882 , 
 n339743 , n339744 , n19885 , n19886 , n339747 , n19888 , n339749 , n19890 , n339751 , n339752 , 
 n339753 , n339754 , n339755 , n339756 , n19897 , n339758 , n339759 , n339760 , n19901 , n339762 , 
 n339763 , n339764 , n339765 , n339766 , n339767 , n339768 , n339769 , n339770 , n19911 , n339772 , 
 n339773 , n19914 , n339775 , n339776 , n339777 , n339778 , n339779 , n19920 , n339781 , n339782 , 
 n19923 , n19924 , n339785 , n339786 , n339787 , n339788 , n339789 , n339790 , n339791 , n19932 , 
 n339793 , n339794 , n339795 , n339796 , n19937 , n19938 , n339799 , n19940 , n19941 , n339802 , 
 n19943 , n339804 , n19945 , n339806 , n339807 , n339808 , n339809 , n339810 , n339811 , n339812 , 
 n339813 , n339814 , n339815 , n339816 , n339817 , n339818 , n19959 , n339820 , n339821 , n19962 , 
 n339823 , n339824 , n339825 , n339826 , n339827 , n339828 , n339829 , n339830 , n19971 , n19972 , 
 n339833 , n19974 , n19975 , n339836 , n339837 , n339838 , n339839 , n339840 , n339841 , n19982 , 
 n339843 , n19984 , n339845 , n339846 , n339847 , n339848 , n19989 , n339850 , n339851 , n339852 , 
 n339853 , n339854 , n339855 , n339856 , n339857 , n339858 , n339859 , n20000 , n20001 , n20002 , 
 n20003 , n20004 , n339865 , n20006 , n339867 , n339868 , n339869 , n339870 , n339871 , n339872 , 
 n20013 , n339874 , n339875 , n339876 , n339877 , n339878 , n339879 , n339880 , n339881 , n339882 , 
 n339883 , n339884 , n339885 , n339886 , n339887 , n339888 , n20029 , n339890 , n339891 , n339892 , 
 n20033 , n20034 , n339895 , n339896 , n20037 , n339898 , n339899 , n339900 , n339901 , n339902 , 
 n20043 , n339904 , n339905 , n20046 , n339907 , n339908 , n20049 , n339910 , n339911 , n20052 , 
 n20053 , n339914 , n20055 , n339916 , n20057 , n339918 , n339919 , n20060 , n339921 , n20062 , 
 n339923 , n20064 , n339925 , n20066 , n339927 , n339928 , n339929 , n339930 , n339931 , n339932 , 
 n339933 , n339934 , n339935 , n339936 , n20077 , n339938 , n339939 , n20080 , n20081 , n339942 , 
 n339943 , n339944 , n339945 , n339946 , n339947 , n339948 , n339949 , n339950 , n20091 , n20092 , 
 n339953 , n339954 , n20095 , n20096 , n20097 , n339958 , n339959 , n20100 , n339961 , n339962 , 
 n339963 , n339964 , n339965 , n20106 , n339967 , n339968 , n339969 , n339970 , n20111 , n20112 , 
 n339973 , n339974 , n20115 , n20116 , n339977 , n339978 , n339979 , n20120 , n339981 , n339982 , 
 n339983 , n20124 , n339985 , n339986 , n339987 , n339988 , n339989 , n20130 , n339991 , n339992 , 
 n339993 , n20134 , n20135 , n339996 , n20137 , n339998 , n20139 , n340000 , n340001 , n340002 , 
 n340003 , n340004 , n340005 , n340006 , n340007 , n20148 , n340009 , n340010 , n340011 , n20152 , 
 n340013 , n340014 , n340015 , n340016 , n340017 , n340018 , n20159 , n20160 , n340021 , n20162 , 
 n340023 , n20164 , n20165 , n20166 , n20167 , n340028 , n20169 , n20170 , n340031 , n340032 , 
 n20173 , n340034 , n340035 , n20176 , n340037 , n20178 , n340039 , n20180 , n340041 , n340042 , 
 n20183 , n340044 , n20185 , n340046 , n340047 , n340048 , n20189 , n340050 , n340051 , n20192 , 
 n340053 , n340054 , n20195 , n340056 , n340057 , n340058 , n340059 , n340060 , n340061 , n340062 , 
 n340063 , n20204 , n340065 , n340066 , n20207 , n340068 , n340069 , n20210 , n340071 , n340072 , 
 n20213 , n340074 , n340075 , n20216 , n20217 , n340078 , n340079 , n340080 , n340081 , n340082 , 
 n20223 , n340084 , n340085 , n340086 , n340087 , n340088 , n340089 , n340090 , n20231 , n340092 , 
 n340093 , n340094 , n20235 , n340096 , n340097 , n340098 , n340099 , n340100 , n340101 , n340102 , 
 n340103 , n340104 , n340105 , n340106 , n340107 , n340108 , n340109 , n340110 , n340111 , n340112 , 
 n20253 , n340114 , n340115 , n20256 , n340117 , n20258 , n340119 , n340120 , n340121 , n340122 , 
 n340123 , n20264 , n340125 , n340126 , n340127 , n20268 , n340129 , n340130 , n20271 , n340132 , 
 n340133 , n340134 , n340135 , n20276 , n340137 , n340138 , n20279 , n20280 , n340141 , n20282 , 
 n20283 , n340144 , n340145 , n340146 , n340147 , n340148 , n20289 , n20290 , n340151 , n340152 , 
 n340153 , n340154 , n340155 , n20296 , n340157 , n340158 , n340159 , n340160 , n20301 , n340162 , 
 n340163 , n340164 , n340165 , n340166 , n340167 , n340168 , n340169 , n340170 , n340171 , n340172 , 
 n340173 , n340174 , n340175 , n340176 , n340177 , n340178 , n340179 , n20320 , n340181 , n340182 , 
 n340183 , n340184 , n20325 , n340186 , n340187 , n20328 , n340189 , n340190 , n340191 , n340192 , 
 n20333 , n20334 , n20335 , n340196 , n340197 , n20338 , n340199 , n20340 , n340201 , n340202 , 
 n340203 , n20344 , n340205 , n340206 , n340207 , n340208 , n20349 , n20350 , n340211 , n340212 , 
 n20353 , n340214 , n20355 , n340216 , n340217 , n20358 , n340219 , n340220 , n340221 , n340222 , 
 n340223 , n20364 , n20365 , n340226 , n340227 , n340228 , n340229 , n340230 , n340231 , n20372 , 
 n340233 , n340234 , n340235 , n340236 , n20377 , n340238 , n340239 , n340240 , n340241 , n340242 , 
 n340243 , n340244 , n340245 , n340246 , n340247 , n340248 , n20389 , n340250 , n340251 , n20392 , 
 n340253 , n20394 , n340255 , n340256 , n340257 , n340258 , n340259 , n340260 , n340261 , n20402 , 
 n340263 , n340264 , n340265 , n340266 , n340267 , n340268 , n340269 , n340270 , n340271 , n20412 , 
 n340273 , n340274 , n340275 , n340276 , n340277 , n340278 , n340279 , n340280 , n340281 , n340282 , 
 n20423 , n340284 , n340285 , n20426 , n340287 , n20428 , n340289 , n340290 , n20431 , n20432 , 
 n340293 , n340294 , n340295 , n340296 , n340297 , n20438 , n340299 , n20440 , n20441 , n20442 , 
 n20443 , n340304 , n340305 , n340306 , n340307 , n340308 , n340309 , n340310 , n20451 , n340312 , 
 n340313 , n20454 , n20455 , n340316 , n20457 , n340318 , n340319 , n340320 , n20461 , n340322 , 
 n20463 , n20464 , n340325 , n340326 , n340327 , n20468 , n20469 , n20470 , n340331 , n20472 , 
 n340333 , n340334 , n340335 , n340336 , n20477 , n340338 , n20479 , n340340 , n340341 , n20482 , 
 n340343 , n340344 , n20485 , n340346 , n340347 , n340348 , n340349 , n340350 , n20491 , n340352 , 
 n20493 , n340354 , n20495 , n340356 , n20497 , n340358 , n340359 , n340360 , n20501 , n340362 , 
 n340363 , n340364 , n20505 , n20506 , n20507 , n20508 , n20509 , n340370 , n340371 , n340372 , 
 n340373 , n340374 , n340375 , n340376 , n340377 , n340378 , n340379 , n340380 , n340381 , n340382 , 
 n340383 , n20524 , n340385 , n340386 , n20527 , n340388 , n340389 , n340390 , n20531 , n340392 , 
 n340393 , n340394 , n340395 , n340396 , n20537 , n340398 , n340399 , n20540 , n20541 , n20542 , 
 n20543 , n20544 , n340405 , n340406 , n340407 , n20548 , n340409 , n340410 , n340411 , n20552 , 
 n340413 , n340414 , n340415 , n340416 , n340417 , n340418 , n20559 , n340420 , n340421 , n20562 , 
 n340423 , n340424 , n20565 , n20566 , n340427 , n340428 , n340429 , n340430 , n340431 , n20572 , 
 n340433 , n340434 , n20575 , n340436 , n20577 , n340438 , n340439 , n20580 , n340441 , n340442 , 
 n340443 , n340444 , n20585 , n340446 , n20587 , n20588 , n340449 , n340450 , n20591 , n340452 , 
 n340453 , n340454 , n20595 , n20596 , n20597 , n340458 , n340459 , n340460 , n20601 , n340462 , 
 n340463 , n340464 , n340465 , n340466 , n20607 , n340468 , n340469 , n340470 , n20611 , n340472 , 
 n340473 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n340481 , n340482 , 
 n340483 , n340484 , n20625 , n340486 , n20627 , n340488 , n340489 , n340490 , n340491 , n340492 , 
 n340493 , n340494 , n340495 , n340496 , n340497 , n340498 , n340499 , n20640 , n340501 , n340502 , 
 n20643 , n340504 , n340505 , n340506 , n340507 , n340508 , n20649 , n340510 , n340511 , n340512 , 
 n20653 , n340514 , n340515 , n20656 , n340517 , n340518 , n340519 , n340520 , n340521 , n20662 , 
 n340523 , n340524 , n20665 , n340526 , n340527 , n20668 , n20669 , n340530 , n20671 , n340532 , 
 n20673 , n20674 , n340535 , n340536 , n340537 , n340538 , n340539 , n340540 , n340541 , n340542 , 
 n340543 , n340544 , n340545 , n340546 , n340547 , n20688 , n340549 , n340550 , n340551 , n340552 , 
 n340553 , n20694 , n340555 , n340556 , n20697 , n20698 , n20699 , n340560 , n20701 , n20702 , 
 n340563 , n20704 , n340565 , n340566 , n340567 , n340568 , n340569 , n340570 , n340571 , n20712 , 
 n340573 , n340574 , n340575 , n20716 , n340577 , n340578 , n20719 , n340580 , n340581 , n20722 , 
 n340583 , n340584 , n20725 , n340586 , n340587 , n340588 , n340589 , n340590 , n340591 , n340592 , 
 n340593 , n340594 , n340595 , n340596 , n340597 , n340598 , n340599 , n340600 , n20738 , n340602 , 
 n340603 , n340604 , n340605 , n20743 , n20744 , n340608 , n340609 , n340610 , n340611 , n20749 , 
 n340613 , n340614 , n20752 , n340616 , n20754 , n20755 , n340619 , n340620 , n340621 , n340622 , 
 n340623 , n340624 , n20756 , n340626 , n340627 , n340628 , n340629 , n20761 , n340631 , n340632 , 
 n340633 , n340634 , n340635 , n340636 , n340637 , n340638 , n340639 , n340640 , n340641 , n20766 , 
 n340643 , n20768 , n340645 , n340646 , n340647 , n340648 , n340649 , n340650 , n340651 , n340652 , 
 n340653 , n340654 , n340655 , n340656 , n340657 , n340658 , n340659 , n340660 , n340661 , n340662 , 
 n340663 , n340664 , n340665 , n340666 , n340667 , n340668 , n340669 , n340670 , n20785 , n340672 , 
 n340673 , n340674 , n340675 , n340676 , n340677 , n20792 , n20793 , n340680 , n20795 , n340682 , 
 n340683 , n340684 , n20799 , n340686 , n340687 , n340688 , n340689 , n340690 , n340691 , n340692 , 
 n20807 , n340694 , n20809 , n340696 , n20811 , n340698 , n340699 , n20814 , n340701 , n340702 , 
 n340703 , n340704 , n340705 , n340706 , n340707 , n20822 , n340709 , n340710 , n340711 , n340712 , 
 n340713 , n340714 , n340715 , n340716 , n340717 , n20832 , n340719 , n20833 , n340721 , n340722 , 
 n340723 , n340724 , n340725 , n340726 , n340727 , n340728 , n340729 , n340730 , n340731 , n20844 , 
 n340733 , n20846 , n340735 , n340736 , n20849 , n340738 , n340739 , n340740 , n340741 , n340742 , 
 n340743 , n340744 , n340745 , n20858 , n340747 , n20860 , n20861 , n340750 , n20863 , n340752 , 
 n340753 , n340754 , n340755 , n340756 , n340757 , n340758 , n20871 , n340760 , n340761 , n340762 , 
 n340763 , n20876 , n20877 , n340766 , n340767 , n340768 , n340769 , n340770 , n340771 , n340772 , 
 n340773 , n340774 , n340775 , n340776 , n340777 , n340778 , n340779 , n340780 , n340781 , n20894 , 
 n20895 , n340784 , n340785 , n20898 , n340787 , n20900 , n340789 , n340790 , n340791 , n20904 , 
 n340793 , n340794 , n340795 , n20908 , n340797 , n340798 , n340799 , n340800 , n340801 , n20914 , 
 n340803 , n340804 , n20917 , n340806 , n340807 , n340808 , n340809 , n340810 , n340811 , n20924 , 
 n340813 , n20926 , n340815 , n340816 , n340817 , n340818 , n340819 , n340820 , n340821 , n340822 , 
 n20935 , n340824 , n340825 , n340826 , n340827 , n340828 , n340829 , n340830 , n340831 , n20944 , 
 n340833 , n340834 , n340835 , n20948 , n340837 , n340838 , n340839 , n340840 , n340841 , n340842 , 
 n340843 , n20956 , n20957 , n340846 , n340847 , n340848 , n20961 , n340850 , n340851 , n20964 , 
 n340853 , n20966 , n20967 , n340856 , n20969 , n340858 , n340859 , n340860 , n340861 , n20974 , 
 n340863 , n20976 , n340865 , n340866 , n340867 , n340868 , n20981 , n20982 , n340871 , n340872 , 
 n340873 , n20986 , n340875 , n20988 , n340877 , n340878 , n340879 , n340880 , n20993 , n340882 , 
 n340883 , n340884 , n20997 , n340886 , n340887 , n21000 , n340889 , n340890 , n340891 , n340892 , 
 n340893 , n340894 , n340895 , n340896 , n340897 , n21010 , n21011 , n21012 , n340901 , n340902 , 
 n340903 , n340904 , n340905 , n340906 , n21019 , n21020 , n340909 , n340910 , n340911 , n340912 , 
 n340913 , n340914 , n340915 , n21028 , n340917 , n340918 , n21031 , n21032 , n21033 , n340922 , 
 n21035 , n21036 , n340925 , n340926 , n340927 , n21040 , n340929 , n340930 , n340931 , n340932 , 
 n21045 , n340934 , n340935 , n340936 , n340937 , n340938 , n340939 , n21052 , n340941 , n340942 , 
 n340943 , n340944 , n340945 , n340946 , n340947 , n340948 , n340949 , n340950 , n21063 , n21064 , 
 n340953 , n21066 , n340955 , n340956 , n21069 , n21070 , n21071 , n340960 , n340961 , n21074 , 
 n21075 , n340964 , n340965 , n340966 , n21079 , n340968 , n340969 , n340970 , n340971 , n340972 , 
 n340973 , n21086 , n340975 , n340976 , n21089 , n340978 , n21091 , n340980 , n340981 , n21094 , 
 n340983 , n21096 , n340985 , n340986 , n340987 , n21100 , n21101 , n340990 , n340991 , n340992 , 
 n340993 , n340994 , n340995 , n21108 , n340997 , n340998 , n340999 , n341000 , n341001 , n21114 , 
 n341003 , n21116 , n341005 , n341006 , n341007 , n341008 , n341009 , n341010 , n341011 , n341012 , 
 n341013 , n341014 , n21127 , n341016 , n341017 , n21130 , n341019 , n341020 , n341021 , n21134 , 
 n341023 , n341024 , n21137 , n341026 , n341027 , n341028 , n341029 , n341030 , n341031 , n341032 , 
 n21145 , n341034 , n341035 , n341036 , n21149 , n341038 , n341039 , n21152 , n341041 , n341042 , 
 n341043 , n21156 , n341045 , n21158 , n21159 , n341048 , n341049 , n341050 , n341051 , n21164 , 
 n341053 , n341054 , n21167 , n341056 , n341057 , n341058 , n341059 , n341060 , n341061 , n21174 , 
 n341063 , n341064 , n21177 , n21178 , n341067 , n341068 , n341069 , n341070 , n341071 , n341072 , 
 n341073 , n21186 , n341075 , n341076 , n21189 , n341078 , n341079 , n341080 , n341081 , n341082 , 
 n341083 , n341084 , n341085 , n341086 , n341087 , n341088 , n341089 , n341090 , n341091 , n341092 , 
 n341093 , n21206 , n341095 , n341096 , n341097 , n341098 , n341099 , n341100 , n21213 , n21214 , 
 n341103 , n341104 , n21217 , n341106 , n341107 , n341108 , n341109 , n341110 , n341111 , n21224 , 
 n341113 , n341114 , n341115 , n341116 , n341117 , n341118 , n341119 , n341120 , n341121 , n341122 , 
 n341123 , n341124 , n341125 , n341126 , n341127 , n341128 , n341129 , n341130 , n341131 , n341132 , 
 n341133 , n341134 , n21245 , n341136 , n341137 , n341138 , n341139 , n341140 , n21251 , n341142 , 
 n341143 , n341144 , n341145 , n341146 , n341147 , n341148 , n341149 , n341150 , n21261 , n341152 , 
 n341153 , n21264 , n341155 , n341156 , n21267 , n341158 , n341159 , n341160 , n341161 , n341162 , 
 n21272 , n341164 , n341165 , n21275 , n341167 , n341168 , n341169 , n21279 , n341171 , n341172 , 
 n341173 , n341174 , n341175 , n341176 , n341177 , n341178 , n341179 , n341180 , n21290 , n341182 , 
 n341183 , n341184 , n341185 , n341186 , n21296 , n341188 , n21298 , n341190 , n341191 , n21301 , 
 n21302 , n21303 , n341195 , n341196 , n21306 , n21307 , n21308 , n341200 , n341201 , n21311 , 
 n341203 , n21313 , n341205 , n341206 , n21316 , n21317 , n341209 , n21319 , n341211 , n341212 , 
 n341213 , n341214 , n21324 , n341216 , n341217 , n21327 , n341219 , n341220 , n21330 , n21331 , 
 n341223 , n21333 , n341225 , n21335 , n341227 , n21337 , n341229 , n341230 , n21340 , n21341 , 
 n21342 , n341234 , n341235 , n341236 , n341237 , n21347 , n341239 , n341240 , n21350 , n341242 , 
 n21352 , n341244 , n341245 , n341246 , n21356 , n21357 , n341249 , n341250 , n21360 , n341252 , 
 n341253 , n21363 , n21364 , n21365 , n21366 , n341258 , n341259 , n341260 , n341261 , n341262 , 
 n341263 , n341264 , n341265 , n21375 , n341267 , n341268 , n341269 , n341270 , n21380 , n21381 , 
 n341273 , n341274 , n341275 , n341276 , n341277 , n341278 , n21388 , n341280 , n341281 , n341282 , 
 n341283 , n341284 , n341285 , n341286 , n341287 , n341288 , n341289 , n341290 , n341291 , n21399 , 
 n341293 , n21401 , n21402 , n341296 , n21404 , n21405 , n21406 , n341300 , n341301 , n341302 , 
 n341303 , n341304 , n341305 , n341306 , n341307 , n341308 , n341309 , n341310 , n341311 , n341312 , 
 n341313 , n341314 , n21422 , n341316 , n341317 , n341318 , n341319 , n341320 , n21427 , n341322 , 
 n21429 , n341324 , n341325 , n21430 , n341327 , n341328 , n341329 , n21431 , n341331 , n21433 , 
 n21434 , n341334 , n21436 , n341336 , n341337 , n341338 , n21440 , n341340 , n341341 , n341342 , 
 n21444 , n341344 , n341345 , n21447 , n341347 , n341348 , n21448 , n341350 , n341351 , n341352 , 
 n341353 , n341354 , n341355 , n341356 , n341357 , n341358 , n341359 , n341360 , n341361 , n341362 , 
 n341363 , n341364 , n341365 , n341366 , n341367 , n341368 , n341369 , n21466 , n341371 , n341372 , 
 n341373 , n341374 , n341375 , n341376 , n341377 , n341378 , n341379 , n341380 , n341381 , n21478 , 
 n341383 , n341384 , n21481 , n21482 , n21483 , n21484 , n341389 , n341390 , n341391 , n341392 , 
 n21489 , n341394 , n341395 , n21492 , n21493 , n341398 , n21495 , n341400 , n341401 , n341402 , 
 n341403 , n341404 , n341405 , n341406 , n341407 , n21503 , n341409 , n341410 , n341411 , n341412 , 
 n341413 , n341414 , n341415 , n341416 , n341417 , n341418 , n341419 , n341420 , n21515 , n341422 , 
 n21517 , n341424 , n341425 , n21520 , n341427 , n341428 , n21523 , n341430 , n341431 , n341432 , 
 n341433 , n341434 , n341435 , n21530 , n341437 , n341438 , n341439 , n341440 , n341441 , n341442 , 
 n341443 , n341444 , n341445 , n341446 , n341447 , n341448 , n21543 , n341450 , n21545 , n21546 , 
 n21547 , n341454 , n341455 , n341456 , n341457 , n341458 , n341459 , n341460 , n341461 , n341462 , 
 n341463 , n341464 , n341465 , n21560 , n341467 , n341468 , n341469 , n341470 , n341471 , n21566 , 
 n341473 , n341474 , n341475 , n21570 , n341477 , n21572 , n21573 , n21574 , n341481 , n21576 , 
 n341483 , n341484 , n341485 , n341486 , n341487 , n341488 , n341489 , n341490 , n341491 , n21586 , 
 n341493 , n341494 , n341495 , n21590 , n21591 , n341498 , n341499 , n21594 , n341501 , n341502 , 
 n21597 , n341504 , n341505 , n341506 , n21601 , n341508 , n341509 , n341510 , n21605 , n341512 , 
 n341513 , n341514 , n341515 , n21610 , n21611 , n341518 , n21613 , n341520 , n21615 , n341522 , 
 n341523 , n341524 , n21619 , n21620 , n341527 , n341528 , n21623 , n21624 , n21625 , n341532 , 
 n341533 , n21628 , n21629 , n21630 , n341537 , n341538 , n21633 , n341540 , n341541 , n21636 , 
 n21637 , n341544 , n21639 , n21640 , n341547 , n341548 , n341549 , n341550 , n341551 , n341552 , 
 n341553 , n341554 , n21649 , n341556 , n341557 , n341558 , n341559 , n341560 , n341561 , n341562 , 
 n341563 , n21658 , n341565 , n341566 , n21661 , n341568 , n341569 , n341570 , n21665 , n341572 , 
 n341573 , n341574 , n341575 , n21670 , n341577 , n21672 , n341579 , n341580 , n341581 , n341582 , 
 n341583 , n341584 , n341585 , n341586 , n21681 , n341588 , n341589 , n21684 , n341591 , n341592 , 
 n341593 , n21688 , n341595 , n341596 , n21691 , n341598 , n341599 , n341600 , n341601 , n341602 , 
 n341603 , n341604 , n341605 , n341606 , n341607 , n21702 , n21703 , n341610 , n341611 , n21706 , 
 n341613 , n341614 , n21709 , n341616 , n341617 , n21712 , n341619 , n341620 , n341621 , n21716 , 
 n341623 , n21718 , n341625 , n21720 , n21721 , n21722 , n21723 , n341630 , n21725 , n341632 , 
 n341633 , n341634 , n341635 , n21730 , n341637 , n341638 , n341639 , n341640 , n341641 , n21736 , 
 n21737 , n341644 , n21739 , n341646 , n341647 , n341648 , n21743 , n21744 , n341651 , n341652 , 
 n341653 , n341654 , n341655 , n341656 , n341657 , n21752 , n341659 , n341660 , n21755 , n341662 , 
 n341663 , n341664 , n341665 , n341666 , n21761 , n341668 , n341669 , n21764 , n21765 , n341672 , 
 n341673 , n341674 , n341675 , n21770 , n341677 , n341678 , n341679 , n21774 , n21775 , n21776 , 
 n341683 , n341684 , n341685 , n21780 , n341687 , n341688 , n341689 , n341690 , n21785 , n341692 , 
 n341693 , n341694 , n21789 , n341696 , n341697 , n341698 , n341699 , n341700 , n341701 , n341702 , 
 n341703 , n21798 , n341705 , n21800 , n341707 , n341708 , n341709 , n341710 , n341711 , n341712 , 
 n341713 , n341714 , n341715 , n341716 , n341717 , n21812 , n341719 , n341720 , n341721 , n341722 , 
 n341723 , n21818 , n341725 , n341726 , n341727 , n21822 , n341729 , n341730 , n21825 , n341732 , 
 n21827 , n21828 , n21829 , n341736 , n21831 , n21832 , n21833 , n21834 , n341741 , n341742 , 
 n21837 , n341744 , n341745 , n21840 , n21841 , n341748 , n341749 , n21844 , n341751 , n21846 , 
 n21847 , n341754 , n21849 , n341756 , n21851 , n21852 , n341759 , n341760 , n21855 , n341762 , 
 n341763 , n21858 , n341765 , n341766 , n341767 , n341768 , n341769 , n341770 , n21865 , n341772 , 
 n21867 , n341774 , n21869 , n341776 , n341777 , n21872 , n341779 , n341780 , n341781 , n341782 , 
 n341783 , n21878 , n21879 , n21880 , n341787 , n341788 , n341789 , n341790 , n341791 , n341792 , 
 n341793 , n341794 , n341795 , n341796 , n341797 , n341798 , n21893 , n21894 , n341801 , n21896 , 
 n21897 , n341804 , n341805 , n341806 , n341807 , n21902 , n341809 , n341810 , n341811 , n21906 , 
 n341813 , n341814 , n341815 , n21910 , n341817 , n341818 , n21913 , n341820 , n341821 , n341822 , 
 n341823 , n341824 , n341825 , n21920 , n341827 , n341828 , n341829 , n341830 , n341831 , n21926 , 
 n21927 , n21928 , n341835 , n341836 , n21931 , n21932 , n341839 , n21934 , n341841 , n341842 , 
 n341843 , n21938 , n341845 , n21940 , n341847 , n21942 , n21943 , n21944 , n341851 , n341852 , 
 n21947 , n21948 , n21949 , n341856 , n341857 , n21952 , n21953 , n341860 , n341861 , n341862 , 
 n21957 , n21958 , n21959 , n341866 , n341867 , n21962 , n341869 , n21964 , n341871 , n21966 , 
 n21967 , n21968 , n341875 , n21970 , n341877 , n21972 , n341879 , n341880 , n341881 , n341882 , 
 n341883 , n341884 , n341885 , n341886 , n341887 , n21982 , n341889 , n341890 , n341891 , n341892 , 
 n341893 , n341894 , n341895 , n21990 , n341897 , n341898 , n341899 , n341900 , n341901 , n21996 , 
 n341903 , n341904 , n21999 , n341906 , n341907 , n22002 , n341909 , n22004 , n341911 , n341912 , 
 n341913 , n341914 , n341915 , n341916 , n341917 , n341918 , n22011 , n341920 , n22013 , n22014 , 
 n22015 , n22016 , n22017 , n341926 , n341927 , n341928 , n341929 , n341930 , n341931 , n22024 , 
 n341933 , n341934 , n341935 , n341936 , n341937 , n341938 , n341939 , n22031 , n341941 , n22033 , 
 n22034 , n341944 , n22036 , n341946 , n341947 , n22037 , n341949 , n341950 , n341951 , n341952 , 
 n341953 , n22040 , n341955 , n341956 , n341957 , n22044 , n341959 , n341960 , n341961 , n341962 , 
 n341963 , n341964 , n341965 , n341966 , n341967 , n22054 , n341969 , n22056 , n341971 , n341972 , 
 n341973 , n341974 , n341975 , n341976 , n341977 , n341978 , n341979 , n341980 , n341981 , n22063 , 
 n341983 , n341984 , n341985 , n341986 , n341987 , n341988 , n22070 , n341990 , n341991 , n22073 , 
 n341993 , n22075 , n341995 , n22077 , n22078 , n341998 , n341999 , n22081 , n342001 , n342002 , 
 n342003 , n342004 , n342005 , n342006 , n342007 , n342008 , n342009 , n342010 , n342011 , n342012 , 
 n342013 , n342014 , n342015 , n22097 , n342017 , n342018 , n342019 , n342020 , n342021 , n342022 , 
 n342023 , n342024 , n342025 , n22107 , n22108 , n22109 , n342029 , n342030 , n342031 , n22112 , 
 n342033 , n342034 , n342035 , n342036 , n342037 , n342038 , n342039 , n22119 , n22120 , n342042 , 
 n342043 , n22123 , n342045 , n22125 , n342047 , n342048 , n22128 , n342050 , n342051 , n342052 , 
 n22132 , n342054 , n342055 , n342056 , n342057 , n342058 , n342059 , n342060 , n342061 , n342062 , 
 n342063 , n22143 , n342065 , n342066 , n342067 , n342068 , n342069 , n22149 , n22150 , n342072 , 
 n342073 , n342074 , n342075 , n342076 , n342077 , n342078 , n342079 , n342080 , n342081 , n342082 , 
 n22162 , n342084 , n342085 , n342086 , n342087 , n22167 , n342089 , n22169 , n342091 , n342092 , 
 n342093 , n342094 , n22174 , n342096 , n342097 , n22177 , n342099 , n342100 , n22180 , n342102 , 
 n342103 , n342104 , n342105 , n342106 , n22186 , n342108 , n342109 , n22189 , n342111 , n342112 , 
 n342113 , n22193 , n342115 , n342116 , n22196 , n342118 , n342119 , n22199 , n342121 , n22201 , 
 n22202 , n342124 , n342125 , n22205 , n342127 , n22207 , n342129 , n342130 , n342131 , n22211 , 
 n342133 , n342134 , n342135 , n342136 , n342137 , n342138 , n22218 , n342140 , n342141 , n342142 , 
 n22222 , n22223 , n342145 , n342146 , n342147 , n342148 , n342149 , n22229 , n342151 , n342152 , 
 n342153 , n342154 , n342155 , n342156 , n342157 , n342158 , n342159 , n22239 , n342161 , n342162 , 
 n22242 , n342164 , n342165 , n22245 , n342167 , n342168 , n342169 , n342170 , n342171 , n342172 , 
 n342173 , n342174 , n342175 , n342176 , n342177 , n22257 , n342179 , n342180 , n342181 , n342182 , 
 n22262 , n22263 , n342185 , n342186 , n22266 , n342188 , n342189 , n22269 , n342191 , n342192 , 
 n342193 , n22273 , n342195 , n342196 , n342197 , n342198 , n342199 , n342200 , n22280 , n342202 , 
 n342203 , n22283 , n342205 , n342206 , n342207 , n342208 , n342209 , n342210 , n342211 , n22291 , 
 n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n342222 , 
 n342223 , n342224 , n342225 , n342226 , n22306 , n342228 , n342229 , n22309 , n342231 , n22311 , 
 n342233 , n22313 , n342235 , n22315 , n342237 , n342238 , n22318 , n342240 , n342241 , n342242 , 
 n22322 , n342244 , n342245 , n22325 , n22326 , n342248 , n22328 , n342250 , n342251 , n342252 , 
 n22332 , n342254 , n342255 , n342256 , n342257 , n342258 , n22338 , n342260 , n342261 , n22341 , 
 n342263 , n22343 , n342265 , n342266 , n22346 , n22347 , n22348 , n342270 , n342271 , n22351 , 
 n342273 , n342274 , n342275 , n342276 , n22356 , n22357 , n22358 , n342280 , n22360 , n22361 , 
 n22362 , n22363 , n342285 , n342286 , n22366 , n22367 , n22368 , n22369 , n342291 , n342292 , 
 n22372 , n342294 , n342295 , n342296 , n22376 , n342298 , n342299 , n22379 , n342301 , n342302 , 
 n342303 , n342304 , n22384 , n342306 , n22386 , n342308 , n342309 , n22389 , n342311 , n342312 , 
 n342313 , n342314 , n342315 , n342316 , n342317 , n342318 , n22398 , n342320 , n22400 , n22401 , 
 n22402 , n22403 , n22404 , n22405 , n342327 , n342328 , n22408 , n342330 , n342331 , n22411 , 
 n342333 , n342334 , n342335 , n342336 , n342337 , n342338 , n342339 , n342340 , n22420 , n342342 , 
 n22422 , n22423 , n342345 , n342346 , n342347 , n342348 , n342349 , n22429 , n342351 , n342352 , 
 n342353 , n22433 , n342355 , n342356 , n22436 , n342358 , n342359 , n22439 , n342361 , n342362 , 
 n22442 , n22443 , n342365 , n342366 , n342367 , n342368 , n342369 , n342370 , n342371 , n22449 , 
 n22450 , n22451 , n342375 , n342376 , n342377 , n22455 , n22456 , n22457 , n22458 , n342382 , 
 n342383 , n342384 , n342385 , n342386 , n342387 , n342388 , n342389 , n342390 , n342391 , n342392 , 
 n342393 , n342394 , n342395 , n342396 , n22465 , n342398 , n342399 , n342400 , n22469 , n342402 , 
 n342403 , n22472 , n342405 , n342406 , n22473 , n342408 , n342409 , n342410 , n22474 , n342412 , 
 n22476 , n342414 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n342422 , 
 n22486 , n342424 , n342425 , n342426 , n22490 , n342428 , n22492 , n342430 , n342431 , n342432 , 
 n342433 , n342434 , n342435 , n342436 , n342437 , n342438 , n342439 , n342440 , n342441 , n342442 , 
 n342443 , n22499 , n342445 , n342446 , n342447 , n22503 , n342449 , n342450 , n22506 , n342452 , 
 n342453 , n342454 , n342455 , n342456 , n342457 , n22513 , n22514 , n342460 , n342461 , n22517 , 
 n342463 , n342464 , n342465 , n342466 , n342467 , n342468 , n342469 , n22525 , n342471 , n342472 , 
 n22528 , n22529 , n342475 , n342476 , n342477 , n22533 , n342479 , n22535 , n342481 , n342482 , 
 n22538 , n342484 , n22540 , n342486 , n342487 , n342488 , n22544 , n22545 , n342491 , n22547 , 
 n22548 , n342494 , n342495 , n342496 , n342497 , n22552 , n342499 , n342500 , n22555 , n342502 , 
 n22556 , n342504 , n342505 , n22559 , n342507 , n22560 , n342509 , n342510 , n342511 , n342512 , 
 n342513 , n342514 , n22567 , n342516 , n342517 , n342518 , n342519 , n342520 , n22573 , n22574 , 
 n22575 , n22576 , n342525 , n342526 , n342527 , n342528 , n342529 , n22582 , n342531 , n342532 , 
 n22585 , n342534 , n342535 , n22588 , n342537 , n342538 , n342539 , n342540 , n22593 , n342542 , 
 n22595 , n342544 , n342545 , n342546 , n22599 , n22600 , n342549 , n342550 , n22603 , n22604 , 
 n22605 , n342554 , n342555 , n22608 , n342557 , n22610 , n342559 , n342560 , n22613 , n22614 , 
 n22615 , n342564 , n22617 , n22618 , n22619 , n342568 , n22621 , n342570 , n342571 , n22624 , 
 n342573 , n22626 , n22627 , n342576 , n342577 , n342578 , n342579 , n22632 , n22633 , n342582 , 
 n22635 , n342584 , n22637 , n342586 , n342587 , n22640 , n342589 , n342590 , n342591 , n342592 , 
 n342593 , n342594 , n22647 , n22648 , n22649 , n22650 , n342599 , n342600 , n342601 , n22654 , 
 n342603 , n22656 , n342605 , n22658 , n342607 , n342608 , n342609 , n22662 , n342611 , n342612 , 
 n22665 , n342614 , n22667 , n342616 , n342617 , n342618 , n342619 , n22672 , n342621 , n342622 , 
 n22675 , n22676 , n342625 , n342626 , n342627 , n342628 , n342629 , n342630 , n22683 , n342632 , 
 n342633 , n22686 , n342635 , n342636 , n22689 , n342638 , n342639 , n22692 , n342641 , n342642 , 
 n22695 , n342644 , n342645 , n22698 , n342647 , n22700 , n342649 , n342650 , n22703 , n22704 , 
 n342653 , n342654 , n22707 , n342656 , n342657 , n22710 , n342659 , n342660 , n342661 , n342662 , 
 n342663 , n342664 , n22717 , n342666 , n342667 , n342668 , n342669 , n22722 , n342671 , n342672 , 
 n342673 , n22726 , n342675 , n22728 , n342677 , n22730 , n342679 , n342680 , n342681 , n342682 , 
 n342683 , n342684 , n342685 , n342686 , n342687 , n342688 , n342689 , n22742 , n22743 , n342692 , 
 n22745 , n22746 , n22747 , n22748 , n342697 , n342698 , n342699 , n342700 , n342701 , n22754 , 
 n342703 , n22756 , n342705 , n342706 , n22759 , n342708 , n342709 , n22762 , n342711 , n342712 , 
 n22765 , n342714 , n342715 , n22768 , n22769 , n342718 , n342719 , n22772 , n342721 , n22774 , 
 n342723 , n342724 , n22777 , n342726 , n342727 , n22780 , n342729 , n342730 , n342731 , n342732 , 
 n342733 , n342734 , n342735 , n342736 , n342737 , n22790 , n342739 , n342740 , n342741 , n342742 , 
 n342743 , n22796 , n342745 , n342746 , n342747 , n22800 , n342749 , n22802 , n342751 , n342752 , 
 n22805 , n342754 , n22807 , n342756 , n22809 , n22810 , n342759 , n342760 , n342761 , n342762 , 
 n342763 , n22816 , n342765 , n342766 , n342767 , n342768 , n342769 , n22822 , n342771 , n342772 , 
 n342773 , n342774 , n342775 , n22828 , n342777 , n342778 , n342779 , n342780 , n342781 , n342782 , 
 n342783 , n342784 , n342785 , n342786 , n342787 , n342788 , n342789 , n342790 , n342791 , n342792 , 
 n342793 , n342794 , n342795 , n342796 , n342797 , n342798 , n342799 , n342800 , n342801 , n22854 , 
 n342803 , n342804 , n342805 , n22858 , n342807 , n22860 , n342809 , n342810 , n22863 , n342812 , 
 n342813 , n342814 , n342815 , n342816 , n22869 , n342818 , n22871 , n342820 , n342821 , n22874 , 
 n342823 , n342824 , n342825 , n342826 , n22879 , n342828 , n342829 , n342830 , n342831 , n22884 , 
 n22885 , n22886 , n342835 , n342836 , n342837 , n22890 , n22891 , n342840 , n22893 , n342842 , 
 n22895 , n22896 , n342845 , n342846 , n22899 , n342848 , n342849 , n22902 , n342851 , n342852 , 
 n342853 , n342854 , n342855 , n342856 , n22909 , n342858 , n342859 , n342860 , n342861 , n342862 , 
 n342863 , n342864 , n342865 , n22916 , n342867 , n342868 , n22919 , n342870 , n342871 , n342872 , 
 n342873 , n342874 , n342875 , n342876 , n342877 , n342878 , n342879 , n22930 , n342881 , n342882 , 
 n342883 , n22934 , n342885 , n342886 , n342887 , n342888 , n342889 , n342890 , n342891 , n22941 , 
 n342893 , n22943 , n22944 , n342896 , n22946 , n22947 , n22948 , n22949 , n342901 , n342902 , 
 n22952 , n342904 , n22954 , n22955 , n22956 , n342908 , n342909 , n22959 , n22960 , n22961 , 
 n342913 , n342914 , n342915 , n342916 , n22966 , n342918 , n342919 , n22969 , n342921 , n342922 , 
 n342923 , n342924 , n342925 , n342926 , n22976 , n342928 , n342929 , n342930 , n342931 , n342932 , 
 n342933 , n342934 , n342935 , n342936 , n342937 , n22985 , n342939 , n342940 , n342941 , n342942 , 
 n342943 , n342944 , n342945 , n342946 , n342947 , n22995 , n22996 , n22997 , n342951 , n22999 , 
 n23000 , n342954 , n342955 , n23003 , n23004 , n342958 , n23006 , n342960 , n23008 , n23009 , 
 n342963 , n342964 , n342965 , n342966 , n342967 , n342968 , n342969 , n342970 , n342971 , n342972 , 
 n23013 , n342974 , n23015 , n342976 , n342977 , n23016 , n342979 , n342980 , n342981 , n342982 , 
 n342983 , n23019 , n342985 , n342986 , n23022 , n342988 , n342989 , n342990 , n342991 , n342992 , 
 n342993 , n342994 , n23027 , n342996 , n342997 , n23030 , n342999 , n23032 , n343001 , n23034 , 
 n343003 , n23036 , n23037 , n343006 , n343007 , n343008 , n23041 , n343010 , n343011 , n343012 , 
 n343013 , n343014 , n343015 , n343016 , n343017 , n343018 , n343019 , n343020 , n343021 , n343022 , 
 n343023 , n343024 , n23057 , n23058 , n23059 , n343028 , n343029 , n23062 , n343031 , n343032 , 
 n343033 , n343034 , n343035 , n343036 , n23069 , n343038 , n343039 , n343040 , n23073 , n343042 , 
 n343043 , n343044 , n343045 , n23078 , n343047 , n23080 , n23081 , n343050 , n343051 , n23084 , 
 n343053 , n343054 , n343055 , n343056 , n343057 , n23090 , n343059 , n23091 , n343061 , n343062 , 
 n23094 , n343064 , n343065 , n343066 , n343067 , n23098 , n23099 , n343070 , n343071 , n23102 , 
 n343073 , n23104 , n343075 , n23106 , n23107 , n23108 , n343079 , n343080 , n23111 , n343082 , 
 n343083 , n343084 , n343085 , n343086 , n343087 , n343088 , n343089 , n343090 , n343091 , n23122 , 
 n343093 , n343094 , n23125 , n343096 , n343097 , n343098 , n23129 , n343100 , n343101 , n343102 , 
 n23133 , n23134 , n343105 , n343106 , n343107 , n23138 , n343109 , n343110 , n23141 , n343112 , 
 n343113 , n343114 , n343115 , n343116 , n343117 , n343118 , n343119 , n343120 , n343121 , n343122 , 
 n343123 , n343124 , n343125 , n23156 , n343127 , n343128 , n343129 , n343130 , n343131 , n343132 , 
 n343133 , n343134 , n343135 , n23166 , n343137 , n343138 , n343139 , n343140 , n343141 , n23170 , 
 n343143 , n343144 , n343145 , n343146 , n343147 , n343148 , n343149 , n343150 , n343151 , n343152 , 
 n343153 , n343154 , n343155 , n23184 , n343157 , n343158 , n23187 , n343160 , n343161 , n23190 , 
 n343163 , n343164 , n23193 , n343166 , n343167 , n343168 , n343169 , n343170 , n343171 , n343172 , 
 n343173 , n343174 , n23203 , n343176 , n23205 , n23206 , n343179 , n343180 , n23208 , n343182 , 
 n343183 , n343184 , n343185 , n343186 , n343187 , n23213 , n343189 , n343190 , n23215 , n343192 , 
 n343193 , n343194 , n343195 , n343196 , n343197 , n343198 , n343199 , n23219 , n343201 , n343202 , 
 n23222 , n343204 , n343205 , n343206 , n23226 , n343208 , n343209 , n343210 , n23230 , n23231 , 
 n23232 , n343214 , n23234 , n23235 , n343217 , n343218 , n343219 , n343220 , n23240 , n343222 , 
 n343223 , n343224 , n23244 , n23245 , n343227 , n343228 , n343229 , n343230 , n343231 , n343232 , 
 n343233 , n343234 , n343235 , n343236 , n343237 , n343238 , n343239 , n343240 , n343241 , n343242 , 
 n343243 , n343244 , n23264 , n343246 , n343247 , n343248 , n23268 , n23269 , n343251 , n343252 , 
 n343253 , n23271 , n23272 , n343256 , n343257 , n343258 , n343259 , n23277 , n343261 , n23278 , 
 n343263 , n343264 , n343265 , n343266 , n23282 , n343268 , n343269 , n343270 , n343271 , n343272 , 
 n23288 , n343274 , n343275 , n23291 , n343277 , n343278 , n343279 , n343280 , n343281 , n23297 , 
 n343283 , n343284 , n343285 , n23301 , n343287 , n343288 , n343289 , n343290 , n343291 , n23307 , 
 n343293 , n343294 , n343295 , n343296 , n343297 , n343298 , n343299 , n343300 , n343301 , n343302 , 
 n343303 , n343304 , n343305 , n343306 , n343307 , n343308 , n23322 , n343310 , n343311 , n23325 , 
 n343313 , n343314 , n343315 , n343316 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , 
 n23336 , n23337 , n23338 , n23339 , n23340 , n343328 , n343329 , n343330 , n343331 , n23345 , 
 n23346 , n23347 , n343335 , n343336 , n343337 , n23351 , n23352 , n343340 , n343341 , n343342 , 
 n23356 , n23357 , n343345 , n343346 , n343347 , n23361 , n343349 , n343350 , n23364 , n343352 , 
 n343353 , n343354 , n23368 , n343356 , n343357 , n23371 , n343359 , n343360 , n23374 , n343362 , 
 n343363 , n343364 , n23378 , n343366 , n343367 , n343368 , n23382 , n343370 , n343371 , n23385 , 
 n23386 , n343374 , n343375 , n343376 , n343377 , n343378 , n343379 , n343380 , n343381 , n23395 , 
 n343383 , n343384 , n23398 , n343386 , n343387 , n343388 , n343389 , n343390 , n343391 , n23405 , 
 n23406 , n23407 , n343395 , n343396 , n23410 , n343398 , n343399 , n23413 , n343401 , n343402 , 
 n23416 , n23417 , n343405 , n343406 , n23420 , n343408 , n343409 , n23423 , n343411 , n23424 , 
 n343413 , n343414 , n343415 , n343416 , n343417 , n343418 , n343419 , n23430 , n23431 , n343422 , 
 n343423 , n343424 , n343425 , n343426 , n343427 , n343428 , n343429 , n343430 , n343431 , n23440 , 
 n343433 , n343434 , n343435 , n343436 , n343437 , n343438 , n343439 , n343440 , n23448 , n343442 , 
 n343443 , n343444 , n23452 , n343446 , n343447 , n343448 , n343449 , n343450 , n343451 , n343452 , 
 n343453 , n23459 , n23460 , n343456 , n23462 , n23463 , n23464 , n343460 , n343461 , n343462 , 
 n343463 , n343464 , n343465 , n23471 , n343467 , n343468 , n23474 , n23475 , n343471 , n23477 , 
 n343473 , n23479 , n343475 , n343476 , n343477 , n343478 , n343479 , n23485 , n343481 , n343482 , 
 n23488 , n23489 , n343485 , n343486 , n343487 , n343488 , n343489 , n343490 , n343491 , n343492 , 
 n343493 , n343494 , n343495 , n23499 , n343497 , n343498 , n23502 , n343500 , n343501 , n343502 , 
 n343503 , n343504 , n343505 , n343506 , n343507 , n343508 , n343509 , n343510 , n343511 , n343512 , 
 n343513 , n343514 , n23518 , n23519 , n343517 , n343518 , n23522 , n343520 , n343521 , n23525 , 
 n23526 , n343524 , n343525 , n23529 , n23530 , n343528 , n23532 , n343530 , n343531 , n343532 , 
 n343533 , n343534 , n343535 , n343536 , n343537 , n343538 , n23540 , n343540 , n23542 , n343542 , 
 n343543 , n23545 , n343545 , n343546 , n343547 , n343548 , n23550 , n23551 , n23552 , n343552 , 
 n343553 , n343554 , n23553 , n23554 , n343557 , n23556 , n23557 , n343560 , n23559 , n343562 , 
 n343563 , n343564 , n343565 , n343566 , n343567 , n343568 , n343569 , n343570 , n343571 , n343572 , 
 n343573 , n343574 , n343575 , n343576 , n343577 , n343578 , n343579 , n343580 , n343581 , n343582 , 
 n343583 , n343584 , n343585 , n343586 , n343587 , n23575 , n343589 , n343590 , n343591 , n343592 , 
 n343593 , n343594 , n343595 , n343596 , n343597 , n343598 , n343599 , n343600 , n343601 , n343602 , 
 n23590 , n343604 , n343605 , n23593 , n343607 , n343608 , n23596 , n343610 , n23598 , n343612 , 
 n343613 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n343620 , n23608 , n343622 , 
 n343623 , n343624 , n343625 , n343626 , n343627 , n343628 , n343629 , n343630 , n343631 , n343632 , 
 n343633 , n343634 , n343635 , n23612 , n23613 , n23614 , n343639 , n23615 , n23616 , n343642 , 
 n23618 , n343644 , n23620 , n23621 , n23622 , n343648 , n343649 , n343650 , n343651 , n343652 , 
 n23626 , n343654 , n343655 , n23629 , n23630 , n343658 , n23632 , n23633 , n343661 , n343662 , 
 n23636 , n23637 , n343665 , n343666 , n23640 , n343668 , n343669 , n23643 , n343671 , n343672 , 
 n343673 , n23647 , n343675 , n343676 , n23649 , n343678 , n343679 , n23652 , n343681 , n343682 , 
 n343683 , n23656 , n343685 , n343686 , n23659 , n343688 , n343689 , n343690 , n343691 , n23664 , 
 n343693 , n343694 , n23667 , n343696 , n343697 , n23670 , n343699 , n23672 , n343701 , n23674 , 
 n343703 , n343704 , n343705 , n343706 , n343707 , n23680 , n23681 , n343710 , n343711 , n23684 , 
 n343713 , n343714 , n23687 , n343716 , n343717 , n343718 , n343719 , n343720 , n343721 , n23692 , 
 n343723 , n23694 , n343725 , n23696 , n343727 , n343728 , n343729 , n343730 , n343731 , n343732 , 
 n23703 , n343734 , n343735 , n343736 , n343737 , n343738 , n343739 , n343740 , n343741 , n343742 , 
 n23713 , n343744 , n343745 , n343746 , n343747 , n343748 , n343749 , n343750 , n343751 , n343752 , 
 n343753 , n23723 , n343755 , n343756 , n343757 , n343758 , n343759 , n343760 , n23730 , n343762 , 
 n343763 , n23733 , n343765 , n23735 , n343767 , n343768 , n343769 , n343770 , n343771 , n343772 , 
 n343773 , n343774 , n343775 , n343776 , n343777 , n343778 , n343779 , n343780 , n343781 , n23750 , 
 n23751 , n343784 , n343785 , n23754 , n23755 , n343788 , n23757 , n23758 , n343791 , n23760 , 
 n343793 , n343794 , n23763 , n23764 , n343797 , n343798 , n23766 , n343800 , n343801 , n343802 , 
 n343803 , n343804 , n23772 , n343806 , n23774 , n343808 , n23776 , n23777 , n343811 , n343812 , 
 n23780 , n343814 , n343815 , n23783 , n343817 , n343818 , n23786 , n343820 , n23788 , n343822 , 
 n23790 , n23791 , n343825 , n343826 , n23794 , n23795 , n343829 , n23797 , n23798 , n343832 , 
 n23800 , n23801 , n343835 , n343836 , n343837 , n343838 , n343839 , n343840 , n343841 , n343842 , 
 n343843 , n343844 , n343845 , n343846 , n343847 , n343848 , n343849 , n343850 , n343851 , n343852 , 
 n343853 , n343854 , n343855 , n23823 , n343857 , n343858 , n23826 , n343860 , n343861 , n343862 , 
 n343863 , n343864 , n343865 , n343866 , n23834 , n343868 , n343869 , n343870 , n343871 , n343872 , 
 n343873 , n23841 , n343875 , n343876 , n23844 , n343878 , n343879 , n343880 , n343881 , n343882 , 
 n343883 , n343884 , n343885 , n343886 , n23854 , n343888 , n343889 , n343890 , n343891 , n23859 , 
 n23860 , n23861 , n343895 , n343896 , n23864 , n343898 , n343899 , n23867 , n23868 , n23869 , 
 n23870 , n343904 , n343905 , n343906 , n343907 , n343908 , n343909 , n343910 , n343911 , n23879 , 
 n343913 , n23881 , n343915 , n23883 , n343917 , n23885 , n343919 , n23887 , n343921 , n23889 , 
 n343923 , n23891 , n343925 , n343926 , n343927 , n343928 , n343929 , n343930 , n23898 , n343932 , 
 n343933 , n343934 , n23902 , n343936 , n343937 , n23905 , n23906 , n343940 , n23908 , n343942 , 
 n23910 , n23911 , n343945 , n343946 , n343947 , n343948 , n343949 , n23917 , n343951 , n23919 , 
 n343953 , n23921 , n343955 , n23923 , n343957 , n23925 , n343959 , n343960 , n23928 , n343962 , 
 n23930 , n343964 , n23932 , n343966 , n23934 , n343968 , n343969 , n343970 , n343971 , n343972 , 
 n343973 , n23941 , n343975 , n343976 , n343977 , n23945 , n343979 , n23947 , n23948 , n343982 , 
 n343983 , n23951 , n343985 , n343986 , n23954 , n23955 , n343989 , n23957 , n343991 , n343992 , 
 n343993 , n343994 , n343995 , n343996 , n343997 , n343998 , n343999 , n344000 , n344001 , n344002 , 
 n344003 , n23971 , n23972 , n344006 , n23974 , n344008 , n344009 , n23977 , n344011 , n344012 , 
 n23980 , n344014 , n344015 , n23983 , n344017 , n344018 , n344019 , n344020 , n344021 , n23989 , 
 n344023 , n23991 , n344025 , n23993 , n344027 , n23995 , n23996 , n344030 , n344031 , n344032 , 
 n344033 , n344034 , n344035 , n24003 , n24004 , n24005 , n24006 , n344040 , n24008 , n24009 , 
 n344043 , n344044 , n24012 , n344046 , n24014 , n24015 , n24016 , n24017 , n344051 , n24019 , 
 n344053 , n344054 , n344055 , n344056 , n344057 , n344058 , n24026 , n344060 , n344061 , n344062 , 
 n24030 , n344064 , n344065 , n344066 , n344067 , n344068 , n344069 , n344070 , n344071 , n344072 , 
 n344073 , n344074 , n344075 , n344076 , n24044 , n344078 , n344079 , n24047 , n344081 , n344082 , 
 n344083 , n24051 , n344085 , n344086 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , 
 n344093 , n24061 , n24062 , n344096 , n344097 , n24065 , n344099 , n344100 , n24068 , n344102 , 
 n344103 , n344104 , n24072 , n344106 , n344107 , n24075 , n344109 , n344110 , n24078 , n344112 , 
 n344113 , n344114 , n24082 , n344116 , n344117 , n24085 , n344119 , n24087 , n24088 , n24089 , 
 n24090 , n24091 , n24092 , n344126 , n344127 , n24095 , n344129 , n344130 , n24098 , n344132 , 
 n344133 , n344134 , n344135 , n344136 , n344137 , n24105 , n24106 , n344140 , n24108 , n24109 , 
 n24110 , n344144 , n24112 , n344146 , n24114 , n344148 , n344149 , n24117 , n344151 , n344152 , 
 n24120 , n344154 , n344155 , n344156 , n24124 , n344158 , n24126 , n344160 , n344161 , n344162 , 
 n344163 , n344164 , n344165 , n344166 , n344167 , n344168 , n344169 , n24137 , n344171 , n24139 , 
 n344173 , n344174 , n344175 , n344176 , n344177 , n344178 , n344179 , n24147 , n344181 , n24149 , 
 n24150 , n344184 , n344185 , n24153 , n344187 , n344188 , n344189 , n344190 , n344191 , n344192 , 
 n344193 , n344194 , n24162 , n344196 , n344197 , n24165 , n344199 , n24167 , n344201 , n24169 , 
 n344203 , n344204 , n24172 , n344206 , n344207 , n24175 , n24176 , n24177 , n344211 , n24179 , 
 n24180 , n344214 , n24182 , n24183 , n344217 , n24185 , n344219 , n344220 , n344221 , n344222 , 
 n344223 , n344224 , n344225 , n344226 , n24194 , n24195 , n344229 , n344230 , n344231 , n344232 , 
 n24200 , n344234 , n344235 , n24203 , n344237 , n344238 , n344239 , n344240 , n344241 , n344242 , 
 n344243 , n344244 , n344245 , n344246 , n344247 , n344248 , n24216 , n344250 , n24218 , n344252 , 
 n24220 , n24221 , n344255 , n344256 , n24224 , n344258 , n344259 , n344260 , n344261 , n344262 , 
 n344263 , n344264 , n344265 , n344266 , n344267 , n344268 , n344269 , n24237 , n344271 , n344272 , 
 n344273 , n344274 , n24242 , n24243 , n344277 , n344278 , n24246 , n344280 , n344281 , n344282 , 
 n24250 , n344284 , n344285 , n24253 , n24254 , n344288 , n344289 , n344290 , n344291 , n24259 , 
 n24260 , n24261 , n344295 , n344296 , n24264 , n24265 , n344299 , n344300 , n344301 , n344302 , 
 n344303 , n24271 , n344305 , n344306 , n24274 , n344308 , n344309 , n24277 , n24278 , n344312 , 
 n24280 , n344314 , n24282 , n24283 , n24284 , n344318 , n24286 , n24287 , n344321 , n344322 , 
 n24290 , n344324 , n344325 , n24293 , n24294 , n24295 , n24296 , n24297 , n344331 , n344332 , 
 n24300 , n344334 , n344335 , n344336 , n344337 , n344338 , n344339 , n344340 , n344341 , n344342 , 
 n344343 , n24311 , n344345 , n344346 , n24314 , n344348 , n344349 , n344350 , n344351 , n344352 , 
 n344353 , n344354 , n344355 , n24323 , n344357 , n344358 , n24326 , n344360 , n344361 , n344362 , 
 n24330 , n344364 , n344365 , n344366 , n344367 , n344368 , n24336 , n344370 , n344371 , n24339 , 
 n24340 , n24341 , n24342 , n24343 , n344377 , n24345 , n24346 , n344380 , n24348 , n24349 , 
 n344383 , n344384 , n24352 , n344386 , n344387 , n344388 , n344389 , n344390 , n344391 , n344392 , 
 n24360 , n344394 , n344395 , n24363 , n344397 , n24365 , n24366 , n344400 , n344401 , n24369 , 
 n344403 , n344404 , n24372 , n344406 , n24374 , n24375 , n24376 , n24377 , n24378 , n344412 , 
 n344413 , n344414 , n24382 , n24383 , n24384 , n344418 , n344419 , n24387 , n24388 , n24389 , 
 n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n344429 , n344430 , n24398 , n344432 , 
 n24400 , n24401 , n344435 , n344436 , n24404 , n344438 , n344439 , n24407 , n24408 , n344442 , 
 n344443 , n24411 , n344445 , n344446 , n24414 , n344448 , n344449 , n344450 , n344451 , n344452 , 
 n24420 , n344454 , n344455 , n344456 , n24424 , n344458 , n344459 , n24427 , n344461 , n344462 , 
 n344463 , n24431 , n24432 , n344466 , n344467 , n24435 , n344469 , n344470 , n24438 , n24439 , 
 n344473 , n344474 , n344475 , n24443 , n344477 , n344478 , n344479 , n344480 , n344481 , n344482 , 
 n344483 , n344484 , n24452 , n344486 , n344487 , n344488 , n344489 , n24457 , n344491 , n344492 , 
 n344493 , n344494 , n344495 , n24463 , n24464 , n24465 , n344499 , n344500 , n344501 , n344502 , 
 n344503 , n344504 , n344505 , n344506 , n344507 , n344508 , n344509 , n344510 , n344511 , n344512 , 
 n344513 , n344514 , n344515 , n24483 , n24484 , n24485 , n344519 , n344520 , n344521 , n344522 , 
 n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n344532 , 
 n344533 , n24501 , n344535 , n24503 , n344537 , n24505 , n344539 , n344540 , n24508 , n344542 , 
 n344543 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n344550 , n344551 , n344552 , 
 n344553 , n344554 , n344555 , n24523 , n344557 , n344558 , n344559 , n344560 , n24528 , n344562 , 
 n344563 , n24531 , n344565 , n344566 , n344567 , n344568 , n344569 , n344570 , n344571 , n344572 , 
 n24540 , n24541 , n24542 , n24543 , n344577 , n344578 , n24546 , n24547 , n344581 , n344582 , 
 n344583 , n24551 , n344585 , n24553 , n344587 , n344588 , n344589 , n344590 , n344591 , n344592 , 
 n344593 , n344594 , n344595 , n344596 , n344597 , n344598 , n344599 , n344600 , n24568 , n344602 , 
 n344603 , n344604 , n344605 , n24573 , n24574 , n344608 , n344609 , n24577 , n24578 , n24579 , 
 n344613 , n344614 , n24582 , n344616 , n344617 , n344618 , n24586 , n344620 , n24588 , n344622 , 
 n344623 , n24591 , n344625 , n344626 , n24594 , n24595 , n344629 , n24597 , n344631 , n344632 , 
 n24600 , n24601 , n344635 , n344636 , n24604 , n344638 , n24606 , n344640 , n344641 , n24609 , 
 n24610 , n24611 , n24612 , n344646 , n344647 , n344648 , n344649 , n344650 , n344651 , n344652 , 
 n344653 , n344654 , n344655 , n24623 , n344657 , n24625 , n24626 , n344660 , n24628 , n24629 , 
 n24630 , n24631 , n344665 , n24633 , n344667 , n344668 , n24636 , n344670 , n24638 , n344672 , 
 n344673 , n344674 , n344675 , n344676 , n344677 , n24645 , n344679 , n344680 , n344681 , n344682 , 
 n24650 , n344684 , n344685 , n344686 , n344687 , n344688 , n344689 , n344690 , n344691 , n24659 , 
 n24660 , n344694 , n344695 , n24663 , n344697 , n344698 , n344699 , n24667 , n24668 , n344702 , 
 n344703 , n344704 , n344705 , n344706 , n24674 , n344708 , n344709 , n344710 , n344711 , n344712 , 
 n344713 , n24681 , n344715 , n344716 , n344717 , n344718 , n344719 , n24687 , n344721 , n344722 , 
 n344723 , n24691 , n344725 , n344726 , n344727 , n24695 , n344729 , n24697 , n344731 , n24699 , 
 n24700 , n24701 , n344735 , n344736 , n344737 , n344738 , n344739 , n24707 , n24708 , n344742 , 
 n344743 , n24711 , n344745 , n344746 , n24714 , n344748 , n344749 , n24717 , n344751 , n344752 , 
 n24720 , n344754 , n344755 , n344756 , n344757 , n344758 , n344759 , n24727 , n344761 , n24729 , 
 n344763 , n24731 , n344765 , n24733 , n24734 , n24735 , n24736 , n344770 , n24738 , n344772 , 
 n344773 , n24741 , n344775 , n24743 , n344777 , n344778 , n24746 , n24747 , n344781 , n24749 , 
 n344783 , n344784 , n24752 , n24753 , n344787 , n344788 , n24756 , n344790 , n344791 , n344792 , 
 n24760 , n24761 , n344795 , n344796 , n344797 , n344798 , n344799 , n344800 , n344801 , n24769 , 
 n24770 , n24771 , n344805 , n24773 , n344807 , n344808 , n344809 , n344810 , n344811 , n344812 , 
 n344813 , n344814 , n344815 , n344816 , n344817 , n344818 , n24786 , n344820 , n344821 , n24789 , 
 n344823 , n344824 , n24792 , n344826 , n344827 , n344828 , n344829 , n344830 , n344831 , n24799 , 
 n24800 , n344834 , n24802 , n344836 , n344837 , n344838 , n344839 , n344840 , n344841 , n344842 , 
 n344843 , n344844 , n344845 , n344846 , n24814 , n344848 , n24816 , n24817 , n24818 , n344852 , 
 n344853 , n344854 , n344855 , n344856 , n344857 , n344858 , n344859 , n344860 , n24828 , n24829 , 
 n24830 , n24831 , n344865 , n344866 , n24834 , n344868 , n344869 , n24837 , n344871 , n344872 , 
 n24840 , n24841 , n24842 , n344876 , n344877 , n344878 , n344879 , n344880 , n24848 , n344882 , 
 n344883 , n24851 , n24852 , n24853 , n24854 , n24855 , n344889 , n24857 , n24858 , n344892 , 
 n344893 , n24861 , n344895 , n344896 , n344897 , n24865 , n344899 , n344900 , n344901 , n24869 , 
 n344903 , n344904 , n344905 , n344906 , n24874 , n24875 , n24876 , n24877 , n344911 , n344912 , 
 n24880 , n344914 , n24882 , n344916 , n24884 , n344918 , n344919 , n344920 , n24888 , n344922 , 
 n24890 , n24891 , n344925 , n24893 , n344927 , n344928 , n344929 , n24897 , n344931 , n24899 , 
 n344933 , n24901 , n344935 , n344936 , n344937 , n344938 , n344939 , n344940 , n24908 , n344942 , 
 n344943 , n24911 , n24912 , n344946 , n24914 , n344948 , n24916 , n344950 , n344951 , n344952 , 
 n24920 , n344954 , n344955 , n24923 , n344957 , n344958 , n344959 , n344960 , n344961 , n344962 , 
 n344963 , n344964 , n24932 , n24933 , n24934 , n344968 , n344969 , n344970 , n344971 , n24939 , 
 n24940 , n344974 , n24942 , n344976 , n344977 , n344978 , n24946 , n344980 , n24948 , n344982 , 
 n24950 , n24951 , n344985 , n344986 , n24954 , n344988 , n344989 , n24957 , n344991 , n344992 , 
 n344993 , n344994 , n344995 , n344996 , n24964 , n344998 , n344999 , n345000 , n24968 , n345002 , 
 n24970 , n345004 , n345005 , n345006 , n345007 , n345008 , n345009 , n345010 , n345011 , n345012 , 
 n345013 , n345014 , n345015 , n345016 , n345017 , n24985 , n345019 , n345020 , n345021 , n345022 , 
 n24990 , n345024 , n24992 , n24993 , n24994 , n345028 , n24996 , n24997 , n24998 , n345032 , 
 n345033 , n25001 , n345035 , n25003 , n345037 , n25005 , n345039 , n345040 , n25008 , n345042 , 
 n345043 , n345044 , n345045 , n25013 , n25014 , n345048 , n25016 , n345050 , n25018 , n345052 , 
 n25020 , n25021 , n25022 , n345056 , n25024 , n25025 , n345059 , n25027 , n345061 , n345062 , 
 n25030 , n25031 , n345065 , n25033 , n25034 , n25035 , n25036 , n345070 , n345071 , n345072 , 
 n345073 , n25041 , n345075 , n345076 , n25044 , n345078 , n345079 , n25047 , n345081 , n345082 , 
 n25050 , n345084 , n345085 , n25053 , n345087 , n25055 , n345089 , n25057 , n345091 , n345092 , 
 n345093 , n25061 , n345095 , n345096 , n345097 , n345098 , n345099 , n25067 , n345101 , n345102 , 
 n25070 , n345104 , n345105 , n345106 , n345107 , n345108 , n345109 , n25077 , n345111 , n345112 , 
 n345113 , n345114 , n25082 , n345116 , n25084 , n345118 , n345119 , n25087 , n345121 , n345122 , 
 n345123 , n25091 , n345125 , n25093 , n345127 , n25095 , n25096 , n345130 , n345131 , n345132 , 
 n345133 , n25101 , n345135 , n345136 , n345137 , n25105 , n345139 , n345140 , n345141 , n345142 , 
 n345143 , n345144 , n345145 , n345146 , n345147 , n345148 , n345149 , n25117 , n25118 , n345152 , 
 n345153 , n345154 , n25122 , n345156 , n25124 , n345158 , n345159 , n345160 , n345161 , n345162 , 
 n345163 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , 
 n25140 , n25141 , n345175 , n345176 , n25144 , n345178 , n345179 , n345180 , n345181 , n25149 , 
 n345183 , n25151 , n345185 , n25153 , n25154 , n345188 , n25156 , n345190 , n25158 , n25159 , 
 n25160 , n345194 , n25162 , n345196 , n345197 , n345198 , n345199 , n345200 , n345201 , n345202 , 
 n345203 , n345204 , n345205 , n25173 , n345207 , n25175 , n345209 , n25177 , n345211 , n345212 , 
 n25180 , n345214 , n345215 , n25183 , n25184 , n345218 , n25186 , n25187 , n25188 , n345222 , 
 n345223 , n345224 , n25192 , n345226 , n25194 , n345228 , n345229 , n345230 , n25198 , n345232 , 
 n345233 , n25201 , n345235 , n345236 , n345237 , n345238 , n345239 , n345240 , n345241 , n345242 , 
 n345243 , n345244 , n345245 , n25213 , n345247 , n345248 , n345249 , n345250 , n345251 , n345252 , 
 n345253 , n25221 , n345255 , n345256 , n345257 , n345258 , n25226 , n345260 , n345261 , n345262 , 
 n345263 , n345264 , n25232 , n345266 , n25234 , n25235 , n25236 , n345270 , n345271 , n25239 , 
 n345273 , n345274 , n345275 , n345276 , n345277 , n345278 , n25246 , n345280 , n345281 , n25249 , 
 n345283 , n345284 , n25252 , n25253 , n345287 , n25255 , n345289 , n345290 , n345291 , n25259 , 
 n345293 , n345294 , n345295 , n345296 , n345297 , n25265 , n345299 , n345300 , n25268 , n345302 , 
 n25270 , n345304 , n345305 , n25273 , n25274 , n345308 , n25276 , n345310 , n25278 , n345312 , 
 n345313 , n345314 , n345315 , n25283 , n345317 , n345318 , n25286 , n345320 , n345321 , n345322 , 
 n345323 , n345324 , n25292 , n25293 , n345327 , n25295 , n345329 , n345330 , n345331 , n25299 , 
 n345333 , n345334 , n25302 , n25303 , n345337 , n25305 , n25306 , n25307 , n25308 , n25309 , 
 n345343 , n345344 , n345345 , n345346 , n25314 , n345348 , n345349 , n345350 , n345351 , n345352 , 
 n345353 , n345354 , n25322 , n345356 , n345357 , n25325 , n345359 , n345360 , n345361 , n25329 , 
 n345363 , n345364 , n25332 , n345366 , n25334 , n25335 , n345369 , n25337 , n345371 , n345372 , 
 n345373 , n345374 , n345375 , n345376 , n345377 , n345378 , n345379 , n345380 , n345381 , n25349 , 
 n25350 , n25351 , n25352 , n345386 , n345387 , n345388 , n345389 , n345390 , n345391 , n25359 , 
 n345393 , n345394 , n345395 , n345396 , n345397 , n25365 , n345399 , n25367 , n345401 , n25369 , 
 n345403 , n25371 , n345405 , n345406 , n345407 , n345408 , n25376 , n345410 , n25378 , n345412 , 
 n345413 , n25381 , n345415 , n345416 , n25384 , n25385 , n345419 , n25387 , n345421 , n345422 , 
 n345423 , n345424 , n345425 , n345426 , n345427 , n345428 , n345429 , n25397 , n345431 , n25399 , 
 n345433 , n25401 , n25402 , n25403 , n345437 , n345438 , n25406 , n345440 , n345441 , n345442 , 
 n345443 , n345444 , n345445 , n345446 , n345447 , n345448 , n25416 , n345450 , n345451 , n345452 , 
 n345453 , n345454 , n25422 , n25423 , n25424 , n25425 , n25426 , n345460 , n345461 , n25429 , 
 n345463 , n345464 , n345465 , n25433 , n345467 , n25435 , n345469 , n345470 , n25438 , n345472 , 
 n25440 , n345474 , n345475 , n345476 , n345477 , n345478 , n345479 , n25447 , n345481 , n25449 , 
 n345483 , n345484 , n345485 , n345486 , n25454 , n25455 , n345489 , n25457 , n345491 , n25459 , 
 n345493 , n345494 , n25462 , n345496 , n345497 , n345498 , n345499 , n345500 , n345501 , n345502 , 
 n345503 , n345504 , n345505 , n345506 , n345507 , n25475 , n345509 , n345510 , n345511 , n25479 , 
 n25480 , n345514 , n345515 , n345516 , n345517 , n345518 , n345519 , n345520 , n345521 , n25489 , 
 n345523 , n345524 , n25492 , n25493 , n345527 , n345528 , n345529 , n345530 , n25498 , n345532 , 
 n345533 , n25501 , n345535 , n345536 , n25504 , n345538 , n345539 , n25507 , n345541 , n345542 , 
 n345543 , n25511 , n345545 , n345546 , n345547 , n345548 , n25516 , n345550 , n345551 , n345552 , 
 n345553 , n345554 , n345555 , n25523 , n345557 , n345558 , n345559 , n345560 , n25528 , n25529 , 
 n345563 , n345564 , n345565 , n25533 , n345567 , n345568 , n25536 , n345570 , n345571 , n345572 , 
 n25540 , n345574 , n345575 , n345576 , n345577 , n345578 , n345579 , n25547 , n345581 , n345582 , 
 n345583 , n345584 , n345585 , n345586 , n345587 , n345588 , n345589 , n25557 , n345591 , n345592 , 
 n345593 , n345594 , n345595 , n25563 , n345597 , n345598 , n25566 , n345600 , n345601 , n345602 , 
 n345603 , n345604 , n345605 , n25573 , n345607 , n345608 , n25576 , n345610 , n345611 , n345612 , 
 n345613 , n345614 , n345615 , n345616 , n345617 , n345618 , n345619 , n25587 , n345621 , n345622 , 
 n345623 , n345624 , n25592 , n25593 , n345627 , n345628 , n25596 , n25597 , n345631 , n345632 , 
 n345633 , n345634 , n25602 , n345636 , n345637 , n345638 , n345639 , n25607 , n25608 , n345642 , 
 n345643 , n345644 , n25612 , n25613 , n345647 , n345648 , n25616 , n25617 , n25618 , n345652 , 
 n345653 , n25621 , n25622 , n345656 , n345657 , n345658 , n345659 , n25627 , n345661 , n345662 , 
 n345663 , n25631 , n345665 , n25633 , n345667 , n345668 , n345669 , n25637 , n25638 , n345672 , 
 n345673 , n25641 , n345675 , n345676 , n345677 , n345678 , n25646 , n345680 , n345681 , n345682 , 
 n25650 , n25651 , n25652 , n345686 , n25654 , n345688 , n345689 , n345690 , n345691 , n345692 , 
 n345693 , n345694 , n345695 , n345696 , n25664 , n25665 , n345699 , n25667 , n25668 , n25669 , 
 n345703 , n25671 , n345705 , n345706 , n25674 , n345708 , n345709 , n345710 , n345711 , n25679 , 
 n345713 , n345714 , n345715 , n345716 , n25684 , n345718 , n345719 , n25687 , n345721 , n345722 , 
 n25690 , n25691 , n345725 , n345726 , n345727 , n345728 , n345729 , n25697 , n345731 , n345732 , 
 n345733 , n345734 , n345735 , n345736 , n25704 , n345738 , n25706 , n345740 , n25708 , n25709 , 
 n345743 , n25711 , n345745 , n345746 , n25714 , n345748 , n345749 , n25717 , n345751 , n345752 , 
 n25720 , n345754 , n25722 , n25723 , n345757 , n25725 , n25726 , n345760 , n25728 , n345762 , 
 n345763 , n345764 , n345765 , n345766 , n345767 , n345768 , n345769 , n25737 , n345771 , n345772 , 
 n25740 , n345774 , n345775 , n345776 , n25744 , n345778 , n345779 , n345780 , n345781 , n345782 , 
 n345783 , n345784 , n345785 , n345786 , n345787 , n25755 , n345789 , n345790 , n25758 , n25759 , 
 n345793 , n25761 , n25762 , n25763 , n345797 , n345798 , n345799 , n345800 , n345801 , n345802 , 
 n345803 , n25771 , n345805 , n345806 , n345807 , n345808 , n345809 , n345810 , n345811 , n345812 , 
 n345813 , n345814 , n25782 , n345816 , n345817 , n25785 , n345819 , n345820 , n345821 , n345822 , 
 n345823 , n345824 , n345825 , n345826 , n345827 , n345828 , n345829 , n345830 , n345831 , n25799 , 
 n345833 , n345834 , n25802 , n345836 , n345837 , n345838 , n345839 , n345840 , n345841 , n345842 , 
 n345843 , n345844 , n345845 , n25813 , n25814 , n345848 , n345849 , n345850 , n345851 , n25819 , 
 n345853 , n25821 , n25822 , n345856 , n25824 , n345858 , n345859 , n345860 , n345861 , n345862 , 
 n345863 , n345864 , n345865 , n25833 , n345867 , n25835 , n345869 , n345870 , n345871 , n345872 , 
 n345873 , n25841 , n345875 , n345876 , n25844 , n345878 , n345879 , n345880 , n345881 , n345882 , 
 n345883 , n25851 , n345885 , n345886 , n25854 , n345888 , n345889 , n25857 , n345891 , n345892 , 
 n345893 , n25861 , n345895 , n345896 , n345897 , n345898 , n345899 , n345900 , n345901 , n25869 , 
 n345903 , n345904 , n345905 , n25873 , n25874 , n345908 , n345909 , n25877 , n25878 , n345912 , 
 n345913 , n25881 , n345915 , n345916 , n345917 , n345918 , n345919 , n25887 , n345921 , n345922 , 
 n345923 , n345924 , n25892 , n345926 , n345927 , n25895 , n345929 , n345930 , n25898 , n345932 , 
 n345933 , n345934 , n345935 , n25903 , n345937 , n25905 , n25906 , n345940 , n25908 , n345942 , 
 n345943 , n345944 , n345945 , n345946 , n345947 , n345948 , n345949 , n345950 , n345951 , n25919 , 
 n345953 , n345954 , n345955 , n345956 , n345957 , n345958 , n345959 , n345960 , n25928 , n345962 , 
 n25930 , n345964 , n345965 , n25933 , n345967 , n345968 , n345969 , n345970 , n345971 , n345972 , 
 n25940 , n25941 , n345975 , n25943 , n345977 , n25945 , n345979 , n345980 , n345981 , n345982 , 
 n25950 , n345984 , n345985 , n345986 , n345987 , n345988 , n345989 , n25957 , n345991 , n345992 , 
 n345993 , n345994 , n345995 , n345996 , n345997 , n25965 , n345999 , n346000 , n25968 , n346002 , 
 n25970 , n346004 , n346005 , n346006 , n25974 , n346008 , n25976 , n346010 , n346011 , n25979 , 
 n346013 , n346014 , n25982 , n25983 , n25984 , n25985 , n346019 , n346020 , n346021 , n346022 , 
 n346023 , n25991 , n346025 , n25993 , n25994 , n25995 , n25996 , n25997 , n346031 , n25999 , 
 n26000 , n346034 , n26002 , n26003 , n346037 , n346038 , n346039 , n346040 , n346041 , n346042 , 
 n26010 , n346044 , n346045 , n26013 , n346047 , n346048 , n26016 , n346050 , n26018 , n346052 , 
 n26020 , n26021 , n26022 , n346056 , n346057 , n346058 , n346059 , n346060 , n346061 , n26029 , 
 n346063 , n346064 , n26032 , n26033 , n346067 , n26035 , n346069 , n346070 , n26038 , n346072 , 
 n346073 , n26041 , n346075 , n346076 , n346077 , n346078 , n26046 , n346080 , n346081 , n26049 , 
 n26050 , n346084 , n26052 , n26053 , n346087 , n346088 , n346089 , n346090 , n26058 , n26059 , 
 n346093 , n26061 , n346095 , n346096 , n346097 , n346098 , n346099 , n346100 , n26068 , n346102 , 
 n346103 , n346104 , n346105 , n346106 , n346107 , n346108 , n346109 , n26077 , n346111 , n26079 , 
 n26080 , n346114 , n346115 , n26083 , n346117 , n346118 , n346119 , n346120 , n346121 , n346122 , 
 n346123 , n26091 , n346125 , n346126 , n346127 , n346128 , n346129 , n346130 , n346131 , n346132 , 
 n346133 , n346134 , n346135 , n346136 , n26104 , n346138 , n346139 , n26107 , n346141 , n346142 , 
 n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n346150 , n26118 , n346152 , 
 n346153 , n26121 , n26122 , n346156 , n346157 , n346158 , n346159 , n26127 , n346161 , n346162 , 
 n26130 , n346164 , n346165 , n26133 , n346167 , n346168 , n346169 , n346170 , n346171 , n346172 , 
 n346173 , n346174 , n346175 , n346176 , n26144 , n346178 , n346179 , n346180 , n346181 , n26149 , 
 n26150 , n346184 , n346185 , n346186 , n346187 , n346188 , n26156 , n346190 , n26158 , n26159 , 
 n346193 , n346194 , n26162 , n346196 , n346197 , n26165 , n346199 , n346200 , n26168 , n346202 , 
 n346203 , n26171 , n346205 , n346206 , n346207 , n26175 , n346209 , n346210 , n26178 , n26179 , 
 n346213 , n346214 , n346215 , n346216 , n346217 , n26185 , n26186 , n346220 , n26188 , n346222 , 
 n346223 , n346224 , n26192 , n26193 , n346227 , n346228 , n346229 , n26197 , n346231 , n346232 , 
 n346233 , n346234 , n346235 , n346236 , n346237 , n346238 , n346239 , n26207 , n346241 , n26209 , 
 n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n346249 , n346250 , n26218 , n26219 , 
 n346253 , n346254 , n346255 , n346256 , n346257 , n346258 , n346259 , n346260 , n346261 , n26229 , 
 n346263 , n346264 , n26232 , n26233 , n346267 , n26235 , n346269 , n26237 , n346271 , n26239 , 
 n346273 , n346274 , n346275 , n346276 , n346277 , n346278 , n346279 , n346280 , n346281 , n346282 , 
 n26250 , n346284 , n346285 , n346286 , n26254 , n26255 , n346289 , n346290 , n346291 , n346292 , 
 n346293 , n346294 , n26262 , n346296 , n346297 , n346298 , n346299 , n26267 , n346301 , n346302 , 
 n346303 , n346304 , n346305 , n346306 , n346307 , n346308 , n346309 , n346310 , n346311 , n346312 , 
 n346313 , n346314 , n346315 , n346316 , n346317 , n346318 , n346319 , n26287 , n346321 , n346322 , 
 n346323 , n346324 , n346325 , n26293 , n346327 , n346328 , n26296 , n346330 , n346331 , n346332 , 
 n26300 , n26301 , n346335 , n346336 , n26304 , n346338 , n346339 , n26307 , n346341 , n346342 , 
 n26310 , n346344 , n346345 , n346346 , n26314 , n346348 , n26316 , n346350 , n346351 , n346352 , 
 n26320 , n346354 , n26322 , n346356 , n346357 , n26325 , n26326 , n346360 , n346361 , n346362 , 
 n26330 , n26331 , n346365 , n26333 , n346367 , n346368 , n346369 , n346370 , n346371 , n346372 , 
 n26340 , n346374 , n346375 , n346376 , n346377 , n346378 , n346379 , n346380 , n346381 , n346382 , 
 n346383 , n26351 , n346385 , n346386 , n26354 , n346388 , n346389 , n346390 , n346391 , n346392 , 
 n346393 , n346394 , n346395 , n26363 , n346397 , n346398 , n346399 , n26367 , n346401 , n346402 , 
 n346403 , n346404 , n346405 , n26373 , n26374 , n346408 , n346409 , n346410 , n26378 , n346412 , 
 n26380 , n26381 , n26382 , n346416 , n346417 , n346418 , n346419 , n26387 , n346421 , n346422 , 
 n26390 , n346424 , n346425 , n26393 , n346427 , n346428 , n26396 , n346430 , n346431 , n346432 , 
 n346433 , n26401 , n26402 , n26403 , n26404 , n26405 , n346439 , n346440 , n26408 , n26409 , 
 n26410 , n26411 , n346445 , n26413 , n346447 , n26415 , n26416 , n26417 , n26418 , n26419 , 
 n26420 , n26421 , n26422 , n26423 , n346457 , n26425 , n346459 , n26427 , n346461 , n26429 , 
 n346463 , n346464 , n346465 , n26433 , n346467 , n346468 , n346469 , n26437 , n346471 , n346472 , 
 n346473 , n346474 , n346475 , n346476 , n26444 , n26445 , n346479 , n346480 , n26448 , n346482 , 
 n346483 , n26451 , n346485 , n346486 , n26454 , n346488 , n346489 , n346490 , n346491 , n346492 , 
 n346493 , n346494 , n346495 , n26463 , n346497 , n346498 , n26466 , n346500 , n346501 , n26469 , 
 n346503 , n346504 , n26472 , n346506 , n346507 , n26475 , n346509 , n26477 , n346511 , n346512 , 
 n346513 , n346514 , n26482 , n346516 , n346517 , n26485 , n346519 , n346520 , n26488 , n346522 , 
 n346523 , n346524 , n26492 , n346526 , n346527 , n26495 , n346529 , n346530 , n346531 , n26499 , 
 n346533 , n346534 , n26502 , n346536 , n346537 , n346538 , n346539 , n346540 , n346541 , n346542 , 
 n346543 , n346544 , n346545 , n346546 , n26514 , n346548 , n346549 , n346550 , n346551 , n346552 , 
 n346553 , n346554 , n26522 , n346556 , n346557 , n346558 , n346559 , n346560 , n346561 , n346562 , 
 n26530 , n346564 , n346565 , n346566 , n346567 , n346568 , n26536 , n346570 , n346571 , n346572 , 
 n346573 , n346574 , n346575 , n26543 , n346577 , n346578 , n26546 , n346580 , n346581 , n26549 , 
 n346583 , n346584 , n346585 , n26553 , n346587 , n346588 , n26556 , n346590 , n346591 , n346592 , 
 n346593 , n26561 , n346595 , n346596 , n26564 , n346598 , n346599 , n26567 , n346601 , n346602 , 
 n346603 , n26571 , n26572 , n26573 , n26574 , n26575 , n346609 , n26577 , n346611 , n26579 , 
 n346613 , n26581 , n26582 , n346616 , n26584 , n346618 , n26586 , n26587 , n346621 , n346622 , 
 n26590 , n26591 , n346625 , n26593 , n346627 , n346628 , n346629 , n26597 , n346631 , n346632 , 
 n26600 , n346634 , n346635 , n346636 , n26604 , n26605 , n346639 , n346640 , n26608 , n346642 , 
 n346643 , n346644 , n346645 , n346646 , n26614 , n346648 , n26616 , n26617 , n26618 , n346652 , 
 n26620 , n346654 , n346655 , n346656 , n346657 , n346658 , n346659 , n346660 , n346661 , n346662 , 
 n346663 , n26631 , n26632 , n346666 , n346667 , n346668 , n26636 , n346670 , n26638 , n26639 , 
 n346673 , n26641 , n346675 , n346676 , n26644 , n346678 , n346679 , n346680 , n346681 , n346682 , 
 n346683 , n346684 , n346685 , n346686 , n26654 , n346688 , n346689 , n26657 , n346691 , n346692 , 
 n346693 , n26661 , n346695 , n346696 , n346697 , n26665 , n346699 , n346700 , n346701 , n346702 , 
 n346703 , n26671 , n346705 , n346706 , n346707 , n26675 , n346709 , n346710 , n26678 , n346712 , 
 n346713 , n26681 , n346715 , n346716 , n346717 , n346718 , n346719 , n26687 , n346721 , n346722 , 
 n346723 , n346724 , n26692 , n346726 , n346727 , n26695 , n346729 , n346730 , n346731 , n346732 , 
 n346733 , n346734 , n346735 , n346736 , n346737 , n346738 , n346739 , n346740 , n346741 , n346742 , 
 n346743 , n346744 , n346745 , n26713 , n346747 , n346748 , n26716 , n26717 , n346751 , n26719 , 
 n346753 , n26721 , n346755 , n346756 , n346757 , n346758 , n346759 , n346760 , n346761 , n346762 , 
 n346763 , n346764 , n346765 , n346766 , n346767 , n26735 , n346769 , n346770 , n346771 , n26739 , 
 n26740 , n346774 , n346775 , n346776 , n346777 , n346778 , n346779 , n346780 , n346781 , n26749 , 
 n346783 , n26751 , n346785 , n26753 , n346787 , n346788 , n346789 , n346790 , n26758 , n346792 , 
 n346793 , n346794 , n26762 , n26763 , n346797 , n26765 , n346799 , n346800 , n346801 , n346802 , 
 n26770 , n346804 , n346805 , n26773 , n346807 , n346808 , n26776 , n346810 , n26778 , n346812 , 
 n26780 , n26781 , n346815 , n346816 , n346817 , n26785 , n26786 , n26787 , n346821 , n346822 , 
 n346823 , n346824 , n346825 , n346826 , n346827 , n346828 , n26796 , n26797 , n346831 , n26799 , 
 n346833 , n346834 , n26802 , n346836 , n346837 , n26805 , n346839 , n346840 , n26808 , n26809 , 
 n346843 , n26811 , n346845 , n26813 , n346847 , n346848 , n26816 , n346850 , n346851 , n346852 , 
 n346853 , n346854 , n346855 , n26823 , n346857 , n26825 , n346859 , n26827 , n346861 , n346862 , 
 n26830 , n26831 , n26832 , n346866 , n26834 , n26835 , n346869 , n346870 , n26838 , n346872 , 
 n346873 , n26841 , n346875 , n346876 , n346877 , n26845 , n346879 , n26847 , n26848 , n346882 , 
 n26850 , n26851 , n346885 , n26853 , n346887 , n346888 , n346889 , n346890 , n346891 , n346892 , 
 n26860 , n346894 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n346902 , 
 n346903 , n26871 , n346905 , n346906 , n346907 , n346908 , n26876 , n346910 , n346911 , n346912 , 
 n26880 , n26881 , n26882 , n346916 , n346917 , n346918 , n26886 , n26887 , n346921 , n346922 , 
 n346923 , n346924 , n26892 , n346926 , n346927 , n26895 , n346929 , n346930 , n346931 , n346932 , 
 n346933 , n26901 , n346935 , n26903 , n346937 , n26905 , n346939 , n346940 , n26908 , n346942 , 
 n346943 , n26911 , n346945 , n346946 , n26914 , n346948 , n346949 , n346950 , n346951 , n346952 , 
 n346953 , n26921 , n346955 , n346956 , n26924 , n346958 , n346959 , n346960 , n346961 , n346962 , 
 n346963 , n346964 , n346965 , n346966 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , 
 n346973 , n346974 , n346975 , n26943 , n346977 , n346978 , n346979 , n346980 , n346981 , n346982 , 
 n346983 , n346984 , n346985 , n346986 , n346987 , n346988 , n346989 , n26957 , n346991 , n346992 , 
 n346993 , n26961 , n346995 , n346996 , n26964 , n346998 , n346999 , n347000 , n26968 , n347002 , 
 n26970 , n347004 , n26972 , n26973 , n347007 , n26975 , n347009 , n26977 , n26978 , n347012 , 
 n347013 , n347014 , n347015 , n347016 , n26984 , n347018 , n347019 , n347020 , n26988 , n347022 , 
 n347023 , n26991 , n347025 , n347026 , n26994 , n347028 , n347029 , n26997 , n347031 , n347032 , 
 n347033 , n27001 , n27002 , n27003 , n347037 , n347038 , n347039 , n347040 , n347041 , n347042 , 
 n347043 , n27011 , n347045 , n347046 , n27014 , n347048 , n347049 , n347050 , n347051 , n347052 , 
 n347053 , n27021 , n347055 , n347056 , n347057 , n347058 , n347059 , n347060 , n347061 , n347062 , 
 n347063 , n347064 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n347071 , n347072 , 
 n27040 , n347074 , n27042 , n347076 , n347077 , n347078 , n347079 , n347080 , n347081 , n347082 , 
 n347083 , n347084 , n347085 , n347086 , n347087 , n347088 , n347089 , n347090 , n347091 , n27059 , 
 n347093 , n347094 , n347095 , n347096 , n27064 , n347098 , n347099 , n347100 , n347101 , n347102 , 
 n347103 , n347104 , n347105 , n347106 , n347107 , n347108 , n347109 , n347110 , n347111 , n347112 , 
 n27080 , n347114 , n347115 , n347116 , n347117 , n347118 , n27086 , n347120 , n347121 , n27089 , 
 n347123 , n347124 , n27092 , n347126 , n347127 , n347128 , n347129 , n347130 , n27098 , n27099 , 
 n27100 , n347134 , n347135 , n347136 , n27104 , n347138 , n347139 , n347140 , n27108 , n347142 , 
 n347143 , n27111 , n347145 , n347146 , n347147 , n347148 , n347149 , n347150 , n347151 , n347152 , 
 n347153 , n347154 , n347155 , n347156 , n347157 , n347158 , n27126 , n347160 , n347161 , n347162 , 
 n347163 , n347164 , n347165 , n27133 , n347167 , n347168 , n347169 , n347170 , n347171 , n27139 , 
 n347173 , n347174 , n27142 , n27143 , n347177 , n347178 , n347179 , n347180 , n347181 , n347182 , 
 n347183 , n347184 , n347185 , n347186 , n347187 , n27155 , n27156 , n347190 , n347191 , n347192 , 
 n347193 , n347194 , n27162 , n347196 , n347197 , n27165 , n27166 , n347200 , n347201 , n347202 , 
 n347203 , n27171 , n27172 , n27173 , n347207 , n27175 , n347209 , n27177 , n347211 , n27179 , 
 n347213 , n27181 , n347215 , n347216 , n347217 , n347218 , n27186 , n347220 , n347221 , n27189 , 
 n347223 , n27191 , n347225 , n347226 , n347227 , n347228 , n347229 , n27197 , n347231 , n347232 , 
 n27200 , n347234 , n347235 , n347236 , n347237 , n347238 , n347239 , n347240 , n27208 , n27209 , 
 n347243 , n27211 , n27212 , n27213 , n347247 , n347248 , n27216 , n347250 , n27218 , n347252 , 
 n27220 , n347254 , n347255 , n347256 , n27224 , n347258 , n27226 , n27227 , n347261 , n347262 , 
 n27230 , n27231 , n27232 , n347266 , n27234 , n27235 , n347269 , n27237 , n347271 , n347272 , 
 n27240 , n347274 , n27242 , n347276 , n347277 , n27245 , n27246 , n27247 , n347281 , n347282 , 
 n27250 , n27251 , n347285 , n347286 , n27254 , n347288 , n27256 , n347290 , n27258 , n347292 , 
 n27260 , n27261 , n347295 , n347296 , n27264 , n347298 , n347299 , n27267 , n347301 , n347302 , 
 n27270 , n27271 , n347305 , n347306 , n27274 , n347308 , n347309 , n27277 , n347311 , n347312 , 
 n347313 , n347314 , n347315 , n347316 , n347317 , n27285 , n347319 , n347320 , n347321 , n27289 , 
 n347323 , n347324 , n27292 , n347326 , n347327 , n27295 , n347329 , n347330 , n347331 , n347332 , 
 n347333 , n347334 , n347335 , n347336 , n27304 , n27305 , n347339 , n347340 , n27308 , n347342 , 
 n347343 , n27311 , n347345 , n347346 , n347347 , n347348 , n347349 , n27317 , n347351 , n347352 , 
 n27320 , n347354 , n347355 , n347356 , n347357 , n347358 , n347359 , n27327 , n27328 , n347362 , 
 n347363 , n347364 , n27332 , n347366 , n347367 , n347368 , n347369 , n347370 , n347371 , n347372 , 
 n347373 , n347374 , n27342 , n347376 , n347377 , n27345 , n347379 , n347380 , n347381 , n347382 , 
 n27350 , n27351 , n347385 , n27353 , n347387 , n347388 , n347389 , n347390 , n347391 , n27359 , 
 n347393 , n347394 , n347395 , n347396 , n27364 , n347398 , n27366 , n347400 , n27368 , n347402 , 
 n27370 , n347404 , n347405 , n27373 , n347407 , n347408 , n347409 , n347410 , n347411 , n347412 , 
 n347413 , n347414 , n347415 , n27383 , n27384 , n27385 , n347419 , n27387 , n347421 , n27389 , 
 n347423 , n347424 , n347425 , n347426 , n347427 , n347428 , n27396 , n347430 , n347431 , n347432 , 
 n27400 , n347434 , n347435 , n347436 , n347437 , n347438 , n347439 , n27407 , n27408 , n347442 , 
 n347443 , n347444 , n347445 , n347446 , n27414 , n347448 , n347449 , n27417 , n27418 , n27419 , 
 n347453 , n347454 , n347455 , n27423 , n347457 , n347458 , n347459 , n27427 , n27428 , n27429 , 
 n347463 , n27431 , n347465 , n27433 , n27434 , n347468 , n347469 , n27437 , n347471 , n347472 , 
 n27440 , n347474 , n27442 , n347476 , n347477 , n347478 , n27446 , n347480 , n347481 , n347482 , 
 n347483 , n347484 , n27452 , n347486 , n347487 , n27455 , n347489 , n347490 , n347491 , n27459 , 
 n347493 , n27461 , n347495 , n27463 , n347497 , n27465 , n347499 , n27467 , n347501 , n347502 , 
 n347503 , n347504 , n27472 , n347506 , n347507 , n347508 , n27476 , n347510 , n347511 , n27479 , 
 n347513 , n347514 , n27482 , n27483 , n347517 , n347518 , n347519 , n347520 , n347521 , n27489 , 
 n347523 , n347524 , n347525 , n27493 , n347527 , n27495 , n27496 , n347530 , n347531 , n347532 , 
 n347533 , n347534 , n347535 , n347536 , n347537 , n347538 , n347539 , n347540 , n27508 , n347542 , 
 n347543 , n347544 , n347545 , n347546 , n347547 , n347548 , n347549 , n347550 , n347551 , n27519 , 
 n347553 , n347554 , n347555 , n347556 , n347557 , n27525 , n27526 , n27527 , n347561 , n347562 , 
 n27530 , n347564 , n27532 , n347566 , n347567 , n27535 , n347569 , n347570 , n347571 , n347572 , 
 n347573 , n27541 , n347575 , n347576 , n27544 , n27545 , n347579 , n347580 , n347581 , n347582 , 
 n347583 , n347584 , n347585 , n347586 , n27554 , n27555 , n27556 , n27557 , n27558 , n347592 , 
 n347593 , n27561 , n347595 , n347596 , n347597 , n347598 , n27566 , n347600 , n347601 , n347602 , 
 n27570 , n347604 , n27572 , n347606 , n347607 , n347608 , n27576 , n27577 , n347611 , n347612 , 
 n27580 , n347614 , n347615 , n347616 , n347617 , n347618 , n27586 , n27587 , n347621 , n27589 , 
 n347623 , n27591 , n27592 , n347626 , n347627 , n347628 , n347629 , n347630 , n27598 , n347632 , 
 n347633 , n347634 , n347635 , n347636 , n347637 , n347638 , n347639 , n27607 , n347641 , n347642 , 
 n27610 , n347644 , n347645 , n347646 , n27614 , n347648 , n347649 , n27617 , n347651 , n347652 , 
 n347653 , n347654 , n27622 , n347656 , n347657 , n347658 , n27626 , n347660 , n347661 , n347662 , 
 n27630 , n347664 , n347665 , n347666 , n347667 , n347668 , n347669 , n27637 , n347671 , n347672 , 
 n27640 , n347674 , n27642 , n347676 , n347677 , n347678 , n347679 , n347680 , n347681 , n347682 , 
 n347683 , n347684 , n347685 , n27653 , n347687 , n347688 , n347689 , n347690 , n347691 , n27659 , 
 n347693 , n27661 , n347695 , n27663 , n347697 , n347698 , n27666 , n347700 , n27668 , n27669 , 
 n347703 , n27671 , n347705 , n347706 , n347707 , n27675 , n347709 , n347710 , n27678 , n347712 , 
 n347713 , n27681 , n347715 , n347716 , n27684 , n347718 , n347719 , n27687 , n347721 , n347722 , 
 n347723 , n347724 , n347725 , n347726 , n27694 , n347728 , n347729 , n347730 , n347731 , n347732 , 
 n347733 , n347734 , n347735 , n347736 , n347737 , n347738 , n27706 , n347740 , n347741 , n347742 , 
 n347743 , n347744 , n347745 , n347746 , n347747 , n347748 , n347749 , n347750 , n347751 , n347752 , 
 n347753 , n347754 , n347755 , n27723 , n347757 , n27725 , n347759 , n347760 , n347761 , n347762 , 
 n347763 , n347764 , n347765 , n347766 , n347767 , n347768 , n27736 , n347770 , n347771 , n347772 , 
 n347773 , n347774 , n347775 , n27743 , n347777 , n347778 , n347779 , n347780 , n347781 , n347782 , 
 n347783 , n347784 , n347785 , n347786 , n27754 , n347788 , n347789 , n347790 , n347791 , n27759 , 
 n347793 , n347794 , n27762 , n27763 , n347797 , n347798 , n347799 , n347800 , n27768 , n347802 , 
 n347803 , n347804 , n347805 , n27773 , n347807 , n347808 , n347809 , n347810 , n347811 , n347812 , 
 n347813 , n27781 , n347815 , n27783 , n347817 , n347818 , n27786 , n347820 , n347821 , n27789 , 
 n347823 , n347824 , n347825 , n347826 , n347827 , n347828 , n347829 , n27797 , n27798 , n347832 , 
 n27800 , n347834 , n347835 , n347836 , n347837 , n27805 , n27806 , n347840 , n27808 , n347842 , 
 n347843 , n347844 , n27812 , n347846 , n347847 , n347848 , n347849 , n347850 , n347851 , n347852 , 
 n347853 , n347854 , n347855 , n347856 , n27824 , n347858 , n347859 , n347860 , n347861 , n347862 , 
 n347863 , n347864 , n347865 , n347866 , n347867 , n347868 , n347869 , n347870 , n27838 , n27839 , 
 n27840 , n347874 , n347875 , n347876 , n27844 , n347878 , n347879 , n347880 , n347881 , n27849 , 
 n347883 , n347884 , n347885 , n347886 , n27854 , n347888 , n347889 , n347890 , n347891 , n347892 , 
 n347893 , n347894 , n347895 , n347896 , n347897 , n347898 , n347899 , n347900 , n27868 , n27869 , 
 n27870 , n347904 , n347905 , n27873 , n27874 , n347908 , n347909 , n347910 , n347911 , n347912 , 
 n27880 , n27881 , n347915 , n347916 , n347917 , n347918 , n347919 , n27887 , n347921 , n347922 , 
 n347923 , n347924 , n347925 , n347926 , n347927 , n347928 , n347929 , n347930 , n347931 , n27899 , 
 n27900 , n27901 , n347935 , n347936 , n347937 , n347938 , n347939 , n27907 , n347941 , n347942 , 
 n347943 , n347944 , n27912 , n347946 , n347947 , n347948 , n347949 , n27917 , n347951 , n347952 , 
 n27920 , n27921 , n27922 , n27923 , n347957 , n347958 , n347959 , n347960 , n347961 , n347962 , 
 n347963 , n347964 , n347965 , n347966 , n27934 , n347968 , n347969 , n347970 , n347971 , n27939 , 
 n347973 , n347974 , n27942 , n27943 , n347977 , n347978 , n347979 , n347980 , n27948 , n27949 , 
 n347983 , n27951 , n347985 , n347986 , n347987 , n347988 , n347989 , n27957 , n347991 , n27959 , 
 n347993 , n347994 , n347995 , n27963 , n347997 , n347998 , n347999 , n348000 , n348001 , n348002 , 
 n27970 , n27971 , n348005 , n27973 , n348007 , n27975 , n348009 , n348010 , n348011 , n348012 , 
 n348013 , n348014 , n348015 , n348016 , n348017 , n348018 , n348019 , n348020 , n27988 , n348022 , 
 n348023 , n348024 , n348025 , n348026 , n348027 , n348028 , n348029 , n27997 , n348031 , n348032 , 
 n348033 , n348034 , n348035 , n348036 , n348037 , n348038 , n28006 , n348040 , n348041 , n348042 , 
 n348043 , n28011 , n28012 , n28013 , n348047 , n348048 , n348049 , n348050 , n348051 , n348052 , 
 n348053 , n348054 , n348055 , n348056 , n28024 , n348058 , n348059 , n28027 , n28028 , n348062 , 
 n28030 , n348064 , n28032 , n348066 , n348067 , n28035 , n28036 , n348070 , n28038 , n348072 , 
 n28040 , n348074 , n348075 , n28043 , n348077 , n348078 , n348079 , n28047 , n348081 , n348082 , 
 n348083 , n28051 , n28052 , n28053 , n28054 , n28055 , n348089 , n348090 , n348091 , n348092 , 
 n348093 , n348094 , n348095 , n348096 , n348097 , n348098 , n348099 , n348100 , n348101 , n348102 , 
 n348103 , n348104 , n348105 , n348106 , n348107 , n348108 , n348109 , n28077 , n28078 , n28079 , 
 n28080 , n348114 , n348115 , n28083 , n348117 , n348118 , n348119 , n348120 , n348121 , n348122 , 
 n348123 , n348124 , n28092 , n348126 , n348127 , n348128 , n28096 , n28097 , n348131 , n28099 , 
 n348133 , n28101 , n348135 , n348136 , n348137 , n348138 , n348139 , n348140 , n28108 , n348142 , 
 n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n348150 , n348151 , n348152 , 
 n348153 , n348154 , n28122 , n348156 , n28124 , n348158 , n348159 , n348160 , n28128 , n28129 , 
 n28130 , n28131 , n348165 , n348166 , n28134 , n348168 , n348169 , n348170 , n348171 , n348172 , 
 n348173 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n348180 , n348181 , n348182 , 
 n28150 , n348184 , n348185 , n348186 , n348187 , n348188 , n348189 , n28157 , n348191 , n348192 , 
 n348193 , n28161 , n28162 , n348196 , n28164 , n348198 , n348199 , n348200 , n28168 , n348202 , 
 n348203 , n348204 , n348205 , n348206 , n28174 , n348208 , n28176 , n348210 , n348211 , n348212 , 
 n348213 , n348214 , n348215 , n348216 , n348217 , n348218 , n28186 , n348220 , n348221 , n28189 , 
 n28190 , n348224 , n348225 , n28193 , n348227 , n348228 , n28196 , n28197 , n348231 , n28199 , 
 n348233 , n348234 , n348235 , n28203 , n348237 , n348238 , n28206 , n28207 , n28208 , n348242 , 
 n28210 , n348244 , n348245 , n28213 , n348247 , n348248 , n28216 , n348250 , n348251 , n348252 , 
 n348253 , n348254 , n348255 , n28223 , n348257 , n348258 , n348259 , n348260 , n28228 , n348262 , 
 n348263 , n348264 , n28232 , n28233 , n28234 , n28235 , n348269 , n28237 , n28238 , n28239 , 
 n28240 , n348274 , n28242 , n348276 , n28244 , n28245 , n348279 , n348280 , n28248 , n348282 , 
 n348283 , n348284 , n348285 , n348286 , n348287 , n348288 , n348289 , n348290 , n28258 , n348292 , 
 n348293 , n348294 , n348295 , n28263 , n348297 , n28265 , n348299 , n348300 , n28268 , n348302 , 
 n348303 , n28271 , n348305 , n28273 , n28274 , n28275 , n348309 , n348310 , n348311 , n348312 , 
 n348313 , n348314 , n348315 , n348316 , n348317 , n348318 , n28286 , n28287 , n348321 , n28289 , 
 n348323 , n348324 , n348325 , n348326 , n348327 , n348328 , n348329 , n28297 , n348331 , n348332 , 
 n348333 , n348334 , n28302 , n28303 , n348337 , n348338 , n28306 , n348340 , n28308 , n348342 , 
 n348343 , n28311 , n348345 , n28313 , n348347 , n348348 , n348349 , n28317 , n348351 , n348352 , 
 n348353 , n348354 , n348355 , n348356 , n28324 , n28325 , n348359 , n348360 , n348361 , n28329 , 
 n348363 , n348364 , n28332 , n348366 , n348367 , n348368 , n348369 , n348370 , n348371 , n348372 , 
 n348373 , n348374 , n28342 , n348376 , n348377 , n348378 , n348379 , n348380 , n348381 , n28349 , 
 n348383 , n28351 , n28352 , n348386 , n348387 , n348388 , n348389 , n348390 , n348391 , n28359 , 
 n348393 , n28361 , n348395 , n28363 , n348397 , n348398 , n28366 , n348400 , n28368 , n348402 , 
 n348403 , n28371 , n348405 , n348406 , n28374 , n348408 , n28376 , n348410 , n348411 , n348412 , 
 n348413 , n348414 , n28382 , n348416 , n28384 , n348418 , n348419 , n28387 , n28388 , n28389 , 
 n348423 , n348424 , n348425 , n348426 , n348427 , n348428 , n348429 , n348430 , n348431 , n348432 , 
 n348433 , n348434 , n348435 , n348436 , n28404 , n348438 , n348439 , n348440 , n348441 , n28409 , 
 n348443 , n348444 , n348445 , n28413 , n348447 , n348448 , n28416 , n348450 , n28418 , n28419 , 
 n348453 , n348454 , n348455 , n28423 , n348457 , n348458 , n348459 , n28427 , n348461 , n28429 , 
 n28430 , n348464 , n28432 , n28433 , n348467 , n348468 , n348469 , n28437 , n348471 , n348472 , 
 n348473 , n348474 , n348475 , n28443 , n28444 , n348478 , n348479 , n348480 , n28448 , n348482 , 
 n348483 , n348484 , n28452 , n348486 , n348487 , n348488 , n348489 , n348490 , n28458 , n28459 , 
 n28460 , n28461 , n348495 , n28463 , n28464 , n348498 , n348499 , n28467 , n348501 , n348502 , 
 n348503 , n348504 , n348505 , n348506 , n348507 , n28475 , n348509 , n28477 , n348511 , n28479 , 
 n348513 , n348514 , n348515 , n348516 , n348517 , n348518 , n348519 , n348520 , n348521 , n28489 , 
 n348523 , n348524 , n28492 , n348526 , n28494 , n28495 , n348529 , n348530 , n28498 , n28499 , 
 n348533 , n28501 , n348535 , n348536 , n348537 , n348538 , n348539 , n28507 , n348541 , n348542 , 
 n348543 , n28511 , n28512 , n348546 , n28514 , n28515 , n348549 , n348550 , n348551 , n348552 , 
 n28520 , n348554 , n28522 , n348556 , n28524 , n348558 , n348559 , n348560 , n348561 , n348562 , 
 n348563 , n348564 , n348565 , n348566 , n348567 , n348568 , n28536 , n348570 , n348571 , n348572 , 
 n28540 , n348574 , n348575 , n348576 , n348577 , n348578 , n28546 , n348580 , n348581 , n28549 , 
 n348583 , n348584 , n28552 , n348586 , n348587 , n28555 , n28556 , n348590 , n348591 , n28559 , 
 n348593 , n348594 , n348595 , n28563 , n348597 , n28565 , n28566 , n348600 , n348601 , n28569 , 
 n28570 , n348604 , n348605 , n348606 , n28574 , n348608 , n348609 , n28577 , n348611 , n28579 , 
 n28580 , n348614 , n348615 , n28583 , n348617 , n348618 , n348619 , n348620 , n348621 , n348622 , 
 n348623 , n348624 , n28592 , n28593 , n348627 , n348628 , n348629 , n348630 , n348631 , n28599 , 
 n348633 , n348634 , n348635 , n348636 , n348637 , n348638 , n348639 , n348640 , n28608 , n28609 , 
 n348643 , n348644 , n348645 , n348646 , n28614 , n348648 , n348649 , n28617 , n348651 , n348652 , 
 n348653 , n348654 , n348655 , n348656 , n28624 , n348658 , n348659 , n348660 , n348661 , n348662 , 
 n348663 , n348664 , n348665 , n28633 , n348667 , n348668 , n348669 , n348670 , n348671 , n348672 , 
 n28640 , n348674 , n28642 , n348676 , n348677 , n28645 , n28646 , n28647 , n28648 , n28649 , 
 n28650 , n348684 , n348685 , n28653 , n348687 , n348688 , n28656 , n348690 , n28658 , n348692 , 
 n348693 , n348694 , n28662 , n28663 , n28664 , n348698 , n348699 , n348700 , n348701 , n348702 , 
 n348703 , n348704 , n348705 , n28673 , n348707 , n348708 , n348709 , n348710 , n348711 , n348712 , 
 n348713 , n348714 , n348715 , n348716 , n348717 , n348718 , n348719 , n348720 , n348721 , n348722 , 
 n28690 , n348724 , n28692 , n28693 , n348727 , n348728 , n28696 , n348730 , n348731 , n28699 , 
 n348733 , n28701 , n348735 , n348736 , n348737 , n348738 , n348739 , n348740 , n348741 , n348742 , 
 n348743 , n348744 , n28712 , n28713 , n348747 , n28715 , n348749 , n28717 , n348751 , n28719 , 
 n28720 , n348754 , n348755 , n28723 , n348757 , n348758 , n28726 , n348760 , n28728 , n28729 , 
 n348763 , n348764 , n348765 , n348766 , n348767 , n348768 , n348769 , n348770 , n348771 , n348772 , 
 n348773 , n348774 , n348775 , n348776 , n348777 , n348778 , n28746 , n348780 , n28748 , n348782 , 
 n348783 , n28751 , n28752 , n348786 , n348787 , n28755 , n28756 , n348790 , n348791 , n348792 , 
 n348793 , n348794 , n348795 , n348796 , n348797 , n348798 , n348799 , n348800 , n348801 , n348802 , 
 n348803 , n348804 , n28772 , n28773 , n348807 , n348808 , n348809 , n348810 , n348811 , n348812 , 
 n348813 , n348814 , n348815 , n348816 , n348817 , n28785 , n28786 , n348820 , n348821 , n28789 , 
 n348823 , n28791 , n28792 , n348826 , n348827 , n348828 , n348829 , n348830 , n28798 , n348832 , 
 n28800 , n348834 , n348835 , n28803 , n348837 , n28805 , n348839 , n28807 , n348841 , n348842 , 
 n348843 , n348844 , n348845 , n348846 , n348847 , n348848 , n28816 , n28817 , n28818 , n28819 , 
 n348853 , n28821 , n348855 , n28823 , n348857 , n348858 , n28826 , n28827 , n348861 , n348862 , 
 n348863 , n348864 , n348865 , n348866 , n348867 , n348868 , n348869 , n348870 , n28838 , n28839 , 
 n348873 , n348874 , n348875 , n348876 , n348877 , n28845 , n348879 , n348880 , n348881 , n28849 , 
 n348883 , n348884 , n28852 , n348886 , n348887 , n28855 , n28856 , n348890 , n28858 , n348892 , 
 n348893 , n28861 , n348895 , n348896 , n28864 , n348898 , n348899 , n28867 , n28868 , n348902 , 
 n348903 , n348904 , n348905 , n348906 , n28874 , n348908 , n348909 , n28877 , n348911 , n348912 , 
 n28880 , n28881 , n348915 , n28883 , n348917 , n348918 , n28886 , n348920 , n348921 , n28889 , 
 n348923 , n348924 , n28892 , n348926 , n348927 , n28895 , n348929 , n348930 , n348931 , n28899 , 
 n348933 , n348934 , n28902 , n348936 , n348937 , n348938 , n348939 , n28907 , n348941 , n348942 , 
 n348943 , n28911 , n348945 , n28913 , n28914 , n28915 , n348949 , n28917 , n348951 , n348952 , 
 n28920 , n348954 , n28922 , n28923 , n348957 , n348958 , n348959 , n348960 , n348961 , n348962 , 
 n28930 , n348964 , n348965 , n28933 , n348967 , n348968 , n28936 , n348970 , n348971 , n348972 , 
 n28940 , n348974 , n348975 , n348976 , n348977 , n348978 , n348979 , n348980 , n348981 , n348982 , 
 n348983 , n348984 , n348985 , n348986 , n348987 , n348988 , n348989 , n28957 , n348991 , n348992 , 
 n348993 , n348994 , n348995 , n348996 , n348997 , n348998 , n348999 , n349000 , n349001 , n349002 , 
 n349003 , n28971 , n349005 , n349006 , n349007 , n349008 , n349009 , n349010 , n349011 , n28979 , 
 n349013 , n349014 , n28982 , n349016 , n349017 , n349018 , n349019 , n28987 , n349021 , n28989 , 
 n349023 , n349024 , n349025 , n349026 , n28994 , n349028 , n28996 , n349030 , n349031 , n28999 , 
 n349033 , n349034 , n29002 , n29003 , n349037 , n29005 , n349039 , n349040 , n29008 , n349042 , 
 n29010 , n349044 , n29012 , n29013 , n349047 , n349048 , n29016 , n349050 , n349051 , n29019 , 
 n349053 , n349054 , n29022 , n29023 , n29024 , n349058 , n349059 , n29027 , n349061 , n349062 , 
 n29030 , n349064 , n349065 , n349066 , n349067 , n349068 , n349069 , n349070 , n349071 , n349072 , 
 n349073 , n349074 , n29042 , n29043 , n349077 , n29045 , n349079 , n349080 , n349081 , n349082 , 
 n349083 , n349084 , n349085 , n29053 , n349087 , n29055 , n349089 , n349090 , n29058 , n349092 , 
 n349093 , n349094 , n349095 , n349096 , n349097 , n349098 , n29066 , n349100 , n349101 , n29069 , 
 n349103 , n349104 , n349105 , n29073 , n349107 , n349108 , n29076 , n349110 , n29078 , n29079 , 
 n29080 , n349114 , n349115 , n349116 , n349117 , n349118 , n349119 , n349120 , n349121 , n29089 , 
 n349123 , n349124 , n349125 , n349126 , n349127 , n349128 , n29096 , n29097 , n349131 , n349132 , 
 n29100 , n349134 , n349135 , n29103 , n29104 , n29105 , n349139 , n29107 , n349141 , n349142 , 
 n349143 , n349144 , n349145 , n29113 , n349147 , n349148 , n349149 , n349150 , n29118 , n349152 , 
 n349153 , n29121 , n349155 , n349156 , n349157 , n349158 , n349159 , n349160 , n349161 , n349162 , 
 n349163 , n29131 , n29132 , n349166 , n349167 , n349168 , n349169 , n349170 , n349171 , n349172 , 
 n349173 , n349174 , n349175 , n349176 , n349177 , n349178 , n349179 , n349180 , n29148 , n349182 , 
 n349183 , n349184 , n349185 , n29153 , n349187 , n349188 , n349189 , n349190 , n349191 , n349192 , 
 n29160 , n29161 , n349195 , n29163 , n349197 , n29165 , n29166 , n349200 , n349201 , n349202 , 
 n349203 , n29171 , n349205 , n349206 , n349207 , n349208 , n349209 , n29177 , n349211 , n349212 , 
 n349213 , n349214 , n349215 , n349216 , n349217 , n349218 , n349219 , n29187 , n349221 , n349222 , 
 n349223 , n349224 , n349225 , n349226 , n349227 , n29195 , n29196 , n349230 , n29198 , n349232 , 
 n29200 , n29201 , n349235 , n349236 , n349237 , n349238 , n349239 , n349240 , n349241 , n349242 , 
 n349243 , n349244 , n29212 , n29213 , n349247 , n349248 , n349249 , n349250 , n349251 , n349252 , 
 n349253 , n349254 , n349255 , n349256 , n349257 , n29225 , n349259 , n29227 , n349261 , n349262 , 
 n349263 , n349264 , n349265 , n349266 , n29234 , n349268 , n349269 , n349270 , n29238 , n349272 , 
 n349273 , n29241 , n349275 , n349276 , n29244 , n349278 , n349279 , n29247 , n349281 , n349282 , 
 n349283 , n349284 , n349285 , n29253 , n349287 , n29255 , n349289 , n349290 , n349291 , n349292 , 
 n29260 , n29261 , n29262 , n349296 , n29264 , n349298 , n349299 , n349300 , n29268 , n349302 , 
 n349303 , n349304 , n29272 , n349306 , n349307 , n349308 , n349309 , n349310 , n29278 , n349312 , 
 n349313 , n349314 , n349315 , n29283 , n349317 , n349318 , n29286 , n29287 , n349321 , n29289 , 
 n29290 , n349324 , n349325 , n29293 , n349327 , n349328 , n349329 , n349330 , n349331 , n349332 , 
 n349333 , n349334 , n349335 , n349336 , n349337 , n349338 , n349339 , n349340 , n29308 , n349342 , 
 n349343 , n349344 , n349345 , n29313 , n29314 , n349348 , n29316 , n29317 , n349351 , n349352 , 
 n29320 , n29321 , n349355 , n349356 , n29324 , n29325 , n349359 , n349360 , n349361 , n29329 , 
 n29330 , n349364 , n349365 , n349366 , n349367 , n349368 , n349369 , n349370 , n349371 , n349372 , 
 n349373 , n349374 , n349375 , n29343 , n29344 , n349378 , n29346 , n29347 , n29348 , n29349 , 
 n349383 , n349384 , n349385 , n349386 , n349387 , n349388 , n349389 , n349390 , n349391 , n29359 , 
 n29360 , n349394 , n29362 , n29363 , n349397 , n349398 , n349399 , n349400 , n29368 , n349402 , 
 n349403 , n29371 , n349405 , n349406 , n349407 , n29375 , n349409 , n349410 , n29378 , n29379 , 
 n349413 , n349414 , n29382 , n349416 , n349417 , n29385 , n349419 , n349420 , n349421 , n29389 , 
 n349423 , n29391 , n349425 , n29393 , n349427 , n29395 , n349429 , n29397 , n29398 , n349432 , 
 n349433 , n29401 , n29402 , n349436 , n349437 , n29405 , n349439 , n349440 , n29408 , n29409 , 
 n349443 , n349444 , n29412 , n29413 , n349447 , n29415 , n29416 , n349450 , n29418 , n29419 , 
 n29420 , n349454 , n349455 , n349456 , n349457 , n349458 , n349459 , n349460 , n349461 , n349462 , 
 n29430 , n349464 , n349465 , n349466 , n29434 , n349468 , n349469 , n349470 , n349471 , n29439 , 
 n349473 , n349474 , n29442 , n349476 , n29444 , n29445 , n29446 , n349480 , n29448 , n349482 , 
 n349483 , n29451 , n349485 , n349486 , n29454 , n349488 , n29456 , n349490 , n29458 , n349492 , 
 n29460 , n29461 , n349495 , n349496 , n349497 , n349498 , n349499 , n349500 , n349501 , n349502 , 
 n29470 , n349504 , n349505 , n349506 , n349507 , n349508 , n349509 , n349510 , n349511 , n349512 , 
 n29480 , n349514 , n349515 , n349516 , n349517 , n349518 , n349519 , n349520 , n29488 , n349522 , 
 n349523 , n29491 , n29492 , n349526 , n29494 , n349528 , n349529 , n29497 , n29498 , n349532 , 
 n349533 , n349534 , n349535 , n349536 , n29504 , n349538 , n349539 , n29507 , n29508 , n349542 , 
 n349543 , n349544 , n349545 , n349546 , n29514 , n349548 , n29516 , n349550 , n349551 , n349552 , 
 n349553 , n29521 , n349555 , n349556 , n29524 , n29525 , n349559 , n29527 , n29528 , n349562 , 
 n349563 , n29531 , n349565 , n349566 , n29534 , n29535 , n29536 , n29537 , n29538 , n349572 , 
 n349573 , n29541 , n349575 , n349576 , n349577 , n349578 , n349579 , n349580 , n349581 , n349582 , 
 n349583 , n29551 , n349585 , n29553 , n29554 , n29555 , n349589 , n349590 , n349591 , n349592 , 
 n349593 , n349594 , n349595 , n349596 , n349597 , n349598 , n349599 , n349600 , n349601 , n29569 , 
 n29570 , n349604 , n349605 , n349606 , n29574 , n29575 , n349609 , n349610 , n349611 , n349612 , 
 n29580 , n349614 , n349615 , n349616 , n349617 , n349618 , n349619 , n29587 , n29588 , n349622 , 
 n29590 , n29591 , n349625 , n349626 , n29594 , n349628 , n349629 , n349630 , n29598 , n349632 , 
 n349633 , n349634 , n29602 , n349636 , n349637 , n29605 , n349639 , n349640 , n349641 , n349642 , 
 n349643 , n349644 , n349645 , n29613 , n349647 , n349648 , n29616 , n349650 , n349651 , n29619 , 
 n349653 , n349654 , n29622 , n29623 , n349657 , n349658 , n349659 , n349660 , n349661 , n349662 , 
 n29630 , n29631 , n349665 , n29633 , n349667 , n349668 , n349669 , n349670 , n29638 , n349672 , 
 n349673 , n349674 , n349675 , n349676 , n349677 , n349678 , n349679 , n349680 , n349681 , n349682 , 
 n349683 , n349684 , n29652 , n349686 , n29654 , n349688 , n349689 , n349690 , n349691 , n29659 , 
 n349693 , n349694 , n349695 , n349696 , n29664 , n349698 , n29666 , n349700 , n349701 , n29669 , 
 n349703 , n349704 , n349705 , n349706 , n349707 , n349708 , n349709 , n29677 , n29678 , n349712 , 
 n349713 , n349714 , n349715 , n349716 , n29684 , n349718 , n349719 , n349720 , n29688 , n349722 , 
 n349723 , n349724 , n349725 , n349726 , n349727 , n349728 , n349729 , n349730 , n349731 , n29699 , 
 n29700 , n29701 , n29702 , n29703 , n29704 , n349738 , n29706 , n349740 , n349741 , n349742 , 
 n349743 , n349744 , n349745 , n349746 , n29714 , n29715 , n349749 , n349750 , n349751 , n29719 , 
 n349753 , n349754 , n349755 , n349756 , n349757 , n349758 , n349759 , n349760 , n349761 , n349762 , 
 n29730 , n29731 , n349765 , n349766 , n349767 , n349768 , n29736 , n349770 , n349771 , n29739 , 
 n29740 , n349774 , n349775 , n29743 , n29744 , n349778 , n349779 , n29747 , n29748 , n349782 , 
 n29750 , n349784 , n349785 , n29753 , n349787 , n29755 , n349789 , n349790 , n29758 , n349792 , 
 n349793 , n349794 , n349795 , n349796 , n349797 , n29765 , n29766 , n29767 , n29768 , n29769 , 
 n29770 , n29771 , n349805 , n29773 , n349807 , n29775 , n29776 , n349810 , n29778 , n349812 , 
 n349813 , n349814 , n349815 , n29783 , n29784 , n349818 , n29786 , n349820 , n349821 , n349822 , 
 n29790 , n349824 , n349825 , n349826 , n349827 , n349828 , n349829 , n349830 , n349831 , n349832 , 
 n349833 , n349834 , n349835 , n349836 , n349837 , n349838 , n29806 , n349840 , n349841 , n349842 , 
 n349843 , n29811 , n29812 , n349846 , n29814 , n349848 , n29816 , n349850 , n349851 , n349852 , 
 n349853 , n349854 , n349855 , n349856 , n349857 , n349858 , n349859 , n349860 , n349861 , n349862 , 
 n349863 , n349864 , n349865 , n349866 , n349867 , n349868 , n29836 , n349870 , n349871 , n349872 , 
 n29840 , n349874 , n349875 , n29843 , n349877 , n349878 , n349879 , n349880 , n349881 , n29849 , 
 n349883 , n349884 , n349885 , n29853 , n349887 , n349888 , n349889 , n349890 , n349891 , n29859 , 
 n349893 , n349894 , n349895 , n29863 , n349897 , n349898 , n349899 , n349900 , n349901 , n349902 , 
 n29870 , n349904 , n349905 , n349906 , n29874 , n349908 , n29876 , n29877 , n29878 , n349912 , 
 n29880 , n29881 , n349915 , n29883 , n29884 , n349918 , n29886 , n349920 , n349921 , n349922 , 
 n349923 , n349924 , n349925 , n349926 , n349927 , n349928 , n349929 , n29897 , n349931 , n29899 , 
 n29900 , n349934 , n349935 , n29903 , n349937 , n349938 , n29906 , n349940 , n349941 , n29909 , 
 n349943 , n349944 , n349945 , n29913 , n349947 , n349948 , n349949 , n349950 , n349951 , n349952 , 
 n349953 , n349954 , n349955 , n349956 , n349957 , n29925 , n349959 , n349960 , n349961 , n349962 , 
 n349963 , n349964 , n349965 , n349966 , n349967 , n29935 , n349969 , n349970 , n349971 , n349972 , 
 n29940 , n349974 , n29942 , n349976 , n349977 , n29945 , n349979 , n29947 , n29948 , n29949 , 
 n349983 , n29951 , n349985 , n349986 , n349987 , n349988 , n349989 , n349990 , n349991 , n349992 , 
 n349993 , n349994 , n349995 , n29963 , n349997 , n29965 , n349999 , n29967 , n350001 , n350002 , 
 n29970 , n350004 , n350005 , n350006 , n350007 , n350008 , n29976 , n350010 , n350011 , n29979 , 
 n350013 , n350014 , n29982 , n350016 , n350017 , n350018 , n350019 , n350020 , n350021 , n350022 , 
 n29990 , n350024 , n350025 , n350026 , n350027 , n350028 , n350029 , n29997 , n350031 , n29999 , 
 n350033 , n350034 , n30002 , n350036 , n350037 , n350038 , n30006 , n350040 , n30008 , n350042 , 
 n30010 , n350044 , n350045 , n30013 , n350047 , n350048 , n30016 , n30017 , n30018 , n30019 , 
 n30020 , n350054 , n350055 , n30023 , n350057 , n350058 , n350059 , n350060 , n30028 , n350062 , 
 n350063 , n30031 , n350065 , n350066 , n30034 , n30035 , n350069 , n350070 , n350071 , n30039 , 
 n350073 , n350074 , n350075 , n350076 , n350077 , n350078 , n350079 , n350080 , n350081 , n350082 , 
 n350083 , n350084 , n350085 , n350086 , n30054 , n350088 , n350089 , n30057 , n350091 , n350092 , 
 n30060 , n350094 , n350095 , n30063 , n30064 , n350098 , n350099 , n350100 , n350101 , n350102 , 
 n350103 , n350104 , n350105 , n350106 , n350107 , n30075 , n350109 , n350110 , n350111 , n350112 , 
 n350113 , n350114 , n350115 , n350116 , n350117 , n350118 , n350119 , n30087 , n30088 , n30089 , 
 n30090 , n350124 , n350125 , n350126 , n350127 , n30095 , n350129 , n30097 , n350131 , n350132 , 
 n350133 , n350134 , n350135 , n350136 , n350137 , n350138 , n350139 , n350140 , n350141 , n30109 , 
 n30110 , n30111 , n350145 , n350146 , n350147 , n350148 , n350149 , n350150 , n350151 , n350152 , 
 n30120 , n30121 , n350155 , n350156 , n350157 , n350158 , n350159 , n30127 , n350161 , n350162 , 
 n30130 , n350164 , n350165 , n30133 , n350167 , n30135 , n30136 , n30137 , n350171 , n30139 , 
 n30140 , n350174 , n350175 , n30143 , n350177 , n350178 , n350179 , n350180 , n350181 , n350182 , 
 n30150 , n350184 , n350185 , n30153 , n350187 , n350188 , n350189 , n350190 , n350191 , n30159 , 
 n350193 , n30161 , n30162 , n350196 , n30164 , n350198 , n30166 , n350200 , n350201 , n30169 , 
 n350203 , n350204 , n350205 , n350206 , n350207 , n350208 , n350209 , n350210 , n350211 , n350212 , 
 n350213 , n350214 , n350215 , n30183 , n30184 , n350218 , n350219 , n30187 , n350221 , n350222 , 
 n30190 , n350224 , n350225 , n30193 , n350227 , n350228 , n350229 , n30197 , n30198 , n30199 , 
 n350233 , n350234 , n350235 , n350236 , n350237 , n30205 , n350239 , n350240 , n30208 , n350242 , 
 n350243 , n30211 , n350245 , n350246 , n350247 , n350248 , n350249 , n350250 , n350251 , n350252 , 
 n350253 , n30221 , n350255 , n350256 , n30224 , n350258 , n350259 , n350260 , n350261 , n30229 , 
 n350263 , n350264 , n350265 , n350266 , n350267 , n350268 , n350269 , n350270 , n30238 , n350272 , 
 n350273 , n350274 , n350275 , n350276 , n350277 , n350278 , n350279 , n350280 , n350281 , n350282 , 
 n350283 , n350284 , n350285 , n350286 , n30254 , n350288 , n30256 , n30257 , n30258 , n350292 , 
 n30260 , n350294 , n350295 , n350296 , n30264 , n350298 , n350299 , n30267 , n350301 , n350302 , 
 n30270 , n350304 , n350305 , n350306 , n350307 , n350308 , n30276 , n350310 , n350311 , n30279 , 
 n30280 , n350314 , n350315 , n350316 , n30284 , n30285 , n350319 , n350320 , n350321 , n350322 , 
 n350323 , n350324 , n350325 , n350326 , n30294 , n350328 , n350329 , n350330 , n30298 , n350332 , 
 n350333 , n350334 , n350335 , n350336 , n30304 , n30305 , n30306 , n350340 , n30308 , n30309 , 
 n350343 , n350344 , n350345 , n350346 , n30314 , n30315 , n30316 , n30317 , n30318 , n350352 , 
 n350353 , n350354 , n350355 , n350356 , n350357 , n350358 , n350359 , n350360 , n30328 , n350362 , 
 n350363 , n30331 , n350365 , n350366 , n350367 , n350368 , n30336 , n350370 , n350371 , n350372 , 
 n350373 , n350374 , n30342 , n350376 , n350377 , n30345 , n350379 , n350380 , n350381 , n350382 , 
 n350383 , n350384 , n350385 , n350386 , n350387 , n30355 , n30356 , n30357 , n30358 , n350392 , 
 n350393 , n30361 , n350395 , n350396 , n350397 , n30365 , n350399 , n350400 , n350401 , n30369 , 
 n350403 , n350404 , n350405 , n30373 , n350407 , n350408 , n350409 , n30377 , n350411 , n350412 , 
 n350413 , n350414 , n350415 , n350416 , n350417 , n350418 , n350419 , n350420 , n350421 , n350422 , 
 n350423 , n350424 , n350425 , n350426 , n350427 , n30395 , n30396 , n350430 , n350431 , n350432 , 
 n350433 , n350434 , n30402 , n350436 , n350437 , n350438 , n350439 , n350440 , n350441 , n350442 , 
 n350443 , n350444 , n350445 , n350446 , n30414 , n350448 , n350449 , n30417 , n30418 , n350452 , 
 n350453 , n350454 , n350455 , n30423 , n350457 , n350458 , n350459 , n350460 , n350461 , n350462 , 
 n350463 , n30431 , n30432 , n30433 , n350467 , n350468 , n350469 , n350470 , n350471 , n30439 , 
 n30440 , n350474 , n350475 , n350476 , n350477 , n350478 , n30446 , n30447 , n350481 , n30449 , 
 n30450 , n350484 , n350485 , n350486 , n30454 , n30455 , n350489 , n30457 , n350491 , n30459 , 
 n350493 , n350494 , n30462 , n350496 , n350497 , n350498 , n350499 , n350500 , n350501 , n350502 , 
 n350503 , n350504 , n30472 , n350506 , n30474 , n350508 , n350509 , n30477 , n30478 , n350512 , 
 n350513 , n30481 , n350515 , n350516 , n350517 , n350518 , n350519 , n350520 , n350521 , n30489 , 
 n350523 , n350524 , n350525 , n350526 , n30494 , n350528 , n350529 , n350530 , n350531 , n350532 , 
 n350533 , n350534 , n30502 , n30503 , n350537 , n350538 , n30506 , n350540 , n350541 , n30509 , 
 n30510 , n350544 , n30512 , n350546 , n350547 , n30515 , n350549 , n30517 , n30518 , n30519 , 
 n30520 , n30521 , n30522 , n350556 , n30524 , n350558 , n350559 , n350560 , n30528 , n350562 , 
 n350563 , n350564 , n350565 , n350566 , n30534 , n350568 , n350569 , n350570 , n350571 , n30539 , 
 n350573 , n350574 , n350575 , n350576 , n350577 , n30545 , n350579 , n30547 , n350581 , n350582 , 
 n350583 , n350584 , n350585 , n350586 , n350587 , n350588 , n350589 , n30557 , n350591 , n30559 , 
 n350593 , n30561 , n350595 , n350596 , n30564 , n350598 , n30566 , n350600 , n30568 , n350602 , 
 n350603 , n350604 , n350605 , n350606 , n30574 , n350608 , n30576 , n350610 , n350611 , n350612 , 
 n350613 , n30581 , n30582 , n350616 , n30584 , n350618 , n350619 , n350620 , n350621 , n350622 , 
 n350623 , n350624 , n350625 , n350626 , n350627 , n30595 , n350629 , n30597 , n350631 , n350632 , 
 n350633 , n350634 , n350635 , n350636 , n350637 , n350638 , n350639 , n350640 , n350641 , n350642 , 
 n30610 , n30611 , n350645 , n30613 , n350647 , n30615 , n30616 , n350650 , n350651 , n30619 , 
 n350653 , n350654 , n30622 , n350656 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , 
 n30630 , n30631 , n350665 , n350666 , n350667 , n350668 , n30636 , n30637 , n350671 , n350672 , 
 n30640 , n350674 , n350675 , n30643 , n30644 , n350678 , n30646 , n350680 , n350681 , n350682 , 
 n350683 , n30651 , n350685 , n350686 , n30654 , n30655 , n350689 , n30657 , n350691 , n30659 , 
 n30660 , n350694 , n350695 , n350696 , n350697 , n350698 , n30666 , n350700 , n30668 , n350702 , 
 n30670 , n350704 , n30672 , n350706 , n350707 , n30675 , n350709 , n30677 , n350711 , n350712 , 
 n30680 , n350714 , n30682 , n350716 , n350717 , n350718 , n350719 , n350720 , n350721 , n350722 , 
 n350723 , n350724 , n350725 , n350726 , n350727 , n30695 , n350729 , n350730 , n350731 , n350732 , 
 n350733 , n30701 , n30702 , n350736 , n30704 , n350738 , n350739 , n30707 , n350741 , n350742 , 
 n30710 , n350744 , n350745 , n350746 , n350747 , n350748 , n350749 , n350750 , n350751 , n350752 , 
 n30720 , n350754 , n350755 , n350756 , n350757 , n350758 , n30726 , n350760 , n30728 , n350762 , 
 n350763 , n350764 , n350765 , n350766 , n30734 , n350768 , n350769 , n350770 , n30738 , n350772 , 
 n350773 , n350774 , n30742 , n30743 , n350777 , n350778 , n350779 , n30747 , n350781 , n350782 , 
 n350783 , n30751 , n30752 , n350786 , n350787 , n350788 , n350789 , n350790 , n350791 , n350792 , 
 n350793 , n30761 , n30762 , n350796 , n350797 , n30765 , n350799 , n350800 , n30768 , n350802 , 
 n350803 , n350804 , n350805 , n350806 , n350807 , n350808 , n350809 , n350810 , n350811 , n30779 , 
 n350813 , n350814 , n350815 , n350816 , n350817 , n350818 , n350819 , n350820 , n350821 , n350822 , 
 n350823 , n350824 , n350825 , n350826 , n350827 , n350828 , n30796 , n350830 , n350831 , n350832 , 
 n30800 , n350834 , n30802 , n30803 , n350837 , n350838 , n30806 , n350840 , n350841 , n30809 , 
 n350843 , n350844 , n30812 , n30813 , n350847 , n350848 , n30816 , n350850 , n350851 , n30819 , 
 n30820 , n350854 , n30822 , n350856 , n350857 , n350858 , n350859 , n30827 , n350861 , n30829 , 
 n350863 , n30831 , n30832 , n350866 , n30834 , n350868 , n30836 , n350870 , n350871 , n350872 , 
 n30840 , n350874 , n350875 , n30843 , n350877 , n350878 , n350879 , n30847 , n350881 , n350882 , 
 n30850 , n350884 , n350885 , n350886 , n30854 , n350888 , n350889 , n30857 , n350891 , n350892 , 
 n350893 , n350894 , n350895 , n350896 , n350897 , n30865 , n30866 , n350900 , n350901 , n350902 , 
 n350903 , n350904 , n30872 , n30873 , n350907 , n30875 , n350909 , n30877 , n30878 , n350912 , 
 n350913 , n350914 , n350915 , n350916 , n30884 , n350918 , n350919 , n350920 , n350921 , n350922 , 
 n350923 , n30891 , n30892 , n350926 , n350927 , n30895 , n350929 , n350930 , n350931 , n350932 , 
 n30900 , n350934 , n350935 , n350936 , n350937 , n30905 , n30906 , n350940 , n350941 , n30909 , 
 n350943 , n30911 , n30912 , n350946 , n350947 , n350948 , n350949 , n30917 , n350951 , n350952 , 
 n30920 , n350954 , n350955 , n350956 , n30924 , n350958 , n30926 , n30927 , n350961 , n350962 , 
 n30930 , n30931 , n350965 , n30933 , n30934 , n350968 , n350969 , n30937 , n350971 , n350972 , 
 n350973 , n350974 , n350975 , n350976 , n30944 , n350978 , n350979 , n350980 , n350981 , n30949 , 
 n350983 , n30951 , n350985 , n30953 , n350987 , n350988 , n350989 , n350990 , n350991 , n350992 , 
 n30960 , n350994 , n350995 , n30963 , n350997 , n350998 , n350999 , n351000 , n351001 , n351002 , 
 n30970 , n351004 , n351005 , n351006 , n351007 , n30975 , n351009 , n351010 , n30978 , n30979 , 
 n351013 , n30981 , n30982 , n30983 , n351017 , n351018 , n351019 , n30987 , n30988 , n351022 , 
 n351023 , n351024 , n351025 , n30993 , n351027 , n351028 , n351029 , n30997 , n351031 , n351032 , 
 n31000 , n351034 , n31002 , n351036 , n351037 , n351038 , n351039 , n351040 , n31008 , n31009 , 
 n351043 , n351044 , n351045 , n351046 , n351047 , n351048 , n351049 , n351050 , n351051 , n351052 , 
 n351053 , n351054 , n351055 , n351056 , n31024 , n31025 , n351059 , n351060 , n31028 , n351062 , 
 n351063 , n351064 , n351065 , n351066 , n351067 , n31035 , n351069 , n351070 , n31038 , n351072 , 
 n351073 , n351074 , n351075 , n351076 , n351077 , n351078 , n351079 , n351080 , n351081 , n31049 , 
 n351083 , n31051 , n351085 , n31053 , n31054 , n351088 , n351089 , n31057 , n31058 , n351092 , 
 n351093 , n351094 , n351095 , n351096 , n351097 , n351098 , n351099 , n351100 , n31068 , n351102 , 
 n351103 , n31071 , n31072 , n31073 , n351107 , n351108 , n31076 , n31077 , n351111 , n351112 , 
 n351113 , n31081 , n31082 , n351116 , n351117 , n351118 , n351119 , n351120 , n31088 , n351122 , 
 n351123 , n31091 , n351125 , n31093 , n351127 , n31095 , n31096 , n351130 , n31098 , n351132 , 
 n351133 , n31101 , n351135 , n351136 , n31104 , n351138 , n31106 , n351140 , n31108 , n351142 , 
 n351143 , n351144 , n351145 , n351146 , n31114 , n351148 , n351149 , n351150 , n351151 , n351152 , 
 n351153 , n351154 , n351155 , n351156 , n31124 , n351158 , n31126 , n351160 , n351161 , n351162 , 
 n31130 , n351164 , n351165 , n31133 , n351167 , n351168 , n351169 , n351170 , n351171 , n351172 , 
 n351173 , n351174 , n351175 , n351176 , n31144 , n351178 , n351179 , n351180 , n31148 , n351182 , 
 n351183 , n31151 , n31152 , n351186 , n351187 , n351188 , n351189 , n351190 , n351191 , n351192 , 
 n351193 , n351194 , n351195 , n351196 , n31164 , n31165 , n351199 , n31167 , n31168 , n31169 , 
 n31170 , n351204 , n351205 , n351206 , n351207 , n351208 , n31176 , n351210 , n31178 , n31179 , 
 n31180 , n351214 , n351215 , n351216 , n31184 , n351218 , n351219 , n31187 , n351221 , n31189 , 
 n351223 , n351224 , n31192 , n31193 , n31194 , n351228 , n351229 , n31197 , n351231 , n31199 , 
 n351233 , n351234 , n31202 , n351236 , n31204 , n31205 , n351239 , n351240 , n351241 , n351242 , 
 n31210 , n351244 , n351245 , n31213 , n351247 , n351248 , n31216 , n351250 , n351251 , n31219 , 
 n351253 , n351254 , n351255 , n351256 , n351257 , n31225 , n351259 , n351260 , n31228 , n351262 , 
 n31230 , n31231 , n351265 , n351266 , n351267 , n351268 , n351269 , n351270 , n31238 , n351272 , 
 n351273 , n351274 , n351275 , n351276 , n351277 , n31245 , n351279 , n351280 , n31248 , n31249 , 
 n31250 , n351284 , n31252 , n31253 , n351287 , n351288 , n31256 , n351290 , n351291 , n351292 , 
 n31260 , n351294 , n351295 , n351296 , n351297 , n351298 , n31266 , n351300 , n31268 , n351302 , 
 n351303 , n351304 , n351305 , n31273 , n351307 , n351308 , n31276 , n351310 , n351311 , n31279 , 
 n31280 , n351314 , n351315 , n31283 , n351317 , n351318 , n31286 , n351320 , n31288 , n31289 , 
 n351323 , n351324 , n31292 , n351326 , n351327 , n31295 , n351329 , n351330 , n351331 , n351332 , 
 n351333 , n351334 , n351335 , n351336 , n351337 , n31305 , n351339 , n351340 , n31308 , n351342 , 
 n351343 , n31311 , n351345 , n351346 , n31314 , n351348 , n351349 , n351350 , n31318 , n351352 , 
 n31320 , n351354 , n351355 , n351356 , n351357 , n31325 , n31326 , n351360 , n351361 , n31329 , 
 n351363 , n351364 , n351365 , n351366 , n351367 , n351368 , n31336 , n351370 , n351371 , n31339 , 
 n351373 , n351374 , n351375 , n351376 , n351377 , n351378 , n31346 , n351380 , n351381 , n351382 , 
 n351383 , n351384 , n31352 , n351386 , n351387 , n351388 , n351389 , n31357 , n351391 , n351392 , 
 n351393 , n351394 , n351395 , n31363 , n351397 , n31365 , n31366 , n351400 , n351401 , n351402 , 
 n351403 , n351404 , n351405 , n351406 , n351407 , n351408 , n31376 , n351410 , n351411 , n351412 , 
 n31380 , n351414 , n351415 , n31383 , n351417 , n351418 , n31386 , n351420 , n31388 , n351422 , 
 n31390 , n351424 , n351425 , n31393 , n351427 , n351428 , n351429 , n31397 , n351431 , n351432 , 
 n351433 , n351434 , n351435 , n31403 , n351437 , n351438 , n351439 , n351440 , n351441 , n351442 , 
 n31410 , n351444 , n351445 , n31413 , n351447 , n351448 , n351449 , n351450 , n351451 , n31419 , 
 n351453 , n351454 , n351455 , n351456 , n351457 , n351458 , n351459 , n351460 , n351461 , n31429 , 
 n351463 , n351464 , n351465 , n31433 , n31434 , n351468 , n31436 , n351470 , n351471 , n31439 , 
 n351473 , n351474 , n351475 , n31443 , n31444 , n31445 , n351479 , n351480 , n351481 , n351482 , 
 n31450 , n351484 , n351485 , n31453 , n351487 , n351488 , n31456 , n31457 , n351491 , n31459 , 
 n351493 , n351494 , n351495 , n31463 , n351497 , n351498 , n351499 , n351500 , n351501 , n31469 , 
 n351503 , n351504 , n31472 , n351506 , n351507 , n351508 , n31476 , n351510 , n351511 , n351512 , 
 n351513 , n351514 , n31482 , n351516 , n351517 , n31485 , n351519 , n351520 , n351521 , n31489 , 
 n351523 , n351524 , n351525 , n31493 , n31494 , n351528 , n351529 , n31497 , n31498 , n31499 , 
 n351533 , n351534 , n31502 , n351536 , n351537 , n31505 , n351539 , n31507 , n351541 , n31509 , 
 n351543 , n351544 , n351545 , n351546 , n351547 , n351548 , n351549 , n351550 , n351551 , n31519 , 
 n31520 , n351554 , n351555 , n31523 , n351557 , n351558 , n351559 , n351560 , n351561 , n31529 , 
 n351563 , n351564 , n31532 , n351566 , n31534 , n351568 , n31536 , n351570 , n351571 , n31539 , 
 n351573 , n351574 , n31542 , n31543 , n351577 , n351578 , n351579 , n351580 , n31548 , n31549 , 
 n351583 , n31551 , n31552 , n31553 , n31554 , n351588 , n351589 , n351590 , n351591 , n351592 , 
 n31560 , n31561 , n351595 , n31563 , n31564 , n31565 , n351599 , n351600 , n351601 , n31569 , 
 n31570 , n351604 , n31572 , n351606 , n351607 , n31575 , n351609 , n351610 , n31578 , n31579 , 
 n351613 , n31581 , n351615 , n351616 , n351617 , n351618 , n351619 , n351620 , n31588 , n351622 , 
 n351623 , n351624 , n351625 , n31593 , n351627 , n31595 , n351629 , n351630 , n31598 , n31599 , 
 n351633 , n351634 , n351635 , n351636 , n351637 , n351638 , n351639 , n351640 , n31608 , n351642 , 
 n351643 , n31611 , n351645 , n351646 , n351647 , n351648 , n351649 , n351650 , n31618 , n31619 , 
 n351653 , n351654 , n351655 , n31623 , n351657 , n351658 , n351659 , n351660 , n351661 , n351662 , 
 n31630 , n31631 , n351665 , n351666 , n351667 , n351668 , n31636 , n351670 , n351671 , n351672 , 
 n31640 , n351674 , n351675 , n351676 , n351677 , n351678 , n351679 , n31647 , n351681 , n351682 , 
 n351683 , n31651 , n351685 , n351686 , n31654 , n351688 , n351689 , n351690 , n351691 , n351692 , 
 n351693 , n31661 , n351695 , n31663 , n351697 , n351698 , n351699 , n351700 , n351701 , n351702 , 
 n351703 , n351704 , n31672 , n351706 , n351707 , n351708 , n351709 , n351710 , n351711 , n31679 , 
 n351713 , n351714 , n31682 , n351716 , n351717 , n31685 , n351719 , n31687 , n351721 , n31689 , 
 n351723 , n351724 , n351725 , n351726 , n351727 , n31695 , n31696 , n351730 , n351731 , n351732 , 
 n351733 , n31701 , n351735 , n351736 , n351737 , n351738 , n351739 , n351740 , n31708 , n351742 , 
 n351743 , n351744 , n31712 , n351746 , n31714 , n351748 , n351749 , n351750 , n351751 , n351752 , 
 n351753 , n351754 , n31722 , n351756 , n351757 , n31725 , n31726 , n351760 , n31728 , n351762 , 
 n31730 , n351764 , n351765 , n31733 , n351767 , n31735 , n351769 , n351770 , n351771 , n351772 , 
 n351773 , n351774 , n31742 , n351776 , n351777 , n31745 , n351779 , n351780 , n351781 , n31749 , 
 n351783 , n31751 , n31752 , n31753 , n351787 , n31755 , n351789 , n31757 , n351791 , n351792 , 
 n31760 , n351794 , n31762 , n351796 , n351797 , n351798 , n31766 , n351800 , n351801 , n351802 , 
 n351803 , n31771 , n31772 , n351806 , n351807 , n31775 , n351809 , n31777 , n351811 , n31779 , 
 n351813 , n31781 , n351815 , n351816 , n351817 , n31785 , n351819 , n351820 , n351821 , n351822 , 
 n351823 , n351824 , n31792 , n351826 , n351827 , n31795 , n351829 , n351830 , n351831 , n31799 , 
 n351833 , n351834 , n31802 , n351836 , n351837 , n351838 , n31806 , n31807 , n31808 , n31809 , 
 n31810 , n31811 , n351845 , n351846 , n31814 , n351848 , n351849 , n351850 , n351851 , n351852 , 
 n351853 , n31821 , n351855 , n351856 , n31824 , n351858 , n351859 , n351860 , n351861 , n31829 , 
 n31830 , n31831 , n351865 , n351866 , n31834 , n31835 , n31836 , n351870 , n351871 , n351872 , 
 n351873 , n31841 , n351875 , n351876 , n31844 , n351878 , n31846 , n31847 , n351881 , n351882 , 
 n351883 , n31851 , n31852 , n351886 , n351887 , n351888 , n31856 , n31857 , n351891 , n351892 , 
 n351893 , n31861 , n351895 , n31863 , n351897 , n351898 , n31866 , n351900 , n31868 , n31869 , 
 n351903 , n31871 , n351905 , n31873 , n351907 , n351908 , n351909 , n351910 , n351911 , n31879 , 
 n351913 , n351914 , n351915 , n351916 , n351917 , n31885 , n351919 , n31887 , n351921 , n351922 , 
 n351923 , n351924 , n351925 , n351926 , n351927 , n351928 , n351929 , n351930 , n31898 , n351932 , 
 n351933 , n351934 , n351935 , n351936 , n31904 , n351938 , n351939 , n351940 , n351941 , n351942 , 
 n351943 , n31911 , n351945 , n351946 , n31914 , n31915 , n351949 , n351950 , n351951 , n351952 , 
 n351953 , n351954 , n351955 , n351956 , n351957 , n351958 , n31926 , n351960 , n31928 , n31929 , 
 n351963 , n31931 , n351965 , n31933 , n351967 , n351968 , n351969 , n31937 , n351971 , n351972 , 
 n31940 , n351974 , n31942 , n351976 , n351977 , n351978 , n351979 , n351980 , n351981 , n351982 , 
 n351983 , n351984 , n351985 , n31953 , n351987 , n351988 , n31956 , n351990 , n351991 , n351992 , 
 n351993 , n351994 , n351995 , n351996 , n351997 , n351998 , n351999 , n352000 , n31968 , n352002 , 
 n352003 , n31971 , n352005 , n352006 , n352007 , n352008 , n352009 , n352010 , n352011 , n352012 , 
 n352013 , n352014 , n352015 , n352016 , n352017 , n31985 , n352019 , n352020 , n352021 , n31989 , 
 n31990 , n31991 , n352025 , n352026 , n31994 , n31995 , n31996 , n352030 , n352031 , n31999 , 
 n32000 , n352034 , n32002 , n352036 , n32004 , n32005 , n352039 , n352040 , n352041 , n352042 , 
 n352043 , n352044 , n352045 , n32013 , n352047 , n32015 , n352049 , n32017 , n352051 , n352052 , 
 n32020 , n352054 , n352055 , n32023 , n352057 , n352058 , n352059 , n352060 , n352061 , n352062 , 
 n32030 , n352064 , n352065 , n32033 , n352067 , n352068 , n352069 , n352070 , n32038 , n352072 , 
 n352073 , n32041 , n32042 , n32043 , n352077 , n352078 , n32046 , n352080 , n352081 , n352082 , 
 n352083 , n352084 , n352085 , n352086 , n352087 , n32055 , n352089 , n352090 , n352091 , n352092 , 
 n32060 , n352094 , n352095 , n352096 , n352097 , n32065 , n352099 , n352100 , n352101 , n32069 , 
 n352103 , n352104 , n352105 , n32073 , n32074 , n32075 , n352109 , n352110 , n32078 , n32079 , 
 n32080 , n352114 , n32082 , n32083 , n32084 , n32085 , n352119 , n32087 , n32088 , n352122 , 
 n352123 , n352124 , n352125 , n352126 , n352127 , n352128 , n352129 , n352130 , n352131 , n32099 , 
 n352133 , n352134 , n352135 , n352136 , n32104 , n352138 , n352139 , n32107 , n352141 , n32109 , 
 n352143 , n32111 , n352145 , n352146 , n352147 , n352148 , n352149 , n352150 , n352151 , n352152 , 
 n352153 , n352154 , n352155 , n352156 , n352157 , n352158 , n352159 , n352160 , n352161 , n352162 , 
 n352163 , n352164 , n352165 , n352166 , n352167 , n352168 , n32136 , n352170 , n32138 , n352172 , 
 n352173 , n352174 , n352175 , n352176 , n352177 , n352178 , n352179 , n352180 , n32148 , n352182 , 
 n352183 , n32151 , n352185 , n32153 , n32154 , n352188 , n352189 , n32157 , n352191 , n352192 , 
 n32160 , n352194 , n352195 , n352196 , n32164 , n352198 , n352199 , n352200 , n352201 , n352202 , 
 n352203 , n352204 , n352205 , n32173 , n32174 , n32175 , n352209 , n352210 , n352211 , n352212 , 
 n352213 , n352214 , n352215 , n32183 , n352217 , n352218 , n352219 , n32187 , n352221 , n352222 , 
 n32190 , n352224 , n32192 , n352226 , n352227 , n352228 , n352229 , n32197 , n32198 , n32199 , 
 n352233 , n352234 , n32202 , n352236 , n32204 , n32205 , n32206 , n32207 , n32208 , n352242 , 
 n32210 , n352244 , n352245 , n32213 , n32214 , n32215 , n32216 , n352250 , n352251 , n32219 , 
 n352253 , n352254 , n32222 , n32223 , n32224 , n352258 , n352259 , n32227 , n352261 , n32229 , 
 n352263 , n352264 , n32232 , n352266 , n32234 , n352268 , n352269 , n352270 , n352271 , n352272 , 
 n352273 , n352274 , n352275 , n352276 , n352277 , n352278 , n352279 , n352280 , n352281 , n352282 , 
 n352283 , n352284 , n32252 , n352286 , n352287 , n352288 , n352289 , n32257 , n32258 , n352292 , 
 n352293 , n352294 , n32262 , n352296 , n352297 , n352298 , n352299 , n352300 , n352301 , n32269 , 
 n32270 , n352304 , n352305 , n352306 , n352307 , n352308 , n352309 , n352310 , n352311 , n32279 , 
 n352313 , n352314 , n352315 , n32283 , n32284 , n352318 , n352319 , n352320 , n352321 , n352322 , 
 n352323 , n32291 , n352325 , n352326 , n352327 , n352328 , n352329 , n352330 , n32298 , n352332 , 
 n352333 , n32301 , n352335 , n32303 , n352337 , n352338 , n32306 , n352340 , n32308 , n352342 , 
 n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n352349 , n352350 , n32318 , n352352 , 
 n352353 , n352354 , n32322 , n352356 , n352357 , n352358 , n352359 , n352360 , n352361 , n352362 , 
 n352363 , n352364 , n352365 , n352366 , n32334 , n352368 , n352369 , n32337 , n352371 , n352372 , 
 n352373 , n352374 , n352375 , n352376 , n32344 , n352378 , n352379 , n352380 , n352381 , n352382 , 
 n32350 , n32351 , n352385 , n352386 , n352387 , n32355 , n32356 , n32357 , n32358 , n352392 , 
 n352393 , n352394 , n352395 , n352396 , n352397 , n352398 , n352399 , n32367 , n352401 , n352402 , 
 n32370 , n352404 , n352405 , n352406 , n32374 , n32375 , n352409 , n352410 , n32378 , n352412 , 
 n352413 , n32381 , n352415 , n352416 , n32384 , n352418 , n352419 , n352420 , n352421 , n32389 , 
 n352423 , n352424 , n32392 , n352426 , n352427 , n352428 , n352429 , n352430 , n352431 , n32399 , 
 n352433 , n352434 , n352435 , n32403 , n32404 , n352438 , n352439 , n352440 , n32408 , n352442 , 
 n32410 , n352444 , n352445 , n32413 , n352447 , n352448 , n352449 , n32417 , n352451 , n352452 , 
 n32420 , n352454 , n352455 , n32423 , n352457 , n352458 , n352459 , n352460 , n352461 , n352462 , 
 n352463 , n32431 , n352465 , n352466 , n352467 , n352468 , n32436 , n352470 , n352471 , n352472 , 
 n352473 , n32441 , n352475 , n352476 , n32444 , n32445 , n352479 , n352480 , n352481 , n352482 , 
 n352483 , n352484 , n352485 , n352486 , n352487 , n352488 , n352489 , n352490 , n352491 , n352492 , 
 n352493 , n32461 , n32462 , n352496 , n352497 , n352498 , n352499 , n352500 , n32468 , n352502 , 
 n352503 , n352504 , n32472 , n32473 , n352507 , n352508 , n352509 , n352510 , n352511 , n32479 , 
 n352513 , n352514 , n352515 , n352516 , n352517 , n352518 , n352519 , n352520 , n352521 , n352522 , 
 n32490 , n352524 , n352525 , n352526 , n32494 , n352528 , n352529 , n32497 , n352531 , n352532 , 
 n352533 , n352534 , n352535 , n352536 , n352537 , n352538 , n352539 , n352540 , n352541 , n32509 , 
 n352543 , n352544 , n32512 , n32513 , n352547 , n352548 , n352549 , n352550 , n352551 , n32519 , 
 n352553 , n352554 , n352555 , n352556 , n32524 , n352558 , n32526 , n32527 , n32528 , n32529 , 
 n32530 , n352564 , n32532 , n32533 , n32534 , n352568 , n352569 , n352570 , n352571 , n32539 , 
 n352573 , n352574 , n352575 , n352576 , n352577 , n32545 , n352579 , n352580 , n32548 , n32549 , 
 n32550 , n352584 , n352585 , n32553 , n32554 , n32555 , n352589 , n352590 , n32558 , n32559 , 
 n352593 , n32561 , n352595 , n352596 , n352597 , n352598 , n32566 , n352600 , n352601 , n352602 , 
 n352603 , n352604 , n32572 , n352606 , n352607 , n352608 , n32576 , n352610 , n352611 , n352612 , 
 n352613 , n352614 , n352615 , n32583 , n352617 , n352618 , n32586 , n32587 , n352621 , n352622 , 
 n352623 , n32591 , n352625 , n352626 , n352627 , n352628 , n32596 , n32597 , n352631 , n352632 , 
 n352633 , n32601 , n352635 , n352636 , n352637 , n352638 , n352639 , n32607 , n352641 , n352642 , 
 n352643 , n352644 , n352645 , n352646 , n32614 , n352648 , n352649 , n32617 , n352651 , n352652 , 
 n352653 , n352654 , n352655 , n352656 , n352657 , n352658 , n32626 , n32627 , n32628 , n352662 , 
 n352663 , n352664 , n32632 , n352666 , n32634 , n352668 , n352669 , n32637 , n352671 , n32639 , 
 n352673 , n352674 , n352675 , n352676 , n352677 , n352678 , n32646 , n352680 , n352681 , n32649 , 
 n352683 , n352684 , n352685 , n32653 , n32654 , n32655 , n352689 , n32657 , n352691 , n352692 , 
 n32660 , n352694 , n352695 , n32663 , n32664 , n352698 , n32666 , n352700 , n352701 , n32669 , 
 n352703 , n352704 , n32672 , n32673 , n32674 , n32675 , n32676 , n352710 , n32678 , n32679 , 
 n352713 , n32681 , n32682 , n352716 , n352717 , n352718 , n352719 , n352720 , n32688 , n352722 , 
 n352723 , n352724 , n32692 , n32693 , n32694 , n352728 , n32696 , n32697 , n352731 , n352732 , 
 n352733 , n32701 , n352735 , n352736 , n352737 , n32705 , n352739 , n352740 , n352741 , n352742 , 
 n352743 , n32711 , n352745 , n352746 , n32714 , n352748 , n352749 , n32717 , n352751 , n352752 , 
 n352753 , n352754 , n352755 , n352756 , n352757 , n32725 , n352759 , n352760 , n352761 , n352762 , 
 n352763 , n352764 , n352765 , n32733 , n352767 , n352768 , n352769 , n352770 , n352771 , n352772 , 
 n352773 , n32741 , n352775 , n352776 , n352777 , n32745 , n32746 , n32747 , n352781 , n352782 , 
 n352783 , n352784 , n352785 , n352786 , n32754 , n352788 , n352789 , n32757 , n352791 , n352792 , 
 n32760 , n352794 , n352795 , n32763 , n352797 , n352798 , n352799 , n352800 , n352801 , n32769 , 
 n32770 , n352804 , n32772 , n32773 , n32774 , n352808 , n352809 , n32777 , n352811 , n32779 , 
 n352813 , n352814 , n352815 , n352816 , n32784 , n352818 , n32786 , n352820 , n352821 , n352822 , 
 n32790 , n352824 , n32792 , n352826 , n352827 , n352828 , n352829 , n352830 , n352831 , n352832 , 
 n352833 , n32801 , n352835 , n352836 , n352837 , n352838 , n352839 , n352840 , n352841 , n352842 , 
 n352843 , n32811 , n32812 , n352846 , n352847 , n352848 , n352849 , n352850 , n352851 , n352852 , 
 n352853 , n352854 , n32822 , n352856 , n352857 , n352858 , n32826 , n352860 , n352861 , n32829 , 
 n32830 , n352864 , n352865 , n32833 , n352867 , n352868 , n32836 , n352870 , n352871 , n352872 , 
 n352873 , n32841 , n352875 , n352876 , n352877 , n352878 , n32846 , n32847 , n352881 , n32849 , 
 n32850 , n352884 , n352885 , n32853 , n352887 , n352888 , n32856 , n352890 , n352891 , n352892 , 
 n32860 , n352894 , n352895 , n352896 , n352897 , n352898 , n352899 , n352900 , n352901 , n352902 , 
 n352903 , n352904 , n352905 , n352906 , n352907 , n352908 , n352909 , n352910 , n352911 , n352912 , 
 n352913 , n352914 , n352915 , n352916 , n32884 , n32885 , n352919 , n352920 , n352921 , n352922 , 
 n32890 , n352924 , n32892 , n352926 , n352927 , n352928 , n352929 , n352930 , n352931 , n352932 , 
 n352933 , n352934 , n352935 , n352936 , n352937 , n352938 , n352939 , n352940 , n352941 , n352942 , 
 n352943 , n352944 , n32912 , n352946 , n352947 , n352948 , n352949 , n352950 , n352951 , n32919 , 
 n352953 , n352954 , n32922 , n352956 , n352957 , n352958 , n352959 , n352960 , n352961 , n352962 , 
 n32930 , n32931 , n32932 , n32933 , n352967 , n352968 , n352969 , n352970 , n32938 , n352972 , 
 n352973 , n32941 , n352975 , n32943 , n32944 , n32945 , n352979 , n32947 , n352981 , n32949 , 
 n32950 , n32951 , n352985 , n352986 , n32954 , n352988 , n352989 , n32957 , n352991 , n32959 , 
 n32960 , n352994 , n32962 , n352996 , n352997 , n32965 , n352999 , n353000 , n32968 , n32969 , 
 n353003 , n32971 , n32972 , n353006 , n353007 , n353008 , n353009 , n353010 , n353011 , n353012 , 
 n32980 , n353014 , n353015 , n32983 , n353017 , n32985 , n32986 , n353020 , n32988 , n353022 , 
 n353023 , n32991 , n353025 , n353026 , n353027 , n353028 , n353029 , n353030 , n353031 , n353032 , 
 n353033 , n353034 , n353035 , n33003 , n353037 , n353038 , n33006 , n353040 , n353041 , n353042 , 
 n353043 , n353044 , n353045 , n353046 , n353047 , n353048 , n353049 , n33017 , n353051 , n33019 , 
 n353053 , n353054 , n353055 , n353056 , n33024 , n353058 , n33026 , n353060 , n353061 , n353062 , 
 n353063 , n353064 , n353065 , n353066 , n353067 , n353068 , n33036 , n353070 , n33038 , n353072 , 
 n353073 , n33041 , n33042 , n353076 , n353077 , n353078 , n353079 , n33047 , n33048 , n33049 , 
 n33050 , n33051 , n353085 , n353086 , n353087 , n353088 , n353089 , n33057 , n33058 , n353092 , 
 n33060 , n33061 , n33062 , n33063 , n353097 , n353098 , n353099 , n353100 , n33068 , n353102 , 
 n353103 , n353104 , n33072 , n353106 , n353107 , n33075 , n353109 , n353110 , n353111 , n33079 , 
 n33080 , n353114 , n33082 , n33083 , n353117 , n353118 , n353119 , n353120 , n353121 , n33089 , 
 n353123 , n353124 , n353125 , n353126 , n33094 , n353128 , n353129 , n353130 , n353131 , n353132 , 
 n353133 , n353134 , n353135 , n353136 , n353137 , n353138 , n353139 , n353140 , n353141 , n33109 , 
 n353143 , n353144 , n353145 , n353146 , n353147 , n33115 , n33116 , n353150 , n353151 , n33119 , 
 n353153 , n353154 , n33122 , n353156 , n353157 , n353158 , n353159 , n353160 , n353161 , n353162 , 
 n353163 , n353164 , n353165 , n33133 , n353167 , n33135 , n353169 , n33137 , n33138 , n353172 , 
 n353173 , n33141 , n353175 , n353176 , n33144 , n353178 , n353179 , n33147 , n33148 , n353182 , 
 n33150 , n353184 , n353185 , n353186 , n353187 , n33155 , n33156 , n353190 , n353191 , n33159 , 
 n353193 , n353194 , n33162 , n353196 , n353197 , n353198 , n353199 , n353200 , n353201 , n353202 , 
 n353203 , n353204 , n353205 , n353206 , n353207 , n353208 , n353209 , n353210 , n353211 , n353212 , 
 n33180 , n353214 , n353215 , n353216 , n33184 , n33185 , n353219 , n33187 , n353221 , n33189 , 
 n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n353229 , n353230 , n33198 , n353232 , 
 n353233 , n353234 , n353235 , n353236 , n353237 , n353238 , n353239 , n353240 , n353241 , n353242 , 
 n33210 , n33211 , n353245 , n353246 , n33214 , n353248 , n353249 , n33217 , n353251 , n33219 , 
 n353253 , n353254 , n353255 , n353256 , n353257 , n353258 , n33226 , n353260 , n353261 , n353262 , 
 n353263 , n353264 , n353265 , n33233 , n353267 , n33235 , n353269 , n353270 , n353271 , n353272 , 
 n33240 , n33241 , n353275 , n33243 , n353277 , n353278 , n33246 , n33247 , n353281 , n353282 , 
 n353283 , n33251 , n353285 , n353286 , n353287 , n353288 , n33256 , n353290 , n353291 , n353292 , 
 n33260 , n353294 , n353295 , n33263 , n353297 , n353298 , n353299 , n353300 , n33268 , n353302 , 
 n33270 , n353304 , n353305 , n33273 , n353307 , n353308 , n33276 , n353310 , n33278 , n353312 , 
 n353313 , n33281 , n353315 , n353316 , n33284 , n353318 , n353319 , n33287 , n353321 , n353322 , 
 n33290 , n353324 , n353325 , n353326 , n33294 , n353328 , n353329 , n353330 , n33298 , n353332 , 
 n353333 , n353334 , n33302 , n353336 , n33304 , n353338 , n353339 , n353340 , n353341 , n353342 , 
 n353343 , n353344 , n353345 , n353346 , n33314 , n33315 , n353349 , n33317 , n33318 , n353352 , 
 n353353 , n33321 , n353355 , n353356 , n353357 , n353358 , n353359 , n33327 , n353361 , n353362 , 
 n353363 , n33331 , n353365 , n353366 , n33334 , n353368 , n353369 , n33337 , n353371 , n33339 , 
 n353373 , n33341 , n33342 , n353376 , n353377 , n33345 , n353379 , n33347 , n353381 , n353382 , 
 n353383 , n353384 , n33352 , n353386 , n353387 , n353388 , n353389 , n353390 , n33358 , n353392 , 
 n353393 , n33361 , n353395 , n353396 , n33364 , n353398 , n353399 , n33367 , n33368 , n353402 , 
 n33370 , n353404 , n33372 , n353406 , n353407 , n353408 , n353409 , n33377 , n353411 , n353412 , 
 n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n353419 , n353420 , n353421 , n353422 , 
 n353423 , n353424 , n353425 , n353426 , n353427 , n353428 , n353429 , n353430 , n353431 , n33399 , 
 n353433 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n353441 , n353442 , 
 n33410 , n353444 , n353445 , n353446 , n353447 , n353448 , n353449 , n353450 , n33418 , n353452 , 
 n33420 , n33421 , n353455 , n33423 , n353457 , n353458 , n33426 , n353460 , n353461 , n33429 , 
 n353463 , n353464 , n33432 , n353466 , n353467 , n353468 , n353469 , n353470 , n353471 , n353472 , 
 n353473 , n353474 , n353475 , n353476 , n353477 , n33445 , n353479 , n353480 , n33448 , n353482 , 
 n353483 , n353484 , n33452 , n33453 , n33454 , n33455 , n353489 , n353490 , n353491 , n33459 , 
 n353493 , n353494 , n33462 , n353496 , n353497 , n33465 , n353499 , n353500 , n33468 , n353502 , 
 n353503 , n353504 , n353505 , n353506 , n353507 , n353508 , n33476 , n33477 , n353511 , n33479 , 
 n353513 , n353514 , n353515 , n33483 , n353517 , n33485 , n353519 , n353520 , n33488 , n353522 , 
 n33490 , n353524 , n353525 , n33493 , n353527 , n353528 , n33496 , n353530 , n353531 , n353532 , 
 n353533 , n353534 , n33502 , n353536 , n353537 , n353538 , n353539 , n353540 , n353541 , n353542 , 
 n353543 , n353544 , n33512 , n353546 , n353547 , n353548 , n33516 , n353550 , n353551 , n33519 , 
 n353553 , n353554 , n33522 , n33523 , n353557 , n33525 , n33526 , n353560 , n33528 , n353562 , 
 n353563 , n353564 , n353565 , n353566 , n353567 , n33535 , n33536 , n353570 , n33538 , n353572 , 
 n33540 , n353574 , n353575 , n353576 , n33544 , n33545 , n353579 , n353580 , n33548 , n353582 , 
 n353583 , n353584 , n353585 , n33553 , n353587 , n353588 , n353589 , n353590 , n353591 , n353592 , 
 n353593 , n353594 , n33562 , n353596 , n353597 , n33565 , n353599 , n353600 , n353601 , n353602 , 
 n353603 , n353604 , n353605 , n353606 , n33574 , n353608 , n353609 , n353610 , n353611 , n33579 , 
 n353613 , n33581 , n353615 , n353616 , n33584 , n353618 , n353619 , n353620 , n353621 , n353622 , 
 n33590 , n353624 , n353625 , n353626 , n33594 , n353628 , n353629 , n33597 , n353631 , n33599 , 
 n33600 , n353634 , n353635 , n33603 , n353637 , n353638 , n353639 , n353640 , n353641 , n353642 , 
 n33610 , n353644 , n353645 , n353646 , n353647 , n353648 , n353649 , n33617 , n353651 , n353652 , 
 n353653 , n33621 , n353655 , n33623 , n353657 , n353658 , n33626 , n353660 , n353661 , n33629 , 
 n353663 , n353664 , n353665 , n353666 , n353667 , n353668 , n33636 , n353670 , n353671 , n33639 , 
 n353673 , n33641 , n353675 , n353676 , n33644 , n353678 , n33646 , n353680 , n33648 , n353682 , 
 n33650 , n353684 , n353685 , n33653 , n33654 , n353688 , n353689 , n353690 , n33658 , n353692 , 
 n33660 , n33661 , n33662 , n353696 , n353697 , n353698 , n33666 , n353700 , n353701 , n33669 , 
 n353703 , n353704 , n353705 , n353706 , n33674 , n353708 , n33676 , n353710 , n353711 , n353712 , 
 n353713 , n353714 , n353715 , n353716 , n353717 , n353718 , n353719 , n353720 , n353721 , n33689 , 
 n353723 , n353724 , n33692 , n353726 , n353727 , n33695 , n353729 , n353730 , n353731 , n353732 , 
 n353733 , n353734 , n33702 , n353736 , n353737 , n33705 , n353739 , n33707 , n353741 , n33709 , 
 n33710 , n353744 , n353745 , n353746 , n353747 , n353748 , n353749 , n353750 , n353751 , n353752 , 
 n353753 , n353754 , n353755 , n353756 , n353757 , n353758 , n33726 , n353760 , n33728 , n353762 , 
 n353763 , n353764 , n33732 , n353766 , n33734 , n33735 , n33736 , n353770 , n353771 , n353772 , 
 n353773 , n33741 , n353775 , n33743 , n33744 , n353778 , n353779 , n353780 , n353781 , n33749 , 
 n353783 , n33751 , n33752 , n33753 , n33754 , n353788 , n33756 , n33757 , n33758 , n353792 , 
 n353793 , n33761 , n33762 , n353796 , n353797 , n353798 , n33766 , n33767 , n353801 , n353802 , 
 n353803 , n353804 , n353805 , n353806 , n353807 , n353808 , n353809 , n33777 , n33778 , n33779 , 
 n33780 , n353814 , n353815 , n33783 , n353817 , n33785 , n33786 , n33787 , n353821 , n353822 , 
 n33790 , n33791 , n353825 , n353826 , n353827 , n353828 , n353829 , n353830 , n33798 , n353832 , 
 n353833 , n353834 , n353835 , n353836 , n353837 , n353838 , n33806 , n353840 , n353841 , n33809 , 
 n353843 , n353844 , n353845 , n353846 , n353847 , n33815 , n353849 , n353850 , n353851 , n353852 , 
 n33820 , n33821 , n353855 , n353856 , n33824 , n353858 , n33826 , n33827 , n33828 , n353862 , 
 n353863 , n33831 , n33832 , n353866 , n353867 , n33835 , n33836 , n353870 , n353871 , n353872 , 
 n353873 , n33841 , n353875 , n33843 , n353877 , n353878 , n353879 , n33847 , n353881 , n353882 , 
 n33850 , n353884 , n353885 , n353886 , n353887 , n353888 , n353889 , n353890 , n33858 , n353892 , 
 n353893 , n353894 , n33862 , n353896 , n353897 , n353898 , n33866 , n353900 , n353901 , n33869 , 
 n353903 , n353904 , n353905 , n33873 , n353907 , n353908 , n33876 , n353910 , n353911 , n353912 , 
 n353913 , n353914 , n353915 , n353916 , n33884 , n33885 , n353919 , n353920 , n353921 , n353922 , 
 n353923 , n353924 , n353925 , n353926 , n353927 , n353928 , n33896 , n353930 , n353931 , n353932 , 
 n353933 , n353934 , n353935 , n33903 , n353937 , n33905 , n353939 , n33907 , n33908 , n353942 , 
 n353943 , n33911 , n353945 , n353946 , n33914 , n353948 , n353949 , n353950 , n33918 , n353952 , 
 n353953 , n353954 , n33922 , n33923 , n33924 , n353958 , n33926 , n353960 , n353961 , n33929 , 
 n353963 , n353964 , n353965 , n33933 , n353967 , n353968 , n353969 , n353970 , n33938 , n353972 , 
 n33940 , n353974 , n33942 , n33943 , n353977 , n353978 , n353979 , n353980 , n353981 , n353982 , 
 n353983 , n353984 , n353985 , n33953 , n353987 , n353988 , n33956 , n353990 , n353991 , n33959 , 
 n33960 , n33961 , n353995 , n353996 , n33964 , n353998 , n353999 , n354000 , n354001 , n33969 , 
 n354003 , n33971 , n354005 , n354006 , n33974 , n33975 , n354009 , n354010 , n33978 , n354012 , 
 n33980 , n354014 , n33982 , n33983 , n354017 , n33985 , n354019 , n33987 , n33988 , n354022 , 
 n354023 , n354024 , n354025 , n354026 , n354027 , n354028 , n354029 , n354030 , n33998 , n354032 , 
 n354033 , n354034 , n354035 , n354036 , n354037 , n354038 , n354039 , n354040 , n34008 , n354042 , 
 n34010 , n354044 , n34012 , n34013 , n354047 , n354048 , n34016 , n354050 , n354051 , n34019 , 
 n354053 , n354054 , n354055 , n34023 , n354057 , n354058 , n34026 , n354060 , n354061 , n34029 , 
 n34030 , n34031 , n354065 , n354066 , n34034 , n34035 , n34036 , n354070 , n354071 , n34039 , 
 n34040 , n354074 , n354075 , n354076 , n354077 , n34045 , n34046 , n354080 , n354081 , n34049 , 
 n34050 , n354084 , n354085 , n354086 , n354087 , n34055 , n354089 , n354090 , n354091 , n354092 , 
 n354093 , n354094 , n354095 , n34063 , n34064 , n354098 , n354099 , n354100 , n354101 , n354102 , 
 n354103 , n354104 , n354105 , n354106 , n354107 , n354108 , n34076 , n354110 , n354111 , n354112 , 
 n354113 , n354114 , n354115 , n354116 , n354117 , n354118 , n354119 , n354120 , n354121 , n354122 , 
 n354123 , n354124 , n34092 , n354126 , n354127 , n354128 , n354129 , n354130 , n354131 , n354132 , 
 n354133 , n354134 , n354135 , n354136 , n354137 , n354138 , n34106 , n354140 , n354141 , n354142 , 
 n354143 , n354144 , n34112 , n354146 , n34114 , n34115 , n354149 , n354150 , n354151 , n354152 , 
 n34120 , n354154 , n354155 , n34123 , n354157 , n354158 , n34126 , n354160 , n34128 , n354162 , 
 n34130 , n354164 , n354165 , n354166 , n354167 , n34135 , n354169 , n354170 , n354171 , n354172 , 
 n354173 , n354174 , n354175 , n354176 , n354177 , n354178 , n34146 , n354180 , n354181 , n34149 , 
 n354183 , n354184 , n34152 , n34153 , n34154 , n354188 , n354189 , n34157 , n354191 , n354192 , 
 n34160 , n354194 , n34162 , n34163 , n354197 , n34165 , n354199 , n34167 , n34168 , n354202 , 
 n354203 , n354204 , n354205 , n354206 , n34174 , n354208 , n354209 , n354210 , n34178 , n354212 , 
 n354213 , n34181 , n354215 , n354216 , n34184 , n354218 , n34186 , n34187 , n354221 , n34189 , 
 n354223 , n354224 , n354225 , n354226 , n34194 , n354228 , n354229 , n354230 , n354231 , n34199 , 
 n354233 , n354234 , n34202 , n354236 , n34204 , n354238 , n354239 , n34207 , n354241 , n354242 , 
 n354243 , n354244 , n354245 , n34213 , n354247 , n354248 , n354249 , n354250 , n354251 , n354252 , 
 n354253 , n354254 , n34222 , n354256 , n354257 , n354258 , n354259 , n34227 , n354261 , n354262 , 
 n354263 , n34231 , n354265 , n354266 , n354267 , n354268 , n34236 , n354270 , n354271 , n354272 , 
 n354273 , n354274 , n354275 , n354276 , n354277 , n354278 , n354279 , n354280 , n354281 , n34249 , 
 n354283 , n354284 , n354285 , n354286 , n354287 , n354288 , n34256 , n354290 , n354291 , n34259 , 
 n34260 , n354294 , n354295 , n34263 , n354297 , n354298 , n34266 , n354300 , n354301 , n34269 , 
 n354303 , n34271 , n354305 , n354306 , n34274 , n354308 , n34276 , n354310 , n34278 , n34279 , 
 n354313 , n354314 , n354315 , n354316 , n354317 , n34285 , n354319 , n354320 , n354321 , n354322 , 
 n354323 , n354324 , n354325 , n354326 , n354327 , n34295 , n354329 , n34297 , n354331 , n354332 , 
 n34300 , n354334 , n354335 , n354336 , n354337 , n34305 , n354339 , n354340 , n34308 , n34309 , 
 n354343 , n34311 , n34312 , n354346 , n354347 , n34315 , n354349 , n354350 , n354351 , n354352 , 
 n34320 , n354354 , n354355 , n354356 , n34324 , n354358 , n354359 , n354360 , n354361 , n354362 , 
 n34330 , n354364 , n354365 , n34333 , n354367 , n354368 , n354369 , n354370 , n34338 , n34339 , 
 n34340 , n354374 , n354375 , n34343 , n354377 , n34345 , n354379 , n354380 , n34348 , n354382 , 
 n354383 , n354384 , n34352 , n354386 , n354387 , n34355 , n354389 , n354390 , n354391 , n354392 , 
 n354393 , n354394 , n34362 , n34363 , n34364 , n354398 , n354399 , n354400 , n354401 , n354402 , 
 n354403 , n354404 , n34372 , n34373 , n354407 , n354408 , n34376 , n354410 , n354411 , n34379 , 
 n354413 , n354414 , n34382 , n354416 , n34384 , n354418 , n34386 , n354420 , n354421 , n354422 , 
 n354423 , n354424 , n354425 , n354426 , n354427 , n354428 , n34396 , n354430 , n34398 , n354432 , 
 n354433 , n354434 , n354435 , n354436 , n354437 , n34405 , n354439 , n354440 , n354441 , n354442 , 
 n34410 , n354444 , n34412 , n354446 , n354447 , n354448 , n354449 , n354450 , n34418 , n34419 , 
 n354453 , n354454 , n34422 , n354456 , n354457 , n34425 , n354459 , n354460 , n354461 , n354462 , 
 n354463 , n34431 , n354465 , n354466 , n354467 , n354468 , n354469 , n34437 , n34438 , n354472 , 
 n354473 , n354474 , n354475 , n354476 , n354477 , n354478 , n34446 , n34447 , n34448 , n34449 , 
 n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n354489 , n34457 , n354491 , n34459 , 
 n34460 , n354494 , n354495 , n34463 , n354497 , n34465 , n354499 , n354500 , n34468 , n354502 , 
 n354503 , n34471 , n354505 , n354506 , n34474 , n34475 , n354509 , n354510 , n34478 , n354512 , 
 n354513 , n34481 , n354515 , n354516 , n354517 , n354518 , n354519 , n354520 , n354521 , n354522 , 
 n354523 , n354524 , n354525 , n354526 , n34494 , n354528 , n354529 , n34497 , n354531 , n354532 , 
 n34500 , n354534 , n354535 , n34503 , n34504 , n34505 , n354539 , n354540 , n354541 , n354542 , 
 n34510 , n354544 , n34512 , n34513 , n354547 , n354548 , n34516 , n354550 , n354551 , n34519 , 
 n34520 , n354554 , n34522 , n354556 , n34524 , n354558 , n34526 , n34527 , n354561 , n34529 , 
 n354563 , n354564 , n354565 , n34533 , n354567 , n354568 , n34536 , n354570 , n354571 , n34539 , 
 n34540 , n354574 , n354575 , n34543 , n354577 , n354578 , n34546 , n354580 , n354581 , n354582 , 
 n354583 , n354584 , n354585 , n34553 , n354587 , n34555 , n354589 , n354590 , n34558 , n354592 , 
 n354593 , n34561 , n354595 , n354596 , n34564 , n354598 , n354599 , n354600 , n354601 , n354602 , 
 n354603 , n34571 , n354605 , n354606 , n354607 , n34575 , n34576 , n354610 , n34578 , n354612 , 
 n354613 , n354614 , n354615 , n354616 , n34584 , n354618 , n34586 , n354620 , n354621 , n354622 , 
 n354623 , n354624 , n354625 , n354626 , n354627 , n34595 , n354629 , n354630 , n354631 , n354632 , 
 n354633 , n354634 , n34602 , n354636 , n354637 , n34605 , n354639 , n354640 , n354641 , n34609 , 
 n354643 , n354644 , n354645 , n354646 , n354647 , n354648 , n354649 , n354650 , n354651 , n354652 , 
 n354653 , n34621 , n354655 , n34623 , n354657 , n354658 , n354659 , n354660 , n34628 , n34629 , 
 n354663 , n34631 , n34632 , n354666 , n34634 , n354668 , n354669 , n34637 , n354671 , n354672 , 
 n354673 , n34641 , n354675 , n34643 , n34644 , n354678 , n354679 , n354680 , n354681 , n354682 , 
 n354683 , n34651 , n34652 , n354686 , n34654 , n354688 , n354689 , n34657 , n354691 , n34659 , 
 n34660 , n34661 , n34662 , n354696 , n34664 , n34665 , n34666 , n34667 , n354701 , n354702 , 
 n34670 , n354704 , n354705 , n354706 , n34674 , n354708 , n354709 , n354710 , n354711 , n34679 , 
 n34680 , n354714 , n34682 , n354716 , n34684 , n354718 , n354719 , n354720 , n34688 , n354722 , 
 n354723 , n354724 , n354725 , n354726 , n34694 , n354728 , n354729 , n34697 , n354731 , n34699 , 
 n354733 , n354734 , n354735 , n354736 , n354737 , n354738 , n34706 , n354740 , n34708 , n354742 , 
 n354743 , n34711 , n354745 , n354746 , n34714 , n354748 , n354749 , n34717 , n354751 , n354752 , 
 n354753 , n34721 , n354755 , n354756 , n354757 , n354758 , n354759 , n354760 , n34728 , n354762 , 
 n354763 , n34731 , n354765 , n34733 , n354767 , n354768 , n34736 , n354770 , n354771 , n354772 , 
 n34740 , n354774 , n354775 , n34743 , n354777 , n354778 , n34746 , n354780 , n354781 , n354782 , 
 n354783 , n354784 , n354785 , n354786 , n34754 , n354788 , n354789 , n34757 , n34758 , n354792 , 
 n354793 , n354794 , n354795 , n354796 , n34764 , n354798 , n354799 , n34767 , n354801 , n354802 , 
 n34770 , n354804 , n354805 , n34773 , n354807 , n354808 , n34776 , n34777 , n354811 , n354812 , 
 n354813 , n354814 , n354815 , n34783 , n34784 , n354818 , n34786 , n354820 , n354821 , n354822 , 
 n354823 , n354824 , n34792 , n354826 , n354827 , n354828 , n354829 , n354830 , n354831 , n354832 , 
 n354833 , n34801 , n34802 , n34803 , n354837 , n34805 , n354839 , n354840 , n354841 , n354842 , 
 n354843 , n354844 , n34812 , n354846 , n354847 , n354848 , n354849 , n354850 , n354851 , n34819 , 
 n34820 , n34821 , n354855 , n354856 , n354857 , n354858 , n34826 , n354860 , n354861 , n354862 , 
 n354863 , n34831 , n354865 , n354866 , n354867 , n34835 , n354869 , n354870 , n354871 , n34839 , 
 n354873 , n354874 , n354875 , n34843 , n354877 , n354878 , n354879 , n34847 , n354881 , n354882 , 
 n354883 , n354884 , n354885 , n354886 , n354887 , n354888 , n354889 , n34857 , n354891 , n354892 , 
 n34860 , n354894 , n354895 , n354896 , n354897 , n34865 , n354899 , n354900 , n34868 , n354902 , 
 n354903 , n354904 , n354905 , n354906 , n354907 , n354908 , n354909 , n354910 , n34878 , n354912 , 
 n354913 , n354914 , n34882 , n354916 , n354917 , n34885 , n354919 , n354920 , n34888 , n34889 , 
 n34890 , n34891 , n34892 , n34893 , n354927 , n354928 , n354929 , n354930 , n354931 , n34899 , 
 n354933 , n354934 , n354935 , n354936 , n34904 , n354938 , n354939 , n354940 , n354941 , n34909 , 
 n354943 , n34911 , n354945 , n354946 , n354947 , n34915 , n354949 , n354950 , n354951 , n354952 , 
 n354953 , n354954 , n34922 , n354956 , n354957 , n34925 , n354959 , n354960 , n34928 , n354962 , 
 n354963 , n354964 , n354965 , n34933 , n354967 , n354968 , n34936 , n354970 , n354971 , n354972 , 
 n354973 , n354974 , n34942 , n34943 , n354977 , n354978 , n34946 , n34947 , n34948 , n354982 , 
 n354983 , n34951 , n354985 , n34953 , n354987 , n354988 , n34956 , n354990 , n354991 , n354992 , 
 n34960 , n354994 , n354995 , n34963 , n354997 , n34965 , n354999 , n355000 , n34968 , n355002 , 
 n355003 , n355004 , n355005 , n355006 , n34974 , n355008 , n355009 , n355010 , n34978 , n355012 , 
 n34980 , n355014 , n34982 , n355016 , n355017 , n34985 , n34986 , n34987 , n355021 , n34989 , 
 n355023 , n34991 , n355025 , n355026 , n34994 , n355028 , n355029 , n355030 , n355031 , n355032 , 
 n355033 , n355034 , n355035 , n355036 , n355037 , n355038 , n355039 , n355040 , n355041 , n355042 , 
 n35010 , n35011 , n35012 , n35013 , n355047 , n355048 , n35016 , n355050 , n35018 , n355052 , 
 n35020 , n35021 , n355055 , n355056 , n355057 , n355058 , n355059 , n35027 , n355061 , n35029 , 
 n355063 , n355064 , n35032 , n35033 , n355067 , n355068 , n35036 , n355070 , n35038 , n355072 , 
 n35040 , n355074 , n355075 , n355076 , n355077 , n355078 , n355079 , n355080 , n355081 , n35049 , 
 n355083 , n35051 , n355085 , n355086 , n35054 , n355088 , n355089 , n355090 , n355091 , n355092 , 
 n355093 , n355094 , n35062 , n355096 , n35064 , n355098 , n35066 , n355100 , n35068 , n35069 , 
 n35070 , n355104 , n355105 , n35073 , n35074 , n355108 , n355109 , n35077 , n355111 , n355112 , 
 n355113 , n355114 , n35082 , n355116 , n355117 , n355118 , n35086 , n35087 , n355121 , n355122 , 
 n355123 , n35091 , n355125 , n35093 , n35094 , n355128 , n35096 , n355130 , n35098 , n35099 , 
 n355133 , n355134 , n355135 , n355136 , n355137 , n35105 , n355139 , n355140 , n355141 , n35109 , 
 n355143 , n355144 , n35112 , n355146 , n35114 , n35115 , n355149 , n355150 , n355151 , n355152 , 
 n355153 , n35121 , n35122 , n355156 , n355157 , n35125 , n355159 , n355160 , n35128 , n355162 , 
 n355163 , n35131 , n35132 , n355166 , n355167 , n35135 , n355169 , n355170 , n35138 , n355172 , 
 n355173 , n355174 , n35142 , n35143 , n35144 , n355178 , n35146 , n355180 , n35148 , n355182 , 
 n355183 , n355184 , n355185 , n355186 , n355187 , n355188 , n355189 , n355190 , n355191 , n355192 , 
 n35160 , n355194 , n355195 , n355196 , n35164 , n355198 , n355199 , n355200 , n355201 , n355202 , 
 n355203 , n355204 , n355205 , n355206 , n355207 , n355208 , n355209 , n355210 , n35178 , n355212 , 
 n355213 , n35181 , n355215 , n355216 , n35184 , n355218 , n355219 , n355220 , n355221 , n355222 , 
 n35190 , n35191 , n355225 , n355226 , n355227 , n35195 , n355229 , n355230 , n355231 , n355232 , 
 n355233 , n355234 , n355235 , n355236 , n355237 , n355238 , n355239 , n355240 , n355241 , n35209 , 
 n355243 , n355244 , n35212 , n35213 , n355247 , n35215 , n355249 , n355250 , n355251 , n355252 , 
 n35220 , n35221 , n355255 , n35223 , n355257 , n35225 , n35226 , n35227 , n355261 , n35229 , 
 n355263 , n35231 , n355265 , n35233 , n355267 , n35235 , n355269 , n355270 , n35238 , n355272 , 
 n355273 , n35241 , n355275 , n355276 , n35244 , n355278 , n355279 , n35247 , n355281 , n35249 , 
 n355283 , n355284 , n355285 , n355286 , n355287 , n355288 , n355289 , n35257 , n355291 , n355292 , 
 n35260 , n355294 , n355295 , n355296 , n355297 , n355298 , n355299 , n355300 , n355301 , n35269 , 
 n355303 , n355304 , n35272 , n355306 , n35274 , n355308 , n355309 , n355310 , n355311 , n35279 , 
 n355313 , n355314 , n35282 , n35283 , n35284 , n355318 , n355319 , n355320 , n35288 , n35289 , 
 n355323 , n355324 , n355325 , n355326 , n355327 , n35295 , n355329 , n355330 , n355331 , n35299 , 
 n35300 , n355334 , n355335 , n35303 , n355337 , n355338 , n355339 , n355340 , n355341 , n35309 , 
 n355343 , n35311 , n355345 , n355346 , n355347 , n355348 , n35316 , n355350 , n35318 , n355352 , 
 n35320 , n35321 , n355355 , n355356 , n35324 , n355358 , n35326 , n35327 , n35328 , n355362 , 
 n35330 , n355364 , n355365 , n35333 , n355367 , n35335 , n355369 , n355370 , n35338 , n355372 , 
 n355373 , n35341 , n355375 , n355376 , n355377 , n355378 , n355379 , n355380 , n355381 , n355382 , 
 n355383 , n35351 , n355385 , n355386 , n355387 , n355388 , n355389 , n355390 , n355391 , n35359 , 
 n355393 , n35361 , n355395 , n355396 , n355397 , n355398 , n355399 , n355400 , n35368 , n355402 , 
 n355403 , n35371 , n35372 , n35373 , n355407 , n355408 , n355409 , n35377 , n355411 , n355412 , 
 n35380 , n355414 , n35382 , n355416 , n355417 , n355418 , n355419 , n35387 , n355421 , n355422 , 
 n355423 , n355424 , n355425 , n355426 , n355427 , n35395 , n355429 , n35397 , n35398 , n355432 , 
 n355433 , n35401 , n355435 , n355436 , n355437 , n355438 , n355439 , n355440 , n355441 , n35409 , 
 n355443 , n355444 , n35412 , n355446 , n355447 , n35415 , n35416 , n355450 , n355451 , n35419 , 
 n355453 , n355454 , n355455 , n35423 , n355457 , n355458 , n355459 , n35427 , n355461 , n355462 , 
 n35430 , n35431 , n355465 , n355466 , n35434 , n355468 , n355469 , n35437 , n35438 , n355472 , 
 n35440 , n355474 , n355475 , n35443 , n35444 , n35445 , n355479 , n355480 , n35448 , n35449 , 
 n35450 , n355484 , n355485 , n355486 , n35454 , n355488 , n355489 , n355490 , n35458 , n355492 , 
 n355493 , n355494 , n355495 , n35463 , n355497 , n355498 , n355499 , n355500 , n355501 , n35469 , 
 n355503 , n35471 , n35472 , n355506 , n355507 , n355508 , n35476 , n35477 , n35478 , n355512 , 
 n35480 , n355514 , n355515 , n35483 , n355517 , n35485 , n355519 , n355520 , n355521 , n35489 , 
 n355523 , n355524 , n355525 , n355526 , n35494 , n355528 , n35496 , n355530 , n35498 , n355532 , 
 n355533 , n35501 , n35502 , n355536 , n35504 , n35505 , n35506 , n355540 , n355541 , n35509 , 
 n35510 , n355544 , n355545 , n35513 , n35514 , n35515 , n355549 , n35517 , n35518 , n355552 , 
 n355553 , n355554 , n355555 , n355556 , n355557 , n35525 , n355559 , n355560 , n355561 , n355562 , 
 n35530 , n35531 , n355565 , n355566 , n355567 , n355568 , n35536 , n355570 , n355571 , n35539 , 
 n35540 , n35541 , n355575 , n355576 , n35544 , n355578 , n355579 , n35547 , n35548 , n355582 , 
 n35550 , n355584 , n35552 , n355586 , n355587 , n35555 , n355589 , n35557 , n355591 , n355592 , 
 n355593 , n355594 , n35562 , n355596 , n355597 , n35565 , n355599 , n355600 , n355601 , n35569 , 
 n355603 , n355604 , n35572 , n355606 , n355607 , n355608 , n355609 , n355610 , n35578 , n355612 , 
 n355613 , n355614 , n355615 , n355616 , n35584 , n35585 , n355619 , n35587 , n355621 , n355622 , 
 n35590 , n35591 , n355625 , n355626 , n355627 , n355628 , n35596 , n355630 , n355631 , n355632 , 
 n355633 , n355634 , n355635 , n355636 , n355637 , n355638 , n35606 , n355640 , n355641 , n35609 , 
 n355643 , n355644 , n35612 , n35613 , n35614 , n35615 , n35616 , n355650 , n35618 , n355652 , 
 n355653 , n355654 , n35622 , n355656 , n355657 , n35625 , n355659 , n355660 , n355661 , n355662 , 
 n35630 , n355664 , n355665 , n355666 , n35634 , n355668 , n355669 , n35637 , n35638 , n355672 , 
 n355673 , n35641 , n355675 , n355676 , n35644 , n35645 , n355679 , n35647 , n355681 , n355682 , 
 n35650 , n355684 , n355685 , n355686 , n355687 , n355688 , n355689 , n355690 , n35658 , n35659 , 
 n355693 , n355694 , n355695 , n35663 , n355697 , n355698 , n35666 , n355700 , n35668 , n35669 , 
 n35670 , n355704 , n355705 , n355706 , n355707 , n355708 , n35676 , n355710 , n355711 , n355712 , 
 n355713 , n355714 , n355715 , n35683 , n355717 , n355718 , n355719 , n35687 , n355721 , n355722 , 
 n355723 , n35691 , n355725 , n35693 , n355727 , n35695 , n355729 , n355730 , n355731 , n355732 , 
 n355733 , n355734 , n35702 , n355736 , n355737 , n355738 , n355739 , n35707 , n355741 , n35709 , 
 n355743 , n35711 , n35712 , n35713 , n355747 , n355748 , n355749 , n355750 , n35718 , n355752 , 
 n355753 , n355754 , n355755 , n355756 , n355757 , n355758 , n355759 , n35727 , n35728 , n35729 , 
 n35730 , n355764 , n35732 , n355766 , n355767 , n355768 , n355769 , n355770 , n35738 , n35739 , 
 n355773 , n355774 , n35742 , n355776 , n355777 , n35745 , n355779 , n355780 , n35748 , n35749 , 
 n355783 , n355784 , n35752 , n355786 , n355787 , n35755 , n35756 , n355790 , n35758 , n355792 , 
 n355793 , n35761 , n35762 , n355796 , n355797 , n35765 , n355799 , n355800 , n35768 , n355802 , 
 n355803 , n355804 , n355805 , n355806 , n35774 , n355808 , n355809 , n35777 , n355811 , n355812 , 
 n355813 , n35781 , n355815 , n35783 , n355817 , n355818 , n355819 , n355820 , n355821 , n355822 , 
 n355823 , n355824 , n355825 , n355826 , n355827 , n355828 , n35796 , n355830 , n355831 , n35799 , 
 n355833 , n355834 , n355835 , n355836 , n35804 , n35805 , n355839 , n355840 , n355841 , n355842 , 
 n355843 , n35811 , n355845 , n355846 , n355847 , n355848 , n355849 , n355850 , n355851 , n355852 , 
 n355853 , n355854 , n35822 , n355856 , n355857 , n355858 , n355859 , n355860 , n35828 , n355862 , 
 n355863 , n355864 , n355865 , n355866 , n355867 , n355868 , n35836 , n355870 , n355871 , n35839 , 
 n355873 , n355874 , n355875 , n355876 , n355877 , n355878 , n35846 , n355880 , n355881 , n35849 , 
 n355883 , n355884 , n355885 , n355886 , n355887 , n355888 , n355889 , n355890 , n355891 , n355892 , 
 n355893 , n355894 , n355895 , n35863 , n355897 , n355898 , n355899 , n355900 , n355901 , n35869 , 
 n35870 , n355904 , n355905 , n355906 , n355907 , n355908 , n355909 , n355910 , n355911 , n355912 , 
 n355913 , n355914 , n35879 , n355916 , n355917 , n35882 , n355919 , n355920 , n355921 , n355922 , 
 n355923 , n35888 , n35889 , n355926 , n35891 , n355928 , n35893 , n355930 , n35895 , n355932 , 
 n355933 , n35898 , n355935 , n355936 , n355937 , n355938 , n35903 , n355940 , n35905 , n355942 , 
 n355943 , n355944 , n35909 , n355946 , n355947 , n355948 , n355949 , n355950 , n355951 , n355952 , 
 n35917 , n355954 , n355955 , n355956 , n355957 , n355958 , n355959 , n355960 , n355961 , n355962 , 
 n355963 , n355964 , n355965 , n355966 , n35931 , n355968 , n355969 , n35934 , n355971 , n355972 , 
 n355973 , n355974 , n355975 , n355976 , n355977 , n355978 , n355979 , n355980 , n355981 , n355982 , 
 n355983 , n355984 , n355985 , n355986 , n355987 , n355988 , n355989 , n35954 , n355991 , n355992 , 
 n35957 , n355994 , n355995 , n355996 , n35961 , n355998 , n35963 , n356000 , n356001 , n35966 , 
 n356003 , n356004 , n35969 , n356006 , n356007 , n35972 , n356009 , n35974 , n35975 , n35976 , 
 n35977 , n356014 , n356015 , n356016 , n356017 , n35982 , n35983 , n356020 , n35985 , n356022 , 
 n356023 , n356024 , n35989 , n35990 , n35991 , n356028 , n35993 , n35994 , n356031 , n35996 , 
 n356033 , n35998 , n35999 , n356036 , n356037 , n36002 , n356039 , n356040 , n356041 , n356042 , 
 n356043 , n356044 , n36009 , n356046 , n356047 , n36012 , n356049 , n356050 , n36015 , n356052 , 
 n356053 , n36018 , n356055 , n356056 , n36021 , n36022 , n36023 , n356060 , n36025 , n356062 , 
 n356063 , n356064 , n36029 , n356066 , n356067 , n356068 , n356069 , n356070 , n356071 , n356072 , 
 n356073 , n356074 , n356075 , n356076 , n356077 , n356078 , n356079 , n356080 , n356081 , n356082 , 
 n356083 , n36048 , n356085 , n356086 , n356087 , n356088 , n356089 , n356090 , n356091 , n356092 , 
 n356093 , n356094 , n36059 , n356096 , n356097 , n36062 , n356099 , n356100 , n356101 , n356102 , 
 n36067 , n356104 , n36069 , n356106 , n356107 , n36072 , n356109 , n356110 , n36075 , n356112 , 
 n356113 , n36078 , n356115 , n36080 , n356117 , n356118 , n36083 , n356120 , n356121 , n356122 , 
 n356123 , n356124 , n356125 , n356126 , n36091 , n356128 , n356129 , n36094 , n36095 , n356132 , 
 n36097 , n356134 , n356135 , n36100 , n356137 , n356138 , n36103 , n356140 , n356141 , n36106 , 
 n356143 , n36108 , n36109 , n356146 , n356147 , n356148 , n356149 , n356150 , n356151 , n356152 , 
 n356153 , n356154 , n356155 , n36120 , n36121 , n356158 , n36123 , n356160 , n356161 , n36126 , 
 n356163 , n36128 , n356165 , n36130 , n356167 , n36132 , n356169 , n356170 , n36135 , n356172 , 
 n356173 , n356174 , n36139 , n356176 , n356177 , n356178 , n356179 , n356180 , n356181 , n356182 , 
 n356183 , n356184 , n356185 , n356186 , n356187 , n356188 , n356189 , n356190 , n356191 , n36156 , 
 n36157 , n36158 , n36159 , n356196 , n36161 , n356198 , n356199 , n36164 , n356201 , n356202 , 
 n356203 , n36168 , n356205 , n356206 , n356207 , n356208 , n36173 , n356210 , n356211 , n36176 , 
 n36177 , n36178 , n356215 , n356216 , n356217 , n356218 , n356219 , n356220 , n356221 , n356222 , 
 n356223 , n36188 , n356225 , n36190 , n356227 , n36192 , n356229 , n356230 , n356231 , n356232 , 
 n356233 , n356234 , n356235 , n356236 , n36201 , n356238 , n356239 , n36204 , n36205 , n356242 , 
 n36207 , n356244 , n356245 , n356246 , n356247 , n356248 , n36213 , n356250 , n356251 , n356252 , 
 n36217 , n356254 , n356255 , n356256 , n356257 , n36222 , n356259 , n36224 , n356261 , n36226 , 
 n36227 , n356264 , n356265 , n36230 , n356267 , n356268 , n36233 , n356270 , n36235 , n36236 , 
 n356273 , n356274 , n356275 , n356276 , n356277 , n356278 , n36243 , n356280 , n356281 , n36246 , 
 n356283 , n36248 , n356285 , n356286 , n356287 , n356288 , n356289 , n356290 , n356291 , n356292 , 
 n356293 , n36258 , n36259 , n356296 , n356297 , n356298 , n356299 , n36264 , n356301 , n356302 , 
 n356303 , n36268 , n356305 , n356306 , n36271 , n356308 , n356309 , n36274 , n356311 , n36276 , 
 n36277 , n356314 , n356315 , n356316 , n356317 , n356318 , n36283 , n356320 , n36285 , n356322 , 
 n356323 , n36288 , n356325 , n36290 , n356327 , n356328 , n36293 , n356330 , n36295 , n36296 , 
 n356333 , n36298 , n356335 , n36300 , n356337 , n356338 , n356339 , n356340 , n356341 , n356342 , 
 n356343 , n356344 , n356345 , n356346 , n356347 , n356348 , n356349 , n356350 , n356351 , n356352 , 
 n36317 , n356354 , n356355 , n356356 , n356357 , n356358 , n356359 , n356360 , n356361 , n36326 , 
 n356363 , n356364 , n36329 , n356366 , n356367 , n356368 , n36333 , n356370 , n356371 , n36336 , 
 n356373 , n356374 , n356375 , n356376 , n356377 , n356378 , n36340 , n356380 , n356381 , n36343 , 
 n356383 , n356384 , n36346 , n356386 , n356387 , n356388 , n356389 , n356390 , n36352 , n356392 , 
 n356393 , n356394 , n356395 , n356396 , n356397 , n356398 , n356399 , n356400 , n356401 , n356402 , 
 n356403 , n356404 , n356405 , n356406 , n356407 , n356408 , n36358 , n36359 , n36360 , n36361 , 
 n356413 , n356414 , n356415 , n356416 , n356417 , n36367 , n356419 , n356420 , n356421 , n356422 , 
 n36372 , n356424 , n36374 , n36375 , n356427 , n36377 , n356429 , n36379 , n356431 , n356432 , 
 n356433 , n356434 , n356435 , n36385 , n36386 , n356438 , n356439 , n36389 , n356441 , n356442 , 
 n36392 , n356444 , n356445 , n356446 , n36396 , n356448 , n356449 , n356450 , n356451 , n356452 , 
 n356453 , n356454 , n356455 , n356456 , n356457 , n356458 , n356459 , n356460 , n356461 , n356462 , 
 n356463 , n356464 , n356465 , n356466 , n356467 , n356468 , n356469 , n356470 , n36417 , n356472 , 
 n36419 , n356474 , n356475 , n36422 , n356477 , n36424 , n356479 , n36426 , n356481 , n36428 , 
 n356483 , n356484 , n356485 , n356486 , n36433 , n356488 , n356489 , n356490 , n356491 , n356492 , 
 n36439 , n356494 , n356495 , n356496 , n356497 , n356498 , n356499 , n356500 , n356501 , n356502 , 
 n36449 , n36450 , n36451 , n36452 , n36453 , n356508 , n36455 , n36456 , n356511 , n36458 , 
 n356513 , n356514 , n36461 , n356516 , n356517 , n356518 , n356519 , n356520 , n36467 , n356522 , 
 n36469 , n36470 , n356525 , n356526 , n36473 , n356528 , n356529 , n36476 , n36477 , n356532 , 
 n36479 , n356534 , n356535 , n356536 , n36483 , n356538 , n356539 , n36486 , n36487 , n356542 , 
 n36489 , n356544 , n36491 , n36492 , n356547 , n36494 , n356549 , n356550 , n36497 , n36498 , 
 n356553 , n356554 , n356555 , n356556 , n356557 , n356558 , n36505 , n356560 , n356561 , n36508 , 
 n356563 , n356564 , n356565 , n36512 , n356567 , n356568 , n36515 , n36516 , n356571 , n356572 , 
 n36519 , n356574 , n356575 , n36522 , n356577 , n36524 , n356579 , n36526 , n36527 , n36528 , 
 n356583 , n356584 , n356585 , n36532 , n356587 , n36534 , n36535 , n356590 , n36537 , n356592 , 
 n356593 , n36540 , n36541 , n36542 , n356597 , n36544 , n356599 , n356600 , n356601 , n36548 , 
 n356603 , n356604 , n36551 , n356606 , n36553 , n36554 , n36555 , n356610 , n356611 , n356612 , 
 n356613 , n356614 , n36561 , n356616 , n36563 , n356618 , n356619 , n356620 , n356621 , n356622 , 
 n356623 , n356624 , n36571 , n356626 , n356627 , n356628 , n356629 , n356630 , n36577 , n356632 , 
 n356633 , n36580 , n356635 , n356636 , n36583 , n356638 , n356639 , n356640 , n356641 , n356642 , 
 n36589 , n356644 , n356645 , n36592 , n356647 , n356648 , n36595 , n356650 , n356651 , n356652 , 
 n356653 , n356654 , n356655 , n356656 , n356657 , n36604 , n356659 , n356660 , n36607 , n356662 , 
 n356663 , n36610 , n356665 , n356666 , n356667 , n356668 , n356669 , n356670 , n356671 , n356672 , 
 n36619 , n356674 , n36621 , n356676 , n356677 , n356678 , n356679 , n36626 , n356681 , n356682 , 
 n356683 , n356684 , n356685 , n356686 , n356687 , n356688 , n356689 , n356690 , n356691 , n36638 , 
 n36639 , n36640 , n36641 , n356696 , n356697 , n356698 , n356699 , n356700 , n356701 , n356702 , 
 n356703 , n356704 , n36651 , n356706 , n356707 , n356708 , n356709 , n356710 , n356711 , n356712 , 
 n36659 , n356714 , n356715 , n356716 , n356717 , n356718 , n356719 , n356720 , n36667 , n356722 , 
 n356723 , n356724 , n36671 , n356726 , n36673 , n356728 , n356729 , n356730 , n356731 , n356732 , 
 n356733 , n356734 , n356735 , n36682 , n356737 , n356738 , n356739 , n356740 , n36687 , n356742 , 
 n36689 , n36690 , n36691 , n356746 , n356747 , n356748 , n356749 , n356750 , n36697 , n356752 , 
 n356753 , n36700 , n36701 , n356756 , n356757 , n356758 , n356759 , n356760 , n356761 , n36708 , 
 n356763 , n356764 , n356765 , n356766 , n356767 , n356768 , n356769 , n36714 , n36715 , n36716 , 
 n356773 , n356774 , n356775 , n356776 , n356777 , n356778 , n356779 , n356780 , n356781 , n36720 , 
 n36721 , n356784 , n36723 , n356786 , n356787 , n356788 , n356789 , n36728 , n356791 , n356792 , 
 n36731 , n356794 , n356795 , n356796 , n356797 , n36736 , n356799 , n36738 , n36739 , n356802 , 
 n356803 , n36742 , n356805 , n356806 , n36745 , n356808 , n356809 , n356810 , n356811 , n36750 , 
 n36751 , n356814 , n356815 , n356816 , n356817 , n356818 , n356819 , n36758 , n356821 , n356822 , 
 n36761 , n356824 , n356825 , n356826 , n356827 , n356828 , n356829 , n356830 , n36769 , n356832 , 
 n356833 , n356834 , n356835 , n36774 , n36775 , n356838 , n356839 , n356840 , n356841 , n356842 , 
 n356843 , n356844 , n356845 , n356846 , n356847 , n36783 , n356849 , n356850 , n356851 , n356852 , 
 n356853 , n356854 , n356855 , n356856 , n36792 , n356858 , n356859 , n356860 , n36796 , n356862 , 
 n36798 , n356864 , n356865 , n356866 , n356867 , n36803 , n356869 , n356870 , n36806 , n356872 , 
 n356873 , n36809 , n356875 , n356876 , n356877 , n36813 , n36814 , n356880 , n356881 , n36817 , 
 n36818 , n356884 , n356885 , n36821 , n36822 , n356888 , n36824 , n356890 , n36826 , n356892 , 
 n356893 , n356894 , n356895 , n356896 , n356897 , n356898 , n356899 , n356900 , n356901 , n356902 , 
 n356903 , n356904 , n356905 , n356906 , n356907 , n356908 , n356909 , n356910 , n356911 , n36847 , 
 n356913 , n356914 , n356915 , n36851 , n356917 , n356918 , n356919 , n36855 , n36856 , n356922 , 
 n356923 , n36859 , n356925 , n356926 , n356927 , n356928 , n356929 , n356930 , n356931 , n36867 , 
 n356933 , n356934 , n36870 , n356936 , n356937 , n36873 , n356939 , n356940 , n36876 , n36877 , 
 n356943 , n356944 , n36880 , n356946 , n356947 , n356948 , n356949 , n356950 , n356951 , n36887 , 
 n356953 , n356954 , n36890 , n356956 , n36892 , n356958 , n36894 , n36895 , n36896 , n356962 , 
 n36898 , n356964 , n36900 , n356966 , n36902 , n36903 , n356969 , n356970 , n36906 , n356972 , 
 n356973 , n356974 , n356975 , n356976 , n356977 , n356978 , n356979 , n356980 , n356981 , n356982 , 
 n356983 , n36919 , n36920 , n356986 , n356987 , n356988 , n356989 , n36925 , n356991 , n356992 , 
 n356993 , n356994 , n356995 , n36931 , n356997 , n356998 , n356999 , n357000 , n357001 , n36937 , 
 n357003 , n357004 , n357005 , n357006 , n357007 , n357008 , n36944 , n357010 , n357011 , n36947 , 
 n357013 , n357014 , n36950 , n36951 , n357017 , n357018 , n357019 , n357020 , n36956 , n357022 , 
 n36958 , n357024 , n357025 , n357026 , n36962 , n357028 , n357029 , n357030 , n357031 , n357032 , 
 n36968 , n36969 , n357035 , n357036 , n36972 , n357038 , n357039 , n357040 , n357041 , n357042 , 
 n36978 , n357044 , n357045 , n357046 , n357047 , n357048 , n36984 , n357050 , n357051 , n36987 , 
 n357053 , n357054 , n357055 , n357056 , n357057 , n357058 , n357059 , n357060 , n357061 , n357062 , 
 n357063 , n357064 , n37000 , n357066 , n357067 , n37003 , n357069 , n357070 , n357071 , n37007 , 
 n357073 , n357074 , n37010 , n357076 , n357077 , n357078 , n357079 , n357080 , n37016 , n37017 , 
 n357083 , n37019 , n357085 , n37021 , n357087 , n37023 , n357089 , n357090 , n37026 , n357092 , 
 n357093 , n37029 , n37030 , n357096 , n357097 , n37033 , n357099 , n357100 , n357101 , n357102 , 
 n357103 , n37039 , n357105 , n37041 , n357107 , n357108 , n37044 , n357110 , n357111 , n37047 , 
 n357113 , n357114 , n357115 , n357116 , n357117 , n357118 , n357119 , n357120 , n357121 , n357122 , 
 n357123 , n357124 , n357125 , n357126 , n357127 , n357128 , n357129 , n357130 , n357131 , n357132 , 
 n37068 , n357134 , n37070 , n357136 , n37072 , n357138 , n37074 , n37075 , n357141 , n357142 , 
 n37078 , n357144 , n357145 , n357146 , n357147 , n357148 , n357149 , n357150 , n357151 , n357152 , 
 n357153 , n357154 , n357155 , n357156 , n357157 , n357158 , n357159 , n357160 , n357161 , n357162 , 
 n357163 , n357164 , n357165 , n37100 , n357167 , n357168 , n37103 , n37104 , n37105 , n37106 , 
 n357173 , n357174 , n357175 , n357176 , n37111 , n357178 , n357179 , n357180 , n357181 , n357182 , 
 n37117 , n357184 , n37119 , n37120 , n357187 , n37122 , n357189 , n357190 , n37125 , n357192 , 
 n37127 , n357194 , n37129 , n357196 , n357197 , n37132 , n357199 , n37134 , n357201 , n37136 , 
 n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n357209 , n37144 , n37145 , n37146 , 
 n37147 , n357214 , n357215 , n357216 , n37151 , n37152 , n37153 , n357220 , n357221 , n37156 , 
 n357223 , n357224 , n357225 , n357226 , n357227 , n357228 , n357229 , n357230 , n357231 , n357232 , 
 n357233 , n357234 , n357235 , n37167 , n357237 , n37169 , n357239 , n357240 , n357241 , n37173 , 
 n357243 , n357244 , n357245 , n37177 , n357247 , n37179 , n357249 , n37181 , n37182 , n357252 , 
 n357253 , n357254 , n357255 , n357256 , n357257 , n357258 , n37190 , n37191 , n37192 , n37193 , 
 n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n357269 , n357270 , n357271 , n357272 , 
 n357273 , n357274 , n357275 , n357276 , n357277 , n357278 , n357279 , n357280 , n357281 , n357282 , 
 n357283 , n357284 , n357285 , n357286 , n357287 , n357288 , n37220 , n357290 , n357291 , n357292 , 
 n357293 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , 
 n37234 , n357304 , n357305 , n357306 , n357307 , n357308 , n357309 , n357310 , n357311 , n357312 , 
 n37244 , n357314 , n357315 , n37247 , n37248 , n357318 , n357319 , n357320 , n357321 , n357322 , 
 n357323 , n357324 , n357325 , n357326 , n37258 , n357328 , n37260 , n37261 , n37262 , n37263 , 
 n37264 , n37265 , n357335 , n37267 , n357337 , n357338 , n37270 , n357340 , n357341 , n37273 , 
 n37274 , n357344 , n37276 , n37277 , n357347 , n37279 , n37280 , n357350 , n357351 , n357352 , 
 n357353 , n357354 , n37286 , n357356 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , 
 n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n357370 , n37302 , n357372 , 
 n37304 , n37305 , n37306 , n357376 , n37308 , n357378 , n357379 , n357380 , n357381 , n37313 , 
 n357383 , n357384 , n357385 , n37317 , n357387 , n37319 , n357389 , n37321 , n357391 , n37323 , 
 n357393 , n37325 , n357395 , n357396 , n37328 , n37329 , n357399 , n357400 , n37332 , n357402 , 
 n357403 , n37335 , n357405 , n357406 , n357407 , n357408 , n357409 , n357410 , n37342 , n357412 , 
 n357413 , n357414 , n357415 , n37347 , n357417 , n357418 , n37350 , n357420 , n357421 , n357422 , 
 n357423 , n357424 , n37356 , n357426 , n357427 , n357428 , n357429 , n357430 , n357431 , n357432 , 
 n357433 , n357434 , n37366 , n357436 , n357437 , n357438 , n357439 , n357440 , n357441 , n37373 , 
 n357443 , n37375 , n37376 , n357446 , n357447 , n37379 , n357449 , n37381 , n37382 , n37383 , 
 n37384 , n37385 , n37386 , n357456 , n357457 , n357458 , n357459 , n37391 , n357461 , n357462 , 
 n37394 , n357464 , n357465 , n357466 , n357467 , n37399 , n357469 , n357470 , n37402 , n357472 , 
 n357473 , n37405 , n357475 , n37407 , n37408 , n37409 , n37410 , n357480 , n37412 , n357482 , 
 n37414 , n357484 , n357485 , n357486 , n357487 , n357488 , n357489 , n357490 , n357491 , n37423 , 
 n357493 , n37425 , n37426 , n357496 , n37428 , n357498 , n37430 , n357500 , n37432 , n37433 , 
 n37434 , n357504 , n357505 , n37437 , n357507 , n37439 , n37440 , n357510 , n37442 , n357512 , 
 n357513 , n357514 , n357515 , n357516 , n357517 , n357518 , n357519 , n37451 , n357521 , n37453 , 
 n357523 , n357524 , n357525 , n357526 , n357527 , n357528 , n37460 , n357530 , n37462 , n357532 , 
 n37464 , n37465 , n357535 , n357536 , n37468 , n37469 , n357539 , n357540 , n37472 , n357542 , 
 n357543 , n37475 , n357545 , n37477 , n357547 , n357548 , n37480 , n357550 , n357551 , n37483 , 
 n357553 , n357554 , n357555 , n37487 , n357557 , n37489 , n37490 , n357560 , n357561 , n357562 , 
 n357563 , n357564 , n357565 , n357566 , n357567 , n37499 , n37500 , n357570 , n37502 , n357572 , 
 n37504 , n37505 , n357575 , n357576 , n37508 , n37509 , n357579 , n37511 , n357581 , n357582 , 
 n357583 , n357584 , n357585 , n357586 , n357587 , n37519 , n357589 , n357590 , n37522 , n357592 , 
 n37524 , n37525 , n357595 , n357596 , n37528 , n357598 , n357599 , n37531 , n357601 , n357602 , 
 n357603 , n37535 , n357605 , n357606 , n357607 , n37539 , n357609 , n357610 , n37542 , n357612 , 
 n357613 , n357614 , n357615 , n37547 , n357617 , n357618 , n37550 , n37551 , n357621 , n37553 , 
 n357623 , n357624 , n357625 , n37557 , n357627 , n357628 , n37560 , n357630 , n37562 , n357632 , 
 n357633 , n357634 , n357635 , n357636 , n357637 , n357638 , n357639 , n37571 , n37572 , n357642 , 
 n357643 , n357644 , n37576 , n357646 , n357647 , n37579 , n357649 , n37581 , n357651 , n357652 , 
 n37584 , n357654 , n357655 , n357656 , n357657 , n357658 , n357659 , n357660 , n37592 , n357662 , 
 n37594 , n357664 , n357665 , n357666 , n357667 , n357668 , n357669 , n37601 , n357671 , n357672 , 
 n37604 , n357674 , n357675 , n37607 , n37608 , n357678 , n37610 , n357680 , n357681 , n357682 , 
 n37614 , n357684 , n357685 , n357686 , n357687 , n357688 , n37620 , n357690 , n37622 , n357692 , 
 n37624 , n37625 , n357695 , n357696 , n37628 , n357698 , n37630 , n37631 , n37632 , n357702 , 
 n357703 , n37635 , n357705 , n357706 , n37638 , n357708 , n37640 , n357710 , n37642 , n37643 , 
 n37644 , n37645 , n357715 , n357716 , n357717 , n357718 , n357719 , n37651 , n357721 , n37653 , 
 n37654 , n37655 , n357725 , n357726 , n357727 , n357728 , n357729 , n357730 , n37659 , n37660 , 
 n357733 , n37662 , n37663 , n357736 , n37665 , n357738 , n37667 , n37668 , n357741 , n357742 , 
 n37671 , n357744 , n357745 , n37674 , n357747 , n357748 , n357749 , n357750 , n357751 , n37680 , 
 n357753 , n357754 , n357755 , n357756 , n357757 , n357758 , n357759 , n357760 , n357761 , n357762 , 
 n37691 , n357764 , n357765 , n357766 , n357767 , n357768 , n37697 , n357770 , n37699 , n37700 , 
 n357773 , n357774 , n357775 , n357776 , n357777 , n357778 , n357779 , n357780 , n357781 , n37710 , 
 n357783 , n357784 , n37713 , n37714 , n357787 , n37716 , n37717 , n357790 , n357791 , n37720 , 
 n357793 , n37722 , n357795 , n37724 , n357797 , n357798 , n357799 , n37728 , n37729 , n37730 , 
 n37731 , n37732 , n37733 , n357806 , n357807 , n37736 , n357809 , n37738 , n37739 , n37740 , 
 n357813 , n357814 , n357815 , n37744 , n357817 , n37746 , n357819 , n37748 , n37749 , n37750 , 
 n357823 , n357824 , n357825 , n357826 , n357827 , n37756 , n357829 , n357830 , n37759 , n357832 , 
 n357833 , n37762 , n357835 , n37764 , n37765 , n357838 , n357839 , n37768 , n357841 , n357842 , 
 n37771 , n357844 , n37773 , n357846 , n37775 , n37776 , n357849 , n357850 , n37779 , n37780 , 
 n357853 , n37782 , n37783 , n357856 , n357857 , n357858 , n357859 , n357860 , n357861 , n357862 , 
 n357863 , n357864 , n357865 , n357866 , n357867 , n357868 , n357869 , n37798 , n37799 , n357872 , 
 n37801 , n357874 , n357875 , n357876 , n37802 , n37803 , n357879 , n357880 , n37806 , n357882 , 
 n357883 , n357884 , n357885 , n37811 , n37812 , n357888 , n37814 , n357890 , n37816 , n357892 , 
 n357893 , n357894 , n357895 , n37821 , n37822 , n37823 , n357899 , n37825 , n357901 , n37827 , 
 n357903 , n37829 , n357905 , n357906 , n357907 , n37833 , n357909 , n357910 , n37836 , n357912 , 
 n37838 , n357914 , n37840 , n37841 , n357917 , n37843 , n37844 , n37845 , n37846 , n357922 , 
 n37848 , n357924 , n37850 , n357926 , n357927 , n37853 , n357929 , n357930 , n37856 , n357932 , 
 n37858 , n37859 , n357935 , n37861 , n357937 , n37863 , n37864 , n37865 , n37866 , n37867 , 
 n37868 , n37869 , n37870 , n37871 , n37872 , n357948 , n37874 , n357950 , n357951 , n357952 , 
 n37878 , n37879 , n357955 , n357956 , n37882 , n357958 , n37884 , n357960 , n357961 , n357962 , 
 n357963 , n357964 , n357965 , n357966 , n357967 , n357968 , n357969 , n357970 , n357971 , n357972 , 
 n357973 , n357974 , n357975 , n357976 , n37902 , n357978 , n357979 , n357980 , n357981 , n37907 , 
 n357983 , n357984 , n37910 , n357986 , n357987 , n37913 , n357989 , n357990 , n37916 , n357992 , 
 n37918 , n357994 , n357995 , n37921 , n357997 , n357998 , n37924 , n37925 , n358001 , n37927 , 
 n37928 , n358004 , n358005 , n37931 , n358007 , n358008 , n358009 , n358010 , n37936 , n358012 , 
 n358013 , n358014 , n358015 , n358016 , n358017 , n358018 , n358019 , n358020 , n358021 , n358022 , 
 n358023 , n358024 , n358025 , n358026 , n358027 , n358028 , n358029 , n358030 , n37956 , n358032 , 
 n358033 , n37959 , n358035 , n37961 , n37962 , n358038 , n358039 , n358040 , n358041 , n358042 , 
 n358043 , n37969 , n358045 , n37971 , n358047 , n358048 , n37974 , n358050 , n358051 , n358052 , 
 n358053 , n358054 , n37980 , n358056 , n358057 , n37983 , n37984 , n358060 , n358061 , n358062 , 
 n358063 , n358064 , n358065 , n358066 , n358067 , n37993 , n37994 , n37995 , n37996 , n37997 , 
 n358073 , n358074 , n358075 , n38001 , n358077 , n38003 , n358079 , n358080 , n358081 , n358082 , 
 n38008 , n358084 , n358085 , n358086 , n358087 , n358088 , n358089 , n38015 , n358091 , n358092 , 
 n38018 , n358094 , n38020 , n38021 , n358097 , n358098 , n38024 , n358100 , n358101 , n358102 , 
 n38028 , n38029 , n38030 , n358106 , n38032 , n38033 , n358109 , n38035 , n358111 , n358112 , 
 n38038 , n358114 , n38040 , n358116 , n38042 , n38043 , n358119 , n38045 , n358121 , n38047 , 
 n358123 , n358124 , n38050 , n358126 , n38052 , n38053 , n38054 , n358130 , n38056 , n358132 , 
 n358133 , n358134 , n358135 , n358136 , n358137 , n358138 , n358139 , n358140 , n358141 , n358142 , 
 n358143 , n358144 , n358145 , n358146 , n358147 , n38073 , n358149 , n358150 , n38076 , n358152 , 
 n38078 , n358154 , n358155 , n358156 , n358157 , n358158 , n358159 , n358160 , n358161 , n358162 , 
 n38088 , n358164 , n358165 , n38091 , n358167 , n358168 , n358169 , n358170 , n38096 , n358172 , 
 n38098 , n358174 , n38100 , n358176 , n38102 , n358178 , n358179 , n358180 , n358181 , n358182 , 
 n358183 , n358184 , n38110 , n358186 , n358187 , n358188 , n38114 , n358190 , n38116 , n38117 , 
 n358193 , n358194 , n358195 , n38121 , n358197 , n358198 , n358199 , n358200 , n38126 , n358202 , 
 n358203 , n38129 , n358205 , n358206 , n38132 , n38133 , n358209 , n38135 , n38136 , n358212 , 
 n38138 , n358214 , n358215 , n358216 , n358217 , n358218 , n358219 , n358220 , n38146 , n358222 , 
 n358223 , n38149 , n358225 , n358226 , n38152 , n358228 , n38154 , n358230 , n38156 , n38157 , 
 n358233 , n358234 , n38160 , n358236 , n358237 , n38163 , n38164 , n358240 , n38166 , n38167 , 
 n358243 , n358244 , n358245 , n38171 , n358247 , n38173 , n358249 , n358250 , n358251 , n358252 , 
 n358253 , n358254 , n38180 , n358256 , n358257 , n358258 , n358259 , n358260 , n38186 , n358262 , 
 n358263 , n358264 , n38190 , n358266 , n38192 , n358268 , n38194 , n358270 , n38196 , n38197 , 
 n358273 , n358274 , n358275 , n358276 , n38202 , n358278 , n38204 , n358280 , n358281 , n38207 , 
 n358283 , n38209 , n38210 , n358286 , n358287 , n38213 , n358289 , n38215 , n358291 , n358292 , 
 n38218 , n358294 , n38220 , n358296 , n358297 , n358298 , n38224 , n38225 , n38226 , n38227 , 
 n358303 , n358304 , n38230 , n358306 , n358307 , n38233 , n358309 , n358310 , n38236 , n38237 , 
 n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n358320 , n38246 , n358322 , 
 n358323 , n38249 , n358325 , n358326 , n38252 , n358328 , n358329 , n358330 , n358331 , n358332 , 
 n358333 , n358334 , n358335 , n358336 , n38262 , n358338 , n358339 , n358340 , n358341 , n358342 , 
 n38268 , n358344 , n358345 , n358346 , n38272 , n358348 , n358349 , n358350 , n358351 , n358352 , 
 n358353 , n358354 , n358355 , n358356 , n358357 , n358358 , n358359 , n358360 , n38286 , n38287 , 
 n358363 , n358364 , n358365 , n358366 , n358367 , n358368 , n358369 , n358370 , n358371 , n38297 , 
 n358373 , n358374 , n38300 , n358376 , n358377 , n38303 , n358379 , n38305 , n358381 , n358382 , 
 n358383 , n358384 , n358385 , n358386 , n358387 , n358388 , n358389 , n358390 , n358391 , n358392 , 
 n358393 , n358394 , n358395 , n358396 , n358397 , n38318 , n358399 , n38320 , n38321 , n358402 , 
 n358403 , n38324 , n358405 , n358406 , n358407 , n358408 , n358409 , n38330 , n358411 , n38332 , 
 n358413 , n358414 , n358415 , n358416 , n358417 , n358418 , n358419 , n358420 , n358421 , n358422 , 
 n358423 , n358424 , n358425 , n358426 , n358427 , n358428 , n38349 , n358430 , n38351 , n358432 , 
 n38353 , n358434 , n358435 , n38356 , n358437 , n358438 , n38359 , n358440 , n38361 , n358442 , 
 n38363 , n38364 , n358445 , n358446 , n38367 , n358448 , n358449 , n38370 , n358451 , n358452 , 
 n38373 , n358454 , n358455 , n358456 , n38377 , n358458 , n358459 , n38380 , n358461 , n38382 , 
 n358463 , n358464 , n358465 , n358466 , n358467 , n358468 , n38389 , n358470 , n358471 , n358472 , 
 n358473 , n358474 , n358475 , n358476 , n358477 , n358478 , n358479 , n38400 , n358481 , n358482 , 
 n358483 , n38404 , n358485 , n358486 , n358487 , n358488 , n358489 , n38410 , n358491 , n358492 , 
 n38413 , n358494 , n38415 , n358496 , n358497 , n38418 , n358499 , n358500 , n358501 , n358502 , 
 n358503 , n358504 , n358505 , n358506 , n358507 , n358508 , n358509 , n358510 , n358511 , n38432 , 
 n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n358519 , n38440 , n38441 , n358522 , 
 n38443 , n358524 , n38445 , n38446 , n38447 , n358528 , n358529 , n38450 , n358531 , n358532 , 
 n38453 , n358534 , n358535 , n358536 , n38457 , n358538 , n358539 , n38460 , n358541 , n358542 , 
 n38463 , n38464 , n38465 , n358546 , n358547 , n38468 , n358549 , n38470 , n38471 , n358552 , 
 n38473 , n358554 , n38475 , n38476 , n38477 , n358558 , n38479 , n358560 , n358561 , n358562 , 
 n38483 , n38484 , n358565 , n38486 , n358567 , n358568 , n38489 , n38490 , n358571 , n358572 , 
 n38493 , n358574 , n358575 , n38496 , n358577 , n358578 , n358579 , n358580 , n358581 , n358582 , 
 n358583 , n38504 , n358585 , n358586 , n38507 , n38508 , n358589 , n38510 , n38511 , n358592 , 
 n358593 , n358594 , n358595 , n358596 , n358597 , n38518 , n358599 , n358600 , n38521 , n358602 , 
 n38523 , n358604 , n358605 , n358606 , n38527 , n358608 , n358609 , n358610 , n358611 , n358612 , 
 n38533 , n358614 , n358615 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n358622 , 
 n358623 , n38544 , n358625 , n38546 , n358627 , n358628 , n358629 , n358630 , n358631 , n38552 , 
 n358633 , n38554 , n38555 , n38556 , n358637 , n38558 , n358639 , n358640 , n358641 , n38562 , 
 n358643 , n358644 , n38565 , n358646 , n358647 , n38568 , n358649 , n358650 , n358651 , n358652 , 
 n38573 , n358654 , n358655 , n38576 , n358657 , n358658 , n358659 , n358660 , n358661 , n38582 , 
 n38583 , n38584 , n358665 , n358666 , n358667 , n38588 , n358669 , n358670 , n358671 , n358672 , 
 n38593 , n358674 , n358675 , n358676 , n38597 , n358678 , n358679 , n38600 , n38601 , n358682 , 
 n358683 , n358684 , n358685 , n358686 , n358687 , n38608 , n358689 , n358690 , n358691 , n358692 , 
 n358693 , n38614 , n38615 , n38616 , n358697 , n358698 , n358699 , n358700 , n38621 , n358702 , 
 n38623 , n358704 , n358705 , n358706 , n38627 , n358708 , n358709 , n358710 , n358711 , n358712 , 
 n38630 , n358714 , n358715 , n358716 , n358717 , n38635 , n38636 , n358720 , n38638 , n38639 , 
 n358723 , n38641 , n38642 , n358726 , n358727 , n358728 , n38646 , n358730 , n358731 , n358732 , 
 n358733 , n38651 , n358735 , n358736 , n38654 , n358738 , n358739 , n358740 , n358741 , n358742 , 
 n38660 , n358744 , n358745 , n358746 , n38664 , n358748 , n358749 , n358750 , n358751 , n358752 , 
 n358753 , n358754 , n38672 , n358756 , n358757 , n358758 , n358759 , n38677 , n358761 , n358762 , 
 n38680 , n358764 , n358765 , n38683 , n358767 , n358768 , n38686 , n358770 , n358771 , n358772 , 
 n358773 , n358774 , n358775 , n38693 , n38694 , n38695 , n38696 , n358780 , n38698 , n358782 , 
 n358783 , n38701 , n38702 , n358786 , n358787 , n358788 , n38706 , n38707 , n358791 , n358792 , 
 n358793 , n38711 , n358795 , n358796 , n358797 , n38715 , n38716 , n358800 , n358801 , n38719 , 
 n358803 , n358804 , n358805 , n38723 , n38724 , n358808 , n38726 , n38727 , n358811 , n38729 , 
 n38730 , n358814 , n38732 , n358816 , n38734 , n358818 , n38736 , n358820 , n358821 , n38739 , 
 n38740 , n358824 , n358825 , n38743 , n38744 , n38745 , n358829 , n38747 , n358831 , n358832 , 
 n358833 , n38751 , n358835 , n358836 , n358837 , n358838 , n358839 , n38757 , n358841 , n358842 , 
 n38760 , n358844 , n38762 , n358846 , n358847 , n358848 , n358849 , n38767 , n358851 , n358852 , 
 n38770 , n358854 , n358855 , n38773 , n358857 , n358858 , n358859 , n358860 , n358861 , n358862 , 
 n358863 , n358864 , n358865 , n38783 , n358867 , n358868 , n358869 , n358870 , n358871 , n358872 , 
 n358873 , n358874 , n38792 , n38793 , n358877 , n38795 , n358879 , n358880 , n358881 , n358882 , 
 n358883 , n358884 , n358885 , n358886 , n358887 , n38800 , n38801 , n358890 , n358891 , n38804 , 
 n358893 , n358894 , n358895 , n358896 , n358897 , n358898 , n358899 , n358900 , n358901 , n358902 , 
 n38815 , n38816 , n358905 , n358906 , n38819 , n38820 , n38821 , n358910 , n358911 , n358912 , 
 n358913 , n358914 , n38827 , n358916 , n358917 , n358918 , n358919 , n358920 , n38833 , n358922 , 
 n358923 , n38836 , n358925 , n358926 , n38839 , n358928 , n358929 , n358930 , n358931 , n358932 , 
 n358933 , n38844 , n358935 , n358936 , n358937 , n358938 , n358939 , n358940 , n358941 , n358942 , 
 n358943 , n358944 , n358945 , n358946 , n358947 , n38858 , n38859 , n358950 , n358951 , n358952 , 
 n358953 , n38864 , n358955 , n358956 , n358957 , n358958 , n38869 , n38870 , n358961 , n358962 , 
 n358963 , n358964 , n358965 , n358966 , n358967 , n358968 , n38873 , n358970 , n38875 , n38876 , 
 n38877 , n38878 , n38879 , n358976 , n358977 , n38882 , n358979 , n38884 , n38885 , n358982 , 
 n358983 , n38888 , n358985 , n358986 , n358987 , n358988 , n358989 , n38894 , n358991 , n358992 , 
 n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n358999 , n38904 , n359001 , n38906 , 
 n38907 , n38908 , n38909 , n38910 , n38911 , n359008 , n359009 , n359010 , n359011 , n359012 , 
 n38917 , n359014 , n38919 , n359016 , n359017 , n359018 , n359019 , n359020 , n359021 , n38926 , 
 n359023 , n359024 , n38929 , n359026 , n359027 , n359028 , n359029 , n359030 , n38935 , n359032 , 
 n359033 , n359034 , n359035 , n38940 , n359037 , n359038 , n359039 , n359040 , n38945 , n359042 , 
 n359043 , n359044 , n359045 , n359046 , n38951 , n359048 , n359049 , n359050 , n38955 , n359052 , 
 n359053 , n359054 , n359055 , n38960 , n359057 , n359058 , n38963 , n38964 , n359061 , n38966 , 
 n38967 , n38968 , n359065 , n38970 , n359067 , n359068 , n38973 , n359070 , n359071 , n38976 , 
 n359073 , n38978 , n359075 , n38980 , n38981 , n38982 , n38983 , n359080 , n359081 , n359082 , 
 n359083 , n359084 , n359085 , n359086 , n359087 , n359088 , n359089 , n359090 , n359091 , n359092 , 
 n359093 , n359094 , n359095 , n359096 , n359097 , n359098 , n359099 , n39004 , n359101 , n359102 , 
 n39007 , n359104 , n359105 , n39010 , n39011 , n359108 , n359109 , n359110 , n359111 , n359112 , 
 n39017 , n359114 , n359115 , n39020 , n39021 , n359118 , n39023 , n359120 , n359121 , n39026 , 
 n359123 , n359124 , n39029 , n359126 , n359127 , n359128 , n359129 , n359130 , n359131 , n359132 , 
 n359133 , n359134 , n39039 , n359136 , n359137 , n39042 , n359139 , n39044 , n359141 , n39046 , 
 n39047 , n359144 , n359145 , n39050 , n359147 , n359148 , n359149 , n359150 , n359151 , n359152 , 
 n359153 , n359154 , n359155 , n359156 , n39061 , n359158 , n39063 , n39064 , n359161 , n359162 , 
 n359163 , n359164 , n359165 , n39070 , n359167 , n359168 , n359169 , n359170 , n39075 , n359172 , 
 n39077 , n359174 , n359175 , n359176 , n359177 , n359178 , n39083 , n359180 , n39085 , n359182 , 
 n39087 , n359184 , n359185 , n359186 , n359187 , n39092 , n359189 , n359190 , n359191 , n39096 , 
 n359193 , n359194 , n359195 , n39100 , n39101 , n39102 , n359199 , n359200 , n39105 , n359202 , 
 n359203 , n39108 , n359205 , n359206 , n359207 , n39112 , n359209 , n359210 , n39115 , n359212 , 
 n359213 , n39118 , n359215 , n359216 , n359217 , n359218 , n359219 , n359220 , n359221 , n359222 , 
 n39127 , n359224 , n359225 , n359226 , n39131 , n359228 , n359229 , n359230 , n359231 , n359232 , 
 n359233 , n39138 , n39139 , n359236 , n39141 , n359238 , n359239 , n39144 , n359241 , n359242 , 
 n359243 , n359244 , n359245 , n359246 , n39151 , n359248 , n359249 , n359250 , n359251 , n359252 , 
 n39157 , n359254 , n359255 , n359256 , n39161 , n359258 , n359259 , n359260 , n39165 , n359262 , 
 n359263 , n359264 , n39169 , n359266 , n359267 , n359268 , n359269 , n359270 , n39175 , n359272 , 
 n359273 , n359274 , n359275 , n39180 , n39181 , n359278 , n39183 , n359280 , n39185 , n359282 , 
 n359283 , n39188 , n39189 , n359286 , n359287 , n359288 , n39193 , n359290 , n359291 , n359292 , 
 n39197 , n359294 , n39199 , n359296 , n359297 , n359298 , n39203 , n39204 , n39205 , n359302 , 
 n39207 , n39208 , n359305 , n359306 , n359307 , n359308 , n359309 , n359310 , n359311 , n359312 , 
 n39217 , n39218 , n359315 , n359316 , n359317 , n359318 , n359319 , n359320 , n359321 , n359322 , 
 n39227 , n359324 , n359325 , n359326 , n359327 , n39232 , n359329 , n39234 , n359331 , n359332 , 
 n39237 , n359334 , n39239 , n359336 , n359337 , n39242 , n359339 , n359340 , n359341 , n359342 , 
 n359343 , n359344 , n359345 , n359346 , n359347 , n359348 , n359349 , n359350 , n359351 , n39256 , 
 n39257 , n359354 , n39259 , n39260 , n359357 , n359358 , n359359 , n359360 , n39265 , n359362 , 
 n359363 , n359364 , n359365 , n359366 , n359367 , n359368 , n39273 , n359370 , n359371 , n39276 , 
 n359373 , n359374 , n39279 , n359376 , n359377 , n39282 , n39283 , n359380 , n359381 , n39286 , 
 n359383 , n359384 , n39289 , n359386 , n359387 , n359388 , n39293 , n359390 , n359391 , n359392 , 
 n359393 , n359394 , n359395 , n359396 , n39301 , n359398 , n359399 , n359400 , n359401 , n359402 , 
 n359403 , n359404 , n359405 , n359406 , n359407 , n39312 , n359409 , n359410 , n39315 , n39316 , 
 n359413 , n359414 , n359415 , n359416 , n359417 , n359418 , n359419 , n359420 , n39325 , n359422 , 
 n39327 , n359424 , n359425 , n359426 , n39331 , n39332 , n359429 , n359430 , n359431 , n359432 , 
 n39337 , n359434 , n39339 , n359436 , n359437 , n359438 , n359439 , n359440 , n359441 , n39346 , 
 n359443 , n359444 , n359445 , n39350 , n359447 , n359448 , n359449 , n359450 , n359451 , n359452 , 
 n39357 , n359454 , n359455 , n39360 , n39361 , n359458 , n359459 , n39364 , n359461 , n359462 , 
 n359463 , n359464 , n359465 , n359466 , n39371 , n359468 , n39373 , n359470 , n359471 , n359472 , 
 n359473 , n39378 , n359475 , n359476 , n39381 , n359478 , n359479 , n359480 , n359481 , n359482 , 
 n359483 , n359484 , n359485 , n359486 , n359487 , n359488 , n359489 , n359490 , n359491 , n359492 , 
 n359493 , n359494 , n359495 , n359496 , n359497 , n359498 , n359499 , n359500 , n359501 , n359502 , 
 n39407 , n359504 , n359505 , n39410 , n359507 , n359508 , n359509 , n39414 , n359511 , n359512 , 
 n359513 , n359514 , n359515 , n359516 , n359517 , n359518 , n359519 , n39424 , n39425 , n359522 , 
 n359523 , n359524 , n39429 , n359526 , n359527 , n39432 , n359529 , n359530 , n359531 , n359532 , 
 n39437 , n359534 , n359535 , n359536 , n359537 , n359538 , n39443 , n359540 , n359541 , n359542 , 
 n359543 , n39448 , n39449 , n359546 , n359547 , n39452 , n359549 , n39454 , n39455 , n359552 , 
 n359553 , n39458 , n359555 , n39460 , n359557 , n39462 , n359559 , n359560 , n39465 , n359562 , 
 n39467 , n359564 , n359565 , n359566 , n39471 , n359568 , n39473 , n39474 , n359571 , n359572 , 
 n39477 , n359574 , n359575 , n359576 , n359577 , n359578 , n39483 , n359580 , n359581 , n39486 , 
 n359583 , n359584 , n359585 , n39490 , n359587 , n39492 , n39493 , n359590 , n39495 , n39496 , 
 n359593 , n39498 , n359595 , n359596 , n359597 , n39502 , n359599 , n359600 , n39505 , n359602 , 
 n359603 , n359604 , n39509 , n359606 , n39511 , n39512 , n359609 , n359610 , n39515 , n359612 , 
 n39517 , n359614 , n359615 , n39520 , n39521 , n39522 , n359619 , n359620 , n39525 , n359622 , 
 n359623 , n359624 , n359625 , n359626 , n39531 , n359628 , n359629 , n39534 , n359631 , n359632 , 
 n39537 , n359634 , n39539 , n359636 , n39541 , n39542 , n359639 , n359640 , n359641 , n39546 , 
 n39547 , n359644 , n359645 , n359646 , n359647 , n359648 , n359649 , n39554 , n359651 , n359652 , 
 n39557 , n359654 , n359655 , n39560 , n39561 , n39562 , n359659 , n359660 , n39565 , n39566 , 
 n39567 , n359664 , n359665 , n39570 , n39571 , n359668 , n359669 , n39574 , n359671 , n39576 , 
 n359673 , n39578 , n39579 , n359676 , n39581 , n39582 , n359679 , n359680 , n39585 , n359682 , 
 n359683 , n39588 , n359685 , n359686 , n39591 , n39592 , n359689 , n359690 , n359691 , n359692 , 
 n359693 , n359694 , n359695 , n359696 , n39601 , n359698 , n39603 , n359700 , n39605 , n39606 , 
 n359703 , n359704 , n39609 , n359706 , n359707 , n359708 , n359709 , n359710 , n359711 , n359712 , 
 n359713 , n39618 , n359715 , n39620 , n39621 , n39622 , n359719 , n359720 , n359721 , n359722 , 
 n359723 , n359724 , n359725 , n39630 , n359727 , n359728 , n359729 , n359730 , n359731 , n359732 , 
 n359733 , n39638 , n359735 , n39640 , n39641 , n39642 , n359739 , n39644 , n359741 , n359742 , 
 n359743 , n39648 , n359745 , n359746 , n359747 , n359748 , n359749 , n359750 , n359751 , n359752 , 
 n359753 , n359754 , n359755 , n359756 , n39655 , n359758 , n359759 , n39658 , n39659 , n359762 , 
 n359763 , n39662 , n39663 , n359766 , n359767 , n359768 , n359769 , n359770 , n39666 , n39667 , 
 n359773 , n359774 , n39670 , n39671 , n39672 , n359778 , n359779 , n39675 , n359781 , n359782 , 
 n359783 , n359784 , n359785 , n39681 , n359787 , n359788 , n359789 , n359790 , n359791 , n359792 , 
 n359793 , n359794 , n39690 , n359796 , n359797 , n359798 , n39694 , n359800 , n359801 , n359802 , 
 n359803 , n359804 , n39700 , n39701 , n359807 , n39703 , n359809 , n359810 , n39706 , n39707 , 
 n359813 , n39709 , n359815 , n359816 , n359817 , n359818 , n359819 , n359820 , n359821 , n359822 , 
 n359823 , n359824 , n359825 , n359826 , n359827 , n359828 , n39724 , n359830 , n39726 , n359832 , 
 n39728 , n359834 , n359835 , n359836 , n39732 , n359838 , n359839 , n39735 , n359841 , n359842 , 
 n359843 , n359844 , n359845 , n359846 , n359847 , n359848 , n359849 , n39745 , n359851 , n359852 , 
 n39748 , n39749 , n359855 , n359856 , n359857 , n39753 , n39754 , n359860 , n359861 , n39757 , 
 n39758 , n359864 , n359865 , n359866 , n39762 , n359868 , n359869 , n359870 , n359871 , n359872 , 
 n39768 , n359874 , n359875 , n39771 , n359877 , n359878 , n359879 , n39775 , n359881 , n359882 , 
 n359883 , n39779 , n359885 , n359886 , n39782 , n39783 , n39784 , n359890 , n359891 , n359892 , 
 n359893 , n359894 , n359895 , n359896 , n359897 , n39790 , n359899 , n39792 , n359901 , n359902 , 
 n359903 , n359904 , n359905 , n359906 , n359907 , n359908 , n359909 , n359910 , n359911 , n359912 , 
 n359913 , n359914 , n359915 , n359916 , n359917 , n359918 , n359919 , n359920 , n359921 , n39814 , 
 n39815 , n39816 , n359925 , n359926 , n359927 , n359928 , n39821 , n39822 , n359931 , n39824 , 
 n359933 , n39826 , n359935 , n359936 , n359937 , n39830 , n359939 , n39832 , n39833 , n39834 , 
 n359943 , n359944 , n359945 , n359946 , n359947 , n359948 , n359949 , n359950 , n39843 , n39844 , 
 n359953 , n359954 , n359955 , n39848 , n39849 , n359958 , n359959 , n39852 , n39853 , n39854 , 
 n359963 , n39856 , n39857 , n359966 , n39859 , n39860 , n39861 , n359970 , n39863 , n39864 , 
 n359973 , n359974 , n39867 , n359976 , n359977 , n39870 , n359979 , n359980 , n359981 , n39874 , 
 n359983 , n359984 , n39877 , n39878 , n359987 , n39880 , n39881 , n359990 , n359991 , n359992 , 
 n359993 , n359994 , n359995 , n359996 , n39889 , n39890 , n39891 , n360000 , n39893 , n360002 , 
 n360003 , n39896 , n39897 , n360006 , n39899 , n360008 , n360009 , n360010 , n360011 , n360012 , 
 n360013 , n360014 , n360015 , n360016 , n39909 , n360018 , n360019 , n360020 , n360021 , n360022 , 
 n360023 , n360024 , n360025 , n360026 , n360027 , n39920 , n39921 , n360030 , n39923 , n360032 , 
 n360033 , n39926 , n360035 , n360036 , n39929 , n360038 , n360039 , n39932 , n360041 , n39934 , 
 n360043 , n360044 , n39937 , n360046 , n360047 , n360048 , n360049 , n360050 , n360051 , n360052 , 
 n39945 , n39946 , n360055 , n39948 , n39949 , n39950 , n39951 , n39952 , n360061 , n39954 , 
 n360063 , n360064 , n360065 , n360066 , n360067 , n360068 , n360069 , n39962 , n39963 , n360072 , 
 n39965 , n39966 , n360075 , n39968 , n360077 , n360078 , n39971 , n39972 , n360081 , n39974 , 
 n360083 , n39976 , n39977 , n360086 , n39979 , n39980 , n39981 , n360090 , n360091 , n360092 , 
 n360093 , n360094 , n360095 , n360096 , n360097 , n360098 , n39991 , n360100 , n39993 , n360102 , 
 n360103 , n39996 , n360105 , n39998 , n39999 , n360108 , n40001 , n360110 , n40003 , n40004 , 
 n40005 , n360114 , n40007 , n360116 , n360117 , n40010 , n360119 , n360120 , n360121 , n360122 , 
 n360123 , n40016 , n360125 , n360126 , n360127 , n360128 , n360129 , n360130 , n360131 , n360132 , 
 n360133 , n360134 , n40027 , n360136 , n360137 , n360138 , n360139 , n360140 , n40033 , n360142 , 
 n360143 , n40036 , n360145 , n360146 , n40039 , n360148 , n40041 , n360150 , n40043 , n360152 , 
 n360153 , n360154 , n360155 , n360156 , n360157 , n360158 , n360159 , n360160 , n360161 , n360162 , 
 n40055 , n360164 , n360165 , n40058 , n40059 , n360168 , n40061 , n40062 , n360171 , n360172 , 
 n360173 , n360174 , n360175 , n40068 , n360177 , n40070 , n40071 , n360180 , n40073 , n360182 , 
 n360183 , n360184 , n360185 , n360186 , n360187 , n40080 , n360189 , n360190 , n40083 , n360192 , 
 n360193 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , 
 n360203 , n40096 , n40097 , n360206 , n360207 , n40100 , n360209 , n360210 , n40103 , n360212 , 
 n360213 , n40106 , n360215 , n40108 , n40109 , n360218 , n360219 , n40112 , n360221 , n360222 , 
 n360223 , n360224 , n360225 , n40118 , n360227 , n40120 , n360229 , n360230 , n360231 , n360232 , 
 n360233 , n360234 , n360235 , n360236 , n360237 , n360238 , n360239 , n360240 , n360241 , n360242 , 
 n360243 , n360244 , n360245 , n40138 , n360247 , n360248 , n360249 , n360250 , n360251 , n40144 , 
 n360253 , n360254 , n360255 , n360256 , n360257 , n40150 , n40151 , n360260 , n360261 , n360262 , 
 n360263 , n40156 , n360265 , n360266 , n40159 , n360268 , n360269 , n40162 , n360271 , n360272 , 
 n40165 , n360274 , n360275 , n360276 , n360277 , n360278 , n360279 , n40172 , n360281 , n360282 , 
 n40175 , n360284 , n40177 , n40178 , n360287 , n40180 , n40181 , n40182 , n360291 , n360292 , 
 n360293 , n360294 , n40187 , n360296 , n360297 , n40190 , n360299 , n360300 , n360301 , n360302 , 
 n360303 , n40196 , n360305 , n360306 , n40199 , n360308 , n40201 , n40202 , n40203 , n360312 , 
 n40205 , n360314 , n40207 , n360316 , n40209 , n360318 , n360319 , n360320 , n360321 , n360322 , 
 n360323 , n360324 , n40217 , n360326 , n40219 , n40220 , n360329 , n360330 , n360331 , n360332 , 
 n360333 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n360341 , n360342 , 
 n360343 , n360344 , n360345 , n360346 , n360347 , n360348 , n360349 , n360350 , n360351 , n360352 , 
 n360353 , n360354 , n360355 , n360356 , n360357 , n40235 , n360359 , n360360 , n360361 , n40239 , 
 n360363 , n360364 , n40242 , n360366 , n360367 , n40245 , n360369 , n360370 , n40248 , n360372 , 
 n360373 , n40251 , n40252 , n360376 , n360377 , n40255 , n360379 , n360380 , n360381 , n360382 , 
 n360383 , n360384 , n40262 , n360386 , n360387 , n360388 , n360389 , n40267 , n40268 , n40269 , 
 n40270 , n40271 , n360395 , n40273 , n360397 , n40275 , n360399 , n360400 , n360401 , n360402 , 
 n360403 , n360404 , n360405 , n360406 , n360407 , n360408 , n40286 , n40287 , n40288 , n360412 , 
 n360413 , n40291 , n360415 , n360416 , n360417 , n360418 , n360419 , n360420 , n360421 , n360422 , 
 n360423 , n360424 , n360425 , n360426 , n40304 , n40305 , n40306 , n360430 , n360431 , n360432 , 
 n360433 , n360434 , n360435 , n360436 , n360437 , n360438 , n360439 , n40317 , n360441 , n360442 , 
 n360443 , n360444 , n360445 , n40323 , n40324 , n40325 , n360449 , n40327 , n40328 , n360452 , 
 n360453 , n40331 , n360455 , n360456 , n360457 , n360458 , n360459 , n360460 , n40338 , n40339 , 
 n360463 , n40341 , n360465 , n360466 , n360467 , n360468 , n360469 , n360470 , n360471 , n360472 , 
 n40350 , n360474 , n40352 , n360476 , n40354 , n40355 , n360479 , n40357 , n40358 , n40359 , 
 n360483 , n360484 , n360485 , n40363 , n40364 , n40365 , n40366 , n40367 , n360491 , n360492 , 
 n360493 , n360494 , n40372 , n360496 , n360497 , n360498 , n360499 , n360500 , n40378 , n360502 , 
 n360503 , n40381 , n360505 , n360506 , n360507 , n360508 , n360509 , n360510 , n360511 , n360512 , 
 n360513 , n360514 , n360515 , n360516 , n360517 , n360518 , n360519 , n360520 , n360521 , n360522 , 
 n360523 , n360524 , n360525 , n40403 , n40404 , n40405 , n360529 , n40407 , n40408 , n360532 , 
 n360533 , n40411 , n360535 , n360536 , n40414 , n360538 , n40416 , n360540 , n360541 , n360542 , 
 n360543 , n360544 , n360545 , n40423 , n360547 , n360548 , n40426 , n360550 , n360551 , n360552 , 
 n40430 , n360554 , n40432 , n360556 , n40434 , n40435 , n360559 , n360560 , n40438 , n360562 , 
 n360563 , n40441 , n360565 , n360566 , n40444 , n40445 , n40446 , n360570 , n360571 , n360572 , 
 n360573 , n360574 , n360575 , n360576 , n360577 , n360578 , n40456 , n360580 , n360581 , n360582 , 
 n360583 , n40461 , n360585 , n40463 , n360587 , n40465 , n360589 , n40467 , n360591 , n360592 , 
 n360593 , n40471 , n360595 , n40473 , n40474 , n40475 , n360599 , n360600 , n360601 , n360602 , 
 n360603 , n360604 , n360605 , n360606 , n40484 , n360608 , n360609 , n360610 , n360611 , n40489 , 
 n360613 , n360614 , n360615 , n360616 , n360617 , n360618 , n360619 , n40497 , n360621 , n40499 , 
 n360623 , n360624 , n360625 , n360626 , n360627 , n360628 , n360629 , n360630 , n360631 , n360632 , 
 n360633 , n360634 , n40512 , n360636 , n360637 , n40515 , n40516 , n360640 , n360641 , n360642 , 
 n360643 , n40521 , n360645 , n360646 , n360647 , n360648 , n360649 , n360650 , n360651 , n360652 , 
 n360653 , n360654 , n360655 , n360656 , n360657 , n360658 , n360659 , n360660 , n40538 , n360662 , 
 n40540 , n360664 , n360665 , n360666 , n360667 , n360668 , n360669 , n360670 , n360671 , n360672 , 
 n360673 , n360674 , n360675 , n360676 , n360677 , n40555 , n360679 , n360680 , n40558 , n360682 , 
 n360683 , n360684 , n360685 , n360686 , n360687 , n360688 , n40566 , n360690 , n360691 , n360692 , 
 n40570 , n40571 , n360695 , n40573 , n360697 , n360698 , n40576 , n360700 , n360701 , n40579 , 
 n360703 , n360704 , n360705 , n360706 , n360707 , n360708 , n360709 , n360710 , n360711 , n360712 , 
 n360713 , n360714 , n40589 , n360716 , n40591 , n360718 , n40593 , n360720 , n360721 , n360722 , 
 n360723 , n360724 , n360725 , n40600 , n360727 , n360728 , n40603 , n360730 , n360731 , n40606 , 
 n360733 , n360734 , n40609 , n360736 , n40611 , n40612 , n360739 , n360740 , n360741 , n360742 , 
 n360743 , n360744 , n40619 , n360746 , n360747 , n360748 , n360749 , n360750 , n360751 , n360752 , 
 n360753 , n360754 , n360755 , n40630 , n360757 , n360758 , n360759 , n360760 , n40635 , n360762 , 
 n360763 , n360764 , n360765 , n360766 , n360767 , n360768 , n360769 , n360770 , n360771 , n360772 , 
 n360773 , n360774 , n360775 , n360776 , n360777 , n360778 , n360779 , n360780 , n40653 , n360782 , 
 n360783 , n360784 , n360785 , n360786 , n360787 , n360788 , n40658 , n40659 , n40660 , n360792 , 
 n360793 , n360794 , n360795 , n360796 , n360797 , n360798 , n360799 , n360800 , n360801 , n360802 , 
 n360803 , n360804 , n360805 , n40675 , n360807 , n40677 , n40678 , n40679 , n40680 , n360812 , 
 n40682 , n360814 , n360815 , n40685 , n360817 , n360818 , n360819 , n360820 , n360821 , n360822 , 
 n40692 , n360824 , n360825 , n40695 , n40696 , n40697 , n360829 , n40699 , n40700 , n360832 , 
 n360833 , n40703 , n360835 , n360836 , n360837 , n360838 , n360839 , n40709 , n40710 , n360842 , 
 n360843 , n40713 , n360845 , n360846 , n360847 , n360848 , n360849 , n360850 , n360851 , n360852 , 
 n360853 , n40723 , n360855 , n40725 , n360857 , n360858 , n360859 , n360860 , n360861 , n360862 , 
 n360863 , n360864 , n360865 , n360866 , n40736 , n360868 , n40738 , n40739 , n40740 , n40741 , 
 n40742 , n360874 , n360875 , n360876 , n40746 , n360878 , n360879 , n40749 , n40750 , n360882 , 
 n40752 , n40753 , n360885 , n360886 , n40756 , n360888 , n360889 , n40759 , n360891 , n360892 , 
 n360893 , n360894 , n360895 , n360896 , n360897 , n360898 , n360899 , n360900 , n360901 , n360902 , 
 n360903 , n360904 , n360905 , n360906 , n360907 , n360908 , n360909 , n360910 , n360911 , n360912 , 
 n360913 , n360914 , n360915 , n40782 , n360917 , n360918 , n40785 , n360920 , n360921 , n40788 , 
 n360923 , n360924 , n360925 , n360926 , n360927 , n40794 , n40795 , n360930 , n40797 , n40798 , 
 n360933 , n360934 , n40801 , n360936 , n360937 , n360938 , n360939 , n360940 , n40807 , n40808 , 
 n360943 , n40810 , n360945 , n360946 , n360947 , n360948 , n360949 , n360950 , n360951 , n360952 , 
 n360953 , n360954 , n360955 , n360956 , n40823 , n360958 , n360959 , n360960 , n360961 , n360962 , 
 n40829 , n40830 , n40831 , n360966 , n360967 , n40834 , n360969 , n360970 , n360971 , n40838 , 
 n360973 , n360974 , n40841 , n360976 , n360977 , n40844 , n360979 , n40846 , n40847 , n40848 , 
 n40849 , n40850 , n360985 , n40852 , n360987 , n40854 , n360989 , n40856 , n40857 , n360992 , 
 n360993 , n40860 , n360995 , n360996 , n40863 , n360998 , n360999 , n40866 , n40867 , n361002 , 
 n40869 , n361004 , n40871 , n361006 , n361007 , n40874 , n361009 , n40876 , n361011 , n40878 , 
 n361013 , n361014 , n40881 , n361016 , n361017 , n40884 , n361019 , n40886 , n361021 , n361022 , 
 n361023 , n361024 , n40891 , n361026 , n40893 , n361028 , n40895 , n361030 , n40897 , n361032 , 
 n40899 , n361034 , n361035 , n361036 , n361037 , n361038 , n361039 , n361040 , n361041 , n361042 , 
 n40909 , n361044 , n40911 , n361046 , n361047 , n40914 , n361049 , n361050 , n361051 , n361052 , 
 n361053 , n40920 , n40921 , n361056 , n40923 , n361058 , n40925 , n361060 , n361061 , n40928 , 
 n361063 , n361064 , n361065 , n361066 , n361067 , n40934 , n361069 , n361070 , n361071 , n40938 , 
 n361073 , n361074 , n361075 , n361076 , n40943 , n361078 , n40945 , n361080 , n361081 , n361082 , 
 n361083 , n40950 , n40951 , n361086 , n40953 , n361088 , n361089 , n361090 , n361091 , n40958 , 
 n361093 , n361094 , n361095 , n361096 , n361097 , n361098 , n361099 , n361100 , n361101 , n361102 , 
 n361103 , n361104 , n361105 , n361106 , n361107 , n361108 , n361109 , n40976 , n40977 , n361112 , 
 n361113 , n361114 , n361115 , n361116 , n361117 , n361118 , n361119 , n361120 , n361121 , n361122 , 
 n40989 , n40990 , n361125 , n40992 , n361127 , n361128 , n361129 , n361130 , n361131 , n361132 , 
 n40999 , n361134 , n41001 , n41002 , n361137 , n361138 , n41005 , n361140 , n361141 , n41008 , 
 n361143 , n361144 , n41011 , n41012 , n361147 , n41014 , n361149 , n41016 , n361151 , n361152 , 
 n361153 , n361154 , n361155 , n361156 , n361157 , n361158 , n361159 , n361160 , n361161 , n361162 , 
 n361163 , n361164 , n361165 , n361166 , n41033 , n361168 , n361169 , n361170 , n41037 , n41038 , 
 n361173 , n361174 , n361175 , n361176 , n41043 , n361178 , n361179 , n361180 , n361181 , n361182 , 
 n41049 , n361184 , n361185 , n361186 , n361187 , n361188 , n361189 , n361190 , n361191 , n361192 , 
 n41059 , n361194 , n361195 , n41062 , n361197 , n41064 , n361199 , n361200 , n41067 , n361202 , 
 n361203 , n361204 , n361205 , n361206 , n41073 , n361208 , n361209 , n361210 , n361211 , n41078 , 
 n41079 , n41080 , n361215 , n41082 , n41083 , n361218 , n41085 , n361220 , n361221 , n361222 , 
 n41089 , n361224 , n361225 , n41092 , n361227 , n361228 , n361229 , n361230 , n361231 , n361232 , 
 n41099 , n361234 , n361235 , n361236 , n361237 , n361238 , n361239 , n361240 , n361241 , n41108 , 
 n361243 , n361244 , n361245 , n361246 , n361247 , n361248 , n41115 , n361250 , n361251 , n361252 , 
 n41119 , n361254 , n361255 , n361256 , n361257 , n361258 , n361259 , n361260 , n361261 , n361262 , 
 n361263 , n361264 , n361265 , n361266 , n361267 , n361268 , n361269 , n361270 , n41132 , n41133 , 
 n361273 , n361274 , n361275 , n361276 , n41138 , n361278 , n361279 , n41141 , n361281 , n361282 , 
 n361283 , n361284 , n361285 , n361286 , n361287 , n41149 , n361289 , n361290 , n41152 , n361292 , 
 n361293 , n361294 , n41156 , n361296 , n361297 , n361298 , n361299 , n361300 , n361301 , n361302 , 
 n361303 , n361304 , n361305 , n361306 , n361307 , n361308 , n361309 , n361310 , n361311 , n41173 , 
 n361313 , n41175 , n41176 , n361316 , n41178 , n361318 , n41180 , n361320 , n361321 , n361322 , 
 n361323 , n361324 , n41186 , n361326 , n361327 , n361328 , n361329 , n361330 , n361331 , n41193 , 
 n361333 , n361334 , n361335 , n361336 , n361337 , n41199 , n361339 , n41201 , n361341 , n41203 , 
 n361343 , n361344 , n361345 , n361346 , n361347 , n361348 , n361349 , n361350 , n361351 , n41213 , 
 n41214 , n361354 , n361355 , n41217 , n361357 , n361358 , n41220 , n41221 , n361361 , n41223 , 
 n361363 , n361364 , n41226 , n361366 , n361367 , n41229 , n361369 , n361370 , n361371 , n361372 , 
 n361373 , n361374 , n41236 , n361376 , n361377 , n361378 , n361379 , n361380 , n41242 , n361382 , 
 n361383 , n361384 , n361385 , n361386 , n41248 , n361388 , n361389 , n361390 , n41252 , n41253 , 
 n361393 , n361394 , n361395 , n361396 , n41258 , n361398 , n361399 , n41261 , n361401 , n361402 , 
 n41264 , n41265 , n361405 , n41267 , n41268 , n361408 , n361409 , n41271 , n361411 , n361412 , 
 n41274 , n361414 , n361415 , n41277 , n361417 , n361418 , n41280 , n361420 , n361421 , n361422 , 
 n361423 , n41285 , n361425 , n361426 , n361427 , n361428 , n361429 , n361430 , n361431 , n361432 , 
 n361433 , n41295 , n361435 , n41297 , n361437 , n361438 , n361439 , n361440 , n41302 , n361442 , 
 n41304 , n361444 , n361445 , n41307 , n361447 , n41309 , n361449 , n361450 , n41312 , n41313 , 
 n361453 , n41315 , n361455 , n361456 , n41318 , n361458 , n361459 , n361460 , n361461 , n361462 , 
 n41324 , n41325 , n361465 , n41327 , n361467 , n361468 , n41330 , n361470 , n361471 , n361472 , 
 n361473 , n361474 , n361475 , n361476 , n361477 , n361478 , n361479 , n361480 , n361481 , n361482 , 
 n361483 , n361484 , n41346 , n361486 , n361487 , n361488 , n361489 , n361490 , n361491 , n361492 , 
 n361493 , n361494 , n361495 , n41354 , n361497 , n41356 , n361499 , n361500 , n361501 , n41360 , 
 n361503 , n361504 , n41363 , n361506 , n361507 , n41366 , n361509 , n41368 , n361511 , n41370 , 
 n41371 , n361514 , n361515 , n41374 , n361517 , n361518 , n361519 , n361520 , n361521 , n361522 , 
 n361523 , n361524 , n41383 , n41384 , n41385 , n41386 , n361529 , n361530 , n361531 , n361532 , 
 n361533 , n361534 , n361535 , n361536 , n361537 , n361538 , n361539 , n361540 , n361541 , n361542 , 
 n361543 , n41402 , n361545 , n361546 , n41405 , n41406 , n361549 , n361550 , n361551 , n361552 , 
 n361553 , n361554 , n361555 , n361556 , n361557 , n41416 , n41417 , n41418 , n41419 , n41420 , 
 n361563 , n361564 , n41423 , n361566 , n361567 , n41426 , n41427 , n41428 , n41429 , n41430 , 
 n361573 , n361574 , n41433 , n361576 , n361577 , n41436 , n361579 , n361580 , n361581 , n361582 , 
 n41441 , n361584 , n361585 , n361586 , n41445 , n41446 , n41447 , n41448 , n361591 , n361592 , 
 n41451 , n41452 , n361595 , n41454 , n361597 , n361598 , n41457 , n361600 , n361601 , n361602 , 
 n361603 , n361604 , n361605 , n361606 , n361607 , n361608 , n361609 , n361610 , n361611 , n361612 , 
 n361613 , n41472 , n361615 , n41474 , n361617 , n361618 , n361619 , n361620 , n361621 , n41480 , 
 n41481 , n41482 , n361625 , n361626 , n41485 , n361628 , n361629 , n361630 , n361631 , n361632 , 
 n41491 , n361634 , n361635 , n41494 , n361637 , n361638 , n361639 , n361640 , n361641 , n361642 , 
 n361643 , n361644 , n41503 , n361646 , n361647 , n361648 , n361649 , n41508 , n361651 , n361652 , 
 n361653 , n361654 , n361655 , n361656 , n41515 , n361658 , n41517 , n361660 , n361661 , n361662 , 
 n361663 , n361664 , n361665 , n41524 , n361667 , n361668 , n41527 , n41528 , n361671 , n361672 , 
 n361673 , n361674 , n361675 , n41534 , n361677 , n361678 , n361679 , n361680 , n361681 , n41540 , 
 n361683 , n361684 , n361685 , n361686 , n361687 , n41546 , n41547 , n361690 , n361691 , n361692 , 
 n41551 , n361694 , n41553 , n41554 , n361697 , n361698 , n41557 , n361700 , n361701 , n361702 , 
 n361703 , n361704 , n41563 , n361706 , n41565 , n361708 , n41567 , n361710 , n41569 , n361712 , 
 n361713 , n361714 , n41573 , n361716 , n361717 , n361718 , n361719 , n361720 , n361721 , n361722 , 
 n41581 , n41582 , n361725 , n361726 , n41585 , n361728 , n361729 , n41588 , n41589 , n361732 , 
 n41591 , n361734 , n361735 , n361736 , n41595 , n361738 , n361739 , n41598 , n41599 , n361742 , 
 n41601 , n361744 , n41603 , n361746 , n41605 , n361748 , n41607 , n361750 , n361751 , n361752 , 
 n361753 , n361754 , n41613 , n361756 , n41615 , n41616 , n41617 , n361760 , n361761 , n361762 , 
 n361763 , n41622 , n41623 , n361766 , n41625 , n41626 , n41627 , n41628 , n41629 , n361772 , 
 n41631 , n361774 , n41633 , n361776 , n361777 , n41636 , n361779 , n41638 , n361781 , n41640 , 
 n41641 , n41642 , n361785 , n41644 , n361787 , n41646 , n41647 , n361790 , n361791 , n41650 , 
 n361793 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n361800 , n41659 , n361802 , 
 n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n361809 , n41668 , n361811 , n361812 , 
 n361813 , n361814 , n361815 , n361816 , n361817 , n361818 , n361819 , n361820 , n361821 , n361822 , 
 n361823 , n361824 , n361825 , n361826 , n41685 , n361828 , n361829 , n361830 , n41689 , n361832 , 
 n361833 , n41692 , n361835 , n361836 , n41695 , n361838 , n361839 , n361840 , n361841 , n361842 , 
 n41701 , n41702 , n361845 , n41704 , n361847 , n361848 , n41707 , n361850 , n361851 , n361852 , 
 n361853 , n361854 , n361855 , n41714 , n361857 , n361858 , n361859 , n41718 , n361861 , n361862 , 
 n361863 , n361864 , n361865 , n41724 , n361867 , n41726 , n361869 , n361870 , n41729 , n361872 , 
 n361873 , n361874 , n361875 , n361876 , n41735 , n361878 , n361879 , n361880 , n361881 , n361882 , 
 n361883 , n361884 , n361885 , n361886 , n361887 , n361888 , n361889 , n361890 , n361891 , n361892 , 
 n361893 , n361894 , n361895 , n361896 , n361897 , n361898 , n361899 , n361900 , n361901 , n361902 , 
 n361903 , n361904 , n361905 , n41764 , n361907 , n361908 , n361909 , n361910 , n361911 , n41770 , 
 n41771 , n41772 , n361915 , n41774 , n361917 , n41776 , n41777 , n41778 , n361921 , n361922 , 
 n361923 , n41782 , n41783 , n361926 , n361927 , n361928 , n361929 , n361930 , n361931 , n361932 , 
 n361933 , n361934 , n41793 , n361936 , n41795 , n361938 , n41797 , n41798 , n41799 , n361942 , 
 n41801 , n361944 , n41803 , n41804 , n361947 , n361948 , n41807 , n361950 , n361951 , n41810 , 
 n361953 , n361954 , n361955 , n361956 , n361957 , n41816 , n361959 , n41818 , n41819 , n361962 , 
 n361963 , n361964 , n361965 , n361966 , n361967 , n361968 , n41827 , n361970 , n361971 , n41830 , 
 n41831 , n361974 , n361975 , n41834 , n41835 , n41836 , n361979 , n361980 , n361981 , n361982 , 
 n41841 , n361984 , n361985 , n41844 , n361987 , n361988 , n41847 , n361990 , n361991 , n361992 , 
 n41851 , n361994 , n361995 , n41854 , n361997 , n361998 , n41857 , n41858 , n362001 , n362002 , 
 n41861 , n41862 , n362005 , n41864 , n362007 , n362008 , n41867 , n41868 , n41869 , n362012 , 
 n362013 , n362014 , n362015 , n362016 , n41875 , n362018 , n362019 , n362020 , n362021 , n41880 , 
 n41881 , n41882 , n362025 , n41884 , n362027 , n362028 , n41887 , n362030 , n362031 , n41890 , 
 n362033 , n41892 , n362035 , n41894 , n362037 , n362038 , n362039 , n41898 , n362041 , n41900 , 
 n41901 , n362044 , n362045 , n362046 , n41905 , n362048 , n41907 , n362050 , n362051 , n362052 , 
 n41911 , n362054 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n362061 , n362062 , 
 n362063 , n362064 , n362065 , n362066 , n362067 , n362068 , n362069 , n362070 , n362071 , n362072 , 
 n41931 , n41932 , n362075 , n362076 , n41935 , n362078 , n41937 , n362080 , n362081 , n362082 , 
 n41941 , n362084 , n362085 , n362086 , n41945 , n41946 , n362089 , n362090 , n362091 , n362092 , 
 n362093 , n362094 , n362095 , n362096 , n362097 , n41956 , n362099 , n362100 , n41959 , n362102 , 
 n362103 , n41962 , n362105 , n362106 , n41965 , n362108 , n362109 , n362110 , n362111 , n362112 , 
 n362113 , n41972 , n41973 , n362116 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , 
 n41981 , n41982 , n41983 , n41984 , n362127 , n41986 , n41987 , n362130 , n362131 , n41990 , 
 n362133 , n41992 , n362135 , n362136 , n362137 , n362138 , n362139 , n362140 , n362141 , n41999 , 
 n362143 , n362144 , n362145 , n362146 , n362147 , n362148 , n362149 , n362150 , n362151 , n362152 , 
 n362153 , n362154 , n362155 , n42011 , n42012 , n42013 , n42014 , n362160 , n42016 , n42017 , 
 n362163 , n42019 , n42020 , n362166 , n42022 , n362168 , n362169 , n362170 , n362171 , n362172 , 
 n362173 , n42029 , n362175 , n362176 , n362177 , n362178 , n362179 , n362180 , n42036 , n42037 , 
 n362183 , n362184 , n42040 , n362186 , n362187 , n362188 , n362189 , n362190 , n362191 , n362192 , 
 n362193 , n362194 , n362195 , n362196 , n362197 , n362198 , n362199 , n362200 , n362201 , n362202 , 
 n362203 , n42059 , n362205 , n362206 , n362207 , n362208 , n362209 , n42065 , n362211 , n362212 , 
 n42068 , n362214 , n362215 , n42071 , n42072 , n362218 , n42074 , n42075 , n362221 , n42077 , 
 n42078 , n362224 , n362225 , n42081 , n42082 , n362228 , n42084 , n362230 , n362231 , n362232 , 
 n42088 , n362234 , n362235 , n42091 , n42092 , n362238 , n362239 , n362240 , n362241 , n362242 , 
 n362243 , n362244 , n362245 , n362246 , n362247 , n362248 , n362249 , n362250 , n42106 , n42107 , 
 n362253 , n362254 , n42110 , n362256 , n362257 , n42113 , n42114 , n362260 , n362261 , n362262 , 
 n362263 , n42119 , n362265 , n362266 , n362267 , n362268 , n42124 , n42125 , n362271 , n42127 , 
 n362273 , n42129 , n362275 , n42131 , n42132 , n362278 , n42134 , n362280 , n362281 , n42137 , 
 n362283 , n362284 , n362285 , n362286 , n362287 , n362288 , n362289 , n42145 , n42146 , n42147 , 
 n42148 , n42149 , n42150 , n362296 , n362297 , n362298 , n362299 , n362300 , n362301 , n362302 , 
 n362303 , n42159 , n362305 , n362306 , n362307 , n362308 , n362309 , n362310 , n362311 , n362312 , 
 n362313 , n362314 , n362315 , n42171 , n362317 , n362318 , n362319 , n362320 , n362321 , n362322 , 
 n362323 , n362324 , n362325 , n362326 , n362327 , n362328 , n362329 , n362330 , n362331 , n362332 , 
 n362333 , n362334 , n42190 , n362336 , n362337 , n362338 , n362339 , n362340 , n362341 , n362342 , 
 n362343 , n362344 , n362345 , n42201 , n42202 , n362348 , n42204 , n42205 , n362351 , n42207 , 
 n362353 , n42209 , n362355 , n362356 , n362357 , n42213 , n42214 , n362360 , n362361 , n42217 , 
 n362363 , n362364 , n362365 , n42221 , n362367 , n362368 , n42224 , n362370 , n362371 , n42227 , 
 n42228 , n42229 , n42230 , n362376 , n362377 , n42233 , n362379 , n362380 , n362381 , n42237 , 
 n362383 , n42239 , n362385 , n362386 , n42242 , n362388 , n362389 , n42245 , n362391 , n362392 , 
 n42248 , n362394 , n362395 , n42251 , n362397 , n362398 , n42254 , n362400 , n42256 , n362402 , 
 n362403 , n42259 , n362405 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n362412 , 
 n42268 , n362414 , n362415 , n362416 , n362417 , n362418 , n42274 , n362420 , n362421 , n362422 , 
 n362423 , n362424 , n362425 , n362426 , n362427 , n42283 , n362429 , n362430 , n42286 , n362432 , 
 n362433 , n42289 , n362435 , n362436 , n42292 , n362438 , n362439 , n42295 , n362441 , n362442 , 
 n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n362449 , n362450 , n362451 , n362452 , 
 n362453 , n362454 , n362455 , n362456 , n362457 , n362458 , n362459 , n362460 , n362461 , n362462 , 
 n362463 , n362464 , n362465 , n362466 , n362467 , n362468 , n362469 , n42325 , n362471 , n362472 , 
 n42328 , n362474 , n362475 , n42331 , n362477 , n42333 , n362479 , n362480 , n362481 , n362482 , 
 n42338 , n362484 , n362485 , n362486 , n362487 , n42343 , n362489 , n362490 , n362491 , n362492 , 
 n362493 , n362494 , n362495 , n362496 , n42352 , n362498 , n362499 , n42355 , n362501 , n362502 , 
 n362503 , n42359 , n42360 , n362506 , n362507 , n42363 , n362509 , n362510 , n42366 , n362512 , 
 n362513 , n362514 , n362515 , n362516 , n42372 , n42373 , n362519 , n42375 , n362521 , n362522 , 
 n362523 , n362524 , n42380 , n362526 , n362527 , n42383 , n362529 , n362530 , n42386 , n42387 , 
 n42388 , n362534 , n362535 , n42391 , n362537 , n362538 , n362539 , n362540 , n362541 , n42397 , 
 n362543 , n362544 , n42400 , n42401 , n362547 , n362548 , n362549 , n362550 , n42406 , n362552 , 
 n362553 , n362554 , n362555 , n362556 , n362557 , n362558 , n362559 , n362560 , n362561 , n362562 , 
 n362563 , n362564 , n362565 , n42421 , n362567 , n42423 , n362569 , n362570 , n362571 , n42427 , 
 n362573 , n362574 , n42430 , n42431 , n362577 , n362578 , n362579 , n362580 , n362581 , n362582 , 
 n362583 , n362584 , n362585 , n362586 , n362587 , n362588 , n42444 , n42445 , n362591 , n362592 , 
 n42448 , n362594 , n362595 , n362596 , n362597 , n42453 , n42454 , n42455 , n362601 , n42457 , 
 n362603 , n362604 , n362605 , n362606 , n362607 , n362608 , n42464 , n362610 , n362611 , n42467 , 
 n362613 , n362614 , n42470 , n362616 , n362617 , n42473 , n362619 , n362620 , n42476 , n42477 , 
 n362623 , n42479 , n362625 , n362626 , n42482 , n362628 , n362629 , n362630 , n362631 , n362632 , 
 n42488 , n42489 , n362635 , n362636 , n362637 , n362638 , n362639 , n42495 , n362641 , n362642 , 
 n42498 , n362644 , n362645 , n362646 , n362647 , n362648 , n362649 , n362650 , n362651 , n362652 , 
 n42508 , n362654 , n362655 , n362656 , n362657 , n362658 , n362659 , n362660 , n362661 , n362662 , 
 n362663 , n362664 , n42520 , n362666 , n362667 , n42523 , n362669 , n362670 , n42526 , n362672 , 
 n362673 , n362674 , n362675 , n362676 , n362677 , n362678 , n362679 , n362680 , n362681 , n362682 , 
 n362683 , n362684 , n362685 , n362686 , n362687 , n362688 , n362689 , n362690 , n362691 , n362692 , 
 n362693 , n362694 , n362695 , n42551 , n42552 , n362698 , n362699 , n362700 , n362701 , n362702 , 
 n42558 , n362704 , n362705 , n42561 , n362707 , n362708 , n42564 , n362710 , n362711 , n362712 , 
 n362713 , n362714 , n42570 , n42571 , n362717 , n362718 , n362719 , n362720 , n42576 , n362722 , 
 n362723 , n362724 , n362725 , n362726 , n362727 , n42583 , n362729 , n362730 , n362731 , n362732 , 
 n362733 , n362734 , n42590 , n362736 , n362737 , n42593 , n42594 , n42595 , n362741 , n362742 , 
 n362743 , n42599 , n362745 , n362746 , n362747 , n42603 , n362749 , n362750 , n42606 , n362752 , 
 n362753 , n362754 , n362755 , n362756 , n42612 , n42613 , n362759 , n42615 , n42616 , n362762 , 
 n362763 , n42619 , n362765 , n362766 , n362767 , n362768 , n362769 , n362770 , n362771 , n42627 , 
 n362773 , n362774 , n362775 , n362776 , n362777 , n362778 , n362779 , n362780 , n362781 , n362782 , 
 n362783 , n42639 , n42640 , n362786 , n362787 , n362788 , n362789 , n362790 , n42646 , n362792 , 
 n362793 , n362794 , n42650 , n362796 , n362797 , n42653 , n362799 , n42655 , n362801 , n42657 , 
 n362803 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n362810 , n362811 , n42667 , 
 n362813 , n362814 , n42670 , n362816 , n362817 , n362818 , n362819 , n362820 , n42676 , n362822 , 
 n362823 , n362824 , n362825 , n42681 , n362827 , n362828 , n42684 , n362830 , n362831 , n42687 , 
 n362833 , n362834 , n42690 , n362836 , n362837 , n42693 , n362839 , n362840 , n362841 , n362842 , 
 n362843 , n362844 , n362845 , n362846 , n362847 , n362848 , n362849 , n362850 , n42706 , n42707 , 
 n42708 , n42709 , n362855 , n362856 , n42712 , n362858 , n362859 , n362860 , n362861 , n42717 , 
 n362863 , n362864 , n362865 , n42721 , n362867 , n362868 , n362869 , n42725 , n362871 , n362872 , 
 n362873 , n362874 , n42730 , n362876 , n362877 , n42733 , n362879 , n42735 , n362881 , n362882 , 
 n42738 , n362884 , n362885 , n362886 , n362887 , n362888 , n42744 , n362890 , n362891 , n362892 , 
 n362893 , n362894 , n362895 , n362896 , n362897 , n362898 , n362899 , n362900 , n362901 , n362902 , 
 n362903 , n42759 , n42760 , n362906 , n42762 , n362908 , n362909 , n362910 , n362911 , n362912 , 
 n362913 , n362914 , n362915 , n362916 , n362917 , n362918 , n362919 , n362920 , n362921 , n362922 , 
 n42778 , n362924 , n362925 , n362926 , n42782 , n362928 , n362929 , n42785 , n362931 , n362932 , 
 n362933 , n42789 , n362935 , n362936 , n42792 , n362938 , n362939 , n362940 , n362941 , n362942 , 
 n362943 , n362944 , n362945 , n362946 , n362947 , n362948 , n362949 , n362950 , n362951 , n362952 , 
 n362953 , n362954 , n362955 , n42811 , n362957 , n42813 , n362959 , n42815 , n362961 , n362962 , 
 n42818 , n362964 , n362965 , n42821 , n362967 , n362968 , n42824 , n42825 , n362971 , n42827 , 
 n362973 , n362974 , n42830 , n362976 , n362977 , n42833 , n362979 , n362980 , n42836 , n362982 , 
 n362983 , n362984 , n362985 , n362986 , n362987 , n42843 , n362989 , n42845 , n42846 , n42847 , 
 n42848 , n42849 , n42850 , n42851 , n362997 , n362998 , n362999 , n363000 , n363001 , n363002 , 
 n42852 , n363004 , n363005 , n363006 , n42856 , n363008 , n363009 , n363010 , n363011 , n363012 , 
 n363013 , n363014 , n42864 , n363016 , n363017 , n42867 , n363019 , n42869 , n363021 , n363022 , 
 n363023 , n42873 , n363025 , n363026 , n363027 , n363028 , n42878 , n363030 , n363031 , n363032 , 
 n363033 , n363034 , n363035 , n363036 , n42886 , n363038 , n363039 , n42889 , n363041 , n42891 , 
 n363043 , n42893 , n42894 , n42895 , n42896 , n363048 , n42898 , n363050 , n363051 , n363052 , 
 n363053 , n42903 , n363055 , n363056 , n42906 , n363058 , n42908 , n363060 , n42910 , n42911 , 
 n363063 , n42913 , n363065 , n363066 , n42916 , n363068 , n363069 , n363070 , n363071 , n363072 , 
 n363073 , n363074 , n363075 , n42925 , n42926 , n363078 , n42928 , n42929 , n363081 , n363082 , 
 n363083 , n363084 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n363091 , n363092 , 
 n363093 , n363094 , n42944 , n42945 , n363097 , n42947 , n363099 , n363100 , n363101 , n42951 , 
 n363103 , n363104 , n363105 , n363106 , n363107 , n363108 , n42958 , n363110 , n363111 , n363112 , 
 n363113 , n363114 , n363115 , n363116 , n363117 , n363118 , n363119 , n363120 , n42970 , n363122 , 
 n363123 , n363124 , n363125 , n363126 , n42976 , n363128 , n42978 , n42979 , n42980 , n42981 , 
 n42982 , n42983 , n363135 , n42985 , n42986 , n363138 , n363139 , n42989 , n363141 , n363142 , 
 n42992 , n42993 , n42994 , n363146 , n363147 , n363148 , n363149 , n363150 , n363151 , n363152 , 
 n363153 , n363154 , n363155 , n363156 , n363157 , n363158 , n363159 , n363160 , n363161 , n363162 , 
 n363163 , n363164 , n363165 , n43015 , n363167 , n363168 , n363169 , n43019 , n363171 , n363172 , 
 n363173 , n363174 , n363175 , n363176 , n363177 , n363178 , n363179 , n363180 , n43030 , n43031 , 
 n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , 
 n363193 , n363194 , n43044 , n363196 , n363197 , n363198 , n363199 , n363200 , n363201 , n363202 , 
 n363203 , n363204 , n363205 , n363206 , n43051 , n363208 , n363209 , n363210 , n363211 , n43056 , 
 n363213 , n43058 , n363215 , n363216 , n43061 , n363218 , n43063 , n43064 , n363221 , n43066 , 
 n363223 , n363224 , n363225 , n363226 , n363227 , n363228 , n363229 , n363230 , n363231 , n363232 , 
 n363233 , n363234 , n363235 , n363236 , n43081 , n363238 , n43083 , n363240 , n43085 , n43086 , 
 n363243 , n363244 , n363245 , n363246 , n363247 , n363248 , n363249 , n363250 , n363251 , n363252 , 
 n363253 , n363254 , n363255 , n363256 , n363257 , n363258 , n43103 , n363260 , n363261 , n363262 , 
 n43107 , n363264 , n363265 , n363266 , n363267 , n363268 , n363269 , n363270 , n363271 , n363272 , 
 n43117 , n43118 , n363275 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , 
 n43127 , n363284 , n43129 , n43130 , n43131 , n363288 , n363289 , n43134 , n363291 , n363292 , 
 n363293 , n363294 , n363295 , n43140 , n363297 , n43142 , n43143 , n363300 , n363301 , n363302 , 
 n363303 , n363304 , n363305 , n43150 , n363307 , n363308 , n363309 , n363310 , n363311 , n43156 , 
 n363313 , n363314 , n363315 , n363316 , n363317 , n363318 , n43163 , n43164 , n363321 , n363322 , 
 n43167 , n43168 , n363325 , n363326 , n363327 , n363328 , n363329 , n363330 , n363331 , n363332 , 
 n363333 , n363334 , n43179 , n363336 , n43181 , n363338 , n43183 , n363340 , n363341 , n363342 , 
 n43187 , n363344 , n363345 , n363346 , n363347 , n363348 , n363349 , n43194 , n363351 , n363352 , 
 n43197 , n363354 , n363355 , n363356 , n363357 , n363358 , n363359 , n363360 , n363361 , n363362 , 
 n363363 , n43208 , n363365 , n363366 , n363367 , n363368 , n363369 , n363370 , n43215 , n363372 , 
 n363373 , n363374 , n363375 , n43220 , n363377 , n363378 , n43223 , n363380 , n363381 , n43226 , 
 n363383 , n43228 , n363385 , n363386 , n43231 , n363388 , n43233 , n363390 , n363391 , n363392 , 
 n363393 , n43238 , n363395 , n363396 , n363397 , n363398 , n363399 , n363400 , n363401 , n363402 , 
 n363403 , n363404 , n363405 , n363406 , n363407 , n43252 , n43253 , n363410 , n363411 , n43256 , 
 n363413 , n43258 , n363415 , n363416 , n43261 , n363418 , n363419 , n363420 , n363421 , n363422 , 
 n363423 , n43268 , n363425 , n363426 , n43271 , n363428 , n363429 , n43274 , n363431 , n363432 , 
 n43277 , n363434 , n363435 , n43280 , n363437 , n363438 , n363439 , n363440 , n363441 , n363442 , 
 n363443 , n363444 , n363445 , n363446 , n43282 , n43283 , n363449 , n363450 , n363451 , n363452 , 
 n363453 , n363454 , n363455 , n43291 , n363457 , n363458 , n363459 , n43295 , n363461 , n363462 , 
 n363463 , n363464 , n43300 , n363466 , n363467 , n363468 , n43304 , n43305 , n363471 , n43307 , 
 n363473 , n363474 , n363475 , n363476 , n363477 , n43313 , n363479 , n363480 , n363481 , n43317 , 
 n363483 , n363484 , n363485 , n363486 , n363487 , n43323 , n363489 , n363490 , n43326 , n363492 , 
 n43328 , n363494 , n363495 , n363496 , n363497 , n363498 , n363499 , n363500 , n363501 , n363502 , 
 n363503 , n43339 , n363505 , n43341 , n43342 , n43343 , n43344 , n363510 , n363511 , n363512 , 
 n363513 , n43349 , n43350 , n363516 , n363517 , n43353 , n363519 , n363520 , n43356 , n363522 , 
 n363523 , n363524 , n363525 , n43361 , n363527 , n363528 , n363529 , n363530 , n363531 , n43367 , 
 n363533 , n363534 , n363535 , n363536 , n363537 , n363538 , n363539 , n363540 , n363541 , n43377 , 
 n363543 , n363544 , n43380 , n363546 , n363547 , n363548 , n363549 , n43385 , n43386 , n363552 , 
 n43388 , n43389 , n363555 , n43391 , n363557 , n363558 , n43394 , n363560 , n363561 , n43397 , 
 n363563 , n363564 , n363565 , n363566 , n363567 , n363568 , n363569 , n363570 , n43406 , n363572 , 
 n363573 , n43409 , n363575 , n363576 , n363577 , n363578 , n363579 , n363580 , n363581 , n363582 , 
 n363583 , n363584 , n363585 , n363586 , n363587 , n363588 , n43424 , n363590 , n363591 , n363592 , 
 n43428 , n363594 , n43430 , n363596 , n363597 , n43433 , n363599 , n363600 , n363601 , n363602 , 
 n363603 , n43439 , n363605 , n43441 , n363607 , n363608 , n363609 , n43445 , n363611 , n43447 , 
 n43448 , n43449 , n43450 , n43451 , n43452 , n363618 , n363619 , n43455 , n363621 , n363622 , 
 n363623 , n363624 , n363625 , n43461 , n363627 , n43463 , n363629 , n363630 , n363631 , n363632 , 
 n363633 , n43469 , n363635 , n363636 , n363637 , n43473 , n363639 , n363640 , n363641 , n363642 , 
 n43478 , n43479 , n363645 , n363646 , n363647 , n43483 , n363649 , n363650 , n363651 , n363652 , 
 n363653 , n363654 , n363655 , n43491 , n363657 , n43493 , n363659 , n43495 , n363661 , n43497 , 
 n363663 , n43499 , n363665 , n363666 , n43502 , n363668 , n363669 , n363670 , n363671 , n363672 , 
 n363673 , n43509 , n363675 , n363676 , n43512 , n363678 , n363679 , n363680 , n363681 , n363682 , 
 n43518 , n363684 , n363685 , n363686 , n363687 , n363688 , n363689 , n43525 , n363691 , n363692 , 
 n363693 , n43529 , n363695 , n363696 , n363697 , n363698 , n363699 , n43535 , n363701 , n363702 , 
 n43538 , n363704 , n363705 , n363706 , n43542 , n43543 , n363709 , n43545 , n363711 , n363712 , 
 n43548 , n43549 , n363715 , n363716 , n43552 , n43553 , n363719 , n43555 , n363721 , n363722 , 
 n43558 , n363724 , n363725 , n363726 , n363727 , n363728 , n43564 , n43565 , n363731 , n43567 , 
 n363733 , n363734 , n43570 , n43571 , n43572 , n43573 , n43574 , n363740 , n363741 , n363742 , 
 n363743 , n363744 , n363745 , n363746 , n363747 , n43583 , n363749 , n363750 , n43586 , n363752 , 
 n363753 , n363754 , n363755 , n363756 , n363757 , n363758 , n363759 , n363760 , n363761 , n43597 , 
 n43598 , n363764 , n363765 , n363766 , n363767 , n363768 , n363769 , n363770 , n363771 , n363772 , 
 n363773 , n363774 , n43610 , n363776 , n363777 , n363778 , n363779 , n363780 , n363781 , n43617 , 
 n363783 , n363784 , n363785 , n363786 , n363787 , n363788 , n363789 , n363790 , n363791 , n363792 , 
 n43628 , n363794 , n363795 , n43631 , n363797 , n363798 , n363799 , n363800 , n363801 , n43637 , 
 n363803 , n363804 , n363805 , n363806 , n43642 , n363808 , n363809 , n43645 , n43646 , n363812 , 
 n43648 , n363814 , n363815 , n43651 , n363817 , n363818 , n363819 , n363820 , n363821 , n43657 , 
 n43658 , n363824 , n43660 , n363826 , n363827 , n363828 , n363829 , n363830 , n363831 , n43667 , 
 n363833 , n363834 , n363835 , n43671 , n363837 , n43673 , n363839 , n43675 , n363841 , n363842 , 
 n363843 , n363844 , n363845 , n363846 , n363847 , n363848 , n363849 , n363850 , n363851 , n363852 , 
 n363853 , n363854 , n363855 , n363856 , n363857 , n363858 , n363859 , n363860 , n363861 , n363862 , 
 n363863 , n363864 , n363865 , n363866 , n363867 , n363868 , n363869 , n363870 , n363871 , n363872 , 
 n363873 , n363874 , n43710 , n43711 , n363877 , n43713 , n363879 , n363880 , n363881 , n363882 , 
 n363883 , n363884 , n363885 , n363886 , n363887 , n43723 , n363889 , n363890 , n43726 , n363892 , 
 n363893 , n363894 , n363895 , n43731 , n43732 , n363898 , n43734 , n43735 , n363901 , n363902 , 
 n363903 , n363904 , n363905 , n363906 , n363907 , n363908 , n43744 , n363910 , n363911 , n363912 , 
 n43748 , n363914 , n363915 , n363916 , n363917 , n363918 , n43754 , n363920 , n363921 , n43757 , 
 n363923 , n363924 , n363925 , n43761 , n363927 , n43763 , n363929 , n43765 , n363931 , n363932 , 
 n43768 , n363934 , n363935 , n43771 , n363937 , n363938 , n43774 , n363940 , n363941 , n363942 , 
 n363943 , n43779 , n363945 , n363946 , n363947 , n363948 , n363949 , n43785 , n43786 , n363952 , 
 n363953 , n363954 , n363955 , n363956 , n363957 , n363958 , n363959 , n43795 , n363961 , n43797 , 
 n43798 , n363964 , n43800 , n363966 , n363967 , n363968 , n363969 , n363970 , n363971 , n363972 , 
 n363973 , n363974 , n43810 , n363976 , n43812 , n363978 , n363979 , n363980 , n363981 , n363982 , 
 n363983 , n363984 , n43820 , n43821 , n363987 , n43823 , n363989 , n363990 , n363991 , n363992 , 
 n363993 , n363994 , n363995 , n363996 , n43832 , n363998 , n363999 , n364000 , n364001 , n364002 , 
 n364003 , n43839 , n364005 , n364006 , n364007 , n364008 , n364009 , n43845 , n364011 , n364012 , 
 n43848 , n364014 , n364015 , n364016 , n364017 , n364018 , n364019 , n364020 , n364021 , n364022 , 
 n364023 , n364024 , n364025 , n364026 , n364027 , n364028 , n364029 , n364030 , n364031 , n43867 , 
 n364033 , n43869 , n43870 , n43871 , n43872 , n364038 , n43874 , n364040 , n364041 , n364042 , 
 n364043 , n364044 , n364045 , n364046 , n43882 , n364048 , n43884 , n43885 , n364051 , n364052 , 
 n364053 , n364054 , n364055 , n43891 , n364057 , n364058 , n364059 , n364060 , n43896 , n364062 , 
 n364063 , n364064 , n43900 , n364066 , n43902 , n43903 , n364069 , n43905 , n43906 , n364072 , 
 n43908 , n364074 , n43910 , n364076 , n364077 , n364078 , n364079 , n43915 , n364081 , n364082 , 
 n43918 , n364084 , n364085 , n364086 , n364087 , n43923 , n364089 , n364090 , n364091 , n364092 , 
 n364093 , n43929 , n364095 , n364096 , n43932 , n364098 , n364099 , n364100 , n364101 , n364102 , 
 n364103 , n364104 , n43940 , n364106 , n43942 , n43943 , n364109 , n43945 , n364111 , n364112 , 
 n364113 , n43949 , n364115 , n364116 , n43952 , n43953 , n364119 , n364120 , n364121 , n364122 , 
 n43958 , n364124 , n364125 , n43961 , n364127 , n43963 , n364129 , n43965 , n43966 , n364132 , 
 n43968 , n364134 , n364135 , n364136 , n364137 , n364138 , n43974 , n364140 , n43976 , n43977 , 
 n364143 , n43979 , n364145 , n43981 , n364147 , n364148 , n43984 , n364150 , n364151 , n43987 , 
 n364153 , n364154 , n364155 , n364156 , n364157 , n364158 , n364159 , n43995 , n364161 , n364162 , 
 n364163 , n364164 , n44000 , n364166 , n364167 , n44003 , n44004 , n364170 , n364171 , n364172 , 
 n364173 , n364174 , n44010 , n44011 , n364177 , n44013 , n364179 , n364180 , n364181 , n44017 , 
 n364183 , n364184 , n44020 , n364186 , n44022 , n364188 , n44024 , n364190 , n364191 , n364192 , 
 n44028 , n364194 , n44030 , n364196 , n364197 , n364198 , n364199 , n364200 , n364201 , n364202 , 
 n364203 , n364204 , n364205 , n44041 , n364207 , n364208 , n44044 , n364210 , n364211 , n44047 , 
 n364213 , n44049 , n364215 , n364216 , n364217 , n364218 , n364219 , n364220 , n44056 , n364222 , 
 n364223 , n364224 , n364225 , n364226 , n364227 , n44063 , n44064 , n364230 , n44066 , n364232 , 
 n44068 , n364234 , n44070 , n364236 , n364237 , n364238 , n364239 , n364240 , n364241 , n364242 , 
 n364243 , n364244 , n44080 , n364246 , n364247 , n364248 , n364249 , n364250 , n364251 , n364252 , 
 n44088 , n364254 , n364255 , n44091 , n364257 , n364258 , n364259 , n364260 , n364261 , n364262 , 
 n364263 , n364264 , n364265 , n364266 , n44102 , n44103 , n44104 , n364270 , n44106 , n44107 , 
 n364273 , n44109 , n364275 , n364276 , n44112 , n364278 , n364279 , n364280 , n44116 , n364282 , 
 n364283 , n44119 , n364285 , n364286 , n44122 , n44123 , n364289 , n44125 , n364291 , n364292 , 
 n364293 , n44129 , n364295 , n364296 , n364297 , n364298 , n44134 , n364300 , n44136 , n44137 , 
 n44138 , n364304 , n44140 , n364306 , n364307 , n364308 , n364309 , n364310 , n364311 , n364312 , 
 n364313 , n364314 , n364315 , n44151 , n364317 , n364318 , n44154 , n364320 , n364321 , n364322 , 
 n364323 , n364324 , n44160 , n364326 , n364327 , n364328 , n364329 , n364330 , n364331 , n364332 , 
 n364333 , n44169 , n44170 , n44171 , n364337 , n364338 , n44174 , n44175 , n44176 , n364342 , 
 n44178 , n364344 , n364345 , n44181 , n44182 , n44183 , n44184 , n44185 , n364351 , n364352 , 
 n364353 , n364354 , n364355 , n44191 , n364357 , n44193 , n364359 , n364360 , n44196 , n364362 , 
 n364363 , n364364 , n364365 , n364366 , n44202 , n364368 , n44204 , n364370 , n364371 , n44207 , 
 n364373 , n364374 , n364375 , n364376 , n44212 , n44213 , n364379 , n364380 , n364381 , n364382 , 
 n364383 , n364384 , n364385 , n364386 , n364387 , n44223 , n364389 , n364390 , n364391 , n364392 , 
 n364393 , n44229 , n364395 , n364396 , n364397 , n364398 , n364399 , n364400 , n364401 , n364402 , 
 n364403 , n364404 , n364405 , n364406 , n364407 , n44243 , n364409 , n364410 , n364411 , n364412 , 
 n364413 , n364414 , n364415 , n364416 , n364417 , n364418 , n364419 , n364420 , n364421 , n44257 , 
 n364423 , n364424 , n44260 , n364426 , n364427 , n44263 , n364429 , n364430 , n44266 , n364432 , 
 n364433 , n44269 , n364435 , n44271 , n364437 , n44273 , n44274 , n364440 , n364441 , n44277 , 
 n364443 , n364444 , n364445 , n364446 , n364447 , n44283 , n364449 , n364450 , n364451 , n364452 , 
 n364453 , n364454 , n364455 , n44291 , n364457 , n44293 , n364459 , n364460 , n364461 , n364462 , 
 n364463 , n44299 , n364465 , n364466 , n44302 , n364468 , n364469 , n364470 , n44306 , n364472 , 
 n364473 , n44309 , n364475 , n44311 , n364477 , n364478 , n364479 , n44315 , n364481 , n364482 , 
 n44318 , n364484 , n44320 , n364486 , n364487 , n364488 , n364489 , n364490 , n364491 , n44327 , 
 n364493 , n44329 , n364495 , n364496 , n364497 , n44333 , n364499 , n364500 , n364501 , n364502 , 
 n364503 , n44339 , n44340 , n44341 , n364507 , n364508 , n44344 , n364510 , n364511 , n364512 , 
 n364513 , n364514 , n364515 , n44351 , n364517 , n44353 , n44354 , n364520 , n364521 , n44357 , 
 n364523 , n364524 , n44360 , n364526 , n44362 , n44363 , n364529 , n44365 , n364531 , n364532 , 
 n44368 , n364534 , n44370 , n364536 , n364537 , n44373 , n364539 , n364540 , n364541 , n364542 , 
 n44378 , n364544 , n44380 , n364546 , n364547 , n364548 , n44384 , n364550 , n364551 , n44387 , 
 n364553 , n364554 , n44390 , n44391 , n364557 , n44393 , n364559 , n364560 , n44396 , n364562 , 
 n364563 , n44399 , n44400 , n364566 , n44402 , n364568 , n364569 , n364570 , n364571 , n364572 , 
 n364573 , n364574 , n364575 , n364576 , n44412 , n364578 , n44414 , n364580 , n364581 , n44417 , 
 n364583 , n364584 , n44420 , n364586 , n364587 , n44423 , n364589 , n364590 , n364591 , n364592 , 
 n364593 , n364594 , n364595 , n44431 , n364597 , n364598 , n364599 , n364600 , n364601 , n364602 , 
 n364603 , n364604 , n364605 , n44441 , n364607 , n364608 , n44444 , n364610 , n44446 , n364612 , 
 n44448 , n364614 , n44450 , n364616 , n364617 , n364618 , n364619 , n364620 , n364621 , n364622 , 
 n44458 , n364624 , n364625 , n364626 , n44462 , n364628 , n44464 , n44465 , n364631 , n364632 , 
 n44468 , n364634 , n364635 , n44471 , n364637 , n364638 , n44474 , n364640 , n44476 , n364642 , 
 n364643 , n44479 , n364645 , n44481 , n44482 , n44483 , n364649 , n364650 , n44486 , n364652 , 
 n44488 , n364654 , n364655 , n364656 , n364657 , n364658 , n364659 , n44495 , n364661 , n44497 , 
 n364663 , n364664 , n44500 , n364666 , n364667 , n364668 , n44504 , n44505 , n364671 , n364672 , 
 n44508 , n364674 , n364675 , n44511 , n44512 , n364678 , n364679 , n44515 , n364681 , n364682 , 
 n44518 , n364684 , n364685 , n44521 , n364687 , n364688 , n364689 , n364690 , n44526 , n44527 , 
 n364693 , n44529 , n364695 , n364696 , n44532 , n364698 , n364699 , n44535 , n364701 , n364702 , 
 n364703 , n364704 , n44540 , n44541 , n364707 , n364708 , n364709 , n364710 , n364711 , n364712 , 
 n364713 , n364714 , n364715 , n364716 , n364717 , n44553 , n364719 , n364720 , n364721 , n364722 , 
 n44558 , n44559 , n44560 , n364726 , n44562 , n364728 , n44564 , n364730 , n364731 , n44567 , 
 n44568 , n44569 , n44570 , n364736 , n44572 , n44573 , n364739 , n44575 , n44576 , n364742 , 
 n44578 , n364744 , n364745 , n44581 , n364747 , n364748 , n364749 , n364750 , n364751 , n364752 , 
 n364753 , n364754 , n44590 , n44591 , n364757 , n364758 , n364759 , n364760 , n364761 , n364762 , 
 n364763 , n364764 , n364765 , n364766 , n364767 , n364768 , n44604 , n364770 , n364771 , n364772 , 
 n364773 , n364774 , n364775 , n364776 , n364777 , n364778 , n364779 , n44615 , n364781 , n364782 , 
 n364783 , n364784 , n364785 , n364786 , n364787 , n364788 , n364789 , n364790 , n364791 , n44627 , 
 n364793 , n44629 , n364795 , n364796 , n364797 , n364798 , n44634 , n364800 , n364801 , n44637 , 
 n44638 , n364804 , n364805 , n44641 , n364807 , n364808 , n364809 , n364810 , n364811 , n364812 , 
 n364813 , n364814 , n364815 , n364816 , n364817 , n364818 , n364819 , n44655 , n364821 , n364822 , 
 n44658 , n364824 , n364825 , n44661 , n364827 , n364828 , n44664 , n364830 , n364831 , n364832 , 
 n364833 , n44669 , n364835 , n364836 , n364837 , n44673 , n364839 , n364840 , n364841 , n364842 , 
 n364843 , n364844 , n364845 , n44681 , n364847 , n364848 , n364849 , n364850 , n44686 , n364852 , 
 n364853 , n364854 , n364855 , n364856 , n44692 , n364858 , n364859 , n364860 , n364861 , n44697 , 
 n364863 , n364864 , n364865 , n364866 , n364867 , n364868 , n364869 , n364870 , n44706 , n44707 , 
 n364873 , n364874 , n44710 , n364876 , n364877 , n364878 , n364879 , n44715 , n364881 , n44717 , 
 n364883 , n364884 , n364885 , n364886 , n364887 , n364888 , n364889 , n364890 , n364891 , n44727 , 
 n44728 , n364894 , n364895 , n44731 , n364897 , n364898 , n364899 , n364900 , n364901 , n44737 , 
 n364903 , n44739 , n364905 , n364906 , n364907 , n44743 , n364909 , n364910 , n44746 , n364912 , 
 n364913 , n44749 , n364915 , n364916 , n364917 , n364918 , n364919 , n364920 , n364921 , n364922 , 
 n364923 , n364924 , n364925 , n364926 , n364927 , n44763 , n364929 , n364930 , n44766 , n44767 , 
 n364933 , n364934 , n44770 , n364936 , n364937 , n364938 , n364939 , n44775 , n44776 , n364942 , 
 n364943 , n44779 , n364945 , n364946 , n364947 , n44783 , n364949 , n364950 , n44786 , n364952 , 
 n364953 , n364954 , n44790 , n364956 , n364957 , n364958 , n364959 , n364960 , n44796 , n364962 , 
 n44798 , n364964 , n364965 , n364966 , n364967 , n364968 , n44804 , n44805 , n364971 , n364972 , 
 n44808 , n364974 , n364975 , n364976 , n364977 , n364978 , n364979 , n44815 , n364981 , n364982 , 
 n44818 , n44819 , n364985 , n44821 , n364987 , n364988 , n44824 , n44825 , n44826 , n364992 , 
 n44828 , n364994 , n364995 , n364996 , n364997 , n364998 , n44834 , n365000 , n365001 , n44837 , 
 n365003 , n365004 , n365005 , n44841 , n365007 , n44843 , n44844 , n365010 , n365011 , n365012 , 
 n365013 , n365014 , n44850 , n44851 , n365017 , n44853 , n365019 , n365020 , n365021 , n365022 , 
 n365023 , n365024 , n365025 , n44861 , n44862 , n365028 , n44864 , n365030 , n44866 , n365032 , 
 n365033 , n365034 , n365035 , n365036 , n365037 , n365038 , n365039 , n365040 , n365041 , n365042 , 
 n365043 , n365044 , n44880 , n44881 , n365047 , n365048 , n44884 , n365050 , n365051 , n365052 , 
 n365053 , n44889 , n365055 , n365056 , n44892 , n365058 , n365059 , n365060 , n365061 , n365062 , 
 n44898 , n44899 , n365065 , n365066 , n44902 , n365068 , n44904 , n365070 , n44906 , n365072 , 
 n44908 , n365074 , n365075 , n365076 , n44912 , n44913 , n44914 , n44915 , n365081 , n365082 , 
 n365083 , n365084 , n365085 , n365086 , n365087 , n44923 , n365089 , n44925 , n44926 , n365092 , 
 n365093 , n365094 , n44930 , n365096 , n365097 , n365098 , n365099 , n365100 , n365101 , n44937 , 
 n365103 , n365104 , n365105 , n365106 , n365107 , n365108 , n44944 , n44945 , n44946 , n365112 , 
 n365113 , n365114 , n365115 , n365116 , n365117 , n365118 , n44954 , n365120 , n44956 , n44957 , 
 n365123 , n365124 , n44960 , n365126 , n365127 , n44963 , n365129 , n365130 , n44966 , n365132 , 
 n365133 , n365134 , n365135 , n365136 , n365137 , n365138 , n365139 , n44970 , n365141 , n365142 , 
 n365143 , n365144 , n365145 , n365146 , n365147 , n365148 , n365149 , n365150 , n365151 , n365152 , 
 n365153 , n365154 , n365155 , n44986 , n365157 , n44988 , n365159 , n365160 , n44991 , n365162 , 
 n365163 , n365164 , n365165 , n365166 , n365167 , n365168 , n365169 , n365170 , n365171 , n365172 , 
 n365173 , n365174 , n45005 , n365176 , n365177 , n45008 , n365179 , n45010 , n365181 , n45012 , 
 n365183 , n45014 , n45015 , n365186 , n365187 , n45018 , n365189 , n365190 , n45021 , n365192 , 
 n365193 , n45024 , n365195 , n365196 , n365197 , n45028 , n45029 , n365200 , n45031 , n365202 , 
 n365203 , n45034 , n365205 , n365206 , n365207 , n365208 , n45039 , n365210 , n365211 , n45042 , 
 n365213 , n365214 , n45045 , n45046 , n365217 , n365218 , n45049 , n45050 , n45051 , n45052 , 
 n45053 , n365224 , n45055 , n365226 , n365227 , n45058 , n365229 , n45060 , n45061 , n45062 , 
 n45063 , n365234 , n45065 , n365236 , n365237 , n365238 , n365239 , n365240 , n45071 , n365242 , 
 n45073 , n45074 , n45075 , n45076 , n45077 , n365248 , n45079 , n365250 , n365251 , n365252 , 
 n45083 , n365254 , n45085 , n365256 , n365257 , n365258 , n365259 , n365260 , n45091 , n45092 , 
 n365263 , n365264 , n45095 , n365266 , n365267 , n365268 , n365269 , n365270 , n365271 , n365272 , 
 n45103 , n365274 , n365275 , n365276 , n365277 , n365278 , n365279 , n365280 , n365281 , n365282 , 
 n45113 , n365284 , n365285 , n45116 , n365287 , n45118 , n365289 , n365290 , n365291 , n45122 , 
 n365293 , n365294 , n45125 , n365296 , n365297 , n365298 , n365299 , n365300 , n365301 , n365302 , 
 n365303 , n365304 , n365305 , n365306 , n365307 , n365308 , n365309 , n365310 , n365311 , n365312 , 
 n45143 , n365314 , n365315 , n45146 , n365317 , n365318 , n365319 , n365320 , n365321 , n45152 , 
 n365323 , n45154 , n365325 , n365326 , n45157 , n365328 , n365329 , n365330 , n365331 , n365332 , 
 n365333 , n365334 , n365335 , n45166 , n365337 , n365338 , n45169 , n45170 , n365341 , n45172 , 
 n365343 , n365344 , n365345 , n45176 , n45177 , n365348 , n45179 , n365350 , n45181 , n365352 , 
 n365353 , n365354 , n365355 , n45186 , n365357 , n365358 , n45189 , n365360 , n365361 , n365362 , 
 n365363 , n45194 , n45195 , n45196 , n365367 , n365368 , n45199 , n45200 , n45201 , n365372 , 
 n365373 , n45204 , n365375 , n365376 , n365377 , n45208 , n45209 , n45210 , n365381 , n365382 , 
 n45213 , n365384 , n365385 , n365386 , n365387 , n365388 , n45219 , n365390 , n365391 , n365392 , 
 n365393 , n365394 , n365395 , n365396 , n365397 , n365398 , n365399 , n45230 , n45231 , n365402 , 
 n45233 , n45234 , n365405 , n365406 , n45237 , n365408 , n45239 , n45240 , n45241 , n45242 , 
 n45243 , n45244 , n365415 , n365416 , n365417 , n365418 , n365419 , n365420 , n365421 , n365422 , 
 n365423 , n365424 , n45250 , n365426 , n365427 , n365428 , n365429 , n365430 , n365431 , n365432 , 
 n365433 , n365434 , n365435 , n365436 , n365437 , n365438 , n365439 , n365440 , n45266 , n45267 , 
 n45268 , n45269 , n45270 , n365446 , n365447 , n45273 , n365449 , n45275 , n365451 , n365452 , 
 n365453 , n365454 , n365455 , n365456 , n365457 , n365458 , n45284 , n45285 , n365461 , n45287 , 
 n365463 , n365464 , n45290 , n365466 , n365467 , n365468 , n365469 , n365470 , n365471 , n45297 , 
 n365473 , n365474 , n45300 , n365476 , n365477 , n45303 , n365479 , n365480 , n365481 , n365482 , 
 n365483 , n365484 , n365485 , n365486 , n45312 , n365488 , n365489 , n365490 , n365491 , n45317 , 
 n365493 , n45319 , n365495 , n365496 , n45322 , n365498 , n365499 , n45325 , n365501 , n365502 , 
 n365503 , n365504 , n365505 , n45331 , n365507 , n45333 , n365509 , n45335 , n45336 , n365512 , 
 n45338 , n45339 , n365515 , n45341 , n365517 , n365518 , n365519 , n45345 , n365521 , n365522 , 
 n365523 , n365524 , n365525 , n365526 , n45352 , n365528 , n365529 , n365530 , n45356 , n365532 , 
 n365533 , n365534 , n365535 , n365536 , n45362 , n365538 , n45364 , n365540 , n365541 , n365542 , 
 n365543 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n365552 , 
 n365553 , n45379 , n45380 , n365556 , n365557 , n365558 , n45384 , n365560 , n365561 , n365562 , 
 n365563 , n365564 , n365565 , n45391 , n365567 , n45393 , n365569 , n365570 , n365571 , n45397 , 
 n365573 , n365574 , n45400 , n45401 , n365577 , n45403 , n45404 , n365580 , n45406 , n365582 , 
 n365583 , n365584 , n45410 , n365586 , n45412 , n365588 , n45414 , n365590 , n365591 , n45417 , 
 n365593 , n365594 , n365595 , n365596 , n365597 , n365598 , n365599 , n365600 , n365601 , n365602 , 
 n365603 , n45429 , n365605 , n365606 , n365607 , n365608 , n365609 , n365610 , n365611 , n45437 , 
 n45438 , n365614 , n45440 , n45441 , n365617 , n365618 , n365619 , n365620 , n365621 , n365622 , 
 n365623 , n365624 , n45450 , n365626 , n365627 , n45453 , n45454 , n45455 , n365631 , n45457 , 
 n45458 , n45459 , n365635 , n365636 , n365637 , n365638 , n365639 , n365640 , n365641 , n365642 , 
 n365643 , n365644 , n365645 , n365646 , n365647 , n45473 , n365649 , n365650 , n365651 , n45477 , 
 n45478 , n365654 , n365655 , n365656 , n365657 , n45483 , n45484 , n45485 , n365661 , n45487 , 
 n365663 , n45489 , n365665 , n45491 , n45492 , n45493 , n45494 , n365670 , n365671 , n45497 , 
 n365673 , n365674 , n365675 , n365676 , n365677 , n45503 , n45504 , n365680 , n365681 , n365682 , 
 n45508 , n365684 , n45510 , n365686 , n45512 , n365688 , n365689 , n45515 , n365691 , n365692 , 
 n365693 , n45519 , n45520 , n45521 , n45522 , n45523 , n365699 , n365700 , n45526 , n45527 , 
 n45528 , n365704 , n365705 , n365706 , n365707 , n365708 , n45534 , n365710 , n365711 , n365712 , 
 n365713 , n365714 , n365715 , n365716 , n365717 , n45543 , n45544 , n365720 , n45546 , n365722 , 
 n365723 , n45549 , n365725 , n365726 , n45552 , n45553 , n365729 , n45555 , n45556 , n365732 , 
 n45558 , n365734 , n365735 , n365736 , n365737 , n45563 , n365739 , n45565 , n45566 , n365742 , 
 n365743 , n45569 , n45570 , n365746 , n365747 , n45573 , n365749 , n365750 , n365751 , n365752 , 
 n365753 , n45579 , n365755 , n365756 , n365757 , n365758 , n365759 , n365760 , n45586 , n45587 , 
 n45588 , n45589 , n365765 , n45591 , n45592 , n365768 , n45594 , n45595 , n365771 , n45597 , 
 n365773 , n365774 , n365775 , n365776 , n365777 , n365778 , n365779 , n365780 , n365781 , n365782 , 
 n45608 , n45609 , n365785 , n45611 , n365787 , n365788 , n45614 , n45615 , n365791 , n365792 , 
 n365793 , n365794 , n45620 , n365796 , n365797 , n45623 , n365799 , n365800 , n365801 , n365802 , 
 n365803 , n365804 , n365805 , n45631 , n365807 , n45633 , n365809 , n365810 , n365811 , n45637 , 
 n365813 , n365814 , n45640 , n365816 , n365817 , n365818 , n45644 , n45645 , n365821 , n45647 , 
 n365823 , n45649 , n365825 , n365826 , n45652 , n365828 , n365829 , n365830 , n45656 , n45657 , 
 n365833 , n365834 , n365835 , n365836 , n365837 , n365838 , n365839 , n365840 , n365841 , n365842 , 
 n365843 , n365844 , n45670 , n365846 , n365847 , n365848 , n45674 , n365850 , n365851 , n365852 , 
 n365853 , n365854 , n365855 , n365856 , n365857 , n365858 , n365859 , n365860 , n365861 , n45687 , 
 n365863 , n45689 , n45690 , n45691 , n365867 , n45693 , n45694 , n365870 , n45696 , n365872 , 
 n45698 , n365874 , n45700 , n365876 , n45702 , n365878 , n45704 , n45705 , n45706 , n365882 , 
 n45708 , n45709 , n365885 , n45711 , n365887 , n45713 , n365889 , n45715 , n365891 , n45717 , 
 n45718 , n365894 , n365895 , n365896 , n365897 , n365898 , n365899 , n365900 , n365901 , n365902 , 
 n365903 , n45729 , n365905 , n365906 , n45732 , n45733 , n45734 , n365910 , n365911 , n365912 , 
 n365913 , n45739 , n365915 , n365916 , n45742 , n365918 , n45744 , n45745 , n45746 , n45747 , 
 n365923 , n45749 , n365925 , n45751 , n365927 , n365928 , n365929 , n365930 , n365931 , n365932 , 
 n365933 , n365934 , n365935 , n45761 , n365937 , n365938 , n45764 , n365940 , n365941 , n45767 , 
 n365943 , n365944 , n365945 , n365946 , n365947 , n365948 , n365949 , n365950 , n365951 , n365952 , 
 n45778 , n365954 , n365955 , n45781 , n365957 , n365958 , n365959 , n365960 , n365961 , n45787 , 
 n365963 , n45789 , n45790 , n365966 , n365967 , n365968 , n45794 , n45795 , n365971 , n45797 , 
 n45798 , n365974 , n45800 , n45801 , n45802 , n365978 , n45804 , n365980 , n365981 , n365982 , 
 n365983 , n45809 , n365985 , n365986 , n365987 , n365988 , n365989 , n365990 , n365991 , n365992 , 
 n365993 , n45819 , n365995 , n365996 , n365997 , n365998 , n365999 , n366000 , n366001 , n366002 , 
 n366003 , n366004 , n366005 , n45831 , n366007 , n366008 , n45834 , n366010 , n45836 , n366012 , 
 n366013 , n366014 , n366015 , n366016 , n366017 , n366018 , n366019 , n45845 , n366021 , n366022 , 
 n366023 , n366024 , n366025 , n366026 , n45852 , n366028 , n366029 , n45855 , n366031 , n366032 , 
 n45858 , n45859 , n366035 , n366036 , n366037 , n366038 , n45864 , n366040 , n366041 , n366042 , 
 n366043 , n366044 , n366045 , n366046 , n366047 , n45873 , n45874 , n366050 , n366051 , n45877 , 
 n366053 , n366054 , n45880 , n366056 , n366057 , n366058 , n366059 , n366060 , n45886 , n366062 , 
 n366063 , n366064 , n366065 , n366066 , n366067 , n366068 , n366069 , n366070 , n366071 , n366072 , 
 n366073 , n366074 , n45900 , n45901 , n366077 , n366078 , n366079 , n366080 , n366081 , n45907 , 
 n45908 , n366084 , n45910 , n366086 , n366087 , n366088 , n45914 , n45915 , n45916 , n366092 , 
 n366093 , n366094 , n366095 , n366096 , n366097 , n366098 , n366099 , n366100 , n45926 , n366102 , 
 n366103 , n45929 , n366105 , n366106 , n45932 , n366108 , n45934 , n45935 , n366111 , n45937 , 
 n366113 , n366114 , n366115 , n366116 , n366117 , n366118 , n45944 , n366120 , n366121 , n45947 , 
 n366123 , n45949 , n366125 , n366126 , n366127 , n366128 , n366129 , n366130 , n366131 , n366132 , 
 n366133 , n366134 , n366135 , n366136 , n366137 , n366138 , n366139 , n366140 , n45966 , n366142 , 
 n366143 , n366144 , n366145 , n45971 , n366147 , n366148 , n366149 , n366150 , n366151 , n45977 , 
 n45978 , n366154 , n366155 , n366156 , n366157 , n45983 , n366159 , n45985 , n366161 , n45987 , 
 n45988 , n366164 , n45990 , n366166 , n366167 , n45993 , n366169 , n366170 , n45996 , n45997 , 
 n366173 , n366174 , n366175 , n46001 , n366177 , n366178 , n366179 , n366180 , n366181 , n46007 , 
 n46008 , n366184 , n366185 , n46011 , n366187 , n46013 , n46014 , n366190 , n366191 , n366192 , 
 n366193 , n366194 , n366195 , n366196 , n366197 , n46023 , n366199 , n46025 , n366201 , n366202 , 
 n366203 , n366204 , n46030 , n46031 , n366207 , n46033 , n366209 , n46035 , n46036 , n366212 , 
 n46038 , n46039 , n46040 , n46041 , n366217 , n366218 , n46044 , n366220 , n366221 , n366222 , 
 n46048 , n366224 , n46050 , n366226 , n366227 , n46053 , n366229 , n366230 , n366231 , n366232 , 
 n46058 , n366234 , n366235 , n46061 , n366237 , n46063 , n46064 , n366240 , n366241 , n46067 , 
 n366243 , n46069 , n366245 , n366246 , n46072 , n366248 , n366249 , n46075 , n366251 , n366252 , 
 n366253 , n366254 , n366255 , n366256 , n366257 , n46083 , n46084 , n366260 , n366261 , n46087 , 
 n366263 , n46089 , n46090 , n366266 , n366267 , n366268 , n366269 , n366270 , n366271 , n366272 , 
 n46098 , n46099 , n366275 , n46101 , n366277 , n366278 , n366279 , n46105 , n366281 , n366282 , 
 n46108 , n46109 , n366285 , n46111 , n366287 , n366288 , n46113 , n366290 , n366291 , n366292 , 
 n366293 , n366294 , n366295 , n366296 , n46121 , n366298 , n366299 , n46124 , n46125 , n46126 , 
 n366303 , n46128 , n366305 , n366306 , n366307 , n366308 , n366309 , n366310 , n366311 , n366312 , 
 n366313 , n366314 , n366315 , n46135 , n366317 , n366318 , n46138 , n366320 , n366321 , n366322 , 
 n366323 , n46143 , n46144 , n366326 , n366327 , n46147 , n366329 , n366330 , n46150 , n366332 , 
 n366333 , n46153 , n366335 , n366336 , n46156 , n46157 , n366339 , n46159 , n366341 , n366342 , 
 n46162 , n366344 , n366345 , n366346 , n366347 , n46167 , n46168 , n366350 , n366351 , n46171 , 
 n366353 , n366354 , n46174 , n366356 , n366357 , n46177 , n366359 , n366360 , n366361 , n366362 , 
 n366363 , n366364 , n366365 , n46185 , n366367 , n46187 , n46188 , n46189 , n46190 , n366372 , 
 n46192 , n46193 , n366375 , n366376 , n366377 , n366378 , n46198 , n366380 , n366381 , n46201 , 
 n46202 , n366384 , n46204 , n366386 , n366387 , n46207 , n46208 , n366390 , n366391 , n46211 , 
 n366393 , n366394 , n366395 , n366396 , n366397 , n366398 , n366399 , n366400 , n366401 , n366402 , 
 n366403 , n366404 , n46224 , n46225 , n366407 , n46227 , n366409 , n46229 , n366411 , n366412 , 
 n46232 , n366414 , n366415 , n46235 , n46236 , n366418 , n46238 , n366420 , n366421 , n366422 , 
 n366423 , n366424 , n366425 , n366426 , n366427 , n366428 , n366429 , n366430 , n366431 , n366432 , 
 n366433 , n366434 , n366435 , n46255 , n366437 , n366438 , n366439 , n366440 , n366441 , n46261 , 
 n366443 , n366444 , n46264 , n366446 , n366447 , n366448 , n366449 , n46269 , n46270 , n46271 , 
 n366453 , n46273 , n46274 , n366456 , n46276 , n366458 , n46278 , n366460 , n46280 , n366462 , 
 n366463 , n46283 , n366465 , n366466 , n46286 , n366468 , n366469 , n46289 , n46290 , n366472 , 
 n366473 , n366474 , n366475 , n366476 , n46296 , n366478 , n366479 , n46299 , n366481 , n46301 , 
 n366483 , n46303 , n366485 , n366486 , n366487 , n46307 , n366489 , n366490 , n366491 , n366492 , 
 n366493 , n366494 , n46314 , n46315 , n366497 , n46317 , n366499 , n366500 , n46320 , n366502 , 
 n46322 , n366504 , n46324 , n366506 , n46326 , n366508 , n366509 , n366510 , n46330 , n366512 , 
 n366513 , n46333 , n366515 , n366516 , n46336 , n366518 , n46338 , n46339 , n46340 , n366522 , 
 n46342 , n366524 , n366525 , n366526 , n366527 , n46347 , n366529 , n366530 , n46350 , n366532 , 
 n366533 , n366534 , n366535 , n46355 , n366537 , n366538 , n366539 , n46359 , n366541 , n366542 , 
 n46362 , n366544 , n366545 , n366546 , n366547 , n366548 , n366549 , n366550 , n366551 , n366552 , 
 n366553 , n366554 , n366555 , n366556 , n46376 , n366558 , n366559 , n366560 , n366561 , n366562 , 
 n366563 , n46383 , n46384 , n46385 , n366567 , n366568 , n366569 , n46389 , n46390 , n366572 , 
 n46392 , n46393 , n366575 , n366576 , n46396 , n46397 , n366579 , n46399 , n46400 , n366582 , 
 n366583 , n366584 , n366585 , n366586 , n366587 , n366588 , n366589 , n366590 , n366591 , n46404 , 
 n366593 , n366594 , n46407 , n46408 , n366597 , n46410 , n366599 , n366600 , n366601 , n366602 , 
 n366603 , n366604 , n366605 , n46418 , n366607 , n366608 , n46421 , n366610 , n366611 , n366612 , 
 n366613 , n46426 , n366615 , n46428 , n46429 , n46430 , n366619 , n46432 , n366621 , n366622 , 
 n46435 , n366624 , n46437 , n46438 , n46439 , n366628 , n366629 , n366630 , n366631 , n46444 , 
 n366633 , n366634 , n366635 , n366636 , n366637 , n366638 , n366639 , n366640 , n46453 , n46454 , 
 n366643 , n366644 , n46457 , n366646 , n46459 , n366648 , n366649 , n366650 , n46463 , n366652 , 
 n366653 , n366654 , n366655 , n366656 , n46469 , n366658 , n366659 , n366660 , n46473 , n46474 , 
 n366663 , n46476 , n46477 , n366666 , n46479 , n366668 , n366669 , n366670 , n366671 , n366672 , 
 n366673 , n366674 , n366675 , n366676 , n366677 , n46490 , n46491 , n366680 , n366681 , n46494 , 
 n366683 , n366684 , n366685 , n366686 , n366687 , n46500 , n366689 , n366690 , n366691 , n366692 , 
 n46505 , n366694 , n46507 , n366696 , n46509 , n366698 , n46511 , n366700 , n46513 , n366702 , 
 n366703 , n366704 , n46517 , n366706 , n366707 , n366708 , n46521 , n46522 , n366711 , n366712 , 
 n366713 , n46526 , n366715 , n366716 , n366717 , n366718 , n366719 , n46532 , n366721 , n366722 , 
 n366723 , n366724 , n366725 , n46538 , n366727 , n366728 , n366729 , n366730 , n366731 , n366732 , 
 n46545 , n46546 , n46547 , n46548 , n46549 , n366738 , n366739 , n366740 , n46553 , n366742 , 
 n46555 , n46556 , n46557 , n366746 , n366747 , n366748 , n366749 , n46562 , n366751 , n366752 , 
 n46565 , n366754 , n366755 , n366756 , n366757 , n366758 , n366759 , n366760 , n366761 , n366762 , 
 n366763 , n366764 , n366765 , n366766 , n366767 , n366768 , n46581 , n46582 , n46583 , n366772 , 
 n366773 , n46586 , n46587 , n366776 , n366777 , n46590 , n366779 , n366780 , n46593 , n366782 , 
 n366783 , n366784 , n366785 , n46598 , n366787 , n366788 , n46601 , n46602 , n366791 , n366792 , 
 n46605 , n46606 , n46607 , n366796 , n46609 , n46610 , n46611 , n366800 , n366801 , n46614 , 
 n366803 , n366804 , n366805 , n366806 , n46619 , n46620 , n366809 , n366810 , n366811 , n46624 , 
 n46625 , n366814 , n46627 , n366816 , n46629 , n46630 , n46631 , n366820 , n366821 , n366822 , 
 n366823 , n46636 , n366825 , n366826 , n366827 , n46640 , n46641 , n366830 , n366831 , n46644 , 
 n366833 , n366834 , n366835 , n366836 , n366837 , n46650 , n366839 , n46652 , n46653 , n46654 , 
 n366843 , n366844 , n46657 , n366846 , n366847 , n366848 , n366849 , n46662 , n366851 , n366852 , 
 n46665 , n46666 , n366855 , n366856 , n366857 , n366858 , n46671 , n366860 , n366861 , n366862 , 
 n366863 , n366864 , n46677 , n46678 , n366867 , n46680 , n366869 , n46682 , n366871 , n366872 , 
 n366873 , n46686 , n366875 , n366876 , n366877 , n366878 , n366879 , n366880 , n46693 , n366882 , 
 n366883 , n46696 , n366885 , n366886 , n46699 , n366888 , n46701 , n46702 , n46703 , n366892 , 
 n366893 , n366894 , n366895 , n366896 , n366897 , n366898 , n366899 , n366900 , n366901 , n46714 , 
 n366903 , n366904 , n366905 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , 
 n366913 , n46726 , n366915 , n366916 , n366917 , n366918 , n366919 , n366920 , n366921 , n366922 , 
 n366923 , n366924 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , 
 n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n366940 , n366941 , n46754 , 
 n366943 , n366944 , n366945 , n46758 , n46759 , n366948 , n366949 , n366950 , n366951 , n366952 , 
 n46765 , n366954 , n366955 , n46768 , n366957 , n366958 , n366959 , n366960 , n366961 , n366962 , 
 n366963 , n366964 , n46777 , n366966 , n366967 , n366968 , n46781 , n366970 , n366971 , n366972 , 
 n366973 , n46786 , n366975 , n366976 , n46789 , n366978 , n366979 , n46792 , n366981 , n46794 , 
 n366983 , n366984 , n46797 , n366986 , n366987 , n366988 , n366989 , n366990 , n46803 , n46804 , 
 n366993 , n366994 , n366995 , n366996 , n366997 , n366998 , n366999 , n46812 , n367001 , n367002 , 
 n367003 , n46816 , n367005 , n367006 , n46819 , n367008 , n46821 , n367010 , n367011 , n46824 , 
 n367013 , n367014 , n367015 , n367016 , n46829 , n46830 , n367019 , n367020 , n46833 , n46834 , 
 n367023 , n46836 , n367025 , n367026 , n367027 , n367028 , n367029 , n46842 , n367031 , n367032 , 
 n367033 , n367034 , n46847 , n46848 , n367037 , n46850 , n367039 , n367040 , n367041 , n367042 , 
 n46855 , n367044 , n46857 , n46858 , n46859 , n367048 , n46861 , n46862 , n367051 , n367052 , 
 n367053 , n367054 , n367055 , n46868 , n367057 , n367058 , n367059 , n46872 , n367061 , n367062 , 
 n367063 , n367064 , n367065 , n367066 , n46879 , n46880 , n367069 , n46882 , n46883 , n367072 , 
 n367073 , n367074 , n367075 , n367076 , n46889 , n367078 , n367079 , n367080 , n367081 , n367082 , 
 n46895 , n367084 , n367085 , n46898 , n367087 , n46900 , n367089 , n46902 , n367091 , n46904 , 
 n367093 , n46906 , n367095 , n367096 , n46909 , n46910 , n46911 , n367100 , n367101 , n367102 , 
 n367103 , n367104 , n367105 , n367106 , n367107 , n46920 , n367109 , n367110 , n46923 , n367112 , 
 n367113 , n367114 , n46927 , n367116 , n367117 , n367118 , n46931 , n367120 , n367121 , n46934 , 
 n367123 , n367124 , n46937 , n367126 , n367127 , n367128 , n367129 , n367130 , n367131 , n367132 , 
 n367133 , n367134 , n46947 , n367136 , n367137 , n46950 , n367139 , n367140 , n367141 , n367142 , 
 n367143 , n367144 , n367145 , n46958 , n367147 , n46960 , n46961 , n367150 , n367151 , n46964 , 
 n367153 , n367154 , n46967 , n367156 , n46969 , n367158 , n367159 , n46972 , n367161 , n367162 , 
 n367163 , n46976 , n367165 , n367166 , n367167 , n367168 , n46981 , n46982 , n367171 , n367172 , 
 n46985 , n367174 , n46987 , n367176 , n46989 , n367178 , n367179 , n46992 , n367181 , n367182 , 
 n367183 , n367184 , n46997 , n46998 , n367187 , n47000 , n47001 , n367190 , n367191 , n367192 , 
 n367193 , n367194 , n367195 , n367196 , n367197 , n367198 , n367199 , n367200 , n47013 , n47014 , 
 n367203 , n367204 , n47017 , n367206 , n367207 , n47020 , n367209 , n367210 , n367211 , n47024 , 
 n367213 , n367214 , n47027 , n367216 , n367217 , n47030 , n47031 , n367220 , n367221 , n367222 , 
 n367223 , n47036 , n367225 , n367226 , n47039 , n367228 , n367229 , n47042 , n367231 , n367232 , 
 n367233 , n367234 , n47047 , n367236 , n47049 , n367238 , n367239 , n367240 , n47053 , n367242 , 
 n47055 , n367244 , n367245 , n367246 , n47059 , n367248 , n367249 , n47062 , n47063 , n367252 , 
 n47065 , n367254 , n367255 , n367256 , n367257 , n367258 , n367259 , n47072 , n367261 , n367262 , 
 n47075 , n367264 , n367265 , n47078 , n367267 , n367268 , n367269 , n367270 , n367271 , n367272 , 
 n367273 , n367274 , n367275 , n367276 , n47089 , n367278 , n367279 , n367280 , n367281 , n367282 , 
 n47095 , n367284 , n367285 , n367286 , n367287 , n367288 , n367289 , n367290 , n367291 , n47104 , 
 n367293 , n47106 , n367295 , n367296 , n367297 , n367298 , n367299 , n367300 , n47113 , n367302 , 
 n367303 , n367304 , n367305 , n367306 , n367307 , n367308 , n367309 , n367310 , n367311 , n47124 , 
 n47125 , n47126 , n47127 , n47128 , n47129 , n367318 , n47131 , n367320 , n47133 , n367322 , 
 n47135 , n367324 , n367325 , n367326 , n367327 , n367328 , n367329 , n47142 , n367331 , n367332 , 
 n367333 , n367334 , n367335 , n367336 , n47149 , n367338 , n367339 , n367340 , n367341 , n367342 , 
 n47155 , n367344 , n367345 , n47158 , n367347 , n367348 , n367349 , n367350 , n47163 , n47164 , 
 n47165 , n367354 , n367355 , n367356 , n47169 , n47170 , n367359 , n367360 , n47173 , n47174 , 
 n367363 , n47176 , n367365 , n47178 , n47179 , n367368 , n47181 , n47182 , n367371 , n47184 , 
 n367373 , n47186 , n367375 , n47188 , n47189 , n367378 , n47191 , n47192 , n47193 , n367382 , 
 n47195 , n367384 , n367385 , n367386 , n47199 , n367388 , n47201 , n367390 , n367391 , n47204 , 
 n47205 , n367394 , n47207 , n367396 , n367397 , n47210 , n367399 , n47212 , n47213 , n367402 , 
 n367403 , n47216 , n367405 , n47218 , n367407 , n47220 , n367409 , n47222 , n47223 , n47224 , 
 n367413 , n47226 , n47227 , n367416 , n367417 , n367418 , n367419 , n47232 , n367421 , n367422 , 
 n367423 , n47236 , n367425 , n367426 , n367427 , n367428 , n367429 , n47242 , n367431 , n367432 , 
 n47245 , n47246 , n367435 , n367436 , n47249 , n367438 , n47251 , n367440 , n47253 , n47254 , 
 n47255 , n367444 , n47257 , n367446 , n47259 , n367448 , n47261 , n47262 , n367451 , n47264 , 
 n367453 , n367454 , n367455 , n47268 , n367457 , n367458 , n367459 , n367460 , n367461 , n367462 , 
 n367463 , n367464 , n367465 , n367466 , n367467 , n367468 , n367469 , n367470 , n367471 , n367472 , 
 n367473 , n367474 , n47287 , n367476 , n47289 , n47290 , n367479 , n367480 , n367481 , n367482 , 
 n47295 , n367484 , n367485 , n367486 , n367487 , n367488 , n367489 , n367490 , n367491 , n367492 , 
 n47305 , n367494 , n367495 , n47308 , n367497 , n367498 , n47311 , n367500 , n47313 , n367502 , 
 n367503 , n47316 , n367505 , n47318 , n47319 , n367508 , n47321 , n367510 , n47323 , n367512 , 
 n367513 , n47326 , n367515 , n367516 , n367517 , n47330 , n47331 , n367520 , n47333 , n367522 , 
 n367523 , n367524 , n367525 , n47338 , n367527 , n367528 , n47341 , n367530 , n367531 , n47344 , 
 n47345 , n367534 , n47347 , n367536 , n47349 , n367538 , n367539 , n367540 , n367541 , n367542 , 
 n367543 , n47356 , n367545 , n47358 , n367547 , n47360 , n367549 , n47362 , n47363 , n367552 , 
 n367553 , n47366 , n367555 , n47368 , n47369 , n47370 , n367559 , n47372 , n367561 , n367562 , 
 n367563 , n367564 , n367565 , n367566 , n47379 , n367568 , n47381 , n367570 , n367571 , n367572 , 
 n47385 , n47386 , n367575 , n367576 , n367577 , n367578 , n367579 , n47392 , n367581 , n367582 , 
 n47395 , n47396 , n367585 , n47398 , n367587 , n367588 , n47401 , n367590 , n47403 , n367592 , 
 n367593 , n367594 , n367595 , n47408 , n367597 , n367598 , n47411 , n367600 , n367601 , n47414 , 
 n367603 , n367604 , n367605 , n47418 , n367607 , n367608 , n47421 , n367610 , n367611 , n47424 , 
 n367613 , n367614 , n367615 , n47428 , n47429 , n367618 , n47431 , n47432 , n47433 , n367622 , 
 n367623 , n47436 , n47437 , n367626 , n367627 , n47440 , n367629 , n367630 , n47443 , n367632 , 
 n367633 , n47446 , n367635 , n47448 , n47449 , n47450 , n367639 , n47452 , n367641 , n367642 , 
 n47455 , n367644 , n47457 , n367646 , n47459 , n367648 , n47461 , n47462 , n367651 , n47464 , 
 n367653 , n47466 , n47467 , n367656 , n47469 , n367658 , n47471 , n47472 , n367661 , n367662 , 
 n47475 , n367664 , n367665 , n367666 , n367667 , n47480 , n367669 , n47482 , n367671 , n367672 , 
 n367673 , n47486 , n47487 , n47488 , n47489 , n47490 , n367679 , n367680 , n367681 , n367682 , 
 n47495 , n47496 , n47497 , n367686 , n47499 , n47500 , n367689 , n47502 , n367691 , n47504 , 
 n47505 , n47506 , n47507 , n367696 , n47509 , n367698 , n47511 , n367700 , n367701 , n47514 , 
 n367703 , n47516 , n367705 , n47518 , n367707 , n367708 , n47521 , n367710 , n367711 , n47524 , 
 n367713 , n367714 , n367715 , n367716 , n367717 , n367718 , n47531 , n47532 , n47533 , n47534 , 
 n47535 , n47536 , n47537 , n367726 , n367727 , n367728 , n367729 , n367730 , n367731 , n367732 , 
 n367733 , n367734 , n47547 , n367736 , n367737 , n367738 , n367739 , n47552 , n47553 , n47554 , 
 n367743 , n47556 , n367745 , n47558 , n47559 , n367748 , n367749 , n47562 , n367751 , n367752 , 
 n47565 , n367754 , n367755 , n367756 , n47569 , n367758 , n367759 , n367760 , n47573 , n367762 , 
 n367763 , n367764 , n367765 , n367766 , n367767 , n367768 , n367769 , n367770 , n47583 , n367772 , 
 n367773 , n47586 , n367775 , n47588 , n367777 , n367778 , n47591 , n367780 , n367781 , n47594 , 
 n367783 , n47596 , n367785 , n367786 , n367787 , n367788 , n367789 , n47602 , n367791 , n367792 , 
 n367793 , n367794 , n47607 , n367796 , n367797 , n367798 , n367799 , n367800 , n47613 , n47614 , 
 n47615 , n47616 , n47617 , n47618 , n367807 , n367808 , n367809 , n367810 , n367811 , n367812 , 
 n367813 , n367814 , n367815 , n367816 , n47629 , n367818 , n47631 , n367820 , n367821 , n47634 , 
 n47635 , n47636 , n367825 , n367826 , n367827 , n367828 , n367829 , n367830 , n367831 , n367832 , 
 n367833 , n367834 , n367835 , n367836 , n367837 , n367838 , n367839 , n367840 , n367841 , n47654 , 
 n367843 , n367844 , n47657 , n367846 , n47659 , n47660 , n367849 , n367850 , n47663 , n367852 , 
 n47665 , n47666 , n367855 , n367856 , n47669 , n367858 , n367859 , n367860 , n367861 , n367862 , 
 n367863 , n367864 , n367865 , n367866 , n367867 , n367868 , n47681 , n367870 , n47683 , n47684 , 
 n367873 , n367874 , n367875 , n367876 , n367877 , n47690 , n367879 , n367880 , n47693 , n367882 , 
 n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n367889 , n47702 , n367891 , n367892 , 
 n367893 , n367894 , n367895 , n367896 , n367897 , n47710 , n367899 , n367900 , n367901 , n367902 , 
 n47715 , n367904 , n367905 , n47718 , n367907 , n367908 , n47721 , n367910 , n367911 , n47724 , 
 n367913 , n367914 , n47727 , n367916 , n367917 , n47730 , n47731 , n367920 , n367921 , n367922 , 
 n367923 , n367924 , n367925 , n367926 , n367927 , n47733 , n367929 , n367930 , n367931 , n367932 , 
 n367933 , n367934 , n367935 , n367936 , n47742 , n47743 , n47744 , n367940 , n367941 , n367942 , 
 n47748 , n367944 , n47750 , n367946 , n47752 , n47753 , n47754 , n47755 , n47756 , n367952 , 
 n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , 
 n47768 , n367964 , n47770 , n47771 , n47772 , n367968 , n47774 , n47775 , n367971 , n367972 , 
 n367973 , n367974 , n367975 , n47781 , n47782 , n367978 , n367979 , n47785 , n367981 , n367982 , 
 n47788 , n367984 , n367985 , n47791 , n47792 , n367988 , n367989 , n367990 , n367991 , n367992 , 
 n367993 , n367994 , n367995 , n367996 , n367997 , n367998 , n367999 , n368000 , n368001 , n368002 , 
 n368003 , n47809 , n47810 , n368006 , n47812 , n368008 , n368009 , n368010 , n368011 , n368012 , 
 n368013 , n368014 , n368015 , n368016 , n368017 , n368018 , n47824 , n368020 , n368021 , n47827 , 
 n368023 , n368024 , n47830 , n47831 , n47832 , n47833 , n368029 , n47835 , n368031 , n368032 , 
 n368033 , n47839 , n47840 , n47841 , n47842 , n368038 , n368039 , n47845 , n47846 , n47847 , 
 n47848 , n47849 , n368045 , n368046 , n368047 , n368048 , n47854 , n47855 , n368051 , n47857 , 
 n368053 , n47859 , n368055 , n368056 , n368057 , n368058 , n47864 , n47865 , n47866 , n47867 , 
 n368063 , n368064 , n47870 , n368066 , n47872 , n368068 , n47874 , n47875 , n47876 , n368072 , 
 n47878 , n368074 , n47880 , n368076 , n47882 , n368078 , n368079 , n368080 , n368081 , n47887 , 
 n368083 , n47889 , n368085 , n368086 , n368087 , n368088 , n368089 , n368090 , n368091 , n368092 , 
 n368093 , n368094 , n47900 , n368096 , n368097 , n368098 , n368099 , n368100 , n368101 , n368102 , 
 n368103 , n368104 , n47910 , n368106 , n47912 , n368108 , n368109 , n368110 , n47916 , n368112 , 
 n368113 , n47919 , n368115 , n368116 , n47922 , n368118 , n47924 , n368120 , n368121 , n47927 , 
 n368123 , n47929 , n368125 , n47931 , n368127 , n368128 , n368129 , n47935 , n368131 , n368132 , 
 n47938 , n368134 , n368135 , n368136 , n368137 , n368138 , n368139 , n368140 , n368141 , n368142 , 
 n47948 , n368144 , n368145 , n47951 , n368147 , n47953 , n368149 , n368150 , n368151 , n368152 , 
 n368153 , n368154 , n368155 , n47961 , n368157 , n47963 , n368159 , n368160 , n47966 , n368162 , 
 n368163 , n368164 , n368165 , n368166 , n47972 , n368168 , n368169 , n368170 , n368171 , n368172 , 
 n368173 , n368174 , n368175 , n368176 , n47982 , n368178 , n368179 , n47985 , n368181 , n368182 , 
 n47988 , n47989 , n368185 , n368186 , n368187 , n368188 , n368189 , n368190 , n47996 , n368192 , 
 n368193 , n368194 , n368195 , n368196 , n368197 , n368198 , n368199 , n368200 , n368201 , n368202 , 
 n48008 , n368204 , n368205 , n368206 , n48012 , n368208 , n368209 , n48015 , n368211 , n368212 , 
 n48018 , n48019 , n368215 , n368216 , n368217 , n368218 , n368219 , n368220 , n368221 , n48027 , 
 n368223 , n368224 , n368225 , n368226 , n368227 , n368228 , n368229 , n368230 , n368231 , n368232 , 
 n48038 , n368234 , n368235 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , 
 n368243 , n368244 , n48050 , n368246 , n368247 , n368248 , n48054 , n368250 , n48056 , n48057 , 
 n48058 , n368254 , n368255 , n48061 , n368257 , n368258 , n368259 , n368260 , n48066 , n368262 , 
 n368263 , n368264 , n368265 , n368266 , n368267 , n48073 , n48074 , n48075 , n48076 , n48077 , 
 n48078 , n368274 , n368275 , n368276 , n368277 , n48083 , n48084 , n48085 , n368281 , n48087 , 
 n368283 , n368284 , n368285 , n368286 , n368287 , n368288 , n48094 , n368290 , n368291 , n48097 , 
 n48098 , n368294 , n368295 , n48101 , n368297 , n368298 , n48104 , n368300 , n368301 , n368302 , 
 n368303 , n368304 , n368305 , n368306 , n368307 , n368308 , n368309 , n368310 , n48116 , n48117 , 
 n368313 , n48119 , n368315 , n368316 , n48122 , n48123 , n368319 , n368320 , n48126 , n368322 , 
 n368323 , n368324 , n48130 , n368326 , n48132 , n48133 , n368329 , n368330 , n368331 , n368332 , 
 n368333 , n368334 , n368335 , n48141 , n48142 , n368338 , n48144 , n368340 , n368341 , n368342 , 
 n48148 , n48149 , n368345 , n48151 , n48152 , n368348 , n48154 , n48155 , n368351 , n368352 , 
 n368353 , n368354 , n48160 , n48161 , n368357 , n368358 , n48164 , n368360 , n48166 , n368362 , 
 n48168 , n368364 , n368365 , n368366 , n368367 , n368368 , n368369 , n48175 , n368371 , n368372 , 
 n368373 , n368374 , n368375 , n368376 , n368377 , n48183 , n368379 , n368380 , n368381 , n48187 , 
 n368383 , n368384 , n368385 , n368386 , n48192 , n368388 , n368389 , n368390 , n48196 , n368392 , 
 n48198 , n368394 , n48200 , n48201 , n368397 , n368398 , n368399 , n48205 , n48206 , n48207 , 
 n368403 , n48209 , n48210 , n368406 , n368407 , n48213 , n368409 , n368410 , n48216 , n48217 , 
 n368413 , n368414 , n368415 , n368416 , n368417 , n368418 , n48224 , n48225 , n368421 , n368422 , 
 n368423 , n368424 , n368425 , n368426 , n368427 , n368428 , n368429 , n368430 , n48236 , n368432 , 
 n368433 , n48239 , n368435 , n368436 , n368437 , n368438 , n368439 , n368440 , n368441 , n368442 , 
 n48248 , n48249 , n48250 , n48251 , n48252 , n368448 , n368449 , n368450 , n368451 , n368452 , 
 n368453 , n368454 , n368455 , n368456 , n48262 , n368458 , n368459 , n368460 , n368461 , n368462 , 
 n48268 , n368464 , n368465 , n368466 , n48272 , n48273 , n368469 , n368470 , n48276 , n368472 , 
 n368473 , n368474 , n48280 , n48281 , n368477 , n368478 , n48284 , n48285 , n48286 , n368482 , 
 n368483 , n368484 , n368485 , n368486 , n48292 , n368488 , n48294 , n368490 , n368491 , n368492 , 
 n48298 , n48299 , n48300 , n368496 , n48302 , n48303 , n368499 , n48305 , n368501 , n368502 , 
 n48308 , n48309 , n368505 , n368506 , n48312 , n368508 , n368509 , n368510 , n368511 , n48317 , 
 n368513 , n48319 , n368515 , n368516 , n48322 , n368518 , n368519 , n48325 , n368521 , n368522 , 
 n48328 , n368524 , n368525 , n368526 , n368527 , n368528 , n368529 , n368530 , n368531 , n368532 , 
 n368533 , n368534 , n368535 , n368536 , n368537 , n368538 , n48338 , n368540 , n368541 , n48341 , 
 n368543 , n48343 , n48344 , n48345 , n368547 , n368548 , n368549 , n368550 , n48350 , n368552 , 
 n48352 , n368554 , n48354 , n48355 , n48356 , n368558 , n368559 , n48359 , n368561 , n368562 , 
 n368563 , n368564 , n368565 , n368566 , n368567 , n48367 , n368569 , n368570 , n368571 , n48371 , 
 n368573 , n368574 , n368575 , n368576 , n368577 , n368578 , n368579 , n48379 , n368581 , n368582 , 
 n48382 , n368584 , n368585 , n368586 , n368587 , n368588 , n368589 , n368590 , n368591 , n368592 , 
 n368593 , n368594 , n48394 , n368596 , n48396 , n368598 , n368599 , n368600 , n368601 , n368602 , 
 n368603 , n368604 , n368605 , n368606 , n368607 , n368608 , n368609 , n368610 , n368611 , n368612 , 
 n368613 , n368614 , n368615 , n48415 , n368617 , n48417 , n48418 , n368620 , n368621 , n368622 , 
 n368623 , n368624 , n368625 , n368626 , n368627 , n48427 , n48428 , n368630 , n368631 , n48431 , 
 n368633 , n368634 , n48434 , n368636 , n368637 , n48437 , n368639 , n368640 , n368641 , n368642 , 
 n48442 , n368644 , n368645 , n48445 , n368647 , n368648 , n48448 , n368650 , n368651 , n48451 , 
 n48452 , n368654 , n368655 , n368656 , n368657 , n48457 , n48458 , n48459 , n368661 , n368662 , 
 n368663 , n368664 , n368665 , n368666 , n368667 , n368668 , n48468 , n368670 , n368671 , n368672 , 
 n368673 , n368674 , n368675 , n48475 , n368677 , n368678 , n48478 , n368680 , n368681 , n368682 , 
 n368683 , n368684 , n368685 , n368686 , n368687 , n368688 , n368689 , n368690 , n48490 , n368692 , 
 n48492 , n48493 , n368695 , n368696 , n48496 , n368698 , n368699 , n368700 , n368701 , n368702 , 
 n48502 , n368704 , n368705 , n368706 , n48506 , n368708 , n368709 , n368710 , n368711 , n368712 , 
 n48512 , n368714 , n368715 , n368716 , n48516 , n48517 , n368719 , n368720 , n48520 , n48521 , 
 n368723 , n368724 , n368725 , n368726 , n368727 , n48527 , n368729 , n368730 , n48530 , n48531 , 
 n368733 , n368734 , n48534 , n368736 , n368737 , n368738 , n48538 , n368740 , n368741 , n368742 , 
 n48542 , n368744 , n368745 , n368746 , n368747 , n368748 , n368749 , n48549 , n368751 , n368752 , 
 n48552 , n48553 , n368755 , n368756 , n48556 , n368758 , n48558 , n368760 , n368761 , n48561 , 
 n368763 , n48563 , n368765 , n368766 , n48566 , n48567 , n48568 , n368770 , n48570 , n48571 , 
 n368773 , n48573 , n368775 , n368776 , n368777 , n368778 , n368779 , n48579 , n368781 , n368782 , 
 n48582 , n368784 , n368785 , n48585 , n368787 , n368788 , n368789 , n368790 , n368791 , n368792 , 
 n368793 , n368794 , n368795 , n368796 , n368797 , n48597 , n368799 , n368800 , n48600 , n368802 , 
 n368803 , n48603 , n48604 , n368806 , n48606 , n368808 , n368809 , n48609 , n368811 , n368812 , 
 n368813 , n368814 , n368815 , n368816 , n368817 , n368818 , n368819 , n368820 , n368821 , n368822 , 
 n368823 , n368824 , n48624 , n368826 , n368827 , n368828 , n368829 , n368830 , n48630 , n48631 , 
 n368833 , n368834 , n48634 , n368836 , n368837 , n368838 , n368839 , n368840 , n48640 , n368842 , 
 n48642 , n368844 , n368845 , n368846 , n48646 , n368848 , n48648 , n368850 , n368851 , n368852 , 
 n368853 , n368854 , n48654 , n368856 , n48656 , n368858 , n48658 , n48659 , n368861 , n368862 , 
 n48662 , n368864 , n368865 , n48665 , n368867 , n368868 , n48668 , n48669 , n48670 , n48671 , 
 n48672 , n48673 , n48674 , n368876 , n48676 , n368878 , n368879 , n48679 , n48680 , n368882 , 
 n368883 , n48683 , n48684 , n368886 , n48686 , n368888 , n48688 , n48689 , n368891 , n368892 , 
 n48692 , n368894 , n368895 , n48695 , n368897 , n48697 , n48698 , n48699 , n48700 , n48701 , 
 n48702 , n368904 , n48704 , n368906 , n368907 , n48707 , n368909 , n368910 , n48710 , n368912 , 
 n48712 , n368914 , n368915 , n48715 , n368917 , n368918 , n48718 , n368920 , n368921 , n48721 , 
 n368923 , n368924 , n368925 , n48725 , n368927 , n368928 , n368929 , n368930 , n48730 , n368932 , 
 n368933 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n368940 , n48740 , n368942 , 
 n48742 , n368944 , n368945 , n48745 , n368947 , n368948 , n368949 , n368950 , n368951 , n368952 , 
 n368953 , n368954 , n48754 , n368956 , n368957 , n368958 , n368959 , n368960 , n368961 , n368962 , 
 n368963 , n368964 , n368965 , n368966 , n48766 , n368968 , n48768 , n48769 , n368971 , n48771 , 
 n368973 , n368974 , n48774 , n368976 , n368977 , n48777 , n368979 , n368980 , n48780 , n48781 , 
 n368983 , n368984 , n368985 , n368986 , n368987 , n48787 , n368989 , n368990 , n48790 , n48791 , 
 n48792 , n368994 , n368995 , n48795 , n368997 , n368998 , n368999 , n369000 , n369001 , n48801 , 
 n48802 , n369004 , n369005 , n48805 , n48806 , n369008 , n48808 , n369010 , n48810 , n369012 , 
 n48812 , n48813 , n369015 , n369016 , n369017 , n369018 , n369019 , n369020 , n48820 , n369022 , 
 n369023 , n48823 , n369025 , n369026 , n369027 , n369028 , n369029 , n369030 , n48830 , n48831 , 
 n369033 , n48833 , n369035 , n369036 , n369037 , n369038 , n369039 , n369040 , n369041 , n369042 , 
 n48842 , n369044 , n369045 , n369046 , n48846 , n369048 , n48848 , n369050 , n369051 , n369052 , 
 n369053 , n369054 , n369055 , n369056 , n369057 , n369058 , n369059 , n369060 , n369061 , n48861 , 
 n369063 , n48863 , n369065 , n369066 , n369067 , n48867 , n48868 , n48869 , n48870 , n369072 , 
 n369073 , n369074 , n369075 , n369076 , n48876 , n369078 , n369079 , n369080 , n369081 , n369082 , 
 n369083 , n48883 , n369085 , n369086 , n369087 , n48887 , n369089 , n369090 , n369091 , n369092 , 
 n369093 , n369094 , n369095 , n369096 , n369097 , n369098 , n369099 , n369100 , n369101 , n369102 , 
 n369103 , n369104 , n48904 , n48905 , n369107 , n369108 , n369109 , n369110 , n369111 , n48911 , 
 n369113 , n48913 , n48914 , n48915 , n48916 , n369118 , n48918 , n369120 , n369121 , n369122 , 
 n48922 , n369124 , n48924 , n369126 , n48926 , n369128 , n48928 , n369130 , n48930 , n48931 , 
 n369133 , n48933 , n369135 , n48935 , n48936 , n48937 , n369139 , n48939 , n369141 , n48941 , 
 n48942 , n369144 , n369145 , n48945 , n369147 , n369148 , n48948 , n369150 , n369151 , n48951 , 
 n369153 , n369154 , n48954 , n369156 , n369157 , n369158 , n369159 , n369160 , n369161 , n369162 , 
 n369163 , n369164 , n369165 , n369166 , n369167 , n369168 , n48968 , n48969 , n48970 , n48971 , 
 n48972 , n369174 , n48974 , n369176 , n48976 , n48977 , n369179 , n48979 , n48980 , n369182 , 
 n369183 , n48983 , n369185 , n369186 , n48986 , n369188 , n48988 , n48989 , n369191 , n369192 , 
 n48992 , n48993 , n369195 , n369196 , n48996 , n369198 , n369199 , n48999 , n49000 , n369202 , 
 n369203 , n49003 , n369205 , n369206 , n369207 , n369208 , n369209 , n49009 , n369211 , n49011 , 
 n49012 , n49013 , n369215 , n49015 , n369217 , n369218 , n369219 , n369220 , n369221 , n49021 , 
 n369223 , n369224 , n49024 , n369226 , n49026 , n49027 , n49028 , n369230 , n369231 , n49031 , 
 n369233 , n49033 , n49034 , n369236 , n369237 , n49037 , n369239 , n369240 , n49040 , n369242 , 
 n369243 , n369244 , n49044 , n369246 , n49046 , n49047 , n369249 , n369250 , n49050 , n369252 , 
 n369253 , n369254 , n369255 , n369256 , n49056 , n369258 , n49058 , n369260 , n369261 , n49061 , 
 n49062 , n369264 , n369265 , n49065 , n369267 , n369268 , n49068 , n369270 , n369271 , n49071 , 
 n369273 , n369274 , n369275 , n49075 , n369277 , n369278 , n49078 , n369280 , n49080 , n369282 , 
 n369283 , n49083 , n49084 , n369286 , n369287 , n49087 , n369289 , n369290 , n49090 , n369292 , 
 n369293 , n369294 , n369295 , n369296 , n369297 , n49097 , n369299 , n369300 , n49100 , n49101 , 
 n49102 , n369304 , n369305 , n49105 , n369307 , n49107 , n49108 , n369310 , n49110 , n369312 , 
 n49112 , n369314 , n49114 , n369316 , n369317 , n369318 , n369319 , n369320 , n49120 , n369322 , 
 n49122 , n369324 , n369325 , n49125 , n49126 , n49127 , n369329 , n49129 , n369331 , n49131 , 
 n49132 , n369334 , n49134 , n369336 , n49136 , n369338 , n369339 , n49139 , n369341 , n49141 , 
 n369343 , n369344 , n49144 , n49145 , n369347 , n49147 , n369349 , n369350 , n49150 , n369352 , 
 n369353 , n49153 , n49154 , n369356 , n369357 , n49157 , n369359 , n369360 , n369361 , n49161 , 
 n369363 , n369364 , n369365 , n369366 , n49166 , n49167 , n49168 , n369370 , n369371 , n369372 , 
 n49172 , n369374 , n49174 , n369376 , n49176 , n369378 , n49178 , n369380 , n369381 , n369382 , 
 n49182 , n369384 , n369385 , n369386 , n369387 , n369388 , n49188 , n369390 , n369391 , n369392 , 
 n369393 , n369394 , n369395 , n369396 , n369397 , n369398 , n369399 , n369400 , n49200 , n49201 , 
 n369403 , n49203 , n49204 , n369406 , n369407 , n49207 , n369409 , n49209 , n49210 , n369412 , 
 n369413 , n369414 , n369415 , n369416 , n369417 , n49217 , n369419 , n369420 , n49218 , n369422 , 
 n369423 , n369424 , n369425 , n49223 , n369427 , n369428 , n369429 , n49227 , n369431 , n369432 , 
 n49230 , n49231 , n49232 , n49233 , n369437 , n369438 , n369439 , n49237 , n369441 , n369442 , 
 n369443 , n369444 , n369445 , n49243 , n369447 , n369448 , n369449 , n49247 , n369451 , n49249 , 
 n49250 , n369454 , n369455 , n369456 , n369457 , n369458 , n49256 , n369460 , n369461 , n49259 , 
 n369463 , n369464 , n49262 , n369466 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , 
 n369473 , n369474 , n369475 , n49273 , n369477 , n369478 , n49276 , n369480 , n369481 , n49279 , 
 n369483 , n369484 , n369485 , n369486 , n369487 , n49285 , n369489 , n369490 , n369491 , n369492 , 
 n369493 , n369494 , n369495 , n369496 , n369497 , n369498 , n49296 , n369500 , n369501 , n49299 , 
 n369503 , n369504 , n369505 , n369506 , n369507 , n369508 , n49306 , n369510 , n49308 , n369512 , 
 n49310 , n369514 , n49312 , n49313 , n369517 , n49315 , n49316 , n49317 , n49318 , n49319 , 
 n49320 , n49321 , n369525 , n49323 , n369527 , n369528 , n369529 , n369530 , n369531 , n369532 , 
 n49330 , n49331 , n369535 , n49333 , n369537 , n49335 , n369539 , n369540 , n49338 , n49339 , 
 n369543 , n369544 , n369545 , n369546 , n369547 , n369548 , n369549 , n369550 , n369551 , n49349 , 
 n369553 , n369554 , n369555 , n369556 , n369557 , n49355 , n369559 , n369560 , n369561 , n49359 , 
 n369563 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n369570 , n369571 , n369572 , 
 n369573 , n369574 , n369575 , n369576 , n369577 , n369578 , n369579 , n369580 , n369581 , n369582 , 
 n369583 , n369584 , n369585 , n369586 , n369587 , n369588 , n369589 , n369590 , n49388 , n369592 , 
 n369593 , n369594 , n369595 , n369596 , n369597 , n369598 , n369599 , n369600 , n49398 , n49399 , 
 n369603 , n369604 , n369605 , n49403 , n369607 , n49405 , n49406 , n369610 , n369611 , n49409 , 
 n369613 , n49411 , n369615 , n49413 , n49414 , n369618 , n369619 , n369620 , n369621 , n369622 , 
 n369623 , n369624 , n369625 , n369626 , n369627 , n369628 , n369629 , n369630 , n369631 , n369632 , 
 n369633 , n369634 , n369635 , n369636 , n369637 , n369638 , n369639 , n49437 , n369641 , n369642 , 
 n369643 , n49441 , n49442 , n369646 , n49444 , n369648 , n369649 , n49447 , n369651 , n369652 , 
 n49450 , n369654 , n369655 , n49453 , n49454 , n49455 , n49456 , n49457 , n369661 , n369662 , 
 n49460 , n369664 , n49462 , n369666 , n49464 , n369668 , n369669 , n49467 , n49468 , n49469 , 
 n369673 , n369674 , n49472 , n369676 , n369677 , n369678 , n49476 , n369680 , n369681 , n49479 , 
 n369683 , n49481 , n49482 , n369686 , n369687 , n49485 , n369689 , n369690 , n49488 , n49489 , 
 n369693 , n369694 , n49492 , n369696 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , 
 n369703 , n49501 , n369705 , n49503 , n49504 , n369708 , n369709 , n49507 , n369711 , n369712 , 
 n49510 , n369714 , n49512 , n369716 , n49514 , n369718 , n49516 , n369720 , n49518 , n369722 , 
 n369723 , n369724 , n369725 , n369726 , n369727 , n369728 , n369729 , n369730 , n49528 , n369732 , 
 n369733 , n369734 , n49532 , n369736 , n369737 , n49535 , n369739 , n49537 , n369741 , n369742 , 
 n369743 , n369744 , n49542 , n369746 , n49544 , n369748 , n49546 , n49547 , n369751 , n49549 , 
 n369753 , n49551 , n49552 , n369756 , n49554 , n369758 , n369759 , n49557 , n369761 , n369762 , 
 n369763 , n369764 , n49562 , n369766 , n369767 , n49565 , n369769 , n49567 , n49568 , n49569 , 
 n369773 , n369774 , n369775 , n369776 , n369777 , n369778 , n369779 , n49577 , n49578 , n49579 , 
 n369783 , n49581 , n49582 , n369786 , n49584 , n49585 , n369789 , n369790 , n49588 , n369792 , 
 n369793 , n369794 , n369795 , n369796 , n49594 , n369798 , n49596 , n369800 , n369801 , n369802 , 
 n49600 , n369804 , n369805 , n49603 , n49604 , n49605 , n369809 , n369810 , n49608 , n49609 , 
 n369813 , n369814 , n369815 , n369816 , n369817 , n49615 , n369819 , n369820 , n369821 , n369822 , 
 n369823 , n369824 , n49622 , n369826 , n49624 , n369828 , n369829 , n49627 , n369831 , n369832 , 
 n49630 , n369834 , n369835 , n49633 , n49634 , n369838 , n369839 , n369840 , n369841 , n369842 , 
 n49640 , n49641 , n369845 , n369846 , n369847 , n369848 , n49646 , n49647 , n369851 , n369852 , 
 n49650 , n369854 , n369855 , n49653 , n369857 , n49655 , n49656 , n369860 , n49658 , n49659 , 
 n369863 , n369864 , n49662 , n369866 , n369867 , n369868 , n369869 , n369870 , n369871 , n49669 , 
 n369873 , n49671 , n49672 , n49673 , n369877 , n369878 , n369879 , n369880 , n369881 , n49679 , 
 n369883 , n369884 , n49682 , n369886 , n49684 , n369888 , n49686 , n369890 , n369891 , n49689 , 
 n369893 , n369894 , n49692 , n369896 , n369897 , n369898 , n49696 , n369900 , n369901 , n369902 , 
 n49700 , n369904 , n369905 , n369906 , n369907 , n369908 , n369909 , n369910 , n369911 , n369912 , 
 n369913 , n369914 , n49712 , n369916 , n369917 , n49715 , n369919 , n369920 , n49718 , n369922 , 
 n49720 , n369924 , n369925 , n49723 , n369927 , n49725 , n369929 , n369930 , n369931 , n49729 , 
 n369933 , n49731 , n369935 , n369936 , n369937 , n49735 , n369939 , n369940 , n369941 , n369942 , 
 n369943 , n49741 , n369945 , n49743 , n369947 , n369948 , n49746 , n369950 , n369951 , n369952 , 
 n369953 , n369954 , n369955 , n369956 , n369957 , n369958 , n369959 , n369960 , n369961 , n49759 , 
 n369963 , n369964 , n49762 , n369966 , n369967 , n369968 , n369969 , n369970 , n49768 , n369972 , 
 n369973 , n369974 , n49772 , n369976 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , 
 n369983 , n369984 , n49782 , n369986 , n369987 , n369988 , n369989 , n369990 , n369991 , n49789 , 
 n369993 , n369994 , n369995 , n49793 , n369997 , n369998 , n49796 , n370000 , n370001 , n370002 , 
 n370003 , n370004 , n370005 , n370006 , n370007 , n370008 , n370009 , n370010 , n370011 , n370012 , 
 n49810 , n370014 , n370015 , n370016 , n49814 , n370018 , n370019 , n370020 , n370021 , n370022 , 
 n370023 , n370024 , n370025 , n370026 , n370027 , n370028 , n49826 , n49827 , n49828 , n370032 , 
 n49830 , n370034 , n370035 , n370036 , n49834 , n370038 , n49836 , n370040 , n370041 , n370042 , 
 n370043 , n370044 , n49842 , n370046 , n49844 , n370048 , n49846 , n370050 , n370051 , n49849 , 
 n370053 , n370054 , n49852 , n370056 , n370057 , n49855 , n370059 , n370060 , n49858 , n49859 , 
 n370063 , n370064 , n370065 , n370066 , n370067 , n370068 , n49866 , n370070 , n370071 , n370072 , 
 n370073 , n370074 , n370075 , n370076 , n370077 , n370078 , n370079 , n370080 , n49878 , n370082 , 
 n370083 , n49881 , n370085 , n370086 , n49884 , n49885 , n370089 , n370090 , n370091 , n370092 , 
 n370093 , n370094 , n49892 , n370096 , n370097 , n49895 , n370099 , n370100 , n49898 , n370102 , 
 n49900 , n49901 , n370105 , n370106 , n370107 , n370108 , n49906 , n370110 , n49908 , n370112 , 
 n49910 , n370114 , n49912 , n370116 , n370117 , n370118 , n49916 , n49917 , n370121 , n370122 , 
 n49920 , n370124 , n370125 , n49923 , n370127 , n370128 , n49926 , n49927 , n370131 , n370132 , 
 n49930 , n370134 , n370135 , n370136 , n370137 , n370138 , n370139 , n370140 , n370141 , n49939 , 
 n49940 , n49941 , n49942 , n370146 , n49944 , n370148 , n370149 , n370150 , n370151 , n370152 , 
 n370153 , n370154 , n370155 , n370156 , n370157 , n370158 , n49956 , n370160 , n49958 , n370162 , 
 n370163 , n49961 , n370165 , n370166 , n49964 , n370168 , n370169 , n49967 , n49968 , n370172 , 
 n370173 , n370174 , n370175 , n370176 , n49974 , n49975 , n370179 , n49977 , n370181 , n370182 , 
 n370183 , n370184 , n370185 , n49983 , n370187 , n370188 , n49986 , n49987 , n49988 , n370192 , 
 n49990 , n49991 , n49992 , n49993 , n370197 , n49995 , n370199 , n370200 , n370201 , n370202 , 
 n370203 , n50001 , n50002 , n370206 , n50004 , n370208 , n370209 , n370210 , n370211 , n370212 , 
 n370213 , n370214 , n50012 , n370216 , n370217 , n370218 , n370219 , n370220 , n370221 , n50019 , 
 n370223 , n370224 , n370225 , n50023 , n370227 , n370228 , n50026 , n370230 , n370231 , n370232 , 
 n50030 , n370234 , n370235 , n370236 , n370237 , n370238 , n50036 , n50037 , n50038 , n50039 , 
 n50040 , n50041 , n50042 , n370246 , n370247 , n370248 , n370249 , n50047 , n370251 , n370252 , 
 n370253 , n370254 , n370255 , n50053 , n370257 , n370258 , n50056 , n370260 , n370261 , n50059 , 
 n370263 , n370264 , n50062 , n370266 , n370267 , n50065 , n370269 , n370270 , n370271 , n370272 , 
 n370273 , n370274 , n370275 , n370276 , n370277 , n370278 , n370279 , n370280 , n370281 , n370282 , 
 n370283 , n50076 , n370285 , n370286 , n370287 , n370288 , n370289 , n370290 , n370291 , n50084 , 
 n370293 , n370294 , n50087 , n370296 , n370297 , n50090 , n370299 , n370300 , n50093 , n370302 , 
 n370303 , n370304 , n370305 , n370306 , n50099 , n370308 , n50101 , n370310 , n370311 , n50104 , 
 n370313 , n50106 , n370315 , n370316 , n50109 , n370318 , n370319 , n370320 , n370321 , n370322 , 
 n370323 , n50116 , n370325 , n370326 , n370327 , n50120 , n370329 , n370330 , n370331 , n370332 , 
 n370333 , n370334 , n50127 , n50128 , n370337 , n370338 , n370339 , n370340 , n370341 , n370342 , 
 n370343 , n370344 , n370345 , n370346 , n50139 , n370348 , n370349 , n370350 , n370351 , n370352 , 
 n50145 , n370354 , n50147 , n50148 , n50149 , n50150 , n50151 , n370360 , n370361 , n50154 , 
 n370363 , n370364 , n50157 , n370366 , n370367 , n50160 , n370369 , n370370 , n50163 , n370372 , 
 n370373 , n370374 , n370375 , n50168 , n50169 , n370378 , n50171 , n370380 , n370381 , n370382 , 
 n370383 , n50176 , n370385 , n370386 , n370387 , n370388 , n50181 , n370390 , n370391 , n50184 , 
 n370393 , n370394 , n370395 , n370396 , n370397 , n370398 , n370399 , n370400 , n370401 , n370402 , 
 n370403 , n370404 , n370405 , n50198 , n50199 , n370408 , n370409 , n50202 , n370411 , n370412 , 
 n50205 , n370414 , n370415 , n370416 , n50209 , n370418 , n50211 , n50212 , n370421 , n370422 , 
 n370423 , n50216 , n50217 , n370426 , n370427 , n50220 , n370429 , n370430 , n50223 , n50224 , 
 n370433 , n370434 , n50227 , n370436 , n370437 , n50230 , n370439 , n370440 , n50233 , n370442 , 
 n50235 , n370444 , n370445 , n370446 , n50239 , n50240 , n50241 , n370450 , n370451 , n370452 , 
 n50245 , n370454 , n370455 , n370456 , n370457 , n370458 , n370459 , n370460 , n50253 , n370462 , 
 n370463 , n50256 , n370465 , n370466 , n370467 , n50260 , n370469 , n370470 , n370471 , n370472 , 
 n370473 , n370474 , n50267 , n370476 , n370477 , n370478 , n370479 , n50272 , n370481 , n370482 , 
 n50275 , n370484 , n50277 , n370486 , n370487 , n50280 , n370489 , n50282 , n370491 , n370492 , 
 n50285 , n50286 , n370495 , n370496 , n370497 , n370498 , n370499 , n50292 , n370501 , n50294 , 
 n50295 , n370504 , n370505 , n370506 , n370507 , n370508 , n50301 , n370510 , n370511 , n370512 , 
 n50305 , n370514 , n370515 , n50308 , n370517 , n370518 , n50311 , n370520 , n50313 , n50314 , 
 n370523 , n50316 , n370525 , n370526 , n50319 , n370528 , n50321 , n50322 , n370531 , n370532 , 
 n370533 , n370534 , n50327 , n370536 , n370537 , n370538 , n370539 , n370540 , n370541 , n370542 , 
 n50335 , n370544 , n50337 , n370546 , n370547 , n370548 , n50341 , n370550 , n370551 , n370552 , 
 n370553 , n370554 , n370555 , n50348 , n370557 , n50350 , n50351 , n370560 , n370561 , n50354 , 
 n370563 , n370564 , n50357 , n370566 , n50359 , n370568 , n370569 , n50362 , n370571 , n370572 , 
 n370573 , n370574 , n50367 , n370576 , n50369 , n370578 , n50371 , n370580 , n370581 , n370582 , 
 n370583 , n370584 , n370585 , n370586 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , 
 n370593 , n370594 , n370595 , n370596 , n370597 , n50390 , n370599 , n50392 , n50393 , n50394 , 
 n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n370612 , 
 n370613 , n370614 , n370615 , n370616 , n370617 , n370618 , n370619 , n50412 , n370621 , n50414 , 
 n370623 , n370624 , n50417 , n370626 , n370627 , n370628 , n370629 , n370630 , n50423 , n370632 , 
 n370633 , n370634 , n370635 , n370636 , n370637 , n50430 , n370639 , n370640 , n370641 , n370642 , 
 n370643 , n370644 , n370645 , n370646 , n370647 , n50440 , n370649 , n370650 , n50443 , n370652 , 
 n370653 , n50446 , n370655 , n370656 , n370657 , n50450 , n370659 , n370660 , n370661 , n370662 , 
 n370663 , n370664 , n370665 , n370666 , n50459 , n370668 , n370669 , n50462 , n370671 , n370672 , 
 n370673 , n50466 , n50467 , n370676 , n50469 , n370678 , n370679 , n370680 , n50473 , n370682 , 
 n370683 , n50476 , n370685 , n370686 , n50479 , n370688 , n370689 , n370690 , n370691 , n50484 , 
 n50485 , n370694 , n370695 , n50488 , n370697 , n370698 , n50491 , n50492 , n370701 , n370702 , 
 n50495 , n370704 , n50497 , n50498 , n370707 , n370708 , n370709 , n370710 , n370711 , n50504 , 
 n370713 , n50506 , n50507 , n370716 , n50509 , n370718 , n50511 , n50512 , n50513 , n50514 , 
 n370723 , n370724 , n370725 , n370726 , n370727 , n370728 , n370729 , n370730 , n370731 , n370732 , 
 n370733 , n50526 , n370735 , n370736 , n370737 , n370738 , n370739 , n50532 , n50533 , n370742 , 
 n50535 , n50536 , n370745 , n50538 , n370747 , n370748 , n370749 , n370750 , n370751 , n50544 , 
 n370753 , n370754 , n370755 , n370756 , n370757 , n370758 , n370759 , n50552 , n370761 , n370762 , 
 n50555 , n370764 , n370765 , n50558 , n370767 , n370768 , n50561 , n370770 , n50563 , n370772 , 
 n370773 , n370774 , n370775 , n50568 , n370777 , n50570 , n50571 , n370780 , n370781 , n370782 , 
 n370783 , n370784 , n50577 , n50578 , n370787 , n50580 , n370789 , n370790 , n370791 , n370792 , 
 n370793 , n370794 , n370795 , n370796 , n370797 , n50590 , n370799 , n370800 , n50593 , n370802 , 
 n50595 , n50596 , n370805 , n370806 , n370807 , n370808 , n370809 , n370810 , n370811 , n50604 , 
 n370813 , n370814 , n50607 , n370816 , n50609 , n370818 , n370819 , n370820 , n370821 , n370822 , 
 n50615 , n370824 , n370825 , n370826 , n370827 , n370828 , n50621 , n50622 , n370831 , n370832 , 
 n370833 , n370834 , n370835 , n370836 , n50629 , n370838 , n370839 , n50632 , n370841 , n370842 , 
 n370843 , n370844 , n370845 , n370846 , n370847 , n370848 , n370849 , n370850 , n50643 , n50644 , 
 n50645 , n370854 , n370855 , n370856 , n370857 , n370858 , n370859 , n370860 , n50653 , n370862 , 
 n370863 , n50656 , n370865 , n370866 , n50659 , n370868 , n370869 , n370870 , n370871 , n370872 , 
 n370873 , n370874 , n370875 , n370876 , n370877 , n50670 , n370879 , n370880 , n50673 , n370882 , 
 n370883 , n370884 , n370885 , n370886 , n370887 , n370888 , n370889 , n50682 , n370891 , n370892 , 
 n50685 , n370894 , n370895 , n50688 , n370897 , n370898 , n370899 , n370900 , n50693 , n370902 , 
 n370903 , n370904 , n370905 , n370906 , n50699 , n370908 , n370909 , n370910 , n50703 , n370912 , 
 n370913 , n50706 , n370915 , n370916 , n370917 , n370918 , n50711 , n370920 , n370921 , n50714 , 
 n370923 , n370924 , n370925 , n370926 , n370927 , n370928 , n370929 , n50722 , n50723 , n370932 , 
 n50725 , n370934 , n370935 , n370936 , n370937 , n50730 , n370939 , n370940 , n50733 , n370942 , 
 n370943 , n50736 , n370945 , n370946 , n370947 , n370948 , n370949 , n370950 , n50743 , n50744 , 
 n50745 , n50746 , n370955 , n370956 , n370957 , n370958 , n370959 , n50752 , n370961 , n370962 , 
 n50755 , n370964 , n370965 , n50758 , n370967 , n370968 , n50761 , n50762 , n370971 , n50764 , 
 n370973 , n50766 , n50767 , n370976 , n370977 , n370978 , n370979 , n370980 , n370981 , n370982 , 
 n50775 , n370984 , n50777 , n370986 , n50779 , n50780 , n370989 , n50782 , n370991 , n370992 , 
 n370993 , n370994 , n370995 , n370996 , n50789 , n370998 , n370999 , n50792 , n371001 , n371002 , 
 n371003 , n371004 , n371005 , n371006 , n371007 , n371008 , n371009 , n50802 , n371011 , n50804 , 
 n371013 , n371014 , n50807 , n371016 , n371017 , n50810 , n371019 , n50812 , n50813 , n371022 , 
 n371023 , n371024 , n50817 , n371026 , n371027 , n371028 , n371029 , n371030 , n50823 , n371032 , 
 n371033 , n50826 , n50827 , n371036 , n371037 , n50830 , n371039 , n371040 , n50833 , n371042 , 
 n50835 , n371044 , n50837 , n50838 , n371047 , n50840 , n371049 , n50842 , n371051 , n371052 , 
 n50845 , n371054 , n50847 , n371056 , n371057 , n50850 , n371059 , n371060 , n371061 , n50854 , 
 n371063 , n371064 , n371065 , n371066 , n371067 , n371068 , n50861 , n371070 , n371071 , n371072 , 
 n50865 , n371074 , n50867 , n371076 , n50869 , n50870 , n50871 , n371080 , n371081 , n371082 , 
 n371083 , n50876 , n371085 , n371086 , n371087 , n371088 , n371089 , n50882 , n371091 , n371092 , 
 n371093 , n50886 , n371095 , n371096 , n50889 , n371098 , n371099 , n371100 , n371101 , n371102 , 
 n371103 , n371104 , n50897 , n50898 , n371107 , n50900 , n371109 , n371110 , n50903 , n50904 , 
 n371113 , n371114 , n371115 , n371116 , n371117 , n371118 , n371119 , n50912 , n371121 , n50914 , 
 n50915 , n371124 , n50917 , n371126 , n371127 , n371128 , n50921 , n50922 , n371131 , n50924 , 
 n371133 , n371134 , n50927 , n50928 , n371137 , n371138 , n371139 , n371140 , n371141 , n50934 , 
 n371143 , n371144 , n371145 , n371146 , n371147 , n371148 , n50941 , n371150 , n371151 , n371152 , 
 n371153 , n371154 , n371155 , n50948 , n371157 , n371158 , n371159 , n371160 , n50953 , n371162 , 
 n371163 , n50956 , n50957 , n371166 , n50959 , n371168 , n371169 , n50962 , n371171 , n371172 , 
 n371173 , n371174 , n371175 , n371176 , n50969 , n371178 , n371179 , n371180 , n371181 , n371182 , 
 n371183 , n371184 , n371185 , n371186 , n371187 , n371188 , n50981 , n50982 , n371191 , n50984 , 
 n50985 , n371194 , n50987 , n371196 , n371197 , n371198 , n50991 , n371200 , n371201 , n50994 , 
 n371203 , n371204 , n371205 , n371206 , n371207 , n371208 , n371209 , n371210 , n371211 , n371212 , 
 n371213 , n371214 , n371215 , n51008 , n371217 , n371218 , n371219 , n371220 , n371221 , n371222 , 
 n371223 , n371224 , n371225 , n371226 , n371227 , n371228 , n371229 , n371230 , n371231 , n371232 , 
 n371233 , n371234 , n51022 , n371236 , n371237 , n51025 , n371239 , n51027 , n371241 , n371242 , 
 n371243 , n371244 , n51032 , n371246 , n371247 , n371248 , n371249 , n371250 , n371251 , n371252 , 
 n51040 , n371254 , n371255 , n51043 , n371257 , n371258 , n371259 , n51047 , n371261 , n371262 , 
 n51050 , n371264 , n51052 , n51053 , n51054 , n371268 , n51056 , n371270 , n371271 , n371272 , 
 n371273 , n51061 , n371275 , n371276 , n371277 , n371278 , n371279 , n371280 , n371281 , n51069 , 
 n371283 , n371284 , n371285 , n371286 , n51074 , n51075 , n51076 , n51077 , n371291 , n371292 , 
 n371293 , n371294 , n371295 , n51083 , n371297 , n371298 , n371299 , n371300 , n371301 , n371302 , 
 n371303 , n51091 , n371305 , n371306 , n371307 , n371308 , n371309 , n371310 , n51098 , n371312 , 
 n51100 , n51101 , n371315 , n51103 , n371317 , n51105 , n371319 , n51107 , n371321 , n371322 , 
 n371323 , n371324 , n51112 , n371326 , n51114 , n371328 , n51116 , n371330 , n371331 , n371332 , 
 n51120 , n371334 , n371335 , n371336 , n371337 , n51125 , n371339 , n371340 , n51128 , n371342 , 
 n371343 , n51131 , n371345 , n51133 , n371347 , n51135 , n51136 , n371350 , n371351 , n371352 , 
 n371353 , n371354 , n371355 , n371356 , n371357 , n51145 , n371359 , n371360 , n371361 , n371362 , 
 n51150 , n371364 , n371365 , n51153 , n51154 , n371368 , n51156 , n371370 , n51158 , n371372 , 
 n371373 , n371374 , n371375 , n371376 , n371377 , n371378 , n51166 , n371380 , n371381 , n371382 , 
 n371383 , n371384 , n371385 , n51173 , n371387 , n371388 , n371389 , n371390 , n51178 , n51179 , 
 n51180 , n51181 , n371395 , n371396 , n371397 , n371398 , n371399 , n371400 , n371401 , n371402 , 
 n51190 , n371404 , n371405 , n371406 , n51194 , n51195 , n371409 , n371410 , n371411 , n371412 , 
 n371413 , n371414 , n51202 , n371416 , n51204 , n51205 , n51206 , n51207 , n371421 , n51209 , 
 n51210 , n51211 , n51212 , n51213 , n51214 , n371428 , n371429 , n371430 , n371431 , n51219 , 
 n371433 , n371434 , n371435 , n371436 , n371437 , n371438 , n51226 , n51227 , n371441 , n371442 , 
 n51230 , n51231 , n371445 , n371446 , n371447 , n371448 , n371449 , n371450 , n51238 , n371452 , 
 n371453 , n51241 , n371455 , n371456 , n51244 , n371458 , n371459 , n51247 , n371461 , n371462 , 
 n51250 , n371464 , n371465 , n371466 , n371467 , n371468 , n371469 , n371470 , n371471 , n371472 , 
 n371473 , n371474 , n371475 , n371476 , n371477 , n371478 , n51266 , n51267 , n371481 , n371482 , 
 n51270 , n371484 , n51272 , n371486 , n371487 , n371488 , n51276 , n371490 , n371491 , n371492 , 
 n371493 , n51281 , n371495 , n371496 , n51284 , n371498 , n371499 , n371500 , n371501 , n371502 , 
 n51290 , n371504 , n371505 , n371506 , n51294 , n371508 , n371509 , n51297 , n371511 , n371512 , 
 n371513 , n371514 , n371515 , n371516 , n371517 , n371518 , n371519 , n371520 , n51308 , n371522 , 
 n51310 , n51311 , n371525 , n371526 , n51314 , n371528 , n51316 , n371530 , n371531 , n371532 , 
 n51320 , n51321 , n51322 , n371536 , n371537 , n371538 , n371539 , n51327 , n371541 , n371542 , 
 n371543 , n371544 , n371545 , n51333 , n371547 , n371548 , n371549 , n51337 , n51338 , n371552 , 
 n371553 , n371554 , n371555 , n371556 , n51344 , n371558 , n371559 , n371560 , n371561 , n371562 , 
 n371563 , n371564 , n51352 , n51353 , n51354 , n371568 , n371569 , n371570 , n371571 , n371572 , 
 n51360 , n51361 , n371575 , n51363 , n371577 , n371578 , n51366 , n371580 , n371581 , n51369 , 
 n371583 , n371584 , n371585 , n371586 , n371587 , n371588 , n51376 , n371590 , n371591 , n371592 , 
 n371593 , n371594 , n371595 , n371596 , n371597 , n371598 , n51386 , n371600 , n51388 , n51389 , 
 n371603 , n51391 , n371605 , n51393 , n371607 , n371608 , n371609 , n371610 , n371611 , n371612 , 
 n371613 , n371614 , n371615 , n371616 , n371617 , n371618 , n371619 , n51407 , n371621 , n371622 , 
 n51410 , n371624 , n371625 , n371626 , n371627 , n371628 , n371629 , n51417 , n371631 , n371632 , 
 n371633 , n371634 , n371635 , n371636 , n51424 , n371638 , n371639 , n371640 , n371641 , n371642 , 
 n371643 , n371644 , n51432 , n371646 , n371647 , n371648 , n371649 , n371650 , n371651 , n51439 , 
 n371653 , n371654 , n51442 , n371656 , n371657 , n51445 , n51446 , n371660 , n51448 , n371662 , 
 n371663 , n371664 , n371665 , n51453 , n371667 , n371668 , n371669 , n371670 , n51458 , n51459 , 
 n371673 , n371674 , n371675 , n371676 , n371677 , n371678 , n371679 , n371680 , n371681 , n371682 , 
 n371683 , n371684 , n371685 , n371686 , n371687 , n371688 , n371689 , n371690 , n371691 , n371692 , 
 n371693 , n371694 , n371695 , n371696 , n371697 , n371698 , n371699 , n371700 , n51468 , n371702 , 
 n371703 , n371704 , n371705 , n371706 , n371707 , n51471 , n371709 , n371710 , n51474 , n51475 , 
 n371713 , n51477 , n51478 , n371716 , n51480 , n371718 , n51482 , n51483 , n371721 , n51485 , 
 n371723 , n51487 , n371725 , n371726 , n371727 , n371728 , n371729 , n371730 , n371731 , n371732 , 
 n371733 , n371734 , n371735 , n371736 , n51500 , n371738 , n371739 , n371740 , n371741 , n371742 , 
 n371743 , n51507 , n371745 , n371746 , n51510 , n371748 , n51512 , n51513 , n371751 , n51515 , 
 n371753 , n371754 , n371755 , n371756 , n371757 , n371758 , n371759 , n371760 , n51524 , n371762 , 
 n371763 , n371764 , n371765 , n51529 , n371767 , n371768 , n51532 , n51533 , n371771 , n51535 , 
 n371773 , n371774 , n51538 , n371776 , n51540 , n51541 , n51542 , n51543 , n371781 , n371782 , 
 n371783 , n371784 , n371785 , n51549 , n51550 , n371788 , n51552 , n371790 , n51554 , n371792 , 
 n371793 , n371794 , n51558 , n371796 , n371797 , n371798 , n371799 , n371800 , n371801 , n371802 , 
 n371803 , n371804 , n51568 , n371806 , n371807 , n51571 , n371809 , n371810 , n371811 , n371812 , 
 n371813 , n371814 , n371815 , n371816 , n371817 , n371818 , n51582 , n371820 , n371821 , n371822 , 
 n371823 , n371824 , n371825 , n51589 , n371827 , n371828 , n371829 , n51593 , n371831 , n51595 , 
 n51596 , n371834 , n371835 , n51599 , n51600 , n371838 , n371839 , n371840 , n371841 , n371842 , 
 n51606 , n371844 , n51608 , n371846 , n371847 , n371848 , n371849 , n371850 , n371851 , n371852 , 
 n371853 , n371854 , n51618 , n371856 , n371857 , n51621 , n371859 , n371860 , n51624 , n371862 , 
 n371863 , n51627 , n371865 , n371866 , n51630 , n371868 , n371869 , n51633 , n371871 , n371872 , 
 n371873 , n51637 , n371875 , n371876 , n371877 , n371878 , n371879 , n51643 , n371881 , n51645 , 
 n371883 , n51647 , n371885 , n371886 , n371887 , n371888 , n371889 , n371890 , n371891 , n371892 , 
 n371893 , n371894 , n371895 , n51659 , n371897 , n51661 , n51662 , n51663 , n51664 , n371902 , 
 n51666 , n371904 , n51668 , n371906 , n371907 , n51671 , n371909 , n371910 , n51674 , n371912 , 
 n371913 , n51677 , n371915 , n371916 , n51680 , n371918 , n371919 , n371920 , n51684 , n51685 , 
 n371923 , n51687 , n371925 , n371926 , n371927 , n371928 , n371929 , n371930 , n371931 , n51695 , 
 n371933 , n51697 , n51698 , n51699 , n51700 , n371938 , n51702 , n51703 , n371941 , n51705 , 
 n371943 , n371944 , n371945 , n51709 , n371947 , n371948 , n371949 , n371950 , n371951 , n371952 , 
 n371953 , n51717 , n371955 , n51719 , n371957 , n371958 , n51722 , n371960 , n371961 , n51725 , 
 n371963 , n371964 , n51728 , n371966 , n371967 , n371968 , n51732 , n371970 , n371971 , n51735 , 
 n371973 , n371974 , n51738 , n371976 , n371977 , n371978 , n371979 , n51743 , n371981 , n51745 , 
 n371983 , n51747 , n51748 , n371986 , n371987 , n371988 , n371989 , n51753 , n371991 , n371992 , 
 n371993 , n51757 , n371995 , n51759 , n371997 , n371998 , n371999 , n372000 , n372001 , n372002 , 
 n372003 , n372004 , n51768 , n372006 , n372007 , n372008 , n372009 , n51773 , n51774 , n51775 , 
 n372013 , n51777 , n372015 , n372016 , n51780 , n372018 , n372019 , n372020 , n372021 , n372022 , 
 n51786 , n372024 , n372025 , n51789 , n372027 , n372028 , n372029 , n372030 , n372031 , n51795 , 
 n372033 , n372034 , n372035 , n51799 , n372037 , n372038 , n372039 , n372040 , n372041 , n372042 , 
 n372043 , n372044 , n51808 , n372046 , n372047 , n51811 , n372049 , n372050 , n51814 , n51815 , 
 n372053 , n51817 , n372055 , n372056 , n372057 , n372058 , n51822 , n372060 , n372061 , n372062 , 
 n51826 , n51827 , n372065 , n372066 , n372067 , n372068 , n372069 , n372070 , n372071 , n372072 , 
 n51836 , n372074 , n51838 , n51839 , n372077 , n372078 , n51842 , n372080 , n51844 , n372082 , 
 n372083 , n372084 , n372085 , n372086 , n372087 , n372088 , n372089 , n51853 , n51854 , n372092 , 
 n372093 , n51857 , n372095 , n51859 , n372097 , n51861 , n372099 , n372100 , n372101 , n372102 , 
 n372103 , n372104 , n372105 , n372106 , n372107 , n372108 , n372109 , n372110 , n372111 , n51875 , 
 n372113 , n372114 , n51878 , n372116 , n51880 , n51881 , n372119 , n372120 , n372121 , n372122 , 
 n372123 , n372124 , n372125 , n51889 , n372127 , n372128 , n51892 , n372130 , n372131 , n372132 , 
 n372133 , n372134 , n372135 , n51899 , n51900 , n51901 , n372139 , n372140 , n51904 , n372142 , 
 n372143 , n372144 , n372145 , n372146 , n372147 , n51911 , n372149 , n51913 , n51914 , n372152 , 
 n372153 , n51917 , n372155 , n51919 , n372157 , n372158 , n51922 , n372160 , n51924 , n51925 , 
 n372163 , n372164 , n372165 , n372166 , n372167 , n372168 , n372169 , n372170 , n372171 , n372172 , 
 n51936 , n372174 , n372175 , n372176 , n372177 , n372178 , n372179 , n51943 , n372181 , n372182 , 
 n51946 , n372184 , n51948 , n51949 , n372187 , n372188 , n51952 , n51953 , n51954 , n51955 , 
 n51956 , n372194 , n372195 , n372196 , n372197 , n372198 , n372199 , n51963 , n372201 , n372202 , 
 n51966 , n372204 , n372205 , n51969 , n372207 , n372208 , n51972 , n372210 , n372211 , n51975 , 
 n372213 , n372214 , n372215 , n372216 , n51980 , n372218 , n372219 , n372220 , n51984 , n51985 , 
 n51986 , n372224 , n51988 , n372226 , n372227 , n372228 , n51992 , n372230 , n372231 , n51995 , 
 n51996 , n372234 , n51998 , n51999 , n372237 , n372238 , n52002 , n372240 , n372241 , n372242 , 
 n372243 , n372244 , n52008 , n372246 , n372247 , n372248 , n372249 , n372250 , n372251 , n372252 , 
 n372253 , n372254 , n372255 , n372256 , n372257 , n372258 , n52022 , n372260 , n372261 , n52025 , 
 n372263 , n52027 , n52028 , n52029 , n372267 , n372268 , n52032 , n372270 , n372271 , n52035 , 
 n372273 , n52037 , n372275 , n372276 , n372277 , n372278 , n52042 , n372280 , n372281 , n52045 , 
 n372283 , n52047 , n372285 , n372286 , n372287 , n372288 , n372289 , n372290 , n372291 , n372292 , 
 n372293 , n372294 , n372295 , n372296 , n372297 , n372298 , n372299 , n372300 , n372301 , n52065 , 
 n372303 , n372304 , n52068 , n372306 , n372307 , n52071 , n372309 , n372310 , n52074 , n372312 , 
 n52076 , n372314 , n372315 , n372316 , n372317 , n52081 , n372319 , n372320 , n52084 , n372322 , 
 n372323 , n52087 , n372325 , n372326 , n52090 , n52091 , n372329 , n372330 , n52094 , n372332 , 
 n372333 , n52097 , n372335 , n372336 , n52100 , n372338 , n372339 , n372340 , n372341 , n372342 , 
 n372343 , n372344 , n372345 , n372346 , n372347 , n372348 , n372349 , n372350 , n52108 , n372352 , 
 n52110 , n372354 , n52112 , n372356 , n372357 , n52115 , n372359 , n372360 , n52118 , n52119 , 
 n372363 , n372364 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n372371 , n372372 , 
 n372373 , n372374 , n372375 , n372376 , n372377 , n52135 , n372379 , n372380 , n52138 , n372382 , 
 n52140 , n52141 , n52142 , n372386 , n372387 , n52145 , n372389 , n372390 , n372391 , n372392 , 
 n372393 , n372394 , n372395 , n372396 , n52154 , n372398 , n372399 , n52157 , n372401 , n372402 , 
 n372403 , n372404 , n372405 , n52163 , n372407 , n372408 , n52166 , n372410 , n372411 , n372412 , 
 n372413 , n372414 , n372415 , n372416 , n372417 , n372418 , n372419 , n372420 , n372421 , n372422 , 
 n372423 , n372424 , n372425 , n372426 , n52184 , n372428 , n52186 , n372430 , n372431 , n52189 , 
 n372433 , n372434 , n52192 , n372436 , n372437 , n52195 , n372439 , n372440 , n52198 , n52199 , 
 n372443 , n372444 , n52202 , n372446 , n372447 , n52205 , n52206 , n52207 , n372451 , n372452 , 
 n372453 , n372454 , n52212 , n372456 , n52214 , n372458 , n372459 , n372460 , n52218 , n372462 , 
 n372463 , n52221 , n372465 , n372466 , n372467 , n372468 , n372469 , n372470 , n372471 , n372472 , 
 n372473 , n372474 , n372475 , n372476 , n372477 , n372478 , n372479 , n372480 , n52238 , n52239 , 
 n52240 , n52241 , n372485 , n52243 , n372487 , n52245 , n372489 , n372490 , n372491 , n52249 , 
 n372493 , n372494 , n52252 , n372496 , n372497 , n372498 , n52256 , n52257 , n52258 , n372502 , 
 n372503 , n372504 , n372505 , n372506 , n372507 , n372508 , n372509 , n372510 , n372511 , n372512 , 
 n52270 , n372514 , n372515 , n52273 , n52274 , n372518 , n372519 , n52277 , n372521 , n372522 , 
 n372523 , n372524 , n52282 , n52283 , n52284 , n372528 , n372529 , n52287 , n52288 , n372532 , 
 n52290 , n372534 , n372535 , n372536 , n372537 , n372538 , n372539 , n372540 , n372541 , n52299 , 
 n372543 , n372544 , n372545 , n52303 , n372547 , n372548 , n52306 , n372550 , n52308 , n52309 , 
 n52310 , n52311 , n372555 , n372556 , n372557 , n372558 , n372559 , n372560 , n372561 , n372562 , 
 n52320 , n52321 , n372565 , n372566 , n52324 , n372568 , n372569 , n52327 , n372571 , n372572 , 
 n372573 , n52331 , n372575 , n372576 , n372577 , n372578 , n372579 , n372580 , n372581 , n372582 , 
 n372583 , n372584 , n372585 , n372586 , n52344 , n372588 , n372589 , n372590 , n372591 , n52349 , 
 n372593 , n372594 , n52352 , n52353 , n372597 , n372598 , n372599 , n372600 , n52358 , n372602 , 
 n372603 , n52361 , n372605 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , 
 n372613 , n372614 , n372615 , n372616 , n372617 , n372618 , n372619 , n372620 , n372621 , n372622 , 
 n372623 , n372624 , n372625 , n372626 , n372627 , n372628 , n52386 , n372630 , n372631 , n372632 , 
 n52390 , n372634 , n372635 , n372636 , n372637 , n372638 , n372639 , n372640 , n372641 , n372642 , 
 n52400 , n52401 , n372645 , n52403 , n372647 , n52405 , n52406 , n372650 , n372651 , n52409 , 
 n372653 , n372654 , n52412 , n372656 , n372657 , n372658 , n372659 , n372660 , n372661 , n52419 , 
 n372663 , n372664 , n52422 , n52423 , n52424 , n52425 , n52426 , n372670 , n372671 , n372672 , 
 n372673 , n372674 , n372675 , n52433 , n372677 , n372678 , n372679 , n52437 , n52438 , n372682 , 
 n52440 , n52441 , n372685 , n372686 , n372687 , n372688 , n372689 , n372690 , n372691 , n372692 , 
 n372693 , n372694 , n372695 , n372696 , n52454 , n372698 , n52456 , n372700 , n52458 , n372702 , 
 n372703 , n52461 , n372705 , n372706 , n52464 , n372708 , n52466 , n52467 , n372711 , n372712 , 
 n372713 , n372714 , n372715 , n52473 , n372717 , n372718 , n52476 , n372720 , n372721 , n372722 , 
 n372723 , n372724 , n372725 , n372726 , n372727 , n372728 , n372729 , n372730 , n52488 , n372732 , 
 n372733 , n372734 , n372735 , n372736 , n372737 , n372738 , n52496 , n372740 , n372741 , n372742 , 
 n372743 , n372744 , n52502 , n372746 , n52504 , n372748 , n372749 , n372750 , n372751 , n372752 , 
 n52510 , n372754 , n372755 , n372756 , n372757 , n372758 , n372759 , n372760 , n372761 , n372762 , 
 n372763 , n372764 , n372765 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , 
 n52530 , n52531 , n52532 , n52533 , n52534 , n372778 , n52536 , n372780 , n372781 , n52539 , 
 n372783 , n372784 , n372785 , n372786 , n372787 , n372788 , n372789 , n372790 , n52548 , n372792 , 
 n372793 , n372794 , n372795 , n372796 , n372797 , n52555 , n372799 , n52557 , n372801 , n372802 , 
 n372803 , n372804 , n52562 , n372806 , n372807 , n372808 , n52566 , n372810 , n372811 , n372812 , 
 n372813 , n372814 , n372815 , n372816 , n372817 , n372818 , n372819 , n52577 , n372821 , n372822 , 
 n52580 , n372824 , n372825 , n52583 , n372827 , n372828 , n52586 , n372830 , n372831 , n372832 , 
 n372833 , n52591 , n372835 , n372836 , n52594 , n372838 , n372839 , n52597 , n52598 , n372842 , 
 n372843 , n372844 , n372845 , n372846 , n372847 , n372848 , n52606 , n372850 , n372851 , n372852 , 
 n372853 , n372854 , n372855 , n372856 , n52614 , n372858 , n52616 , n52617 , n372861 , n372862 , 
 n372863 , n372864 , n372865 , n372866 , n372867 , n372868 , n372869 , n52627 , n372871 , n52629 , 
 n372873 , n52631 , n372875 , n52633 , n372877 , n52635 , n372879 , n372880 , n52638 , n372882 , 
 n372883 , n372884 , n372885 , n52643 , n372887 , n52645 , n372889 , n52647 , n372891 , n52649 , 
 n52650 , n372894 , n372895 , n372896 , n372897 , n372898 , n52656 , n52657 , n372901 , n52659 , 
 n372903 , n372904 , n52662 , n372906 , n52664 , n372908 , n372909 , n372910 , n372911 , n372912 , 
 n372913 , n372914 , n372915 , n372916 , n52674 , n52675 , n52676 , n372920 , n372921 , n372922 , 
 n372923 , n372924 , n372925 , n372926 , n52684 , n372928 , n372929 , n372930 , n372931 , n372932 , 
 n52690 , n52691 , n372935 , n372936 , n372937 , n372938 , n372939 , n372940 , n372941 , n372942 , 
 n52700 , n372944 , n372945 , n372946 , n372947 , n372948 , n52706 , n372950 , n372951 , n372952 , 
 n372953 , n372954 , n372955 , n372956 , n372957 , n372958 , n372959 , n52717 , n372961 , n52719 , 
 n372963 , n52721 , n52722 , n52723 , n372967 , n52725 , n372969 , n372970 , n372971 , n372972 , 
 n372973 , n372974 , n372975 , n372976 , n52734 , n52735 , n372979 , n52737 , n372981 , n372982 , 
 n52740 , n52741 , n372985 , n372986 , n372987 , n52745 , n372989 , n372990 , n52748 , n372992 , 
 n372993 , n372994 , n372995 , n52753 , n52754 , n372998 , n372999 , n373000 , n373001 , n373002 , 
 n373003 , n373004 , n373005 , n52763 , n373007 , n373008 , n52766 , n373010 , n373011 , n373012 , 
 n373013 , n373014 , n373015 , n373016 , n52774 , n373018 , n52776 , n373020 , n52778 , n52779 , 
 n373023 , n373024 , n373025 , n373026 , n52784 , n52785 , n373029 , n373030 , n52788 , n373032 , 
 n373033 , n52791 , n373035 , n373036 , n52794 , n52795 , n373039 , n373040 , n373041 , n373042 , 
 n373043 , n373044 , n373045 , n52798 , n373047 , n373048 , n52801 , n373050 , n373051 , n373052 , 
 n373053 , n373054 , n52807 , n373056 , n373057 , n52810 , n52811 , n373060 , n52813 , n373062 , 
 n373063 , n52816 , n373065 , n52818 , n52819 , n373068 , n373069 , n373070 , n373071 , n373072 , 
 n52825 , n373074 , n373075 , n52828 , n373077 , n52830 , n373079 , n373080 , n373081 , n373082 , 
 n373083 , n373084 , n373085 , n52838 , n373087 , n373088 , n52841 , n52842 , n373091 , n373092 , 
 n373093 , n373094 , n373095 , n373096 , n52849 , n373098 , n52851 , n373100 , n373101 , n52854 , 
 n373103 , n52856 , n373105 , n52858 , n52859 , n52860 , n373109 , n373110 , n373111 , n52864 , 
 n373113 , n373114 , n52867 , n52868 , n373117 , n52870 , n373119 , n373120 , n373121 , n373122 , 
 n373123 , n373124 , n52877 , n52878 , n373127 , n52880 , n52881 , n373130 , n52883 , n52884 , 
 n373133 , n52886 , n373135 , n52888 , n373137 , n373138 , n52891 , n373140 , n373141 , n52894 , 
 n373143 , n373144 , n52897 , n373146 , n52899 , n373148 , n52901 , n373150 , n373151 , n373152 , 
 n373153 , n373154 , n373155 , n373156 , n373157 , n52910 , n373159 , n373160 , n373161 , n373162 , 
 n373163 , n373164 , n52917 , n373166 , n373167 , n373168 , n373169 , n373170 , n373171 , n52924 , 
 n373173 , n373174 , n373175 , n52928 , n373177 , n373178 , n373179 , n373180 , n373181 , n373182 , 
 n373183 , n373184 , n373185 , n52938 , n373187 , n52940 , n373189 , n52942 , n373191 , n52944 , 
 n373193 , n52946 , n373195 , n373196 , n373197 , n373198 , n373199 , n52952 , n52953 , n373202 , 
 n373203 , n373204 , n373205 , n373206 , n373207 , n373208 , n373209 , n52962 , n373211 , n373212 , 
 n52965 , n52966 , n373215 , n52968 , n52969 , n373218 , n373219 , n373220 , n373221 , n373222 , 
 n52975 , n373224 , n52977 , n373226 , n373227 , n373228 , n52981 , n373230 , n373231 , n373232 , 
 n373233 , n52986 , n373235 , n373236 , n373237 , n373238 , n52991 , n373240 , n373241 , n373242 , 
 n373243 , n52996 , n373245 , n373246 , n52999 , n373248 , n373249 , n53002 , n373251 , n373252 , 
 n53005 , n373254 , n373255 , n53008 , n53009 , n373258 , n373259 , n373260 , n373261 , n373262 , 
 n53015 , n373264 , n373265 , n373266 , n53019 , n373268 , n373269 , n373270 , n373271 , n53024 , 
 n373273 , n373274 , n373275 , n373276 , n373277 , n373278 , n53031 , n373280 , n53033 , n373282 , 
 n53035 , n373284 , n53037 , n373286 , n373287 , n53040 , n53041 , n373290 , n53043 , n373292 , 
 n373293 , n53046 , n373295 , n373296 , n53049 , n373298 , n373299 , n53052 , n53053 , n53054 , 
 n373303 , n373304 , n53057 , n53058 , n53059 , n373308 , n373309 , n53062 , n373311 , n53064 , 
 n373313 , n373314 , n373315 , n373316 , n373317 , n53070 , n373319 , n53072 , n373321 , n373322 , 
 n373323 , n373324 , n373325 , n373326 , n373327 , n373328 , n373329 , n373330 , n373331 , n373332 , 
 n373333 , n373334 , n53087 , n373336 , n373337 , n53090 , n373339 , n373340 , n53093 , n373342 , 
 n373343 , n373344 , n373345 , n53098 , n373347 , n53100 , n373349 , n53102 , n373351 , n373352 , 
 n373353 , n373354 , n373355 , n373356 , n53109 , n53110 , n373359 , n53112 , n373361 , n53114 , 
 n373363 , n373364 , n53117 , n373366 , n373367 , n53120 , n373369 , n373370 , n53123 , n373372 , 
 n373373 , n373374 , n53127 , n53128 , n53129 , n53130 , n373379 , n53132 , n373381 , n373382 , 
 n373383 , n53136 , n373385 , n373386 , n373387 , n53140 , n373389 , n373390 , n53143 , n373392 , 
 n373393 , n373394 , n373395 , n373396 , n373397 , n373398 , n373399 , n373400 , n373401 , n373402 , 
 n373403 , n53156 , n373405 , n373406 , n373407 , n373408 , n373409 , n373410 , n373411 , n373412 , 
 n373413 , n373414 , n373415 , n373416 , n373417 , n373418 , n373419 , n373420 , n373421 , n373422 , 
 n373423 , n373424 , n373425 , n373426 , n373427 , n373428 , n373429 , n373430 , n373431 , n373432 , 
 n373433 , n373434 , n373435 , n373436 , n373437 , n373438 , n373439 , n373440 , n373441 , n373442 , 
 n373443 , n373444 , n373445 , n373446 , n373447 , n373448 , n373449 , n373450 , n373451 , n373452 , 
 n373453 , n373454 , n373455 , n373456 , n373457 , n373458 , n373459 , n373460 , n373461 , n373462 , 
 n373463 , n373464 , n373465 , n373466 , n373467 , n373468 , n373469 , n373470 , n373471 , n373472 , 
 n373473 , n373474 , n373475 , n373476 , n373477 , n373478 , n373479 , n373480 , n373481 , n373482 , 
 n373483 , n373484 , n53161 , n373486 , n373487 , n373488 , n53162 , n373490 , n373491 , n53165 , 
 n373493 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n373501 , n373502 , 
 n373503 , n373504 , n53178 , n373506 , n373507 , n53181 , n373509 , n373510 , n373511 , n373512 , 
 n373513 , n373514 , n373515 , n373516 , n53190 , n373518 , n373519 , n373520 , n373521 , n53195 , 
 n53196 , n53197 , n53198 , n373526 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , 
 n373533 , n53207 , n373535 , n53209 , n373537 , n53211 , n373539 , n53213 , n373541 , n373542 , 
 n373543 , n373544 , n373545 , n373546 , n373547 , n373548 , n53222 , n373550 , n373551 , n373552 , 
 n373553 , n373554 , n373555 , n373556 , n373557 , n373558 , n373559 , n373560 , n373561 , n53235 , 
 n373563 , n373564 , n53238 , n373566 , n373567 , n53241 , n373569 , n373570 , n53244 , n373572 , 
 n373573 , n53247 , n373575 , n53249 , n53250 , n373578 , n373579 , n53253 , n373581 , n373582 , 
 n373583 , n373584 , n373585 , n373586 , n53260 , n373588 , n373589 , n373590 , n53264 , n373592 , 
 n373593 , n373594 , n373595 , n53269 , n53270 , n373598 , n53272 , n373600 , n53274 , n373602 , 
 n373603 , n373604 , n373605 , n373606 , n373607 , n373608 , n53282 , n373610 , n373611 , n53285 , 
 n373613 , n373614 , n53288 , n373616 , n373617 , n373618 , n373619 , n373620 , n373621 , n373622 , 
 n373623 , n373624 , n373625 , n373626 , n373627 , n373628 , n373629 , n53303 , n53304 , n373632 , 
 n373633 , n373634 , n373635 , n373636 , n53310 , n373638 , n373639 , n53313 , n53314 , n373642 , 
 n373643 , n53317 , n373645 , n373646 , n53320 , n373648 , n53322 , n53323 , n373651 , n373652 , 
 n373653 , n53327 , n373655 , n373656 , n373657 , n53331 , n373659 , n53333 , n373661 , n373662 , 
 n53336 , n373664 , n373665 , n53339 , n373667 , n373668 , n53342 , n373670 , n373671 , n373672 , 
 n53346 , n373674 , n373675 , n53349 , n373677 , n53351 , n373679 , n373680 , n53354 , n373682 , 
 n53356 , n53357 , n373685 , n373686 , n53360 , n53361 , n53362 , n53363 , n373691 , n373692 , 
 n53366 , n373694 , n373695 , n373696 , n373697 , n53371 , n53372 , n373700 , n373701 , n53375 , 
 n53376 , n53377 , n373705 , n53379 , n373707 , n53381 , n53382 , n373710 , n373711 , n53385 , 
 n373713 , n53387 , n53388 , n373716 , n373717 , n53391 , n373719 , n373720 , n373721 , n373722 , 
 n373723 , n53397 , n53398 , n373726 , n373727 , n373728 , n373729 , n373730 , n53404 , n373732 , 
 n373733 , n53407 , n373735 , n373736 , n373737 , n373738 , n53412 , n373740 , n373741 , n373742 , 
 n373743 , n373744 , n373745 , n373746 , n373747 , n373748 , n53422 , n373750 , n373751 , n373752 , 
 n373753 , n373754 , n53428 , n373756 , n53430 , n373758 , n53432 , n53433 , n373761 , n373762 , 
 n53436 , n373764 , n53438 , n53439 , n373767 , n53441 , n373769 , n373770 , n373771 , n373772 , 
 n53446 , n373774 , n373775 , n53449 , n373777 , n53451 , n373779 , n373780 , n373781 , n53455 , 
 n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n373789 , n53463 , n53464 , n373792 , 
 n373793 , n53467 , n373795 , n373796 , n53470 , n373798 , n53472 , n373800 , n53474 , n53475 , 
 n373803 , n373804 , n53478 , n53479 , n373807 , n53481 , n373809 , n373810 , n53484 , n373812 , 
 n53486 , n373814 , n53488 , n53489 , n373817 , n53491 , n373819 , n373820 , n53494 , n373822 , 
 n53496 , n53497 , n373825 , n373826 , n53500 , n373828 , n373829 , n53503 , n53504 , n373832 , 
 n53506 , n53507 , n373835 , n373836 , n373837 , n373838 , n373839 , n53513 , n53514 , n53515 , 
 n373843 , n53517 , n373845 , n53519 , n53520 , n373848 , n373849 , n53523 , n373851 , n373852 , 
 n373853 , n373854 , n373855 , n373856 , n373857 , n373858 , n373859 , n373860 , n53534 , n373862 , 
 n373863 , n373864 , n373865 , n373866 , n53540 , n53541 , n53542 , n53543 , n53544 , n373872 , 
 n373873 , n373874 , n373875 , n373876 , n373877 , n373878 , n373879 , n373880 , n373881 , n373882 , 
 n373883 , n373884 , n373885 , n373886 , n53557 , n373888 , n53559 , n373890 , n53561 , n373892 , 
 n53563 , n53564 , n53565 , n53566 , n373897 , n53568 , n373899 , n53570 , n373901 , n53572 , 
 n373903 , n373904 , n373905 , n373906 , n373907 , n373908 , n53579 , n373910 , n373911 , n53582 , 
 n373913 , n373914 , n373915 , n373916 , n373917 , n373918 , n373919 , n373920 , n373921 , n373922 , 
 n373923 , n373924 , n373925 , n373926 , n373927 , n53598 , n373929 , n373930 , n373931 , n373932 , 
 n373933 , n53604 , n373935 , n373936 , n373937 , n373938 , n373939 , n373940 , n53611 , n53612 , 
 n373943 , n373944 , n373945 , n373946 , n53617 , n373948 , n373949 , n53620 , n53621 , n53622 , 
 n53623 , n53624 , n53625 , n373956 , n53627 , n53628 , n373959 , n53630 , n373961 , n53632 , 
 n373963 , n53634 , n373965 , n373966 , n373967 , n53638 , n373969 , n373970 , n373971 , n373972 , 
 n373973 , n53644 , n373975 , n373976 , n373977 , n373978 , n373979 , n373980 , n53651 , n373982 , 
 n373983 , n53654 , n373985 , n373986 , n373987 , n373988 , n373989 , n373990 , n373991 , n53662 , 
 n373993 , n373994 , n373995 , n373996 , n373997 , n373998 , n53669 , n374000 , n374001 , n53672 , 
 n53673 , n374004 , n374005 , n374006 , n374007 , n374008 , n374009 , n374010 , n53681 , n374012 , 
 n53683 , n374014 , n53685 , n374016 , n374017 , n53688 , n374019 , n374020 , n53691 , n374022 , 
 n374023 , n374024 , n53695 , n374026 , n53697 , n374028 , n374029 , n374030 , n374031 , n374032 , 
 n374033 , n374034 , n374035 , n374036 , n53707 , n53708 , n374039 , n374040 , n53711 , n374042 , 
 n374043 , n374044 , n374045 , n374046 , n374047 , n53718 , n374049 , n374050 , n374051 , n374052 , 
 n374053 , n53724 , n374055 , n374056 , n374057 , n374058 , n53729 , n374060 , n374061 , n53732 , 
 n374063 , n374064 , n374065 , n374066 , n374067 , n374068 , n374069 , n374070 , n374071 , n374072 , 
 n374073 , n374074 , n374075 , n374076 , n374077 , n374078 , n374079 , n53750 , n374081 , n374082 , 
 n53753 , n374084 , n374085 , n374086 , n53757 , n374088 , n374089 , n53760 , n374091 , n53762 , 
 n374093 , n374094 , n374095 , n374096 , n53767 , n374098 , n374099 , n374100 , n374101 , n374102 , 
 n374103 , n53774 , n53775 , n374106 , n374107 , n374108 , n374109 , n374110 , n53781 , n374112 , 
 n374113 , n374114 , n374115 , n53786 , n374117 , n374118 , n374119 , n374120 , n53791 , n374122 , 
 n374123 , n374124 , n374125 , n374126 , n53797 , n374128 , n374129 , n374130 , n374131 , n374132 , 
 n374133 , n53804 , n374135 , n374136 , n53807 , n53808 , n374139 , n53810 , n374141 , n374142 , 
 n374143 , n374144 , n374145 , n374146 , n374147 , n53818 , n374149 , n374150 , n53821 , n53822 , 
 n374153 , n374154 , n374155 , n374156 , n374157 , n374158 , n374159 , n374160 , n374161 , n374162 , 
 n53833 , n374164 , n374165 , n53836 , n374167 , n374168 , n53839 , n374170 , n374171 , n53842 , 
 n374173 , n53844 , n374175 , n374176 , n53847 , n374178 , n374179 , n53850 , n374181 , n374182 , 
 n53853 , n374184 , n53855 , n53856 , n374187 , n53858 , n374189 , n53860 , n374191 , n374192 , 
 n374193 , n53864 , n374195 , n374196 , n53867 , n374198 , n374199 , n53870 , n374201 , n53872 , 
 n374203 , n374204 , n374205 , n53876 , n374207 , n53878 , n374209 , n374210 , n374211 , n374212 , 
 n374213 , n374214 , n53885 , n374216 , n374217 , n374218 , n374219 , n374220 , n374221 , n374222 , 
 n53893 , n374224 , n53895 , n374226 , n374227 , n53898 , n374229 , n374230 , n374231 , n374232 , 
 n374233 , n53904 , n374235 , n374236 , n374237 , n374238 , n53909 , n53910 , n53911 , n374242 , 
 n374243 , n53914 , n374245 , n374246 , n374247 , n53918 , n374249 , n374250 , n53921 , n374252 , 
 n374253 , n53924 , n53925 , n374256 , n53927 , n374258 , n374259 , n374260 , n374261 , n53932 , 
 n53933 , n53934 , n53935 , n374266 , n374267 , n374268 , n53939 , n374270 , n374271 , n374272 , 
 n53943 , n374274 , n374275 , n374276 , n53947 , n53948 , n374279 , n374280 , n53951 , n53952 , 
 n53953 , n374284 , n374285 , n374286 , n374287 , n374288 , n53959 , n53960 , n374291 , n53962 , 
 n374293 , n374294 , n374295 , n374296 , n374297 , n374298 , n374299 , n374300 , n374301 , n374302 , 
 n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , 
 n374313 , n374314 , n53985 , n374316 , n53987 , n374318 , n53989 , n53990 , n53991 , n374322 , 
 n374323 , n53994 , n374325 , n53996 , n374327 , n374328 , n374329 , n374330 , n374331 , n374332 , 
 n374333 , n374334 , n374335 , n54006 , n54007 , n374338 , n374339 , n374340 , n374341 , n374342 , 
 n374343 , n374344 , n374345 , n54016 , n374347 , n374348 , n374349 , n374350 , n374351 , n374352 , 
 n374353 , n374354 , n374355 , n374356 , n374357 , n374358 , n374359 , n54030 , n374361 , n54032 , 
 n374363 , n54034 , n374365 , n54036 , n374367 , n374368 , n374369 , n374370 , n374371 , n374372 , 
 n374373 , n54044 , n374375 , n374376 , n374377 , n374378 , n374379 , n374380 , n54051 , n374382 , 
 n374383 , n54054 , n374385 , n374386 , n374387 , n374388 , n374389 , n54060 , n374391 , n374392 , 
 n54063 , n374394 , n374395 , n374396 , n54067 , n54068 , n374399 , n54070 , n54071 , n374402 , 
 n374403 , n374404 , n374405 , n374406 , n374407 , n374408 , n54079 , n374410 , n374411 , n374412 , 
 n374413 , n374414 , n374415 , n374416 , n374417 , n374418 , n374419 , n374420 , n374421 , n374422 , 
 n374423 , n374424 , n54095 , n374426 , n374427 , n374428 , n374429 , n374430 , n374431 , n54102 , 
 n374433 , n54104 , n374435 , n54106 , n54107 , n374438 , n374439 , n374440 , n374441 , n374442 , 
 n374443 , n374444 , n374445 , n374446 , n54117 , n374448 , n374449 , n374450 , n374451 , n54122 , 
 n54123 , n374454 , n54125 , n374456 , n374457 , n374458 , n54129 , n374460 , n374461 , n374462 , 
 n374463 , n374464 , n374465 , n54136 , n374467 , n374468 , n54139 , n54140 , n374471 , n374472 , 
 n54143 , n54144 , n374475 , n54146 , n54147 , n374478 , n374479 , n374480 , n54151 , n374482 , 
 n374483 , n54154 , n374485 , n374486 , n54157 , n54158 , n54159 , n374490 , n374491 , n54162 , 
 n374493 , n54164 , n374495 , n54166 , n54167 , n374498 , n54169 , n374500 , n54171 , n54172 , 
 n374503 , n374504 , n54175 , n374506 , n374507 , n54178 , n374509 , n374510 , n54181 , n374512 , 
 n374513 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n374521 , n374522 , 
 n54193 , n374524 , n54195 , n54196 , n54197 , n374528 , n54199 , n374530 , n54201 , n54202 , 
 n374533 , n374534 , n54205 , n374536 , n374537 , n54208 , n374539 , n374540 , n54211 , n374542 , 
 n54213 , n54214 , n374545 , n54216 , n374547 , n54218 , n54219 , n54220 , n54221 , n374552 , 
 n374553 , n54224 , n374555 , n374556 , n54227 , n374558 , n54229 , n374560 , n54231 , n374562 , 
 n54233 , n54234 , n54235 , n374566 , n54237 , n374568 , n54239 , n54240 , n54241 , n374572 , 
 n54243 , n374574 , n54245 , n374576 , n54247 , n54248 , n374579 , n374580 , n54251 , n374582 , 
 n374583 , n54254 , n374585 , n374586 , n374587 , n54258 , n374589 , n54260 , n54261 , n374592 , 
 n374593 , n54264 , n374595 , n374596 , n54267 , n374598 , n374599 , n54270 , n374601 , n54272 , 
 n374603 , n54274 , n54275 , n374606 , n374607 , n54278 , n374609 , n374610 , n54281 , n374612 , 
 n374613 , n54284 , n374615 , n374616 , n54287 , n374618 , n374619 , n54290 , n54291 , n54292 , 
 n374623 , n374624 , n54295 , n54296 , n54297 , n54298 , n54299 , n374630 , n54301 , n54302 , 
 n54303 , n54304 , n374635 , n374636 , n54307 , n374638 , n374639 , n54310 , n374641 , n54312 , 
 n374643 , n374644 , n374645 , n54316 , n374647 , n54318 , n374649 , n54320 , n54321 , n374652 , 
 n374653 , n54324 , n374655 , n374656 , n54327 , n374658 , n374659 , n54330 , n54331 , n374662 , 
 n374663 , n54334 , n374665 , n374666 , n54337 , n374668 , n374669 , n54340 , n374671 , n54342 , 
 n374673 , n374674 , n54345 , n374676 , n54347 , n54348 , n374679 , n374680 , n54351 , n374682 , 
 n374683 , n54354 , n374685 , n54356 , n54357 , n54358 , n54359 , n374690 , n54361 , n374692 , 
 n54363 , n54364 , n374695 , n374696 , n54367 , n374698 , n374699 , n54370 , n374701 , n374702 , 
 n374703 , n54374 , n374705 , n54376 , n54377 , n54378 , n54379 , n374710 , n54381 , n54382 , 
 n54383 , n374714 , n374715 , n54386 , n374717 , n374718 , n54389 , n374720 , n374721 , n54392 , 
 n54393 , n374724 , n374725 , n54396 , n374727 , n54398 , n374729 , n54400 , n54401 , n374732 , 
 n374733 , n54404 , n374735 , n374736 , n54407 , n374738 , n374739 , n54410 , n54411 , n54412 , 
 n54413 , n54414 , n54415 , n374746 , n374747 , n54418 , n374749 , n374750 , n54421 , n374752 , 
 n374753 , n54424 , n54425 , n54426 , n374757 , n54428 , n54429 , n54430 , n374761 , n374762 , 
 n374763 , n54434 , n374765 , n54436 , n374767 , n54438 , n54439 , n374770 , n374771 , n54442 , 
 n374773 , n374774 , n54445 , n374776 , n374777 , n54448 , n54449 , n374780 , n374781 , n54452 , 
 n374783 , n374784 , n54455 , n374786 , n54457 , n374788 , n54459 , n374790 , n54461 , n374792 , 
 n54463 , n374794 , n54465 , n54466 , n374797 , n374798 , n54469 , n374800 , n374801 , n54472 , 
 n374803 , n374804 , n54475 , n54476 , n374807 , n54478 , n374809 , n54480 , n374811 , n374812 , 
 n54483 , n374814 , n54485 , n374816 , n54487 , n374818 , n374819 , n54490 , n54491 , n374822 , 
 n54493 , n54494 , n374825 , n54496 , n374827 , n54498 , n374829 , n374830 , n54501 , n374832 , 
 n374833 , n374834 , n54505 , n374836 , n54507 , n374838 , n54509 , n374840 , n374841 , n54512 , 
 n374843 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n374850 , n54521 , n54522 , 
 n374853 , n54524 , n374855 , n374856 , n374857 , n54528 , n374859 , n54530 , n374861 , n54532 , 
 n54533 , n374864 , n374865 , n54536 , n374867 , n54538 , n374869 , n54540 , n54541 , n374872 , 
 n374873 , n54544 , n374875 , n374876 , n54547 , n374878 , n374879 , n54550 , n374881 , n54552 , 
 n374883 , n54554 , n54555 , n374886 , n374887 , n54558 , n374889 , n374890 , n54561 , n374892 , 
 n374893 , n54564 , n54565 , n374896 , n374897 , n54568 , n374899 , n54570 , n374901 , n54572 , 
 n54573 , n374904 , n374905 , n54576 , n374907 , n374908 , n54579 , n374910 , n374911 , n54582 , 
 n374913 , n54584 , n54585 , n54586 , n374917 , n54588 , n374919 , n54590 , n374921 , n54592 , 
 n374923 , n54594 , n54595 , n374926 , n374927 , n54598 , n374929 , n374930 , n54601 , n374932 , 
 n54603 , n374934 , n54605 , n374936 , n374937 , n54608 , n374939 , n374940 , n54611 , n374942 , 
 n374943 , n54614 , n374945 , n374946 , n54617 , n374948 , n54619 , n374950 , n54621 , n54622 , 
 n374953 , n374954 , n54625 , n374956 , n374957 , n54628 , n374959 , n374960 , n374961 , n54632 , 
 n374963 , n54634 , n54635 , n374966 , n374967 , n54638 , n374969 , n374970 , n54641 , n374972 , 
 n54643 , n54644 , n54645 , n374976 , n54647 , n374978 , n54649 , n54650 , n374981 , n54652 , 
 n374983 , n54654 , n374985 , n54656 , n54657 , n374988 , n374989 , n54660 , n374991 , n374992 , 
 n54663 , n374994 , n374995 , n54666 , n54667 , n54668 , n54669 , n375000 , n54671 , n375002 , 
 n54673 , n375004 , n54675 , n54676 , n375007 , n375008 , n54679 , n375010 , n375011 , n54682 , 
 n375013 , n375014 , n54685 , n54686 , n54687 , n375018 , n375019 , n54690 , n375021 , n375022 , 
 n54693 , n54694 , n54695 , n375026 , n375027 , n375028 , n54699 , n375030 , n54701 , n54702 , 
 n375033 , n375034 , n54705 , n375036 , n375037 , n54708 , n375039 , n375040 , n375041 , n54712 , 
 n375043 , n54714 , n54715 , n375046 , n375047 , n54718 , n375049 , n375050 , n54721 , n375052 , 
 n375053 , n54724 , n375055 , n54726 , n375057 , n54728 , n54729 , n375060 , n375061 , n54732 , 
 n375063 , n375064 , n54735 , n375066 , n375067 , n54738 , n375069 , n375070 , n54741 , n54742 , 
 n54743 , n54744 , n375075 , n375076 , n54747 , n54748 , n54749 , n54750 , n54751 , n375082 , 
 n375083 , n54754 , n54755 , n375086 , n375087 , n54758 , n54759 , n54760 , n54761 , n375092 , 
 n54763 , n375094 , n54765 , n54766 , n375097 , n54768 , n375099 , n375100 , n54771 , n375102 , 
 n375103 , n54774 , n54775 , n54776 , n375107 , n375108 , n54779 , n54780 , n375111 , n375112 , 
 n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , 
 n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n375130 , n375131 , n54802 , 
 n375133 , n54804 , n375135 , n375136 , n54807 , n375138 , n54809 , n54810 , n375141 , n54812 , 
 n54813 , n54814 , n375145 , n375146 , n54817 , n54818 , n54819 , n375150 , n375151 , n54822 , 
 n54823 , n54824 , n375155 , n375156 , n54827 , n54828 , n54829 , n375160 , n375161 , n54832 , 
 n375163 , n375164 , n54835 , n375166 , n54837 , n375168 , n54839 , n54840 , n375171 , n375172 , 
 n54843 , n375174 , n375175 , n54846 , n375177 , n375178 , n54849 , n54850 , n375181 , n375182 , 
 n54853 , n375184 , n54855 , n375186 , n54857 , n54858 , n375189 , n375190 , n54861 , n375192 , 
 n375193 , n54864 , n375195 , n375196 , n54867 , n54868 , n54869 , n375200 , n375201 , n54872 , 
 n54873 , n375204 , n375205 , n54876 , n375207 , n54878 , n375209 , n54880 , n54881 , n375212 , 
 n375213 , n54884 , n375215 , n54886 , n375217 , n375218 , n54889 , n375220 , n375221 , n54892 , 
 n375223 , n375224 , n54895 , n375226 , n375227 , n54898 , n375229 , n54900 , n375231 , n375232 , 
 n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n375239 , n54910 , n375241 , n375242 , 
 n375243 , n54914 , n375245 , n375246 , n375247 , n54918 , n375249 , n375250 , n54921 , n375252 , 
 n375253 , n54924 , n54925 , n54926 , n375257 , n375258 , n54929 , n54930 , n375261 , n375262 , 
 n54933 , n54934 , n54935 , n375266 , n375267 , n54938 , n54939 , n54940 , n375271 , n375272 , 
 n54943 , n375274 , n375275 , n54946 , n54947 , n375278 , n54949 , n54950 , n54951 , n375282 , 
 n375283 , n54954 , n375285 , n54956 , n375287 , n375288 , n54959 , n375290 , n54961 , n375292 , 
 n54963 , n54964 , n375295 , n375296 , n54967 , n375298 , n54969 , n54970 , n54971 , n54972 , 
 n54973 , n54974 , n54975 , n54976 , n375307 , n54978 , n375309 , n54980 , n54981 , n375312 , 
 n375313 , n54984 , n54985 , n375316 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , 
 n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n375331 , n375332 , 
 n55003 , n375334 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , 
 n375343 , n375344 , n55015 , n55016 , n375347 , n375348 , n55019 , n375350 , n55021 , n375352 , 
 n375353 , n55024 , n375355 , n55026 , n55027 , n375358 , n55029 , n375360 , n375361 , n375362 , 
 n55033 , n375364 , n55035 , n375366 , n375367 , n55038 , n375369 , n375370 , n55041 , n55042 , 
 n55043 , n375374 , n375375 , n55046 , n55047 , n375378 , n375379 , n55050 , n375381 , n375382 , 
 n55053 , n375384 , n55055 , n375386 , n375387 , n55058 , n55059 , n55060 , n375391 , n55062 , 
 n55063 , n55064 , n55065 , n375396 , n55067 , n375398 , n55069 , n55070 , n375401 , n375402 , 
 n55073 , n375404 , n55075 , n55076 , n375407 , n375408 , n55079 , n375410 , n375411 , n55082 , 
 n375413 , n375414 , n375415 , n55086 , n375417 , n375418 , n55089 , n55090 , n375421 , n55092 , 
 n55093 , n375424 , n375425 , n55096 , n375427 , n375428 , n55099 , n55100 , n55101 , n55102 , 
 n375433 , n55104 , n55105 , n375436 , n375437 , n55108 , n55109 , n55110 , n55111 , n55112 , 
 n375443 , n375444 , n375445 , n375446 , n375447 , n375448 , n375449 , n375450 , n55121 , n375452 , 
 n375453 , n375454 , n375455 , n375456 , n375457 , n375458 , n375459 , n375460 , n55131 , n375462 , 
 n375463 , n375464 , n375465 , n55136 , n375467 , n55138 , n55139 , n375470 , n55141 , n375472 , 
 n375473 , n55144 , n55145 , n55146 , n55147 , n55148 , n375479 , n375480 , n55151 , n55152 , 
 n375483 , n375484 , n375485 , n375486 , n375487 , n375488 , n55159 , n55160 , n375491 , n55162 , 
 n375493 , n375494 , n375495 , n375496 , n375497 , n375498 , n375499 , n375500 , n375501 , n375502 , 
 n375503 , n375504 , n375505 , n55176 , n55177 , n375508 , n55179 , n375510 , n375511 , n375512 , 
 n55183 , n375514 , n375515 , n375516 , n375517 , n375518 , n55189 , n375520 , n375521 , n55192 , 
 n375523 , n55194 , n375525 , n375526 , n55197 , n375528 , n375529 , n55200 , n375531 , n375532 , 
 n375533 , n55204 , n375535 , n375536 , n375537 , n375538 , n375539 , n375540 , n55211 , n55212 , 
 n375543 , n55214 , n375545 , n375546 , n375547 , n55218 , n375549 , n375550 , n375551 , n375552 , 
 n375553 , n375554 , n55225 , n55226 , n55227 , n55228 , n375559 , n375560 , n55231 , n55232 , 
 n55233 , n55234 , n55235 , n375566 , n375567 , n375568 , n55239 , n375570 , n55241 , n55242 , 
 n375573 , n375574 , n55245 , n55246 , n375577 , n55248 , n375579 , n375580 , n375581 , n55252 , 
 n375583 , n375584 , n375585 , n375586 , n375587 , n375588 , n375589 , n375590 , n375591 , n55262 , 
 n375593 , n375594 , n55265 , n375596 , n375597 , n375598 , n55269 , n375600 , n375601 , n375602 , 
 n375603 , n375604 , n375605 , n375606 , n375607 , n55278 , n375609 , n55280 , n375611 , n375612 , 
 n375613 , n55284 , n55285 , n375616 , n375617 , n55288 , n375619 , n375620 , n375621 , n375622 , 
 n55293 , n375624 , n375625 , n375626 , n55297 , n55298 , n375629 , n375630 , n375631 , n375632 , 
 n55303 , n375634 , n375635 , n375636 , n55307 , n375638 , n55309 , n375640 , n375641 , n55312 , 
 n375643 , n55314 , n55315 , n375646 , n375647 , n55318 , n375649 , n375650 , n375651 , n375652 , 
 n55323 , n55324 , n55325 , n55326 , n375657 , n55328 , n55329 , n375660 , n55331 , n375662 , 
 n375663 , n55334 , n375665 , n375666 , n55337 , n55338 , n375669 , n375670 , n375671 , n375672 , 
 n55343 , n375674 , n375675 , n55346 , n375677 , n55348 , n375679 , n375680 , n375681 , n375682 , 
 n375683 , n375684 , n375685 , n55356 , n375687 , n375688 , n55359 , n375690 , n375691 , n55362 , 
 n55363 , n375694 , n375695 , n375696 , n55367 , n375698 , n375699 , n375700 , n375701 , n375702 , 
 n375703 , n55374 , n375705 , n375706 , n375707 , n375708 , n375709 , n375710 , n375711 , n55382 , 
 n375713 , n375714 , n375715 , n375716 , n375717 , n375718 , n55389 , n55390 , n375721 , n55392 , 
 n375723 , n375724 , n375725 , n375726 , n375727 , n375728 , n375729 , n55400 , n375731 , n375732 , 
 n55403 , n55404 , n375735 , n55406 , n55407 , n55408 , n375739 , n375740 , n375741 , n55412 , 
 n375743 , n375744 , n375745 , n375746 , n55417 , n375748 , n375749 , n55420 , n375751 , n375752 , 
 n55423 , n375754 , n375755 , n375756 , n375757 , n55428 , n375759 , n55430 , n375761 , n375762 , 
 n55433 , n375764 , n375765 , n55436 , n375767 , n375768 , n375769 , n375770 , n375771 , n375772 , 
 n375773 , n55444 , n375775 , n375776 , n55447 , n375778 , n375779 , n375780 , n375781 , n375782 , 
 n375783 , n375784 , n55455 , n375786 , n375787 , n55458 , n55459 , n375790 , n55461 , n55462 , 
 n375793 , n375794 , n55465 , n55466 , n375797 , n375798 , n375799 , n55470 , n375801 , n375802 , 
 n375803 , n55474 , n375805 , n55476 , n375807 , n55478 , n55479 , n375810 , n375811 , n55482 , 
 n55483 , n375814 , n55485 , n375816 , n375817 , n55488 , n375819 , n375820 , n375821 , n55492 , 
 n375823 , n55494 , n375825 , n375826 , n55497 , n375828 , n375829 , n375830 , n375831 , n55502 , 
 n375833 , n375834 , n55505 , n375836 , n375837 , n375838 , n55509 , n375840 , n55511 , n55512 , 
 n375843 , n375844 , n375845 , n375846 , n375847 , n375848 , n375849 , n55520 , n55521 , n375852 , 
 n375853 , n375854 , n55525 , n375856 , n55527 , n375858 , n55529 , n375860 , n375861 , n375862 , 
 n375863 , n375864 , n375865 , n55536 , n375867 , n375868 , n55539 , n375870 , n55541 , n375872 , 
 n375873 , n375874 , n375875 , n375876 , n375877 , n375878 , n375879 , n375880 , n375881 , n375882 , 
 n375883 , n375884 , n375885 , n375886 , n375887 , n375888 , n375889 , n375890 , n375891 , n375892 , 
 n375893 , n375894 , n375895 , n375896 , n375897 , n375898 , n375899 , n375900 , n375901 , n375902 , 
 n375903 , n375904 , n375905 , n375906 , n375907 , n375908 , n375909 , n55551 , n375911 , n375912 , 
 n375913 , n375914 , n55556 , n375916 , n55558 , n375918 , n55560 , n375920 , n375921 , n375922 , 
 n55564 , n55565 , n375925 , n55567 , n375927 , n375928 , n375929 , n55571 , n375931 , n375932 , 
 n55574 , n375934 , n375935 , n55577 , n375937 , n55578 , n375939 , n375940 , n55581 , n55582 , 
 n55583 , n375944 , n55585 , n55586 , n55587 , n375948 , n375949 , n375950 , n375951 , n375952 , 
 n375953 , n55594 , n375955 , n375956 , n55597 , n55598 , n375959 , n375960 , n55601 , n55602 , 
 n375963 , n375964 , n55605 , n55606 , n55607 , n375968 , n375969 , n55610 , n55611 , n55612 , 
 n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , 
 n55623 , n375984 , n55625 , n55626 , n55627 , n375988 , n55629 , n375990 , n55631 , n55632 , 
 n55633 , n55634 , n55635 , n375996 , n55637 , n375998 , n55639 , n55640 , n376001 , n376002 , 
 n55643 , n376004 , n376005 , n55646 , n376007 , n376008 , n376009 , n55650 , n376011 , n55652 , 
 n376013 , n376014 , n55655 , n376016 , n55657 , n55658 , n55659 , n376020 , n55661 , n376022 , 
 n55663 , n376024 , n376025 , n55666 , n376027 , n376028 , n55669 , n376030 , n376031 , n55672 , 
 n376033 , n55674 , n376035 , n55676 , n55677 , n55678 , n55679 , n55680 , n376041 , n55682 , 
 n376043 , n55684 , n55685 , n376046 , n376047 , n55688 , n376049 , n376050 , n55691 , n376052 , 
 n376053 , n376054 , n55695 , n376056 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , 
 n55703 , n55704 , n55705 , n55706 , n376067 , n55708 , n55709 , n55710 , n55711 , n55712 , 
 n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n376079 , n55720 , n376081 , n376082 , 
 n55723 , n376084 , n55725 , n376086 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , 
 n376093 , n376094 , n55735 , n376096 , n55737 , n55738 , n55739 , n55740 , n376101 , n55742 , 
 n55743 , n376104 , n55745 , n55746 , n376107 , n376108 , n55749 , n376110 , n376111 , n55752 , 
 n376113 , n376114 , n55755 , n376116 , n55757 , n55758 , n376119 , n376120 , n55761 , n376122 , 
 n376123 , n55764 , n376125 , n55766 , n55767 , n55768 , n376129 , n55770 , n55771 , n55772 , 
 n376133 , n55774 , n55775 , n376136 , n55777 , n55778 , n55779 , n376140 , n376141 , n55782 , 
 n376143 , n55784 , n376145 , n55786 , n55787 , n55788 , n376149 , n376150 , n55791 , n55792 , 
 n55793 , n376154 , n376155 , n55796 , n55797 , n376158 , n376159 , n55800 , n376161 , n55802 , 
 n376163 , n55804 , n55805 , n376166 , n55807 , n376168 , n55809 , n55810 , n376171 , n55812 , 
 n376173 , n376174 , n376175 , n55816 , n376177 , n376178 , n55819 , n376180 , n376181 , n376182 , 
 n55823 , n376184 , n376185 , n55826 , n376187 , n376188 , n55829 , n55830 , n376191 , n376192 , 
 n55833 , n55834 , n376195 , n376196 , n55837 , n376198 , n55839 , n55840 , n55841 , n376202 , 
 n55843 , n376204 , n55845 , n55846 , n376207 , n376208 , n55849 , n376210 , n376211 , n55852 , 
 n376213 , n376214 , n376215 , n376216 , n376217 , n376218 , n376219 , n376220 , n55856 , n376222 , 
 n376223 , n55859 , n376225 , n376226 , n55862 , n376228 , n55864 , n376230 , n55866 , n376232 , 
 n55868 , n55869 , n376235 , n376236 , n55872 , n376238 , n376239 , n55875 , n376241 , n376242 , 
 n55878 , n376244 , n55880 , n376246 , n376247 , n55883 , n55884 , n376250 , n376251 , n55887 , 
 n376253 , n376254 , n55890 , n376256 , n376257 , n55893 , n376259 , n55895 , n55896 , n376262 , 
 n376263 , n55899 , n376265 , n376266 , n55902 , n376268 , n55904 , n55905 , n376271 , n376272 , 
 n55908 , n376274 , n376275 , n55911 , n376277 , n55913 , n55914 , n55915 , n376281 , n376282 , 
 n55918 , n376284 , n55920 , n55921 , n55922 , n55923 , n376289 , n55925 , n55926 , n55927 , 
 n376293 , n376294 , n55930 , n376296 , n376297 , n55933 , n55934 , n55935 , n55936 , n55937 , 
 n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n376310 , n55946 , n376312 , 
 n376313 , n55949 , n376315 , n376316 , n376317 , n55953 , n376319 , n55955 , n376321 , n376322 , 
 n55958 , n376324 , n376325 , n55961 , n376327 , n376328 , n55964 , n376330 , n376331 , n55967 , 
 n55968 , n55969 , n376335 , n376336 , n55972 , n55973 , n376339 , n376340 , n55976 , n55977 , 
 n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n376352 , 
 n55988 , n376354 , n376355 , n55991 , n55992 , n55993 , n55994 , n55995 , n376361 , n55997 , 
 n55998 , n376364 , n56000 , n376366 , n56002 , n56003 , n376369 , n376370 , n376371 , n376372 , 
 n376373 , n376374 , n376375 , n376376 , n376377 , n376378 , n376379 , n376380 , n376381 , n376382 , 
 n376383 , n376384 , n376385 , n376386 , n376387 , n376388 , n376389 , n376390 , n376391 , n376392 , 
 n376393 , n376394 , n376395 , n376396 , n376397 , n376398 , n376399 , n376400 , n376401 , n376402 , 
 n376403 , n376404 , n56005 , n56006 , n56007 , n376408 , n376409 , n56010 , n376411 , n56012 , 
 n376413 , n56014 , n376415 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , 
 n56023 , n376424 , n376425 , n56026 , n376427 , n56028 , n56029 , n376430 , n376431 , n56032 , 
 n376433 , n376434 , n56035 , n376436 , n376437 , n56038 , n376439 , n56040 , n56041 , n376442 , 
 n376443 , n56044 , n376445 , n376446 , n56047 , n376448 , n56049 , n56050 , n56051 , n56052 , 
 n56053 , n56054 , n56055 , n56056 , n56057 , n376458 , n56059 , n376460 , n376461 , n56062 , 
 n376463 , n376464 , n56065 , n376466 , n376467 , n56068 , n376469 , n376470 , n56071 , n56072 , 
 n56073 , n376474 , n376475 , n56076 , n56077 , n56078 , n376479 , n376480 , n56081 , n56082 , 
 n376483 , n56084 , n376485 , n376486 , n56087 , n376488 , n56089 , n376490 , n376491 , n56092 , 
 n56093 , n56094 , n56095 , n376496 , n56097 , n56098 , n376499 , n56100 , n376501 , n376502 , 
 n56103 , n56104 , n56105 , n56106 , n56107 , n376508 , n376509 , n56110 , n376511 , n376512 , 
 n56113 , n376514 , n376515 , n376516 , n56117 , n376518 , n56119 , n56120 , n56121 , n56122 , 
 n56123 , n56124 , n56125 , n376526 , n376527 , n56128 , n376529 , n376530 , n56131 , n376532 , 
 n376533 , n56134 , n56135 , n56136 , n376537 , n376538 , n56139 , n56140 , n56141 , n56142 , 
 n56143 , n376544 , n56145 , n376546 , n376547 , n56148 , n376549 , n56150 , n376551 , n56152 , 
 n56153 , n376554 , n376555 , n56156 , n376557 , n376558 , n56159 , n376560 , n376561 , n56162 , 
 n376563 , n56164 , n56165 , n376566 , n376567 , n56168 , n376569 , n376570 , n56171 , n376572 , 
 n376573 , n56174 , n56175 , n56176 , n376577 , n56178 , n376579 , n56180 , n376581 , n56182 , 
 n56183 , n376584 , n56185 , n376586 , n56187 , n56188 , n376589 , n376590 , n56191 , n376592 , 
 n376593 , n56194 , n376595 , n376596 , n376597 , n56198 , n56199 , n376600 , n376601 , n56202 , 
 n376603 , n56204 , n56205 , n376606 , n376607 , n56208 , n376609 , n376610 , n56211 , n376612 , 
 n376613 , n56214 , n376615 , n56216 , n56217 , n376618 , n376619 , n56220 , n376621 , n376622 , 
 n56223 , n376624 , n56225 , n56226 , n56227 , n56228 , n376629 , n376630 , n56231 , n376632 , 
 n376633 , n56234 , n376635 , n56236 , n56237 , n376638 , n56239 , n376640 , n376641 , n56242 , 
 n56243 , n376644 , n376645 , n56246 , n376647 , n376648 , n56249 , n376650 , n376651 , n56252 , 
 n376653 , n376654 , n56255 , n376656 , n376657 , n56258 , n56259 , n376660 , n376661 , n56262 , 
 n56263 , n376664 , n56265 , n376666 , n376667 , n56268 , n376669 , n56270 , n56271 , n376672 , 
 n376673 , n56274 , n56275 , n376676 , n376677 , n56278 , n376679 , n56280 , n56281 , n376682 , 
 n376683 , n56284 , n56285 , n376686 , n376687 , n56288 , n56289 , n376690 , n56291 , n376692 , 
 n56293 , n56294 , n376695 , n376696 , n56297 , n376698 , n376699 , n56300 , n376701 , n376702 , 
 n56303 , n376704 , n56305 , n56306 , n376707 , n376708 , n56309 , n376710 , n376711 , n56312 , 
 n376713 , n376714 , n56315 , n376716 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , 
 n376723 , n376724 , n376725 , n376726 , n376727 , n376728 , n56324 , n376730 , n376731 , n376732 , 
 n376733 , n376734 , n376735 , n56326 , n56327 , n56328 , n56329 , n376740 , n376741 , n56332 , 
 n376743 , n376744 , n56335 , n376746 , n56337 , n56338 , n376749 , n376750 , n56341 , n376752 , 
 n376753 , n56344 , n376755 , n376756 , n56347 , n376758 , n376759 , n56350 , n376761 , n56352 , 
 n56353 , n376764 , n56355 , n376766 , n56357 , n376768 , n376769 , n56360 , n376771 , n376772 , 
 n376773 , n56364 , n376775 , n56366 , n56367 , n376778 , n376779 , n56370 , n376781 , n376782 , 
 n56373 , n376784 , n376785 , n56376 , n376787 , n56378 , n56379 , n376790 , n56381 , n376792 , 
 n56383 , n376794 , n376795 , n56386 , n376797 , n376798 , n56389 , n376800 , n56391 , n56392 , 
 n56393 , n56394 , n56395 , n56396 , n376807 , n56398 , n56399 , n376810 , n376811 , n56402 , 
 n376813 , n376814 , n56405 , n376816 , n376817 , n56408 , n56409 , n56410 , n376821 , n56412 , 
 n56413 , n376824 , n56415 , n56416 , n376827 , n56418 , n376829 , n56420 , n56421 , n376832 , 
 n376833 , n56424 , n376835 , n376836 , n56427 , n376838 , n376839 , n56430 , n376841 , n56432 , 
 n56433 , n56434 , n376845 , n56436 , n376847 , n56438 , n56439 , n56440 , n56441 , n56442 , 
 n376853 , n56444 , n376855 , n56446 , n56447 , n376858 , n376859 , n56450 , n376861 , n376862 , 
 n56453 , n376864 , n56455 , n376866 , n376867 , n376868 , n376869 , n376870 , n376871 , n376872 , 
 n376873 , n56464 , n376875 , n376876 , n56467 , n376878 , n376879 , n376880 , n376881 , n376882 , 
 n56473 , n376884 , n376885 , n56476 , n376887 , n376888 , n376889 , n376890 , n376891 , n376892 , 
 n56483 , n376894 , n376895 , n56486 , n376897 , n56488 , n56489 , n376900 , n56491 , n376902 , 
 n376903 , n376904 , n56495 , n376906 , n376907 , n376908 , n376909 , n376910 , n376911 , n376912 , 
 n56503 , n376914 , n376915 , n56506 , n376917 , n376918 , n376919 , n376920 , n376921 , n376922 , 
 n376923 , n376924 , n376925 , n376926 , n56517 , n376928 , n376929 , n56520 , n376931 , n376932 , 
 n376933 , n376934 , n376935 , n376936 , n376937 , n376938 , n376939 , n376940 , n56531 , n376942 , 
 n376943 , n56534 , n376945 , n376946 , n56537 , n56538 , n56539 , n376950 , n376951 , n56542 , 
 n376953 , n56544 , n376955 , n376956 , n56547 , n376958 , n376959 , n56550 , n376961 , n56552 , 
 n56553 , n376964 , n56555 , n376966 , n56557 , n376968 , n376969 , n56560 , n376971 , n376972 , 
 n56563 , n376974 , n56565 , n56566 , n56567 , n376978 , n376979 , n56570 , n376981 , n376982 , 
 n56573 , n376984 , n376985 , n56576 , n376987 , n376988 , n56579 , n376990 , n376991 , n56582 , 
 n376993 , n376994 , n376995 , n376996 , n376997 , n376998 , n376999 , n377000 , n377001 , n377002 , 
 n377003 , n377004 , n377005 , n377006 , n377007 , n377008 , n377009 , n377010 , n377011 , n377012 , 
 n56603 , n377014 , n377015 , n56606 , n377017 , n56608 , n377019 , n377020 , n56611 , n377022 , 
 n56613 , n377024 , n377025 , n377026 , n377027 , n377028 , n377029 , n377030 , n377031 , n56622 , 
 n56623 , n377034 , n377035 , n377036 , n377037 , n377038 , n377039 , n377040 , n377041 , n377042 , 
 n377043 , n377044 , n377045 , n377046 , n377047 , n56638 , n56639 , n56640 , n56641 , n377052 , 
 n377053 , n377054 , n377055 , n377056 , n377057 , n377058 , n377059 , n377060 , n377061 , n377062 , 
 n377063 , n56654 , n377065 , n377066 , n377067 , n377068 , n377069 , n377070 , n377071 , n377072 , 
 n56663 , n377074 , n377075 , n377076 , n377077 , n377078 , n56669 , n377080 , n377081 , n56672 , 
 n56673 , n377084 , n56675 , n377086 , n377087 , n56678 , n56679 , n56680 , n377091 , n377092 , 
 n377093 , n377094 , n377095 , n56686 , n56687 , n377098 , n56689 , n377100 , n377101 , n56692 , 
 n377103 , n377104 , n56695 , n377106 , n377107 , n377108 , n377109 , n377110 , n377111 , n377112 , 
 n56703 , n377114 , n56705 , n377116 , n56707 , n56708 , n377119 , n377120 , n56711 , n377122 , 
 n377123 , n377124 , n56715 , n56716 , n377127 , n56718 , n56719 , n377130 , n377131 , n377132 , 
 n56723 , n377134 , n377135 , n377136 , n56727 , n377138 , n377139 , n377140 , n377141 , n56732 , 
 n377143 , n377144 , n377145 , n377146 , n377147 , n377148 , n56739 , n377150 , n56741 , n377152 , 
 n377153 , n377154 , n56745 , n377156 , n377157 , n56748 , n377159 , n377160 , n377161 , n377162 , 
 n377163 , n377164 , n56755 , n377166 , n377167 , n377168 , n377169 , n377170 , n377171 , n56762 , 
 n377173 , n377174 , n56765 , n377176 , n377177 , n377178 , n377179 , n377180 , n377181 , n377182 , 
 n56773 , n56774 , n377185 , n377186 , n56777 , n377188 , n56779 , n377190 , n377191 , n56782 , 
 n377193 , n377194 , n377195 , n377196 , n377197 , n56788 , n56789 , n377200 , n56791 , n377202 , 
 n56793 , n56794 , n377205 , n377206 , n377207 , n56798 , n377209 , n56800 , n377211 , n377212 , 
 n56803 , n377214 , n377215 , n56806 , n377217 , n377218 , n377219 , n56810 , n377221 , n377222 , 
 n377223 , n56814 , n377225 , n377226 , n56817 , n377228 , n377229 , n377230 , n377231 , n377232 , 
 n377233 , n377234 , n377235 , n56826 , n56827 , n377238 , n377239 , n377240 , n56831 , n377242 , 
 n377243 , n377244 , n56835 , n377246 , n377247 , n56838 , n377249 , n377250 , n377251 , n377252 , 
 n377253 , n377254 , n377255 , n377256 , n56847 , n56848 , n56849 , n377260 , n56851 , n377262 , 
 n377263 , n56854 , n56855 , n377266 , n377267 , n377268 , n377269 , n377270 , n377271 , n56862 , 
 n377273 , n377274 , n377275 , n377276 , n377277 , n377278 , n377279 , n377280 , n56871 , n377282 , 
 n377283 , n377284 , n56875 , n377286 , n56877 , n377288 , n377289 , n377290 , n377291 , n377292 , 
 n377293 , n377294 , n377295 , n56886 , n377297 , n377298 , n56889 , n377300 , n377301 , n377302 , 
 n377303 , n377304 , n377305 , n377306 , n56897 , n377308 , n377309 , n377310 , n377311 , n377312 , 
 n377313 , n377314 , n377315 , n377316 , n377317 , n377318 , n56909 , n377320 , n56911 , n56912 , 
 n56913 , n377324 , n56915 , n56916 , n56917 , n377328 , n377329 , n56920 , n56921 , n377332 , 
 n56923 , n377334 , n377335 , n377336 , n56927 , n377338 , n377339 , n56930 , n56931 , n377342 , 
 n377343 , n56934 , n377345 , n56936 , n377347 , n56938 , n377349 , n56940 , n377351 , n377352 , 
 n377353 , n377354 , n56945 , n377356 , n377357 , n56948 , n377359 , n377360 , n56951 , n377362 , 
 n377363 , n56954 , n377365 , n377366 , n56957 , n377368 , n377369 , n377370 , n377371 , n377372 , 
 n377373 , n56964 , n377375 , n377376 , n56967 , n377378 , n377379 , n56970 , n377381 , n377382 , 
 n377383 , n377384 , n56975 , n377386 , n377387 , n56978 , n377389 , n377390 , n377391 , n377392 , 
 n377393 , n56984 , n377395 , n377396 , n377397 , n56988 , n377399 , n377400 , n377401 , n377402 , 
 n377403 , n56994 , n377405 , n377406 , n377407 , n377408 , n377409 , n377410 , n377411 , n377412 , 
 n377413 , n377414 , n57005 , n57006 , n377417 , n57008 , n377419 , n377420 , n57011 , n57012 , 
 n377423 , n377424 , n377425 , n377426 , n57017 , n377428 , n377429 , n377430 , n57021 , n57022 , 
 n377433 , n377434 , n57025 , n57026 , n57027 , n377438 , n57029 , n377440 , n57031 , n57032 , 
 n377443 , n377444 , n57035 , n377446 , n57037 , n57038 , n377449 , n377450 , n57041 , n377452 , 
 n377453 , n57044 , n377455 , n377456 , n377457 , n377458 , n377459 , n377460 , n377461 , n377462 , 
 n377463 , n377464 , n377465 , n377466 , n377467 , n377468 , n377469 , n377470 , n377471 , n377472 , 
 n377473 , n377474 , n377475 , n377476 , n377477 , n377478 , n377479 , n377480 , n57051 , n377482 , 
 n57053 , n377484 , n377485 , n377486 , n377487 , n377488 , n377489 , n377490 , n377491 , n377492 , 
 n57063 , n377494 , n377495 , n377496 , n57067 , n57068 , n377499 , n377500 , n377501 , n377502 , 
 n377503 , n377504 , n377505 , n377506 , n377507 , n377508 , n377509 , n377510 , n377511 , n57082 , 
 n377513 , n377514 , n377515 , n57086 , n377517 , n377518 , n377519 , n377520 , n377521 , n377522 , 
 n377523 , n57093 , n377525 , n377526 , n57096 , n377528 , n377529 , n377530 , n57100 , n57101 , 
 n377533 , n57103 , n57104 , n377536 , n377537 , n57107 , n377539 , n377540 , n57110 , n377542 , 
 n57112 , n377544 , n57114 , n57115 , n377547 , n377548 , n57118 , n377550 , n377551 , n57121 , 
 n377553 , n57123 , n377555 , n377556 , n377557 , n57127 , n377559 , n377560 , n57130 , n57131 , 
 n377563 , n377564 , n377565 , n377566 , n377567 , n57137 , n377569 , n377570 , n377571 , n57141 , 
 n377573 , n377574 , n57144 , n57145 , n57146 , n57147 , n377579 , n377580 , n377581 , n377582 , 
 n377583 , n377584 , n377585 , n377586 , n377587 , n377588 , n377589 , n377590 , n377591 , n377592 , 
 n377593 , n377594 , n377595 , n377596 , n57150 , n377598 , n377599 , n57153 , n57154 , n57155 , 
 n57156 , n57157 , n57158 , n377606 , n377607 , n57161 , n57162 , n377610 , n377611 , n377612 , 
 n377613 , n57167 , n377615 , n377616 , n57170 , n377618 , n377619 , n57173 , n377621 , n377622 , 
 n57176 , n377624 , n377625 , n377626 , n377627 , n377628 , n377629 , n57183 , n377631 , n377632 , 
 n377633 , n377634 , n377635 , n377636 , n377637 , n377638 , n377639 , n377640 , n57194 , n377642 , 
 n377643 , n57197 , n377645 , n377646 , n377647 , n377648 , n377649 , n57203 , n377651 , n377652 , 
 n377653 , n377654 , n377655 , n377656 , n57210 , n377658 , n377659 , n57213 , n377661 , n377662 , 
 n377663 , n377664 , n377665 , n57219 , n377667 , n57221 , n377669 , n57223 , n377671 , n377672 , 
 n57226 , n377674 , n57228 , n377676 , n57230 , n377678 , n57232 , n57233 , n57234 , n57235 , 
 n377683 , n377684 , n377685 , n377686 , n377687 , n377688 , n57242 , n377690 , n377691 , n377692 , 
 n377693 , n377694 , n57248 , n377696 , n57250 , n57251 , n377699 , n377700 , n57254 , n377702 , 
 n377703 , n57257 , n377705 , n57259 , n57260 , n57261 , n377709 , n377710 , n377711 , n377712 , 
 n377713 , n57267 , n377715 , n57269 , n57270 , n377718 , n377719 , n57273 , n377721 , n377722 , 
 n57276 , n57277 , n377725 , n377726 , n57280 , n377728 , n377729 , n57283 , n377731 , n377732 , 
 n57286 , n377734 , n377735 , n377736 , n377737 , n57291 , n377739 , n377740 , n377741 , n377742 , 
 n377743 , n57297 , n377745 , n57299 , n57300 , n57301 , n57302 , n377750 , n57304 , n377752 , 
 n57306 , n377754 , n377755 , n57309 , n377757 , n377758 , n377759 , n377760 , n57314 , n377762 , 
 n57316 , n57317 , n377765 , n377766 , n57320 , n57321 , n377769 , n57323 , n377771 , n57325 , 
 n57326 , n377774 , n57328 , n377776 , n377777 , n377778 , n377779 , n377780 , n57334 , n377782 , 
 n57336 , n377784 , n57338 , n57339 , n377787 , n377788 , n377789 , n377790 , n377791 , n57345 , 
 n377793 , n377794 , n377795 , n377796 , n57350 , n377798 , n377799 , n377800 , n377801 , n377802 , 
 n377803 , n377804 , n377805 , n57359 , n377807 , n57361 , n377809 , n377810 , n377811 , n377812 , 
 n57366 , n57367 , n377815 , n377816 , n57370 , n57371 , n377819 , n57373 , n57374 , n377822 , 
 n57376 , n377824 , n377825 , n57379 , n377827 , n57381 , n377829 , n57383 , n377831 , n377832 , 
 n377833 , n377834 , n377835 , n377836 , n377837 , n377838 , n377839 , n377840 , n57394 , n377842 , 
 n57396 , n57397 , n377845 , n377846 , n57400 , n377848 , n377849 , n377850 , n377851 , n377852 , 
 n377853 , n377854 , n377855 , n377856 , n377857 , n57411 , n377859 , n377860 , n57414 , n377862 , 
 n377863 , n377864 , n57418 , n377866 , n377867 , n57421 , n377869 , n377870 , n57424 , n377872 , 
 n377873 , n57427 , n377875 , n57429 , n57430 , n377878 , n57432 , n57433 , n377881 , n377882 , 
 n57436 , n377884 , n57438 , n57439 , n57440 , n57441 , n377889 , n57443 , n377891 , n377892 , 
 n377893 , n377894 , n377895 , n57449 , n377897 , n377898 , n377899 , n377900 , n377901 , n377902 , 
 n57456 , n377904 , n57458 , n57459 , n377907 , n57461 , n57462 , n57463 , n377911 , n57465 , 
 n377913 , n377914 , n57468 , n377916 , n377917 , n57471 , n377919 , n377920 , n57474 , n377922 , 
 n377923 , n57477 , n377925 , n377926 , n377927 , n57481 , n377929 , n377930 , n57484 , n377932 , 
 n377933 , n377934 , n377935 , n377936 , n377937 , n377938 , n377939 , n377940 , n377941 , n377942 , 
 n377943 , n377944 , n377945 , n377946 , n377947 , n377948 , n57485 , n377950 , n57487 , n377952 , 
 n377953 , n377954 , n57489 , n57490 , n377957 , n57492 , n377959 , n57494 , n377961 , n377962 , 
 n57497 , n57498 , n377965 , n377966 , n377967 , n377968 , n377969 , n57504 , n377971 , n377972 , 
 n377973 , n377974 , n377975 , n377976 , n57511 , n377978 , n377979 , n377980 , n57515 , n57516 , 
 n377983 , n377984 , n377985 , n57520 , n377987 , n377988 , n57523 , n377990 , n377991 , n377992 , 
 n57527 , n377994 , n57529 , n57530 , n377997 , n57532 , n57533 , n378000 , n57535 , n378002 , 
 n378003 , n57538 , n378005 , n378006 , n57541 , n378008 , n378009 , n57544 , n378011 , n378012 , 
 n57547 , n378014 , n378015 , n57550 , n378017 , n57552 , n378019 , n378020 , n378021 , n378022 , 
 n378023 , n378024 , n378025 , n378026 , n57561 , n57562 , n57563 , n378030 , n57565 , n378032 , 
 n378033 , n378034 , n57569 , n378036 , n378037 , n57572 , n378039 , n378040 , n378041 , n378042 , 
 n378043 , n57578 , n378045 , n378046 , n57581 , n57582 , n57583 , n378050 , n57585 , n378052 , 
 n378053 , n57588 , n378055 , n378056 , n378057 , n378058 , n378059 , n57594 , n378061 , n378062 , 
 n57597 , n378064 , n57599 , n378066 , n57601 , n378068 , n57603 , n57604 , n57605 , n378072 , 
 n378073 , n57608 , n378075 , n378076 , n57611 , n378078 , n378079 , n57614 , n378081 , n57616 , 
 n57617 , n378084 , n57619 , n378086 , n378087 , n57622 , n378089 , n57624 , n57625 , n57626 , 
 n378093 , n378094 , n378095 , n378096 , n57631 , n378098 , n378099 , n57634 , n378101 , n378102 , 
 n378103 , n378104 , n378105 , n378106 , n378107 , n57642 , n57643 , n378110 , n378111 , n57646 , 
 n378113 , n378114 , n57649 , n378116 , n378117 , n378118 , n378119 , n378120 , n378121 , n378122 , 
 n378123 , n378124 , n57659 , n378126 , n378127 , n57662 , n378129 , n57664 , n378131 , n57666 , 
 n378133 , n378134 , n378135 , n378136 , n378137 , n378138 , n57673 , n378140 , n378141 , n57676 , 
 n378143 , n378144 , n378145 , n378146 , n378147 , n378148 , n378149 , n378150 , n57685 , n378152 , 
 n378153 , n57688 , n378155 , n378156 , n378157 , n378158 , n378159 , n378160 , n378161 , n378162 , 
 n57697 , n378164 , n378165 , n378166 , n57701 , n378168 , n378169 , n378170 , n378171 , n57706 , 
 n378173 , n378174 , n57709 , n378176 , n378177 , n378178 , n378179 , n378180 , n57715 , n378182 , 
 n378183 , n378184 , n378185 , n378186 , n378187 , n57722 , n57723 , n57724 , n378191 , n378192 , 
 n57727 , n378194 , n57729 , n57730 , n378197 , n57732 , n378199 , n57734 , n57735 , n378202 , 
 n378203 , n57738 , n378205 , n378206 , n57741 , n378208 , n378209 , n57744 , n378211 , n57746 , 
 n57747 , n378214 , n378215 , n378216 , n378217 , n378218 , n57753 , n57754 , n378221 , n378222 , 
 n57757 , n378224 , n57759 , n57760 , n378227 , n57762 , n57763 , n57764 , n378231 , n378232 , 
 n57767 , n57768 , n378235 , n378236 , n57771 , n57772 , n57773 , n57774 , n378241 , n57776 , 
 n378243 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n378250 , n57785 , n57786 , 
 n378253 , n378254 , n57789 , n378256 , n57791 , n378258 , n378259 , n378260 , n57795 , n378262 , 
 n57797 , n378264 , n57799 , n57800 , n378267 , n378268 , n378269 , n378270 , n378271 , n57806 , 
 n378273 , n378274 , n57809 , n378276 , n378277 , n378278 , n378279 , n378280 , n378281 , n378282 , 
 n57817 , n378284 , n378285 , n378286 , n378287 , n378288 , n378289 , n57824 , n378291 , n378292 , 
 n378293 , n57828 , n378295 , n378296 , n378297 , n378298 , n378299 , n57834 , n57835 , n57836 , 
 n378303 , n378304 , n378305 , n57840 , n378307 , n378308 , n378309 , n57844 , n378311 , n378312 , 
 n57847 , n378314 , n378315 , n57850 , n378317 , n57852 , n378319 , n378320 , n57855 , n378322 , 
 n378323 , n57858 , n378325 , n57860 , n378327 , n378328 , n57863 , n378330 , n378331 , n57866 , 
 n378333 , n378334 , n57869 , n57870 , n378337 , n378338 , n378339 , n57874 , n378341 , n378342 , 
 n57877 , n378344 , n57879 , n378346 , n378347 , n378348 , n57883 , n378350 , n57885 , n378352 , 
 n378353 , n57888 , n57889 , n57890 , n378357 , n57892 , n57893 , n57894 , n57895 , n57896 , 
 n57897 , n57898 , n57899 , n57900 , n57901 , n378368 , n378369 , n378370 , n378371 , n378372 , 
 n378373 , n378374 , n378375 , n378376 , n57911 , n57912 , n57913 , n57914 , n378381 , n57916 , 
 n378383 , n57918 , n378385 , n378386 , n378387 , n57922 , n378389 , n57924 , n57925 , n57926 , 
 n378393 , n378394 , n57929 , n378396 , n378397 , n57932 , n57933 , n378400 , n378401 , n378402 , 
 n378403 , n378404 , n378405 , n57940 , n57941 , n378408 , n57943 , n378410 , n378411 , n378412 , 
 n378413 , n378414 , n57949 , n57950 , n378417 , n378418 , n378419 , n57954 , n378421 , n57956 , 
 n57957 , n378424 , n378425 , n378426 , n57961 , n378428 , n378429 , n57964 , n378431 , n57966 , 
 n378433 , n57968 , n57969 , n57970 , n378437 , n57972 , n57973 , n57974 , n57975 , n57976 , 
 n378443 , n57978 , n378445 , n57980 , n378447 , n57982 , n57983 , n378450 , n378451 , n57986 , 
 n378453 , n378454 , n378455 , n378456 , n378457 , n378458 , n378459 , n378460 , n378461 , n378462 , 
 n57997 , n378464 , n378465 , n378466 , n378467 , n378468 , n378469 , n378470 , n378471 , n58006 , 
 n378473 , n378474 , n58009 , n378476 , n378477 , n378478 , n58013 , n378480 , n58015 , n378482 , 
 n378483 , n378484 , n378485 , n378486 , n378487 , n378488 , n378489 , n378490 , n58025 , n378492 , 
 n378493 , n378494 , n58029 , n58030 , n378497 , n378498 , n378499 , n378500 , n378501 , n58036 , 
 n378503 , n378504 , n378505 , n378506 , n58041 , n378508 , n378509 , n378510 , n58045 , n58046 , 
 n378513 , n378514 , n58049 , n378516 , n378517 , n378518 , n378519 , n378520 , n58055 , n58056 , 
 n378523 , n378524 , n58059 , n378526 , n378527 , n58062 , n378529 , n378530 , n378531 , n58066 , 
 n58067 , n378534 , n58069 , n378536 , n58071 , n378538 , n58073 , n378540 , n378541 , n58076 , 
 n378543 , n378544 , n58079 , n378546 , n378547 , n378548 , n378549 , n378550 , n58085 , n378552 , 
 n378553 , n58088 , n378555 , n58090 , n378557 , n58092 , n58093 , n378560 , n378561 , n58096 , 
 n378563 , n378564 , n378565 , n378566 , n378567 , n378568 , n58103 , n378570 , n378571 , n58106 , 
 n58107 , n378574 , n58109 , n378576 , n58111 , n58112 , n58113 , n378580 , n58115 , n378582 , 
 n378583 , n378584 , n378585 , n378586 , n378587 , n58122 , n58123 , n58124 , n378591 , n378592 , 
 n378593 , n378594 , n378595 , n378596 , n58131 , n378598 , n378599 , n378600 , n378601 , n58136 , 
 n378603 , n58138 , n378605 , n378606 , n58141 , n378608 , n378609 , n58144 , n378611 , n378612 , 
 n378613 , n378614 , n378615 , n58150 , n378617 , n58152 , n378619 , n378620 , n58155 , n378622 , 
 n58157 , n378624 , n378625 , n58160 , n378627 , n378628 , n58163 , n58164 , n58165 , n58166 , 
 n58167 , n378634 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n378642 , 
 n378643 , n378644 , n58179 , n378646 , n378647 , n58182 , n378649 , n58184 , n58185 , n58186 , 
 n378653 , n378654 , n378655 , n378656 , n378657 , n378658 , n58193 , n378660 , n378661 , n58196 , 
 n378663 , n58198 , n378665 , n378666 , n58201 , n378668 , n378669 , n58204 , n378671 , n378672 , 
 n58207 , n378674 , n378675 , n58210 , n378677 , n58212 , n58213 , n58214 , n58215 , n58216 , 
 n58217 , n378684 , n378685 , n378686 , n378687 , n378688 , n378689 , n58224 , n378691 , n378692 , 
 n58227 , n378694 , n378695 , n378696 , n58231 , n378698 , n378699 , n58234 , n378701 , n378702 , 
 n58237 , n378704 , n378705 , n58240 , n378707 , n378708 , n58243 , n58244 , n378711 , n58246 , 
 n378713 , n378714 , n378715 , n378716 , n378717 , n378718 , n378719 , n378720 , n378721 , n378722 , 
 n378723 , n378724 , n378725 , n378726 , n378727 , n378728 , n378729 , n378730 , n378731 , n58266 , 
 n378733 , n378734 , n378735 , n378736 , n378737 , n378738 , n378739 , n378740 , n58275 , n378742 , 
 n378743 , n378744 , n378745 , n378746 , n378747 , n378748 , n378749 , n378750 , n378751 , n378752 , 
 n378753 , n58288 , n58289 , n378756 , n58291 , n378758 , n378759 , n58294 , n378761 , n378762 , 
 n58297 , n378764 , n58299 , n58300 , n378767 , n378768 , n378769 , n378770 , n378771 , n378772 , 
 n378773 , n58308 , n58309 , n378776 , n58311 , n58312 , n378779 , n58314 , n378781 , n378782 , 
 n378783 , n378784 , n58319 , n378786 , n378787 , n58322 , n378789 , n58324 , n378791 , n58326 , 
 n58327 , n378794 , n378795 , n378796 , n378797 , n378798 , n378799 , n378800 , n58335 , n378802 , 
 n378803 , n378804 , n378805 , n378806 , n378807 , n58342 , n378809 , n58344 , n58345 , n378812 , 
 n58347 , n378814 , n378815 , n58350 , n58351 , n378818 , n378819 , n58354 , n378821 , n378822 , 
 n58357 , n378824 , n58359 , n58360 , n378827 , n378828 , n58363 , n378830 , n378831 , n378832 , 
 n378833 , n378834 , n58369 , n378836 , n378837 , n58372 , n378839 , n378840 , n378841 , n378842 , 
 n378843 , n58378 , n378845 , n58380 , n378847 , n378848 , n58383 , n378850 , n58385 , n378852 , 
 n378853 , n378854 , n58389 , n378856 , n378857 , n58392 , n378859 , n378860 , n378861 , n378862 , 
 n378863 , n58398 , n378865 , n378866 , n58401 , n378868 , n58403 , n378870 , n378871 , n378872 , 
 n378873 , n378874 , n378875 , n58410 , n58411 , n378878 , n58413 , n378880 , n378881 , n58416 , 
 n378883 , n378884 , n378885 , n378886 , n378887 , n58422 , n378889 , n378890 , n58425 , n58426 , 
 n378893 , n378894 , n58429 , n378896 , n378897 , n58432 , n378899 , n58434 , n58435 , n378902 , 
 n378903 , n378904 , n378905 , n378906 , n378907 , n378908 , n378909 , n378910 , n378911 , n378912 , 
 n378913 , n58436 , n378915 , n378916 , n58439 , n378918 , n378919 , n378920 , n378921 , n378922 , 
 n378923 , n58442 , n378925 , n58444 , n378927 , n58446 , n58447 , n58448 , n378931 , n378932 , 
 n378933 , n378934 , n58453 , n378936 , n378937 , n58456 , n58457 , n378940 , n378941 , n378942 , 
 n378943 , n378944 , n378945 , n378946 , n378947 , n58462 , n58463 , n378950 , n58465 , n378952 , 
 n378953 , n58468 , n378955 , n378956 , n58471 , n378958 , n58473 , n378960 , n378961 , n58475 , 
 n378963 , n378964 , n378965 , n378966 , n58478 , n58479 , n378969 , n378970 , n58482 , n378972 , 
 n378973 , n378974 , n378975 , n58487 , n58488 , n378978 , n58490 , n58491 , n378981 , n58493 , 
 n378983 , n58495 , n58496 , n58497 , n378987 , n58499 , n378989 , n58501 , n58502 , n378992 , 
 n378993 , n378994 , n378995 , n58507 , n378997 , n378998 , n58510 , n379000 , n379001 , n58513 , 
 n58514 , n379004 , n379005 , n379006 , n379007 , n379008 , n58520 , n379010 , n379011 , n58523 , 
 n379013 , n379014 , n58526 , n379016 , n58528 , n379018 , n58530 , n379020 , n58532 , n379022 , 
 n58534 , n58535 , n379025 , n379026 , n58538 , n379028 , n379029 , n58541 , n379031 , n58543 , 
 n58544 , n58545 , n58546 , n58547 , n379037 , n379038 , n379039 , n379040 , n379041 , n379042 , 
 n58554 , n379044 , n58556 , n58557 , n58558 , n379048 , n58560 , n379050 , n58562 , n379052 , 
 n379053 , n379054 , n58566 , n379056 , n379057 , n58569 , n379059 , n379060 , n58572 , n379062 , 
 n379063 , n58575 , n379065 , n379066 , n58578 , n379068 , n379069 , n379070 , n58582 , n379072 , 
 n379073 , n379074 , n379075 , n58587 , n379077 , n379078 , n58590 , n379080 , n379081 , n379082 , 
 n58594 , n379084 , n58596 , n379086 , n58598 , n379088 , n58600 , n379090 , n379091 , n58603 , 
 n379093 , n379094 , n58606 , n379096 , n379097 , n58609 , n58610 , n379100 , n58612 , n58613 , 
 n379103 , n58615 , n379105 , n379106 , n379107 , n379108 , n379109 , n379110 , n58622 , n379112 , 
 n379113 , n58625 , n379115 , n379116 , n58628 , n379118 , n379119 , n58631 , n58632 , n379122 , 
 n379123 , n379124 , n379125 , n58637 , n379127 , n58639 , n58640 , n58641 , n58642 , n58643 , 
 n58644 , n379134 , n58646 , n379136 , n379137 , n58649 , n58650 , n58651 , n58652 , n58653 , 
 n379143 , n379144 , n58656 , n379146 , n58658 , n58659 , n379149 , n58661 , n379151 , n379152 , 
 n379153 , n58665 , n58666 , n379156 , n58668 , n379158 , n379159 , n58671 , n379161 , n379162 , 
 n379163 , n379164 , n379165 , n379166 , n379167 , n379168 , n379169 , n379170 , n379171 , n379172 , 
 n58684 , n379174 , n379175 , n58687 , n58688 , n379178 , n58690 , n58691 , n58692 , n58693 , 
 n58694 , n58695 , n379185 , n379186 , n58698 , n58699 , n379189 , n379190 , n58702 , n379192 , 
 n379193 , n379194 , n58706 , n379196 , n379197 , n379198 , n379199 , n379200 , n379201 , n58713 , 
 n58714 , n379204 , n379205 , n379206 , n379207 , n379208 , n379209 , n379210 , n379211 , n379212 , 
 n379213 , n379214 , n58726 , n58727 , n379217 , n379218 , n379219 , n58731 , n379221 , n58733 , 
 n379223 , n379224 , n58736 , n379226 , n379227 , n379228 , n58740 , n379230 , n58742 , n58743 , 
 n58744 , n58745 , n58746 , n58747 , n379237 , n379238 , n58750 , n379240 , n379241 , n379242 , 
 n58754 , n379244 , n379245 , n379246 , n379247 , n379248 , n379249 , n379250 , n379251 , n58763 , 
 n379253 , n379254 , n379255 , n58767 , n379257 , n379258 , n58770 , n379260 , n379261 , n58773 , 
 n379263 , n379264 , n379265 , n379266 , n58778 , n379268 , n58780 , n379270 , n379271 , n379272 , 
 n379273 , n379274 , n379275 , n379276 , n58788 , n379278 , n379279 , n58791 , n58792 , n379282 , 
 n379283 , n58795 , n379285 , n379286 , n379287 , n58799 , n379289 , n379290 , n379291 , n379292 , 
 n379293 , n379294 , n379295 , n379296 , n379297 , n58809 , n379299 , n379300 , n379301 , n379302 , 
 n379303 , n58815 , n379305 , n379306 , n58818 , n379308 , n379309 , n58821 , n379311 , n379312 , 
 n379313 , n379314 , n379315 , n379316 , n379317 , n379318 , n379319 , n379320 , n379321 , n379322 , 
 n379323 , n58835 , n379325 , n379326 , n58838 , n379328 , n379329 , n379330 , n379331 , n379332 , 
 n379333 , n379334 , n379335 , n379336 , n379337 , n379338 , n379339 , n379340 , n379341 , n58853 , 
 n379343 , n379344 , n58856 , n58857 , n379347 , n379348 , n379349 , n379350 , n379351 , n379352 , 
 n379353 , n379354 , n58866 , n58867 , n379357 , n58869 , n379359 , n58871 , n379361 , n58873 , 
 n379363 , n58875 , n379365 , n379366 , n58878 , n379368 , n379369 , n379370 , n379371 , n379372 , 
 n379373 , n379374 , n58886 , n379376 , n58888 , n379378 , n379379 , n379380 , n379381 , n58893 , 
 n58894 , n379384 , n58896 , n58897 , n379387 , n58899 , n379389 , n379390 , n58902 , n379392 , 
 n379393 , n58905 , n379395 , n379396 , n58908 , n379398 , n379399 , n379400 , n58912 , n58913 , 
 n379403 , n58915 , n58916 , n58917 , n379407 , n58919 , n58920 , n379410 , n58922 , n58923 , 
 n379413 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , 
 n58934 , n379424 , n58936 , n58937 , n379427 , n379428 , n379429 , n379430 , n379431 , n58943 , 
 n379433 , n58945 , n379435 , n379436 , n58948 , n379438 , n379439 , n379440 , n379441 , n58953 , 
 n379443 , n379444 , n379445 , n379446 , n379447 , n379448 , n379449 , n58961 , n379451 , n379452 , 
 n379453 , n379454 , n379455 , n379456 , n379457 , n379458 , n379459 , n379460 , n379461 , n58973 , 
 n379463 , n379464 , n379465 , n379466 , n379467 , n379468 , n379469 , n58981 , n379471 , n379472 , 
 n58984 , n379474 , n379475 , n379476 , n58988 , n379478 , n379479 , n379480 , n379481 , n379482 , 
 n379483 , n58995 , n58996 , n379486 , n58998 , n58999 , n379489 , n379490 , n379491 , n379492 , 
 n379493 , n379494 , n379495 , n379496 , n379497 , n59009 , n379499 , n379500 , n59012 , n379502 , 
 n379503 , n59015 , n59016 , n379506 , n59018 , n59019 , n59020 , n379510 , n379511 , n59023 , 
 n379513 , n379514 , n379515 , n379516 , n379517 , n59029 , n379519 , n379520 , n59032 , n59033 , 
 n379523 , n379524 , n379525 , n379526 , n379527 , n379528 , n59040 , n379530 , n379531 , n379532 , 
 n379533 , n379534 , n379535 , n379536 , n379537 , n59049 , n379539 , n379540 , n379541 , n379542 , 
 n379543 , n379544 , n59056 , n59057 , n59058 , n59059 , n59060 , n379550 , n59062 , n379552 , 
 n59064 , n379554 , n379555 , n59067 , n59068 , n379558 , n379559 , n59071 , n379561 , n379562 , 
 n379563 , n379564 , n379565 , n379566 , n59078 , n59079 , n379569 , n59081 , n379571 , n379572 , 
 n379573 , n379574 , n379575 , n379576 , n59088 , n59089 , n379579 , n379580 , n379581 , n59093 , 
 n379583 , n379584 , n59096 , n379586 , n379587 , n59099 , n379589 , n379590 , n379591 , n379592 , 
 n59104 , n379594 , n379595 , n59107 , n379597 , n59109 , n59110 , n379600 , n379601 , n59113 , 
 n379603 , n379604 , n59116 , n379606 , n59118 , n59119 , n379609 , n59121 , n379611 , n379612 , 
 n59124 , n379614 , n379615 , n59127 , n379617 , n59129 , n59130 , n379620 , n59132 , n379622 , 
 n379623 , n59135 , n379625 , n59137 , n59138 , n379628 , n379629 , n59141 , n379631 , n379632 , 
 n59144 , n59145 , n379635 , n59147 , n379637 , n379638 , n59150 , n59151 , n379641 , n59153 , 
 n379643 , n379644 , n379645 , n379646 , n379647 , n379648 , n59160 , n379650 , n379651 , n59163 , 
 n379653 , n379654 , n379655 , n379656 , n59168 , n379658 , n379659 , n379660 , n379661 , n379662 , 
 n59174 , n379664 , n379665 , n59177 , n379667 , n59179 , n379669 , n379670 , n379671 , n379672 , 
 n379673 , n379674 , n379675 , n379676 , n379677 , n379678 , n379679 , n379680 , n379681 , n379682 , 
 n379683 , n59195 , n379685 , n59197 , n59198 , n379688 , n379689 , n59201 , n379691 , n379692 , 
 n379693 , n379694 , n379695 , n379696 , n379697 , n59209 , n59210 , n379700 , n379701 , n59213 , 
 n379703 , n379704 , n59216 , n379706 , n379707 , n379708 , n379709 , n379710 , n59222 , n379712 , 
 n379713 , n59225 , n379715 , n379716 , n59228 , n379718 , n59230 , n379720 , n379721 , n59233 , 
 n379723 , n59235 , n59236 , n59237 , n59238 , n379728 , n379729 , n379730 , n379731 , n379732 , 
 n379733 , n379734 , n59246 , n379736 , n379737 , n379738 , n379739 , n379740 , n379741 , n379742 , 
 n379743 , n379744 , n379745 , n59257 , n379747 , n379748 , n59260 , n379750 , n379751 , n379752 , 
 n379753 , n59265 , n379755 , n59267 , n379757 , n59269 , n379759 , n379760 , n59272 , n379762 , 
 n379763 , n59275 , n379765 , n379766 , n59278 , n59279 , n379769 , n59281 , n379771 , n379772 , 
 n379773 , n379774 , n379775 , n379776 , n59288 , n59289 , n59290 , n59291 , n379781 , n379782 , 
 n59294 , n379784 , n379785 , n379786 , n379787 , n379788 , n379789 , n59301 , n379791 , n59303 , 
 n59304 , n379794 , n59306 , n379796 , n59308 , n379798 , n379799 , n59311 , n379801 , n379802 , 
 n379803 , n59315 , n379805 , n379806 , n59318 , n379808 , n59320 , n59321 , n379811 , n379812 , 
 n59324 , n379814 , n379815 , n379816 , n379817 , n59329 , n59330 , n59331 , n59332 , n59333 , 
 n59334 , n59335 , n59336 , n59337 , n379827 , n59339 , n379829 , n379830 , n59342 , n379832 , 
 n379833 , n379834 , n379835 , n379836 , n59348 , n379838 , n59350 , n379840 , n379841 , n379842 , 
 n379843 , n379844 , n379845 , n379846 , n379847 , n379848 , n59360 , n59361 , n379851 , n379852 , 
 n59364 , n379854 , n379855 , n379856 , n379857 , n379858 , n379859 , n379860 , n379861 , n379862 , 
 n379863 , n379864 , n379865 , n379866 , n379867 , n379868 , n379869 , n379870 , n379871 , n59383 , 
 n379873 , n59385 , n59386 , n379876 , n379877 , n59389 , n379879 , n59391 , n379881 , n379882 , 
 n379883 , n379884 , n379885 , n59397 , n379887 , n379888 , n59400 , n379890 , n379891 , n379892 , 
 n379893 , n379894 , n379895 , n59407 , n379897 , n379898 , n379899 , n59411 , n379901 , n379902 , 
 n379903 , n379904 , n379905 , n379906 , n59418 , n59419 , n59420 , n59421 , n379911 , n379912 , 
 n59424 , n379914 , n59426 , n379916 , n379917 , n59429 , n59430 , n379920 , n59432 , n59433 , 
 n59434 , n59435 , n59436 , n379926 , n59438 , n379928 , n59440 , n59441 , n379931 , n379932 , 
 n59444 , n379934 , n59446 , n59447 , n59448 , n59449 , n379939 , n59451 , n59452 , n379942 , 
 n379943 , n379944 , n59456 , n379946 , n379947 , n379948 , n379949 , n379950 , n379951 , n379952 , 
 n59464 , n379954 , n379955 , n59467 , n59468 , n59469 , n59470 , n379960 , n59472 , n379962 , 
 n59474 , n59475 , n379965 , n379966 , n379967 , n379968 , n379969 , n59481 , n379971 , n379972 , 
 n59484 , n379974 , n379975 , n379976 , n379977 , n59489 , n379979 , n379980 , n59492 , n379982 , 
 n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n379989 , n59501 , n379991 , n59503 , 
 n59504 , n379994 , n379995 , n379996 , n379997 , n379998 , n379999 , n380000 , n59512 , n59513 , 
 n380003 , n380004 , n380005 , n380006 , n59518 , n380008 , n380009 , n59521 , n380011 , n380012 , 
 n380013 , n380014 , n59526 , n380016 , n380017 , n380018 , n380019 , n59531 , n380021 , n380022 , 
 n59534 , n380024 , n380025 , n380026 , n380027 , n59539 , n380029 , n59541 , n380031 , n380032 , 
 n59544 , n380034 , n59546 , n380036 , n59548 , n380038 , n59550 , n380040 , n380041 , n380042 , 
 n380043 , n380044 , n380045 , n380046 , n380047 , n380048 , n380049 , n380050 , n380051 , n380052 , 
 n380053 , n380054 , n380055 , n380056 , n380057 , n380058 , n380059 , n380060 , n380061 , n380062 , 
 n380063 , n380064 , n380065 , n380066 , n380067 , n380068 , n380069 , n380070 , n380071 , n380072 , 
 n380073 , n380074 , n380075 , n59564 , n380077 , n380078 , n380079 , n59568 , n380081 , n380082 , 
 n59571 , n380084 , n380085 , n380086 , n380087 , n380088 , n380089 , n380090 , n380091 , n380092 , 
 n380093 , n380094 , n380095 , n380096 , n380097 , n380098 , n59587 , n59588 , n380101 , n59590 , 
 n59591 , n59592 , n380105 , n380106 , n380107 , n380108 , n380109 , n380110 , n380111 , n380112 , 
 n59601 , n59602 , n59603 , n380116 , n59605 , n59606 , n380119 , n59608 , n380121 , n380122 , 
 n380123 , n380124 , n59612 , n380126 , n59614 , n380128 , n59616 , n380130 , n59618 , n380132 , 
 n380133 , n59621 , n380135 , n380136 , n380137 , n380138 , n59626 , n380140 , n380141 , n59629 , 
 n59630 , n380144 , n380145 , n380146 , n380147 , n59635 , n380149 , n380150 , n59638 , n380152 , 
 n380153 , n59641 , n380155 , n380156 , n380157 , n380158 , n380159 , n59647 , n59648 , n59649 , 
 n380163 , n380164 , n59652 , n380166 , n380167 , n380168 , n380169 , n59657 , n380171 , n380172 , 
 n59660 , n59661 , n380175 , n380176 , n380177 , n380178 , n380179 , n380180 , n380181 , n59669 , 
 n380183 , n380184 , n59672 , n380186 , n380187 , n380188 , n380189 , n59677 , n380191 , n380192 , 
 n380193 , n59681 , n380195 , n380196 , n380197 , n380198 , n380199 , n380200 , n380201 , n380202 , 
 n59690 , n380204 , n380205 , n380206 , n380207 , n380208 , n380209 , n380210 , n380211 , n380212 , 
 n380213 , n380214 , n380215 , n380216 , n59704 , n380218 , n380219 , n59707 , n380221 , n380222 , 
 n380223 , n59711 , n380225 , n380226 , n59714 , n380228 , n380229 , n59717 , n59718 , n59719 , 
 n380233 , n380234 , n59722 , n380236 , n59724 , n380238 , n380239 , n380240 , n380241 , n59729 , 
 n380243 , n380244 , n380245 , n380246 , n59734 , n59735 , n380249 , n380250 , n59738 , n380252 , 
 n380253 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n380261 , n59749 , 
 n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n380270 , n59758 , n59759 , 
 n380273 , n380274 , n59762 , n59763 , n59764 , n59765 , n59766 , n380280 , n380281 , n380282 , 
 n59770 , n380284 , n59772 , n59773 , n380287 , n380288 , n380289 , n380290 , n380291 , n59779 , 
 n59780 , n380294 , n380295 , n59783 , n59784 , n380298 , n59786 , n59787 , n59788 , n59789 , 
 n380303 , n59791 , n59792 , n59793 , n59794 , n380308 , n380309 , n380310 , n380311 , n59799 , 
 n380313 , n380314 , n59802 , n59803 , n380317 , n59805 , n380319 , n380320 , n59808 , n380322 , 
 n59810 , n59811 , n59812 , n59813 , n59814 , n380328 , n380329 , n380330 , n380331 , n380332 , 
 n380333 , n380334 , n380335 , n380336 , n59824 , n380338 , n380339 , n59827 , n59828 , n380342 , 
 n59830 , n380344 , n59832 , n59833 , n59834 , n59835 , n380349 , n59837 , n380351 , n380352 , 
 n380353 , n380354 , n380355 , n380356 , n380357 , n380358 , n380359 , n380360 , n380361 , n380362 , 
 n380363 , n380364 , n380365 , n59853 , n380367 , n380368 , n380369 , n380370 , n380371 , n59859 , 
 n59860 , n380374 , n59862 , n59863 , n380377 , n59865 , n59866 , n59867 , n380381 , n59869 , 
 n380383 , n380384 , n59872 , n59873 , n380387 , n59875 , n380389 , n59877 , n59878 , n380392 , 
 n380393 , n380394 , n380395 , n380396 , n380397 , n380398 , n380399 , n380400 , n380401 , n380402 , 
 n380403 , n380404 , n380405 , n380406 , n380407 , n380408 , n380409 , n380410 , n380411 , n380412 , 
 n380413 , n380414 , n380415 , n380416 , n59904 , n380418 , n380419 , n380420 , n380421 , n380422 , 
 n59910 , n380424 , n59912 , n380426 , n59914 , n380428 , n380429 , n59917 , n59918 , n380432 , 
 n380433 , n380434 , n59922 , n380436 , n59924 , n380438 , n380439 , n380440 , n380441 , n380442 , 
 n380443 , n380444 , n380445 , n380446 , n380447 , n380448 , n380449 , n380450 , n380451 , n380452 , 
 n59940 , n59941 , n59942 , n59943 , n59944 , n380458 , n59946 , n380460 , n380461 , n380462 , 
 n380463 , n59951 , n380465 , n59953 , n59954 , n59955 , n380469 , n380470 , n59958 , n380472 , 
 n380473 , n59961 , n380475 , n380476 , n380477 , n380478 , n380479 , n380480 , n380481 , n380482 , 
 n59970 , n59971 , n380485 , n380486 , n380487 , n59975 , n380489 , n380490 , n380491 , n59979 , 
 n380493 , n380494 , n380495 , n380496 , n380497 , n380498 , n59986 , n380500 , n380501 , n380502 , 
 n380503 , n380504 , n59992 , n380506 , n380507 , n59995 , n59996 , n380510 , n380511 , n380512 , 
 n380513 , n380514 , n380515 , n380516 , n380517 , n380518 , n380519 , n60007 , n380521 , n380522 , 
 n380523 , n380524 , n380525 , n380526 , n60014 , n60015 , n380529 , n380530 , n380531 , n380532 , 
 n380533 , n380534 , n60022 , n380536 , n380537 , n380538 , n380539 , n60027 , n380541 , n380542 , 
 n60030 , n380544 , n60032 , n380546 , n60034 , n380548 , n380549 , n380550 , n60038 , n380552 , 
 n380553 , n380554 , n60042 , n380556 , n380557 , n380558 , n60046 , n380560 , n380561 , n60049 , 
 n60050 , n380564 , n380565 , n380566 , n60054 , n380568 , n380569 , n380570 , n380571 , n60059 , 
 n380573 , n380574 , n60062 , n60063 , n380577 , n380578 , n380579 , n60067 , n380581 , n380582 , 
 n60070 , n380584 , n380585 , n380586 , n380587 , n380588 , n380589 , n380590 , n380591 , n380592 , 
 n60080 , n60081 , n380595 , n380596 , n60084 , n380598 , n60086 , n380600 , n380601 , n60089 , 
 n60090 , n380604 , n380605 , n60093 , n60094 , n380608 , n380609 , n60097 , n380611 , n60099 , 
 n380613 , n60101 , n60102 , n380616 , n380617 , n380618 , n380619 , n60107 , n380621 , n380622 , 
 n60110 , n380624 , n380625 , n380626 , n380627 , n380628 , n380629 , n380630 , n380631 , n380632 , 
 n380633 , n380634 , n380635 , n380636 , n380637 , n380638 , n380639 , n380640 , n380641 , n60129 , 
 n60130 , n60131 , n380645 , n380646 , n380647 , n60135 , n380649 , n60137 , n380651 , n380652 , 
 n380653 , n380654 , n380655 , n60143 , n380657 , n380658 , n380659 , n60147 , n380661 , n380662 , 
 n380663 , n380664 , n380665 , n380666 , n60154 , n60155 , n380669 , n380670 , n380671 , n380672 , 
 n60160 , n380674 , n380675 , n60163 , n60164 , n380678 , n380679 , n380680 , n380681 , n380682 , 
 n380683 , n60171 , n380685 , n380686 , n380687 , n380688 , n380689 , n380690 , n380691 , n380692 , 
 n380693 , n60181 , n60182 , n380696 , n380697 , n380698 , n60186 , n380700 , n380701 , n60189 , 
 n60190 , n380704 , n380705 , n60193 , n60194 , n60195 , n380709 , n380710 , n60198 , n60199 , 
 n60200 , n380714 , n60202 , n60203 , n60204 , n380718 , n380719 , n60207 , n380721 , n380722 , 
 n60210 , n60211 , n380725 , n380726 , n60214 , n380728 , n380729 , n380730 , n380731 , n380732 , 
 n380733 , n380734 , n380735 , n380736 , n380737 , n60225 , n60226 , n60227 , n380741 , n380742 , 
 n380743 , n380744 , n380745 , n380746 , n380747 , n380748 , n60236 , n380750 , n380751 , n60239 , 
 n380753 , n380754 , n60242 , n60243 , n380757 , n380758 , n380759 , n380760 , n380761 , n380762 , 
 n60250 , n380764 , n380765 , n380766 , n60254 , n380768 , n380769 , n380770 , n380771 , n380772 , 
 n380773 , n60261 , n380775 , n60263 , n380777 , n380778 , n380779 , n380780 , n380781 , n380782 , 
 n380783 , n380784 , n60272 , n380786 , n380787 , n380788 , n60276 , n380790 , n380791 , n60279 , 
 n380793 , n380794 , n380795 , n380796 , n380797 , n380798 , n380799 , n380800 , n380801 , n380802 , 
 n380803 , n380804 , n380805 , n60293 , n380807 , n380808 , n60296 , n60297 , n380811 , n380812 , 
 n60300 , n380814 , n380815 , n380816 , n380817 , n380818 , n60306 , n380820 , n380821 , n60309 , 
 n60310 , n380824 , n380825 , n60313 , n380827 , n60315 , n380829 , n60317 , n380831 , n380832 , 
 n380833 , n380834 , n60322 , n380836 , n60324 , n380838 , n380839 , n380840 , n380841 , n380842 , 
 n380843 , n380844 , n380845 , n380846 , n380847 , n380848 , n60336 , n380850 , n380851 , n60339 , 
 n380853 , n380854 , n380855 , n60343 , n60344 , n380858 , n380859 , n60347 , n380861 , n380862 , 
 n60350 , n380864 , n380865 , n380866 , n60354 , n60355 , n380869 , n380870 , n60358 , n60359 , 
 n380873 , n60361 , n380875 , n60363 , n380877 , n60365 , n60366 , n380880 , n380881 , n60369 , 
 n380883 , n380884 , n60372 , n380886 , n380887 , n60375 , n380889 , n380890 , n380891 , n380892 , 
 n60380 , n380894 , n380895 , n380896 , n380897 , n380898 , n380899 , n380900 , n380901 , n380902 , 
 n380903 , n380904 , n380905 , n380906 , n60394 , n380908 , n380909 , n380910 , n60398 , n380912 , 
 n60400 , n380914 , n380915 , n60403 , n380917 , n60405 , n380919 , n380920 , n380921 , n380922 , 
 n380923 , n380924 , n60412 , n380926 , n380927 , n380928 , n380929 , n380930 , n380931 , n60419 , 
 n380933 , n380934 , n380935 , n380936 , n380937 , n380938 , n380939 , n380940 , n380941 , n60429 , 
 n380943 , n380944 , n380945 , n380946 , n380947 , n380948 , n60436 , n60437 , n380951 , n60439 , 
 n380953 , n60441 , n380955 , n380956 , n380957 , n60445 , n380959 , n380960 , n380961 , n380962 , 
 n60450 , n60451 , n60452 , n380966 , n380967 , n380968 , n380969 , n380970 , n380971 , n380972 , 
 n60460 , n380974 , n380975 , n380976 , n380977 , n380978 , n380979 , n60467 , n380981 , n60469 , 
 n380983 , n380984 , n380985 , n380986 , n380987 , n380988 , n380989 , n380990 , n380991 , n380992 , 
 n380993 , n380994 , n60482 , n60483 , n60484 , n380998 , n60486 , n60487 , n60488 , n60489 , 
 n60490 , n381004 , n60492 , n60493 , n381007 , n60495 , n60496 , n60497 , n60498 , n60499 , 
 n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , 
 n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n381030 , n60517 , n381032 , 
 n381033 , n381034 , n381035 , n381036 , n60520 , n381038 , n381039 , n60523 , n381041 , n381042 , 
 n60526 , n381044 , n60528 , n381046 , n381047 , n381048 , n381049 , n381050 , n381051 , n381052 , 
 n60536 , n381054 , n381055 , n60539 , n381057 , n381058 , n381059 , n60543 , n381061 , n60545 , 
 n381063 , n60547 , n60548 , n381066 , n60550 , n60551 , n381069 , n381070 , n381071 , n381072 , 
 n381073 , n381074 , n381075 , n381076 , n381077 , n381078 , n381079 , n381080 , n381081 , n381082 , 
 n381083 , n381084 , n381085 , n381086 , n381087 , n381088 , n381089 , n381090 , n381091 , n381092 , 
 n381093 , n381094 , n381095 , n381096 , n381097 , n60559 , n381099 , n381100 , n381101 , n60563 , 
 n381103 , n381104 , n60566 , n381106 , n381107 , n60569 , n381109 , n381110 , n381111 , n381112 , 
 n381113 , n381114 , n381115 , n381116 , n60578 , n60579 , n60580 , n60581 , n60582 , n381122 , 
 n381123 , n60585 , n381125 , n381126 , n381127 , n381128 , n60590 , n381130 , n381131 , n381132 , 
 n381133 , n381134 , n381135 , n381136 , n381137 , n381138 , n381139 , n381140 , n60602 , n381142 , 
 n381143 , n381144 , n381145 , n60607 , n60608 , n60609 , n381149 , n60611 , n381151 , n381152 , 
 n60614 , n381154 , n381155 , n60617 , n381157 , n381158 , n381159 , n381160 , n60621 , n381162 , 
 n381163 , n381164 , n381165 , n381166 , n381167 , n381168 , n60627 , n381170 , n381171 , n381172 , 
 n381173 , n60632 , n381175 , n381176 , n381177 , n60636 , n60637 , n381180 , n381181 , n381182 , 
 n381183 , n381184 , n60643 , n381186 , n381187 , n60646 , n381189 , n381190 , n60649 , n381192 , 
 n381193 , n60652 , n60653 , n60654 , n60655 , n381198 , n381199 , n60658 , n381201 , n381202 , 
 n381203 , n381204 , n381205 , n60664 , n381207 , n381208 , n381209 , n381210 , n381211 , n60670 , 
 n60671 , n60672 , n60673 , n381216 , n60675 , n381218 , n381219 , n381220 , n381221 , n381222 , 
 n381223 , n60682 , n381225 , n60684 , n60685 , n381228 , n381229 , n60688 , n381231 , n381232 , 
 n381233 , n60692 , n381235 , n60694 , n381237 , n381238 , n381239 , n60698 , n381241 , n381242 , 
 n381243 , n381244 , n381245 , n60704 , n381247 , n381248 , n60707 , n381250 , n381251 , n60710 , 
 n381253 , n381254 , n60713 , n381256 , n60715 , n381258 , n60717 , n381260 , n381261 , n60720 , 
 n381263 , n381264 , n60723 , n381266 , n381267 , n60726 , n381269 , n381270 , n60729 , n381272 , 
 n381273 , n60732 , n381275 , n381276 , n381277 , n381278 , n381279 , n381280 , n60739 , n381282 , 
 n381283 , n381284 , n60743 , n381286 , n381287 , n60746 , n381289 , n381290 , n381291 , n60750 , 
 n60751 , n60752 , n60753 , n381296 , n381297 , n381298 , n381299 , n381300 , n60759 , n381302 , 
 n60761 , n381304 , n381305 , n60764 , n381307 , n60766 , n381309 , n381310 , n381311 , n381312 , 
 n381313 , n381314 , n60773 , n381316 , n381317 , n60776 , n381319 , n381320 , n381321 , n381322 , 
 n60781 , n60782 , n60783 , n381326 , n60785 , n381328 , n60787 , n60788 , n381331 , n60790 , 
 n381333 , n381334 , n381335 , n381336 , n381337 , n381338 , n60797 , n381340 , n60799 , n381342 , 
 n381343 , n381344 , n381345 , n60804 , n381347 , n381348 , n381349 , n381350 , n381351 , n60810 , 
 n381353 , n381354 , n381355 , n60814 , n381357 , n381358 , n60817 , n381360 , n381361 , n60820 , 
 n381363 , n381364 , n60823 , n381366 , n381367 , n381368 , n381369 , n381370 , n60829 , n381372 , 
 n381373 , n381374 , n381375 , n381376 , n381377 , n381378 , n381379 , n60838 , n60839 , n60840 , 
 n381383 , n381384 , n381385 , n381386 , n381387 , n381388 , n381389 , n381390 , n381391 , n381392 , 
 n381393 , n381394 , n381395 , n381396 , n381397 , n381398 , n381399 , n381400 , n381401 , n381402 , 
 n381403 , n60843 , n381405 , n60845 , n381407 , n60847 , n381409 , n381410 , n60850 , n381412 , 
 n60852 , n60853 , n60854 , n381416 , n381417 , n381418 , n381419 , n381420 , n381421 , n381422 , 
 n381423 , n381424 , n60864 , n381426 , n381427 , n60867 , n381429 , n60869 , n381431 , n381432 , 
 n60872 , n381434 , n60874 , n60875 , n381437 , n381438 , n381439 , n381440 , n381441 , n381442 , 
 n381443 , n381444 , n381445 , n381446 , n381447 , n381448 , n381449 , n381450 , n381451 , n60891 , 
 n381453 , n60893 , n60894 , n381456 , n381457 , n60897 , n381459 , n381460 , n60900 , n60901 , 
 n381463 , n381464 , n60904 , n60905 , n60906 , n381468 , n381469 , n60909 , n381471 , n60911 , 
 n381473 , n381474 , n381475 , n381476 , n381477 , n381478 , n381479 , n381480 , n381481 , n60921 , 
 n381483 , n381484 , n381485 , n381486 , n381487 , n381488 , n60928 , n381490 , n381491 , n381492 , 
 n381493 , n60933 , n381495 , n381496 , n381497 , n381498 , n381499 , n381500 , n60940 , n381502 , 
 n60942 , n60943 , n381505 , n60945 , n381507 , n381508 , n60948 , n60949 , n60950 , n60951 , 
 n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n381521 , n60961 , 
 n381523 , n60963 , n60964 , n381526 , n381527 , n60967 , n381529 , n60969 , n60970 , n60971 , 
 n381533 , n60973 , n381535 , n381536 , n381537 , n60977 , n381539 , n381540 , n381541 , n60981 , 
 n381543 , n381544 , n381545 , n381546 , n381547 , n381548 , n381549 , n60989 , n60990 , n381552 , 
 n60992 , n381554 , n381555 , n381556 , n381557 , n60997 , n60998 , n381560 , n381561 , n381562 , 
 n381563 , n381564 , n381565 , n381566 , n381567 , n61007 , n381569 , n381570 , n381571 , n381572 , 
 n381573 , n381574 , n61014 , n381576 , n381577 , n381578 , n381579 , n381580 , n381581 , n61021 , 
 n381583 , n61023 , n61024 , n381586 , n381587 , n61027 , n381589 , n381590 , n61030 , n381592 , 
 n381593 , n381594 , n381595 , n381596 , n381597 , n61037 , n381599 , n381600 , n61040 , n381602 , 
 n381603 , n61043 , n381605 , n381606 , n381607 , n61047 , n61048 , n381610 , n381611 , n61051 , 
 n381613 , n381614 , n61054 , n381616 , n61056 , n381618 , n61058 , n381620 , n381621 , n61061 , 
 n381623 , n61063 , n61064 , n381626 , n61066 , n381628 , n61068 , n381630 , n381631 , n381632 , 
 n61072 , n381634 , n381635 , n381636 , n381637 , n381638 , n381639 , n61079 , n381641 , n381642 , 
 n381643 , n381644 , n381645 , n381646 , n61086 , n381648 , n381649 , n61089 , n381651 , n381652 , 
 n61092 , n381654 , n381655 , n381656 , n61096 , n381658 , n381659 , n61099 , n61100 , n381662 , 
 n61102 , n61103 , n381665 , n61105 , n381667 , n381668 , n381669 , n381670 , n381671 , n381672 , 
 n381673 , n61113 , n381675 , n381676 , n61116 , n381678 , n381679 , n61119 , n381681 , n381682 , 
 n61122 , n381684 , n381685 , n61125 , n381687 , n381688 , n61128 , n381690 , n61130 , n61131 , 
 n381693 , n381694 , n381695 , n381696 , n381697 , n61137 , n381699 , n381700 , n381701 , n381702 , 
 n61142 , n381704 , n381705 , n61145 , n61146 , n381708 , n381709 , n61149 , n381711 , n61151 , 
 n381713 , n381714 , n381715 , n381716 , n381717 , n381718 , n381719 , n381720 , n61160 , n61161 , 
 n61162 , n381724 , n61164 , n61165 , n381727 , n381728 , n381729 , n381730 , n381731 , n61171 , 
 n61172 , n381734 , n61174 , n381736 , n381737 , n381738 , n381739 , n381740 , n61180 , n381742 , 
 n381743 , n61183 , n381745 , n381746 , n61186 , n61187 , n61188 , n61189 , n61190 , n381752 , 
 n61192 , n381754 , n381755 , n381756 , n381757 , n61197 , n381759 , n381760 , n381761 , n381762 , 
 n61199 , n381764 , n381765 , n61202 , n381767 , n381768 , n61205 , n61206 , n381771 , n381772 , 
 n381773 , n61210 , n381775 , n61212 , n61213 , n381778 , n381779 , n381780 , n381781 , n61218 , 
 n381783 , n381784 , n61221 , n381786 , n381787 , n381788 , n381789 , n381790 , n381791 , n381792 , 
 n381793 , n381794 , n61231 , n61232 , n381797 , n61234 , n61235 , n381800 , n381801 , n381802 , 
 n381803 , n381804 , n381805 , n381806 , n381807 , n381808 , n381809 , n61246 , n61247 , n61248 , 
 n61249 , n381814 , n381815 , n61252 , n381817 , n61254 , n61255 , n381820 , n381821 , n381822 , 
 n381823 , n61260 , n381825 , n61262 , n381827 , n61264 , n381829 , n381830 , n61267 , n381832 , 
 n61269 , n381834 , n381835 , n381836 , n381837 , n381838 , n381839 , n381840 , n381841 , n61278 , 
 n381843 , n381844 , n61281 , n381846 , n61283 , n381848 , n381849 , n61286 , n381851 , n381852 , 
 n61289 , n381854 , n381855 , n381856 , n381857 , n381858 , n381859 , n61296 , n381861 , n381862 , 
 n381863 , n381864 , n381865 , n381866 , n61303 , n381868 , n381869 , n381870 , n381871 , n381872 , 
 n381873 , n381874 , n381875 , n381876 , n381877 , n381878 , n61315 , n381880 , n381881 , n381882 , 
 n381883 , n381884 , n381885 , n381886 , n381887 , n381888 , n61325 , n381890 , n381891 , n61328 , 
 n381893 , n61330 , n381895 , n61332 , n381897 , n381898 , n381899 , n381900 , n381901 , n381902 , 
 n381903 , n381904 , n381905 , n381906 , n381907 , n61344 , n381909 , n381910 , n61347 , n381912 , 
 n381913 , n61350 , n61351 , n381916 , n61353 , n381918 , n381919 , n381920 , n381921 , n61358 , 
 n381923 , n381924 , n381925 , n381926 , n381927 , n381928 , n381929 , n381930 , n381931 , n381932 , 
 n61369 , n381934 , n61371 , n61372 , n381937 , n381938 , n381939 , n381940 , n381941 , n61378 , 
 n381943 , n381944 , n61381 , n381946 , n61383 , n381948 , n381949 , n381950 , n381951 , n381952 , 
 n381953 , n61390 , n61391 , n381956 , n61393 , n381958 , n381959 , n381960 , n381961 , n381962 , 
 n381963 , n61400 , n381965 , n61402 , n381967 , n381968 , n381969 , n61406 , n381971 , n381972 , 
 n381973 , n381974 , n381975 , n381976 , n381977 , n381978 , n381979 , n61416 , n61417 , n381982 , 
 n61419 , n381984 , n381985 , n381986 , n381987 , n381988 , n61425 , n381990 , n381991 , n381992 , 
 n381993 , n381994 , n61431 , n381996 , n61433 , n381998 , n381999 , n61436 , n382001 , n382002 , 
 n382003 , n382004 , n382005 , n382006 , n61443 , n382008 , n61445 , n382010 , n382011 , n382012 , 
 n382013 , n382014 , n382015 , n382016 , n382017 , n382018 , n382019 , n382020 , n382021 , n382022 , 
 n61459 , n382024 , n382025 , n61462 , n382027 , n382028 , n61465 , n382030 , n382031 , n61468 , 
 n61469 , n382034 , n382035 , n61472 , n382037 , n61474 , n61475 , n382040 , n382041 , n382042 , 
 n382043 , n382044 , n382045 , n382046 , n382047 , n382048 , n382049 , n61486 , n382051 , n61488 , 
 n61489 , n382054 , n382055 , n61492 , n382057 , n382058 , n61495 , n382060 , n382061 , n61498 , 
 n382063 , n382064 , n61501 , n61502 , n61503 , n382068 , n382069 , n61506 , n61507 , n61508 , 
 n382073 , n382074 , n61511 , n61512 , n61513 , n382078 , n382079 , n61516 , n61517 , n61518 , 
 n61519 , n382084 , n382085 , n61520 , n382087 , n382088 , n382089 , n382090 , n61525 , n382092 , 
 n382093 , n382094 , n382095 , n382096 , n382097 , n382098 , n382099 , n61534 , n382101 , n382102 , 
 n382103 , n61538 , n382105 , n382106 , n61541 , n61542 , n382109 , n61544 , n382111 , n61546 , 
 n382113 , n382114 , n382115 , n382116 , n382117 , n382118 , n382119 , n382120 , n382121 , n382122 , 
 n382123 , n382124 , n382125 , n382126 , n382127 , n382128 , n382129 , n382130 , n382131 , n382132 , 
 n382133 , n382134 , n382135 , n382136 , n382137 , n382138 , n382139 , n382140 , n382141 , n382142 , 
 n382143 , n382144 , n382145 , n382146 , n382147 , n382148 , n382149 , n382150 , n382151 , n382152 , 
 n61557 , n61558 , n382155 , n61560 , n61561 , n61562 , n61563 , n382160 , n61565 , n382162 , 
 n61567 , n382164 , n61569 , n382166 , n61571 , n61572 , n61573 , n382170 , n382171 , n382172 , 
 n61577 , n61578 , n382175 , n61580 , n382177 , n382178 , n61583 , n61584 , n382181 , n382182 , 
 n382183 , n382184 , n382185 , n61590 , n382187 , n61592 , n61593 , n382190 , n382191 , n61596 , 
 n382193 , n382194 , n61599 , n382196 , n61601 , n382198 , n61603 , n382200 , n382201 , n61606 , 
 n382203 , n382204 , n382205 , n61610 , n382207 , n61612 , n382209 , n382210 , n61613 , n61614 , 
 n61615 , n61616 , n61617 , n61618 , n382217 , n382218 , n382219 , n382220 , n61623 , n382222 , 
 n382223 , n61626 , n382225 , n382226 , n61629 , n382228 , n382229 , n61632 , n61633 , n61634 , 
 n382233 , n61636 , n382235 , n382236 , n382237 , n61640 , n382239 , n61642 , n61643 , n382242 , 
 n382243 , n61646 , n382245 , n382246 , n61649 , n382248 , n382249 , n61652 , n382251 , n382252 , 
 n382253 , n382254 , n382255 , n382256 , n382257 , n61660 , n382259 , n382260 , n61663 , n382262 , 
 n382263 , n61666 , n382265 , n382266 , n382267 , n382268 , n382269 , n382270 , n382271 , n61674 , 
 n382273 , n382274 , n382275 , n382276 , n382277 , n382278 , n61681 , n382280 , n382281 , n61684 , 
 n382283 , n382284 , n61687 , n61688 , n61689 , n61690 , n382289 , n382290 , n61693 , n382292 , 
 n382293 , n61696 , n61697 , n61698 , n382297 , n382298 , n61701 , n382300 , n382301 , n61704 , 
 n382303 , n61706 , n382305 , n382306 , n382307 , n61710 , n382309 , n382310 , n61713 , n382312 , 
 n382313 , n382314 , n382315 , n382316 , n61719 , n61720 , n61721 , n61722 , n61723 , n382322 , 
 n382323 , n61726 , n382325 , n382326 , n382327 , n382328 , n382329 , n382330 , n61733 , n382332 , 
 n382333 , n382334 , n382335 , n61738 , n382337 , n382338 , n61741 , n382340 , n382341 , n61744 , 
 n382343 , n382344 , n61747 , n382346 , n382347 , n382348 , n382349 , n61752 , n382351 , n61754 , 
 n382353 , n382354 , n382355 , n382356 , n61759 , n61760 , n382359 , n382360 , n382361 , n382362 , 
 n382363 , n61766 , n382365 , n382366 , n382367 , n61770 , n382369 , n382370 , n382371 , n382372 , 
 n382373 , n61776 , n382375 , n61778 , n382377 , n382378 , n61781 , n382380 , n382381 , n61784 , 
 n382383 , n61786 , n382385 , n382386 , n382387 , n61790 , n382389 , n61792 , n382391 , n382392 , 
 n61795 , n382394 , n382395 , n61798 , n61799 , n382398 , n61801 , n382400 , n382401 , n382402 , 
 n382403 , n61806 , n382405 , n382406 , n382407 , n382408 , n382409 , n61812 , n382411 , n382412 , 
 n61815 , n382414 , n61817 , n61818 , n382417 , n382418 , n61821 , n61822 , n382421 , n61824 , 
 n382423 , n382424 , n61827 , n61828 , n61829 , n382428 , n382429 , n61832 , n382431 , n61834 , 
 n382433 , n382434 , n61837 , n382436 , n382437 , n382438 , n382439 , n382440 , n61843 , n382442 , 
 n382443 , n382444 , n382445 , n382446 , n61849 , n382448 , n382449 , n61852 , n61853 , n382452 , 
 n382453 , n382454 , n382455 , n382456 , n382457 , n382458 , n382459 , n382460 , n382461 , n382462 , 
 n382463 , n382464 , n382465 , n61868 , n382467 , n382468 , n382469 , n382470 , n61873 , n382472 , 
 n382473 , n61876 , n382475 , n382476 , n382477 , n382478 , n382479 , n382480 , n61883 , n382482 , 
 n382483 , n61886 , n382485 , n382486 , n382487 , n382488 , n382489 , n382490 , n61893 , n382492 , 
 n382493 , n382494 , n382495 , n382496 , n382497 , n61900 , n382499 , n382500 , n61903 , n382502 , 
 n382503 , n382504 , n382505 , n382506 , n382507 , n382508 , n382509 , n61912 , n382511 , n382512 , 
 n61915 , n382514 , n382515 , n61918 , n382517 , n382518 , n61921 , n382520 , n382521 , n382522 , 
 n382523 , n382524 , n382525 , n382526 , n382527 , n382528 , n382529 , n382530 , n382531 , n382532 , 
 n61935 , n382534 , n382535 , n382536 , n61939 , n382538 , n382539 , n382540 , n382541 , n382542 , 
 n382543 , n382544 , n382545 , n61948 , n61949 , n382548 , n382549 , n382550 , n382551 , n382552 , 
 n382553 , n382554 , n382555 , n382556 , n382557 , n382558 , n382559 , n382560 , n382561 , n382562 , 
 n61965 , n382564 , n382565 , n382566 , n382567 , n61970 , n382569 , n382570 , n61973 , n61974 , 
 n382573 , n382574 , n61977 , n61978 , n61979 , n382578 , n382579 , n61982 , n382581 , n382582 , 
 n382583 , n61986 , n382585 , n382586 , n61989 , n382588 , n382589 , n61992 , n382591 , n382592 , 
 n382593 , n382594 , n61997 , n382596 , n382597 , n382598 , n62001 , n382600 , n62003 , n382602 , 
 n62005 , n62006 , n62007 , n382606 , n382607 , n382608 , n62011 , n382610 , n382611 , n62014 , 
 n62015 , n62016 , n62017 , n382616 , n62019 , n382618 , n62021 , n62022 , n62023 , n62024 , 
 n382623 , n62026 , n382625 , n62028 , n382627 , n382628 , n382629 , n382630 , n382631 , n382632 , 
 n382633 , n382634 , n382635 , n382636 , n382637 , n382638 , n382639 , n382640 , n62043 , n382642 , 
 n382643 , n62046 , n382645 , n62048 , n382647 , n382648 , n382649 , n382650 , n382651 , n382652 , 
 n382653 , n62056 , n382655 , n382656 , n382657 , n62060 , n382659 , n382660 , n382661 , n62064 , 
 n382663 , n382664 , n382665 , n62068 , n382667 , n382668 , n382669 , n382670 , n382671 , n382672 , 
 n382673 , n382674 , n382675 , n382676 , n382677 , n62080 , n62081 , n382680 , n382681 , n62084 , 
 n382683 , n382684 , n382685 , n62088 , n382687 , n382688 , n62091 , n382690 , n62093 , n382692 , 
 n62095 , n382694 , n62097 , n62098 , n382697 , n62100 , n62101 , n382700 , n62103 , n382702 , 
 n382703 , n62106 , n382705 , n382706 , n382707 , n382708 , n382709 , n382710 , n382711 , n382712 , 
 n382713 , n382714 , n382715 , n62118 , n382717 , n382718 , n382719 , n382720 , n62123 , n382722 , 
 n382723 , n382724 , n62127 , n382726 , n382727 , n382728 , n62131 , n382730 , n382731 , n62134 , 
 n382733 , n382734 , n382735 , n382736 , n382737 , n382738 , n382739 , n382740 , n382741 , n382742 , 
 n382743 , n382744 , n62147 , n62148 , n382747 , n382748 , n382749 , n62152 , n382751 , n382752 , 
 n382753 , n382754 , n382755 , n382756 , n62159 , n62160 , n382759 , n382760 , n382761 , n382762 , 
 n382763 , n62166 , n382765 , n382766 , n382767 , n62170 , n382769 , n382770 , n62173 , n382772 , 
 n382773 , n62176 , n62177 , n382776 , n382777 , n382778 , n382779 , n382780 , n382781 , n62184 , 
 n62185 , n382784 , n382785 , n382786 , n62189 , n62190 , n382789 , n382790 , n62193 , n382792 , 
 n382793 , n62196 , n382795 , n382796 , n382797 , n382798 , n62201 , n62202 , n62203 , n382802 , 
 n382803 , n382804 , n382805 , n62208 , n382807 , n382808 , n382809 , n382810 , n382811 , n382812 , 
 n382813 , n62216 , n62217 , n382816 , n382817 , n62220 , n382819 , n382820 , n62223 , n382822 , 
 n382823 , n382824 , n382825 , n382826 , n382827 , n382828 , n62231 , n62232 , n382831 , n382832 , 
 n382833 , n382834 , n382835 , n382836 , n382837 , n382838 , n382839 , n62242 , n62243 , n382842 , 
 n62245 , n382844 , n382845 , n382846 , n382847 , n62250 , n382849 , n382850 , n62253 , n382852 , 
 n382853 , n382854 , n382855 , n382856 , n382857 , n382858 , n382859 , n382860 , n382861 , n62264 , 
 n382863 , n382864 , n382865 , n62268 , n382867 , n382868 , n62271 , n382870 , n382871 , n62274 , 
 n62275 , n62276 , n382875 , n382876 , n62279 , n382878 , n382879 , n62282 , n382881 , n382882 , 
 n62285 , n62286 , n382885 , n382886 , n62289 , n62290 , n62291 , n382890 , n382891 , n62294 , 
 n62295 , n62296 , n382895 , n382896 , n62299 , n382898 , n382899 , n62302 , n382901 , n62304 , 
 n382903 , n382904 , n382905 , n382906 , n62309 , n382908 , n382909 , n62312 , n382911 , n382912 , 
 n62314 , n382914 , n382915 , n62317 , n382917 , n382918 , n62319 , n382920 , n382921 , n62322 , 
 n382923 , n382924 , n62325 , n382926 , n62327 , n62328 , n62329 , n62330 , n62331 , n382932 , 
 n62333 , n382934 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , 
 n62343 , n382944 , n62345 , n382946 , n62347 , n382948 , n62349 , n382950 , n382951 , n62352 , 
 n382953 , n382954 , n62355 , n382956 , n382957 , n382958 , n382959 , n382960 , n382961 , n382962 , 
 n382963 , n382964 , n382965 , n382966 , n382967 , n382968 , n382969 , n382970 , n382971 , n382972 , 
 n382973 , n382974 , n62358 , n382976 , n62360 , n382978 , n382979 , n382980 , n62364 , n382982 , 
 n382983 , n382984 , n382985 , n382986 , n62370 , n62371 , n382989 , n382990 , n382991 , n62375 , 
 n382993 , n382994 , n382995 , n62379 , n62380 , n382998 , n382999 , n383000 , n383001 , n383002 , 
 n383003 , n383004 , n383005 , n383006 , n383007 , n62391 , n383009 , n62393 , n383011 , n383012 , 
 n383013 , n383014 , n383015 , n62399 , n383017 , n383018 , n383019 , n383020 , n62404 , n62405 , 
 n62406 , n383024 , n383025 , n62409 , n62410 , n383028 , n62412 , n62413 , n383031 , n383032 , 
 n383033 , n62417 , n383035 , n383036 , n383037 , n383038 , n383039 , n383040 , n62424 , n383042 , 
 n383043 , n383044 , n383045 , n62429 , n383047 , n383048 , n383049 , n383050 , n383051 , n383052 , 
 n383053 , n383054 , n383055 , n383056 , n383057 , n383058 , n383059 , n383060 , n383061 , n383062 , 
 n383063 , n383064 , n383065 , n383066 , n383067 , n383068 , n383069 , n383070 , n383071 , n383072 , 
 n383073 , n383074 , n62456 , n383076 , n383077 , n383078 , n383079 , n62461 , n383081 , n383082 , 
 n383083 , n383084 , n62466 , n383086 , n62468 , n383088 , n62470 , n62471 , n383091 , n62473 , 
 n383093 , n383094 , n62476 , n383096 , n62478 , n383098 , n62480 , n62481 , n383101 , n62483 , 
 n383103 , n383104 , n62486 , n383106 , n62488 , n383108 , n62490 , n383110 , n62492 , n62493 , 
 n383113 , n383114 , n383115 , n383116 , n383117 , n383118 , n383119 , n383120 , n383121 , n383122 , 
 n383123 , n383124 , n383125 , n383126 , n383127 , n383128 , n383129 , n383130 , n383131 , n383132 , 
 n383133 , n383134 , n383135 , n383136 , n383137 , n383138 , n383139 , n383140 , n383141 , n383142 , 
 n383143 , n383144 , n383145 , n383146 , n62505 , n383148 , n383149 , n62508 , n383151 , n62510 , 
 n383153 , n383154 , n383155 , n383156 , n383157 , n383158 , n383159 , n383160 , n383161 , n383162 , 
 n383163 , n383164 , n62523 , n383166 , n383167 , n62526 , n383169 , n62528 , n383171 , n383172 , 
 n62531 , n383174 , n383175 , n62534 , n383177 , n383178 , n62537 , n383180 , n383181 , n62540 , 
 n383183 , n383184 , n62543 , n383186 , n383187 , n62546 , n383189 , n383190 , n383191 , n383192 , 
 n383193 , n383194 , n383195 , n383196 , n62555 , n383198 , n383199 , n62558 , n383201 , n383202 , 
 n62561 , n383204 , n383205 , n62564 , n383207 , n383208 , n383209 , n383210 , n383211 , n383212 , 
 n383213 , n383214 , n383215 , n383216 , n62575 , n383218 , n383219 , n383220 , n62579 , n383222 , 
 n62581 , n383224 , n383225 , n383226 , n62585 , n383228 , n383229 , n383230 , n383231 , n62590 , 
 n62591 , n62592 , n62593 , n62594 , n62595 , n383238 , n62597 , n62598 , n383241 , n62600 , 
 n62601 , n383244 , n62603 , n383246 , n383247 , n383248 , n383249 , n62608 , n383251 , n62610 , 
 n383253 , n383254 , n383255 , n383256 , n383257 , n383258 , n62617 , n383260 , n383261 , n383262 , 
 n62621 , n383264 , n383265 , n383266 , n383267 , n383268 , n383269 , n383270 , n383271 , n383272 , 
 n383273 , n383274 , n383275 , n383276 , n383277 , n62636 , n62637 , n62638 , n383281 , n62640 , 
 n383283 , n383284 , n62643 , n383286 , n62645 , n383288 , n383289 , n383290 , n383291 , n383292 , 
 n62651 , n383294 , n383295 , n383296 , n383297 , n383298 , n383299 , n383300 , n62659 , n383302 , 
 n62661 , n383304 , n62663 , n383306 , n62665 , n383308 , n383309 , n62668 , n383311 , n383312 , 
 n62671 , n62672 , n383315 , n62674 , n62675 , n383318 , n383319 , n383320 , n383321 , n62680 , 
 n62681 , n383324 , n383325 , n383326 , n383327 , n62686 , n383329 , n383330 , n62689 , n62690 , 
 n383333 , n383334 , n383335 , n62694 , n383337 , n62696 , n62697 , n383340 , n383341 , n383342 , 
 n383343 , n383344 , n383345 , n383346 , n383347 , n62706 , n62707 , n383350 , n383351 , n383352 , 
 n383353 , n383354 , n383355 , n383356 , n62715 , n383358 , n383359 , n62718 , n62719 , n62720 , 
 n383363 , n383364 , n62723 , n383366 , n62725 , n383368 , n62727 , n62728 , n62729 , n383372 , 
 n62731 , n383374 , n383375 , n62734 , n383377 , n62736 , n383379 , n383380 , n62739 , n383382 , 
 n383383 , n383384 , n383385 , n383386 , n383387 , n383388 , n62747 , n383390 , n383391 , n383392 , 
 n62751 , n383394 , n383395 , n383396 , n62755 , n383398 , n383399 , n383400 , n383401 , n62760 , 
 n383403 , n383404 , n383405 , n383406 , n383407 , n383408 , n62767 , n383410 , n383411 , n383412 , 
 n383413 , n383414 , n62773 , n383416 , n383417 , n383418 , n62777 , n62778 , n383421 , n383422 , 
 n62781 , n62782 , n383425 , n383426 , n383427 , n383428 , n383429 , n62788 , n62789 , n383432 , 
 n62791 , n62792 , n62793 , n383436 , n62795 , n383438 , n383439 , n62798 , n383441 , n383442 , 
 n62801 , n383444 , n383445 , n383446 , n383447 , n62806 , n383449 , n383450 , n62809 , n383452 , 
 n383453 , n383454 , n383455 , n383456 , n383457 , n383458 , n383459 , n383460 , n62819 , n383462 , 
 n383463 , n383464 , n62823 , n383466 , n62825 , n383468 , n383469 , n383470 , n383471 , n383472 , 
 n383473 , n383474 , n383475 , n62834 , n62835 , n383478 , n383479 , n383480 , n383481 , n383482 , 
 n383483 , n62842 , n62843 , n383486 , n383487 , n383488 , n383489 , n62848 , n383491 , n383492 , 
 n383493 , n383494 , n383495 , n383496 , n383497 , n62856 , n383499 , n383500 , n62859 , n383502 , 
 n62861 , n383504 , n62863 , n383506 , n62865 , n62866 , n383509 , n383510 , n62869 , n383512 , 
 n383513 , n383514 , n383515 , n383516 , n383517 , n62876 , n383519 , n383520 , n383521 , n383522 , 
 n383523 , n383524 , n383525 , n62884 , n383527 , n383528 , n383529 , n383530 , n62889 , n383532 , 
 n383533 , n62892 , n383535 , n383536 , n383537 , n383538 , n62897 , n383540 , n383541 , n62900 , 
 n62901 , n383544 , n383545 , n383546 , n383547 , n62906 , n383549 , n383550 , n383551 , n62910 , 
 n62911 , n383554 , n383555 , n383556 , n383557 , n383558 , n383559 , n62918 , n383561 , n383562 , 
 n383563 , n62922 , n383565 , n383566 , n383567 , n383568 , n383569 , n383570 , n62929 , n62930 , 
 n383573 , n383574 , n383575 , n62934 , n383577 , n383578 , n383579 , n383580 , n383581 , n383582 , 
 n383583 , n383584 , n383585 , n62944 , n383587 , n383588 , n62947 , n383590 , n383591 , n383592 , 
 n383593 , n383594 , n383595 , n383596 , n383597 , n62956 , n383599 , n383600 , n383601 , n62960 , 
 n383603 , n383604 , n62963 , n383606 , n383607 , n62966 , n383609 , n383610 , n62969 , n383612 , 
 n383613 , n383614 , n383615 , n383616 , n383617 , n383618 , n62977 , n383620 , n62979 , n383622 , 
 n383623 , n383624 , n62983 , n383626 , n383627 , n383628 , n383629 , n383630 , n62989 , n383632 , 
 n383633 , n62992 , n383635 , n383636 , n62995 , n62996 , n383639 , n383640 , n62999 , n383642 , 
 n63001 , n383644 , n383645 , n383646 , n383647 , n383648 , n383649 , n383650 , n383651 , n383652 , 
 n383653 , n383654 , n383655 , n383656 , n63015 , n383658 , n383659 , n383660 , n383661 , n383662 , 
 n383663 , n383664 , n383665 , n383666 , n383667 , n383668 , n383669 , n63028 , n383671 , n383672 , 
 n63031 , n383674 , n383675 , n63034 , n383677 , n383678 , n63037 , n383680 , n383681 , n383682 , 
 n383683 , n383684 , n383685 , n383686 , n383687 , n63046 , n63047 , n383690 , n63049 , n383692 , 
 n383693 , n383694 , n383695 , n383696 , n63055 , n63056 , n383699 , n383700 , n63059 , n63060 , 
 n63061 , n383704 , n383705 , n63064 , n63065 , n383708 , n383709 , n63068 , n383711 , n383712 , 
 n383713 , n383714 , n63073 , n383716 , n383717 , n383718 , n63077 , n383720 , n63079 , n383722 , 
 n383723 , n63082 , n383725 , n383726 , n63085 , n383728 , n383729 , n63088 , n383731 , n383732 , 
 n383733 , n383734 , n383735 , n383736 , n383737 , n383738 , n383739 , n383740 , n383741 , n383742 , 
 n63101 , n383744 , n63103 , n383746 , n63105 , n63106 , n63107 , n383750 , n383751 , n63110 , 
 n383753 , n383754 , n383755 , n383756 , n63115 , n383758 , n383759 , n63118 , n383761 , n383762 , 
 n63121 , n383764 , n383765 , n383766 , n383767 , n383768 , n63127 , n383770 , n63129 , n63130 , 
 n383773 , n383774 , n383775 , n383776 , n383777 , n383778 , n383779 , n383780 , n383781 , n63140 , 
 n383783 , n383784 , n63143 , n383786 , n383787 , n63146 , n63147 , n383790 , n63149 , n383792 , 
 n383793 , n383794 , n383795 , n383796 , n383797 , n63156 , n63157 , n63158 , n383801 , n63160 , 
 n63161 , n383804 , n63163 , n63164 , n383807 , n63166 , n383809 , n383810 , n383811 , n383812 , 
 n383813 , n383814 , n383815 , n63174 , n383817 , n63176 , n383819 , n383820 , n383821 , n63180 , 
 n63181 , n383824 , n383825 , n63184 , n383827 , n383828 , n383829 , n63188 , n63189 , n383832 , 
 n383833 , n383834 , n383835 , n383836 , n63195 , n383838 , n383839 , n63198 , n383841 , n63200 , 
 n63201 , n63202 , n63203 , n63204 , n383847 , n383848 , n383849 , n383850 , n383851 , n383852 , 
 n383853 , n383854 , n383855 , n383856 , n63215 , n383858 , n63217 , n63218 , n63219 , n63220 , 
 n63221 , n63222 , n63223 , n383866 , n63225 , n383868 , n383869 , n383870 , n383871 , n383872 , 
 n383873 , n383874 , n63233 , n383876 , n383877 , n383878 , n383879 , n383880 , n63239 , n383882 , 
 n383883 , n383884 , n383885 , n383886 , n383887 , n383888 , n383889 , n63248 , n383891 , n383892 , 
 n383893 , n63252 , n383895 , n383896 , n383897 , n383898 , n63257 , n383900 , n383901 , n383902 , 
 n383903 , n63262 , n383905 , n383906 , n383907 , n383908 , n383909 , n383910 , n383911 , n383912 , 
 n63271 , n383914 , n383915 , n383916 , n63275 , n383918 , n383919 , n383920 , n383921 , n383922 , 
 n383923 , n383924 , n383925 , n383926 , n383927 , n383928 , n63287 , n383930 , n383931 , n63290 , 
 n383933 , n63292 , n63293 , n383936 , n63295 , n383938 , n63297 , n383940 , n383941 , n63300 , 
 n383943 , n383944 , n383945 , n383946 , n63305 , n63306 , n383949 , n383950 , n63309 , n63310 , 
 n383953 , n383954 , n63313 , n383956 , n383957 , n63316 , n383959 , n383960 , n383961 , n383962 , 
 n63321 , n383964 , n383965 , n383966 , n383967 , n383968 , n383969 , n383970 , n383971 , n383972 , 
 n383973 , n383974 , n383975 , n383976 , n383977 , n63336 , n63337 , n383980 , n383981 , n63340 , 
 n383983 , n383984 , n63343 , n63344 , n63345 , n383988 , n383989 , n383990 , n63349 , n383992 , 
 n383993 , n383994 , n383995 , n63354 , n63355 , n383998 , n383999 , n63358 , n384001 , n63360 , 
 n384003 , n384004 , n63363 , n384006 , n384007 , n63366 , n63367 , n63368 , n384011 , n63370 , 
 n384013 , n384014 , n63373 , n63374 , n384017 , n63376 , n384019 , n384020 , n63379 , n384022 , 
 n63381 , n63382 , n384025 , n384026 , n384027 , n384028 , n384029 , n384030 , n63389 , n384032 , 
 n384033 , n384034 , n63393 , n384036 , n384037 , n384038 , n63397 , n384040 , n384041 , n63400 , 
 n63401 , n384044 , n63403 , n63404 , n384047 , n63406 , n384049 , n384050 , n63409 , n63410 , 
 n384053 , n384054 , n384055 , n384056 , n63415 , n384058 , n384059 , n384060 , n384061 , n63420 , 
 n384063 , n63422 , n384065 , n384066 , n63425 , n384068 , n384069 , n384070 , n384071 , n384072 , 
 n384073 , n384074 , n384075 , n63434 , n384077 , n63436 , n384079 , n384080 , n63439 , n384082 , 
 n384083 , n63442 , n384085 , n384086 , n384087 , n63446 , n384089 , n384090 , n384091 , n384092 , 
 n384093 , n384094 , n384095 , n384096 , n384097 , n384098 , n63457 , n384100 , n63459 , n63460 , 
 n384103 , n384104 , n63463 , n384106 , n384107 , n63466 , n384109 , n384110 , n384111 , n384112 , 
 n63471 , n384114 , n384115 , n384116 , n63475 , n63476 , n384119 , n63478 , n384121 , n63480 , 
 n384123 , n384124 , n63483 , n384126 , n63485 , n384128 , n63487 , n384130 , n384131 , n63490 , 
 n384133 , n384134 , n63493 , n384136 , n63495 , n63496 , n63497 , n63498 , n384141 , n63500 , 
 n384143 , n384144 , n384145 , n384146 , n384147 , n63506 , n63507 , n384150 , n384151 , n384152 , 
 n384153 , n384154 , n384155 , n63514 , n384157 , n384158 , n384159 , n63518 , n63519 , n384162 , 
 n384163 , n384164 , n63523 , n384166 , n384167 , n384168 , n63527 , n384170 , n384171 , n384172 , 
 n63531 , n384174 , n384175 , n63534 , n63535 , n384178 , n384179 , n63538 , n384181 , n384182 , 
 n63541 , n384184 , n63543 , n384186 , n384187 , n384188 , n63547 , n384190 , n63549 , n384192 , 
 n384193 , n63552 , n384195 , n384196 , n63555 , n384198 , n384199 , n384200 , n384201 , n384202 , 
 n384203 , n63562 , n384205 , n384206 , n384207 , n384208 , n384209 , n384210 , n384211 , n384212 , 
 n384213 , n384214 , n384215 , n63574 , n384217 , n384218 , n384219 , n384220 , n63579 , n384222 , 
 n384223 , n63582 , n384225 , n384226 , n384227 , n384228 , n384229 , n63588 , n384231 , n384232 , 
 n384233 , n63592 , n384235 , n384236 , n63595 , n384238 , n384239 , n384240 , n63599 , n384242 , 
 n384243 , n384244 , n63603 , n384246 , n384247 , n63606 , n384249 , n384250 , n384251 , n384252 , 
 n384253 , n384254 , n384255 , n384256 , n384257 , n384258 , n384259 , n384260 , n384261 , n63620 , 
 n384263 , n384264 , n63623 , n63624 , n384267 , n384268 , n384269 , n63628 , n63629 , n384272 , 
 n384273 , n63632 , n384275 , n384276 , n384277 , n384278 , n384279 , n63638 , n384281 , n384282 , 
 n63641 , n384284 , n63643 , n384286 , n384287 , n384288 , n384289 , n384290 , n384291 , n63650 , 
 n63651 , n384294 , n384295 , n63654 , n384297 , n384298 , n63657 , n63658 , n384301 , n384302 , 
 n384303 , n384304 , n384305 , n63664 , n384307 , n384308 , n63667 , n63668 , n384311 , n384312 , 
 n384313 , n384314 , n384315 , n384316 , n384317 , n384318 , n384319 , n384320 , n384321 , n384322 , 
 n384323 , n384324 , n63683 , n384326 , n384327 , n384328 , n384329 , n63688 , n384331 , n384332 , 
 n384333 , n63692 , n384335 , n63694 , n63695 , n384338 , n384339 , n384340 , n384341 , n63700 , 
 n384343 , n384344 , n63703 , n384346 , n384347 , n63706 , n384349 , n384350 , n384351 , n384352 , 
 n384353 , n384354 , n384355 , n384356 , n384357 , n63716 , n384359 , n384360 , n384361 , n384362 , 
 n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n384369 , n384370 , n384371 , n384372 , 
 n384373 , n384374 , n63733 , n384376 , n384377 , n384378 , n63737 , n384380 , n384381 , n384382 , 
 n384383 , n384384 , n63743 , n384386 , n384387 , n384388 , n384389 , n384390 , n384391 , n384392 , 
 n384393 , n63752 , n384395 , n63754 , n384397 , n384398 , n384399 , n384400 , n384401 , n63760 , 
 n63761 , n63762 , n384405 , n384406 , n63765 , n384408 , n384409 , n63768 , n384411 , n63770 , 
 n63771 , n384414 , n384415 , n63774 , n384417 , n63776 , n384419 , n63778 , n384421 , n384422 , 
 n384423 , n384424 , n384425 , n384426 , n384427 , n63786 , n384429 , n384430 , n384431 , n384432 , 
 n384433 , n63792 , n384435 , n384436 , n384437 , n384438 , n384439 , n384440 , n63799 , n63800 , 
 n384443 , n384444 , n384445 , n384446 , n384447 , n63806 , n63807 , n384450 , n384451 , n63810 , 
 n384453 , n384454 , n384455 , n384456 , n384457 , n63816 , n384459 , n384460 , n384461 , n384462 , 
 n384463 , n63822 , n384465 , n384466 , n63825 , n384468 , n384469 , n384470 , n63829 , n63830 , 
 n384473 , n384474 , n63833 , n384476 , n63835 , n63836 , n384479 , n384480 , n63839 , n384482 , 
 n384483 , n63842 , n384485 , n63844 , n63845 , n63846 , n384489 , n63848 , n63849 , n384492 , 
 n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n384500 , n384501 , n384502 , 
 n384503 , n63862 , n384505 , n63864 , n384507 , n63866 , n384509 , n384510 , n63869 , n384512 , 
 n384513 , n63872 , n63873 , n384516 , n384517 , n384518 , n384519 , n63878 , n384521 , n63880 , 
 n63881 , n384524 , n384525 , n384526 , n384527 , n63886 , n384529 , n384530 , n384531 , n384532 , 
 n384533 , n384534 , n384535 , n384536 , n63895 , n63896 , n384539 , n384540 , n384541 , n384542 , 
 n384543 , n384544 , n384545 , n384546 , n63905 , n384548 , n384549 , n63908 , n384551 , n384552 , 
 n384553 , n384554 , n384555 , n384556 , n384557 , n384558 , n384559 , n384560 , n384561 , n63920 , 
 n384563 , n384564 , n384565 , n384566 , n384567 , n384568 , n384569 , n384570 , n63929 , n384572 , 
 n63931 , n384574 , n384575 , n384576 , n63935 , n384578 , n384579 , n384580 , n384581 , n384582 , 
 n384583 , n384584 , n63943 , n63944 , n384587 , n384588 , n63947 , n384590 , n63949 , n63950 , 
 n63951 , n384594 , n63953 , n384596 , n63955 , n384598 , n63957 , n384600 , n384601 , n384602 , 
 n63961 , n384604 , n384605 , n63964 , n63965 , n63966 , n384609 , n384610 , n63969 , n384612 , 
 n384613 , n63972 , n384615 , n384616 , n384617 , n384618 , n384619 , n384620 , n384621 , n384622 , 
 n63981 , n63982 , n384625 , n384626 , n63985 , n384628 , n384629 , n384630 , n63989 , n384632 , 
 n384633 , n384634 , n384635 , n384636 , n384637 , n384638 , n384639 , n384640 , n384641 , n384642 , 
 n384643 , n64002 , n384645 , n384646 , n384647 , n64006 , n384649 , n64008 , n384651 , n64010 , 
 n384653 , n384654 , n384655 , n64014 , n384657 , n64016 , n384659 , n384660 , n384661 , n384662 , 
 n384663 , n384664 , n384665 , n384666 , n384667 , n384668 , n384669 , n384670 , n384671 , n64030 , 
 n384673 , n384674 , n64033 , n64034 , n384677 , n384678 , n384679 , n384680 , n384681 , n384682 , 
 n384683 , n384684 , n384685 , n384686 , n384687 , n64046 , n384689 , n384690 , n384691 , n384692 , 
 n384693 , n64052 , n384695 , n384696 , n384697 , n384698 , n384699 , n384700 , n384701 , n384702 , 
 n384703 , n64062 , n384705 , n384706 , n64065 , n384708 , n384709 , n64068 , n384711 , n384712 , 
 n384713 , n64072 , n384715 , n384716 , n384717 , n64076 , n64077 , n384720 , n64079 , n64080 , 
 n384723 , n384724 , n384725 , n384726 , n64085 , n384728 , n384729 , n384730 , n64089 , n64090 , 
 n384733 , n384734 , n384735 , n384736 , n384737 , n64096 , n64097 , n384740 , n384741 , n384742 , 
 n64101 , n64102 , n384745 , n384746 , n384747 , n64106 , n64107 , n384750 , n384751 , n64110 , 
 n384753 , n64112 , n384755 , n64114 , n384757 , n384758 , n384759 , n64118 , n384761 , n384762 , 
 n64121 , n384764 , n384765 , n384766 , n64125 , n384768 , n64127 , n384770 , n384771 , n384772 , 
 n64131 , n384774 , n384775 , n384776 , n384777 , n384778 , n384779 , n384780 , n384781 , n64140 , 
 n384783 , n384784 , n64143 , n384786 , n384787 , n384788 , n384789 , n384790 , n384791 , n384792 , 
 n384793 , n384794 , n64153 , n64154 , n384797 , n384798 , n384799 , n384800 , n64159 , n384802 , 
 n384803 , n384804 , n384805 , n384806 , n64165 , n384808 , n384809 , n384810 , n384811 , n384812 , 
 n384813 , n64172 , n64173 , n384816 , n384817 , n64176 , n384819 , n384820 , n384821 , n64180 , 
 n384823 , n384824 , n384825 , n384826 , n64185 , n384828 , n384829 , n384830 , n64189 , n384832 , 
 n384833 , n64192 , n384835 , n384836 , n64195 , n384838 , n384839 , n64198 , n384841 , n384842 , 
 n384843 , n384844 , n64203 , n384846 , n384847 , n64206 , n384849 , n384850 , n384851 , n64210 , 
 n64211 , n384854 , n384855 , n64214 , n384857 , n384858 , n64217 , n384860 , n384861 , n384862 , 
 n384863 , n384864 , n384865 , n384866 , n384867 , n384868 , n384869 , n384870 , n384871 , n384872 , 
 n384873 , n384874 , n384875 , n64234 , n384877 , n64236 , n64237 , n384880 , n384881 , n384882 , 
 n384883 , n384884 , n384885 , n384886 , n384887 , n384888 , n64247 , n384890 , n64249 , n384892 , 
 n384893 , n384894 , n384895 , n64254 , n384897 , n384898 , n64257 , n64258 , n384901 , n384902 , 
 n64261 , n64262 , n64263 , n384906 , n384907 , n64266 , n64267 , n64268 , n384911 , n64270 , 
 n64271 , n64272 , n64273 , n384916 , n384917 , n64276 , n384919 , n384920 , n64279 , n384922 , 
 n64281 , n64282 , n384925 , n384926 , n384927 , n64286 , n384929 , n384930 , n64289 , n64290 , 
 n384933 , n384934 , n384935 , n384936 , n384937 , n384938 , n64297 , n384940 , n384941 , n384942 , 
 n384943 , n384944 , n384945 , n64304 , n384947 , n384948 , n384949 , n384950 , n384951 , n384952 , 
 n384953 , n64312 , n64313 , n384956 , n384957 , n384958 , n64317 , n384960 , n384961 , n64320 , 
 n64321 , n384964 , n384965 , n384966 , n384967 , n384968 , n384969 , n384970 , n64329 , n64330 , 
 n384973 , n384974 , n384975 , n384976 , n384977 , n384978 , n64337 , n64338 , n384981 , n384982 , 
 n64341 , n384984 , n384985 , n384986 , n384987 , n384988 , n64347 , n64348 , n384991 , n384992 , 
 n384993 , n64352 , n384995 , n384996 , n64355 , n384998 , n384999 , n385000 , n385001 , n64360 , 
 n385003 , n385004 , n64363 , n385006 , n385007 , n64366 , n64367 , n64368 , n385011 , n385012 , 
 n64371 , n385014 , n385015 , n64374 , n385017 , n64376 , n385019 , n64378 , n385021 , n385022 , 
 n64381 , n385024 , n385025 , n385026 , n64385 , n385028 , n64387 , n385030 , n64389 , n385032 , 
 n385033 , n64392 , n385035 , n385036 , n64395 , n385038 , n385039 , n385040 , n64399 , n64400 , 
 n385043 , n385044 , n64403 , n385046 , n385047 , n64406 , n385049 , n385050 , n64409 , n64410 , 
 n385053 , n385054 , n385055 , n385056 , n385057 , n64416 , n385059 , n64418 , n64419 , n385062 , 
 n385063 , n385064 , n385065 , n385066 , n64425 , n385068 , n64427 , n385070 , n385071 , n64430 , 
 n385073 , n385074 , n64433 , n385076 , n64435 , n385078 , n385079 , n385080 , n64439 , n385082 , 
 n64441 , n385084 , n64443 , n64444 , n385087 , n385088 , n385089 , n385090 , n64449 , n385092 , 
 n385093 , n64452 , n64453 , n385096 , n385097 , n385098 , n385099 , n385100 , n64459 , n385102 , 
 n385103 , n385104 , n64463 , n385106 , n385107 , n385108 , n64467 , n64468 , n385111 , n64470 , 
 n385113 , n64472 , n385115 , n64474 , n385117 , n385118 , n385119 , n385120 , n64479 , n385122 , 
 n385123 , n64482 , n64483 , n385126 , n64485 , n385128 , n385129 , n64488 , n385131 , n385132 , 
 n385133 , n385134 , n385135 , n64494 , n385137 , n385138 , n385139 , n64498 , n64499 , n385142 , 
 n64501 , n385144 , n64503 , n64504 , n64505 , n385148 , n64507 , n385150 , n64509 , n64510 , 
 n64511 , n64512 , n385155 , n64514 , n385157 , n385158 , n64517 , n385160 , n64519 , n385162 , 
 n385163 , n64522 , n385165 , n64524 , n385167 , n385168 , n385169 , n385170 , n385171 , n385172 , 
 n64531 , n64532 , n64533 , n385176 , n385177 , n385178 , n64537 , n64538 , n385181 , n385182 , 
 n64541 , n385184 , n385185 , n64544 , n385187 , n64546 , n385189 , n385190 , n385191 , n385192 , 
 n64551 , n385194 , n64553 , n385196 , n385197 , n64556 , n64557 , n64558 , n385201 , n385202 , 
 n64561 , n385204 , n64563 , n64564 , n385207 , n385208 , n385209 , n385210 , n385211 , n385212 , 
 n64571 , n385214 , n385215 , n385216 , n385217 , n385218 , n64577 , n385220 , n385221 , n64580 , 
 n385223 , n385224 , n64583 , n385226 , n385227 , n64586 , n64587 , n64588 , n64589 , n385232 , 
 n64591 , n385234 , n385235 , n385236 , n385237 , n385238 , n385239 , n64598 , n385241 , n385242 , 
 n385243 , n64602 , n385245 , n385246 , n64605 , n64606 , n385249 , n64608 , n64609 , n385252 , 
 n385253 , n385254 , n385255 , n385256 , n385257 , n385258 , n385259 , n385260 , n385261 , n385262 , 
 n385263 , n385264 , n385265 , n385266 , n385267 , n385268 , n385269 , n385270 , n385271 , n385272 , 
 n385273 , n385274 , n385275 , n385276 , n385277 , n385278 , n385279 , n385280 , n64615 , n64616 , 
 n385283 , n385284 , n385285 , n385286 , n64621 , n385288 , n385289 , n64624 , n385291 , n385292 , 
 n64627 , n64628 , n385295 , n64630 , n385297 , n385298 , n64633 , n385300 , n64635 , n64636 , 
 n385303 , n385304 , n64639 , n385306 , n385307 , n385308 , n385309 , n385310 , n64645 , n385312 , 
 n385313 , n385314 , n385315 , n385316 , n385317 , n385318 , n385319 , n385320 , n385321 , n385322 , 
 n385323 , n385324 , n385325 , n64660 , n64661 , n385328 , n64663 , n64664 , n385331 , n385332 , 
 n64667 , n385334 , n64669 , n385336 , n64671 , n64672 , n385339 , n64674 , n64675 , n385342 , 
 n64677 , n385344 , n64679 , n64680 , n385347 , n385348 , n64683 , n385350 , n385351 , n385352 , 
 n385353 , n385354 , n64689 , n64690 , n385357 , n385358 , n385359 , n385360 , n385361 , n64696 , 
 n385363 , n64698 , n385365 , n64700 , n385367 , n64702 , n385369 , n385370 , n385371 , n385372 , 
 n64707 , n385374 , n385375 , n385376 , n385377 , n385378 , n385379 , n385380 , n385381 , n385382 , 
 n385383 , n385384 , n385385 , n385386 , n64721 , n385388 , n385389 , n385390 , n385391 , n385392 , 
 n64727 , n64728 , n385395 , n385396 , n385397 , n385398 , n385399 , n385400 , n385401 , n385402 , 
 n385403 , n385404 , n385405 , n385406 , n385407 , n64742 , n385409 , n64744 , n385411 , n385412 , 
 n64747 , n64748 , n385415 , n385416 , n64751 , n385418 , n64753 , n385420 , n385421 , n385422 , 
 n64757 , n64758 , n385425 , n64760 , n385427 , n64762 , n385429 , n64764 , n385431 , n385432 , 
 n64767 , n64768 , n64769 , n385436 , n64771 , n385438 , n64773 , n64774 , n385441 , n64776 , 
 n385443 , n64778 , n385445 , n385446 , n385447 , n64782 , n385449 , n385450 , n385451 , n385452 , 
 n385453 , n385454 , n64789 , n385456 , n385457 , n64792 , n385459 , n385460 , n64795 , n385462 , 
 n64797 , n385464 , n64799 , n385466 , n64801 , n64802 , n385469 , n385470 , n385471 , n385472 , 
 n385473 , n64808 , n385475 , n385476 , n64811 , n385478 , n385479 , n385480 , n385481 , n385482 , 
 n385483 , n64818 , n385485 , n385486 , n385487 , n385488 , n64823 , n385490 , n385491 , n385492 , 
 n385493 , n64828 , n385495 , n385496 , n385497 , n64832 , n385499 , n385500 , n64835 , n385502 , 
 n385503 , n385504 , n385505 , n385506 , n64841 , n385508 , n385509 , n64844 , n385511 , n385512 , 
 n385513 , n385514 , n64849 , n385516 , n64851 , n64852 , n64853 , n64854 , n64855 , n385522 , 
 n385523 , n385524 , n64859 , n385526 , n64861 , n385528 , n385529 , n64864 , n64865 , n385532 , 
 n385533 , n385534 , n385535 , n385536 , n385537 , n64872 , n385539 , n385540 , n64875 , n385542 , 
 n385543 , n64878 , n64879 , n385546 , n64881 , n385548 , n385549 , n64884 , n64885 , n64886 , 
 n385553 , n385554 , n385555 , n64890 , n385557 , n385558 , n385559 , n385560 , n385561 , n64896 , 
 n64897 , n385564 , n385565 , n385566 , n385567 , n385568 , n64902 , n385570 , n385571 , n64905 , 
 n385573 , n385574 , n385575 , n385576 , n385577 , n385578 , n385579 , n64913 , n64914 , n64915 , 
 n385583 , n385584 , n64918 , n385586 , n64920 , n64921 , n385589 , n64923 , n385591 , n64925 , 
 n64926 , n385594 , n385595 , n385596 , n385597 , n385598 , n385599 , n385600 , n385601 , n385602 , 
 n385603 , n385604 , n385605 , n385606 , n385607 , n385608 , n385609 , n385610 , n385611 , n385612 , 
 n385613 , n385614 , n385615 , n385616 , n385617 , n385618 , n385619 , n64930 , n385621 , n385622 , 
 n385623 , n64934 , n385625 , n385626 , n64937 , n385628 , n385629 , n64940 , n385631 , n385632 , 
 n64943 , n64944 , n64945 , n385636 , n385637 , n64948 , n385639 , n385640 , n385641 , n385642 , 
 n385643 , n385644 , n385645 , n64956 , n385647 , n385648 , n64959 , n385650 , n385651 , n64962 , 
 n385653 , n64964 , n385655 , n385656 , n385657 , n385658 , n385659 , n385660 , n385661 , n385662 , 
 n385663 , n385664 , n385665 , n64976 , n385667 , n64978 , n64979 , n385670 , n385671 , n385672 , 
 n385673 , n385674 , n385675 , n64986 , n385677 , n64988 , n385679 , n385680 , n385681 , n385682 , 
 n64993 , n385684 , n385685 , n64996 , n385687 , n385688 , n385689 , n385690 , n385691 , n65002 , 
 n385693 , n385694 , n65005 , n385696 , n65007 , n385698 , n65009 , n385700 , n385701 , n65012 , 
 n385703 , n385704 , n65015 , n385706 , n385707 , n65018 , n385709 , n385710 , n385711 , n385712 , 
 n385713 , n65024 , n385715 , n385716 , n65027 , n385718 , n385719 , n65030 , n385721 , n385722 , 
 n65033 , n65034 , n385725 , n65036 , n385727 , n385728 , n385729 , n385730 , n385731 , n385732 , 
 n65043 , n65044 , n385735 , n65046 , n65047 , n385738 , n65049 , n385740 , n65051 , n385742 , 
 n385743 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n385750 , n65061 , n385752 , 
 n385753 , n65064 , n385755 , n385756 , n65067 , n385758 , n385759 , n385760 , n385761 , n385762 , 
 n65073 , n385764 , n385765 , n65076 , n385767 , n385768 , n385769 , n385770 , n385771 , n385772 , 
 n385773 , n385774 , n385775 , n65086 , n385777 , n385778 , n65089 , n385780 , n385781 , n385782 , 
 n385783 , n385784 , n385785 , n385786 , n65097 , n385788 , n385789 , n65100 , n65101 , n385792 , 
 n385793 , n65104 , n385795 , n385796 , n385797 , n65108 , n65109 , n385800 , n385801 , n385802 , 
 n385803 , n385804 , n385805 , n385806 , n65117 , n385808 , n385809 , n385810 , n385811 , n385812 , 
 n385813 , n65124 , n385815 , n385816 , n385817 , n385818 , n65129 , n65130 , n65131 , n65132 , 
 n65133 , n385824 , n385825 , n385826 , n385827 , n385828 , n385829 , n385830 , n65141 , n385832 , 
 n65143 , n385834 , n385835 , n65146 , n385837 , n385838 , n385839 , n385840 , n385841 , n385842 , 
 n385843 , n385844 , n385845 , n385846 , n385847 , n385848 , n65159 , n385850 , n385851 , n385852 , 
 n385853 , n385854 , n385855 , n65166 , n65167 , n65168 , n65169 , n65170 , n385861 , n65172 , 
 n385863 , n65174 , n385865 , n385866 , n385867 , n385868 , n385869 , n385870 , n385871 , n65182 , 
 n65183 , n65184 , n385875 , n65186 , n385877 , n65188 , n385879 , n385880 , n65191 , n385882 , 
 n65193 , n385884 , n65195 , n385886 , n385887 , n65198 , n65199 , n65200 , n385891 , n385892 , 
 n385893 , n385894 , n385895 , n385896 , n385897 , n385898 , n385899 , n385900 , n65211 , n385902 , 
 n65213 , n385904 , n385905 , n385906 , n385907 , n385908 , n385909 , n385910 , n385911 , n385912 , 
 n385913 , n385914 , n65225 , n385916 , n65227 , n65228 , n385919 , n385920 , n385921 , n385922 , 
 n385923 , n65234 , n385925 , n65236 , n385927 , n65238 , n385929 , n65240 , n65241 , n385932 , 
 n385933 , n385934 , n385935 , n65246 , n385937 , n385938 , n65249 , n385940 , n65251 , n385942 , 
 n385943 , n385944 , n385945 , n385946 , n385947 , n385948 , n385949 , n385950 , n385951 , n385952 , 
 n65263 , n385954 , n385955 , n65266 , n385957 , n65268 , n385959 , n385960 , n65271 , n385962 , 
 n385963 , n385964 , n65275 , n385966 , n385967 , n385968 , n385969 , n65280 , n65281 , n385972 , 
 n385973 , n385974 , n385975 , n385976 , n385977 , n385978 , n65289 , n385980 , n385981 , n385982 , 
 n385983 , n385984 , n65295 , n65296 , n65297 , n65298 , n65299 , n385990 , n385991 , n65302 , 
 n385993 , n385994 , n65305 , n385996 , n385997 , n385998 , n65309 , n386000 , n386001 , n386002 , 
 n386003 , n386004 , n386005 , n386006 , n386007 , n386008 , n386009 , n65320 , n65321 , n386012 , 
 n386013 , n65324 , n386015 , n386016 , n65327 , n386018 , n386019 , n386020 , n65331 , n65332 , 
 n65333 , n386024 , n386025 , n65336 , n386027 , n386028 , n386029 , n386030 , n386031 , n386032 , 
 n65343 , n386034 , n386035 , n386036 , n386037 , n386038 , n65349 , n386040 , n65351 , n386042 , 
 n386043 , n65354 , n386045 , n65356 , n386047 , n386048 , n386049 , n65360 , n386051 , n386052 , 
 n65363 , n386054 , n65365 , n65366 , n386057 , n386058 , n386059 , n386060 , n386061 , n386062 , 
 n386063 , n386064 , n386065 , n386066 , n386067 , n386068 , n386069 , n386070 , n386071 , n386072 , 
 n386073 , n386074 , n386075 , n386076 , n386077 , n386078 , n386079 , n386080 , n386081 , n386082 , 
 n386083 , n386084 , n386085 , n386086 , n386087 , n386088 , n386089 , n386090 , n386091 , n386092 , 
 n386093 , n386094 , n386095 , n386096 , n65372 , n386098 , n386099 , n386100 , n386101 , n386102 , 
 n386103 , n386104 , n386105 , n386106 , n65382 , n386108 , n386109 , n65385 , n386111 , n386112 , 
 n386113 , n386114 , n386115 , n386116 , n65392 , n386118 , n386119 , n386120 , n65396 , n386122 , 
 n386123 , n386124 , n386125 , n386126 , n386127 , n386128 , n386129 , n386130 , n386131 , n386132 , 
 n386133 , n386134 , n386135 , n386136 , n386137 , n65413 , n386139 , n65415 , n386141 , n65417 , 
 n386143 , n386144 , n65420 , n386146 , n386147 , n386148 , n386149 , n386150 , n386151 , n386152 , 
 n65428 , n386154 , n65430 , n386156 , n65432 , n386158 , n386159 , n65435 , n386161 , n386162 , 
 n386163 , n386164 , n386165 , n386166 , n386167 , n386168 , n386169 , n386170 , n386171 , n65441 , 
 n386173 , n386174 , n65444 , n386176 , n386177 , n386178 , n386179 , n386180 , n386181 , n386182 , 
 n386183 , n386184 , n386185 , n386186 , n386187 , n386188 , n386189 , n386190 , n386191 , n386192 , 
 n386193 , n386194 , n386195 , n386196 , n65466 , n386198 , n65468 , n386200 , n386201 , n386202 , 
 n65472 , n386204 , n386205 , n386206 , n386207 , n386208 , n65478 , n386210 , n386211 , n65481 , 
 n386213 , n386214 , n65484 , n386216 , n386217 , n386218 , n386219 , n386220 , n386221 , n386222 , 
 n386223 , n386224 , n386225 , n65495 , n386227 , n386228 , n386229 , n386230 , n386231 , n386232 , 
 n386233 , n386234 , n386235 , n386236 , n65506 , n386238 , n65508 , n386240 , n65510 , n386242 , 
 n65512 , n386244 , n386245 , n65515 , n386247 , n65517 , n386249 , n386250 , n65520 , n65521 , 
 n65522 , n65523 , n65524 , n65525 , n65526 , n386258 , n65528 , n65529 , n386261 , n65531 , 
 n386263 , n386264 , n386265 , n65535 , n386267 , n386268 , n65538 , n386270 , n65540 , n386272 , 
 n65542 , n386274 , n386275 , n386276 , n386277 , n386278 , n386279 , n386280 , n386281 , n65551 , 
 n65552 , n65553 , n386285 , n386286 , n65556 , n386288 , n386289 , n386290 , n386291 , n386292 , 
 n386293 , n386294 , n386295 , n386296 , n386297 , n386298 , n386299 , n386300 , n386301 , n386302 , 
 n386303 , n386304 , n386305 , n386306 , n386307 , n386308 , n386309 , n65557 , n386311 , n386312 , 
 n386313 , n386314 , n386315 , n386316 , n65559 , n386318 , n386319 , n65562 , n386321 , n65564 , 
 n65565 , n386324 , n386325 , n386326 , n386327 , n386328 , n386329 , n65572 , n386331 , n65574 , 
 n65575 , n386334 , n386335 , n65578 , n386337 , n386338 , n386339 , n386340 , n386341 , n386342 , 
 n386343 , n386344 , n386345 , n386346 , n386347 , n65590 , n386349 , n386350 , n386351 , n65594 , 
 n386353 , n386354 , n386355 , n386356 , n386357 , n386358 , n386359 , n386360 , n386361 , n386362 , 
 n386363 , n386364 , n386365 , n386366 , n386367 , n386368 , n386369 , n386370 , n386371 , n386372 , 
 n386373 , n386374 , n386375 , n386376 , n386377 , n386378 , n386379 , n386380 , n386381 , n386382 , 
 n386383 , n65613 , n386385 , n386386 , n386387 , n386388 , n386389 , n386390 , n386391 , n386392 , 
 n65619 , n386394 , n65621 , n65622 , n65623 , n386398 , n65625 , n386400 , n386401 , n386402 , 
 n386403 , n386404 , n386405 , n65632 , n386407 , n386408 , n386409 , n386410 , n386411 , n386412 , 
 n386413 , n386414 , n386415 , n386416 , n65643 , n386418 , n386419 , n65646 , n386421 , n386422 , 
 n386423 , n65650 , n386425 , n386426 , n386427 , n65654 , n386429 , n386430 , n65657 , n65658 , 
 n65659 , n386434 , n386435 , n65662 , n386437 , n386438 , n386439 , n65666 , n386441 , n65668 , 
 n386443 , n65670 , n386445 , n386446 , n386447 , n65674 , n386449 , n386450 , n65677 , n386452 , 
 n386453 , n65680 , n386455 , n386456 , n65683 , n386458 , n386459 , n65686 , n386461 , n386462 , 
 n386463 , n386464 , n386465 , n386466 , n386467 , n65694 , n386469 , n386470 , n65697 , n386472 , 
 n386473 , n386474 , n65701 , n386476 , n386477 , n65704 , n386479 , n386480 , n65707 , n386482 , 
 n65709 , n65710 , n65711 , n386486 , n65713 , n386488 , n65715 , n65716 , n386491 , n65718 , 
 n386493 , n386494 , n65721 , n386496 , n386497 , n65724 , n386499 , n65726 , n386501 , n65728 , 
 n65729 , n386504 , n386505 , n386506 , n386507 , n386508 , n386509 , n386510 , n386511 , n386512 , 
 n386513 , n386514 , n386515 , n386516 , n386517 , n386518 , n386519 , n386520 , n386521 , n386522 , 
 n386523 , n386524 , n386525 , n386526 , n386527 , n386528 , n386529 , n386530 , n386531 , n65738 , 
 n65739 , n386534 , n386535 , n386536 , n65743 , n65744 , n65745 , n386540 , n386541 , n386542 , 
 n386543 , n386544 , n386545 , n386546 , n386547 , n386548 , n386549 , n386550 , n65757 , n386552 , 
 n386553 , n65760 , n386555 , n386556 , n386557 , n386558 , n386559 , n386560 , n386561 , n386562 , 
 n65769 , n65770 , n386565 , n65772 , n386567 , n386568 , n386569 , n386570 , n386571 , n386572 , 
 n386573 , n386574 , n386575 , n386576 , n386577 , n386578 , n386579 , n65773 , n65774 , n386582 , 
 n386583 , n386584 , n386585 , n386586 , n386587 , n65781 , n386589 , n386590 , n386591 , n386592 , 
 n386593 , n65783 , n386595 , n65785 , n386597 , n65787 , n386599 , n65789 , n65790 , n386602 , 
 n386603 , n65793 , n386605 , n386606 , n65796 , n386608 , n386609 , n65799 , n65800 , n386612 , 
 n386613 , n65803 , n386615 , n386616 , n65806 , n386618 , n386619 , n386620 , n65810 , n386622 , 
 n65812 , n65813 , n386625 , n65815 , n386627 , n386628 , n386629 , n386630 , n65820 , n386632 , 
 n386633 , n65823 , n386635 , n386636 , n65826 , n386638 , n386639 , n386640 , n386641 , n386642 , 
 n386643 , n386644 , n65834 , n386646 , n65836 , n386648 , n386649 , n65839 , n386651 , n386652 , 
 n65842 , n386654 , n386655 , n65844 , n386657 , n386658 , n65847 , n65848 , n386661 , n386662 , 
 n386663 , n386664 , n386665 , n386666 , n386667 , n386668 , n386669 , n386670 , n386671 , n386672 , 
 n386673 , n386674 , n386675 , n386676 , n386677 , n386678 , n386679 , n65865 , n65866 , n65867 , 
 n65868 , n65869 , n386685 , n386686 , n65872 , n386688 , n65874 , n65875 , n386691 , n65877 , 
 n386693 , n65879 , n386695 , n65881 , n386697 , n65883 , n386699 , n386700 , n386701 , n386702 , 
 n65888 , n65889 , n65890 , n386706 , n386707 , n386708 , n386709 , n65895 , n386711 , n386712 , 
 n65898 , n386714 , n386715 , n65901 , n65902 , n65903 , n386719 , n65905 , n386721 , n386722 , 
 n65908 , n386724 , n386725 , n386726 , n65912 , n65913 , n386729 , n65915 , n386731 , n386732 , 
 n386733 , n386734 , n386735 , n65921 , n386737 , n386738 , n65924 , n386740 , n386741 , n386742 , 
 n65928 , n386744 , n386745 , n65931 , n386747 , n386748 , n65934 , n386750 , n65936 , n386752 , 
 n65938 , n65939 , n386755 , n65941 , n386757 , n386758 , n65944 , n65945 , n386761 , n386762 , 
 n65948 , n386764 , n65950 , n65951 , n386767 , n65953 , n386769 , n386770 , n65956 , n65957 , 
 n386773 , n65959 , n386775 , n65961 , n386777 , n386778 , n386779 , n386780 , n386781 , n65967 , 
 n65968 , n386784 , n65970 , n386786 , n65972 , n386788 , n65974 , n386790 , n65976 , n65977 , 
 n386793 , n386794 , n65980 , n386796 , n65982 , n386798 , n386799 , n65985 , n386801 , n386802 , 
 n386803 , n65989 , n65990 , n386806 , n386807 , n65993 , n386809 , n386810 , n386811 , n386812 , 
 n65998 , n386814 , n386815 , n66001 , n66002 , n386818 , n386819 , n386820 , n386821 , n386822 , 
 n66008 , n386824 , n66010 , n66011 , n66012 , n66013 , n386829 , n386830 , n386831 , n66017 , 
 n386833 , n386834 , n386835 , n66021 , n386837 , n386838 , n66024 , n386840 , n386841 , n386842 , 
 n386843 , n66029 , n66030 , n66031 , n386847 , n386848 , n386849 , n66035 , n386851 , n386852 , 
 n66038 , n386854 , n66040 , n386856 , n386857 , n386858 , n66044 , n66045 , n386861 , n66047 , 
 n386863 , n386864 , n386865 , n386866 , n386867 , n386868 , n66054 , n386870 , n66056 , n386872 , 
 n386873 , n66059 , n386875 , n386876 , n66062 , n66063 , n66064 , n386880 , n66066 , n66067 , 
 n66068 , n386884 , n66070 , n386886 , n66072 , n386888 , n66074 , n66075 , n66076 , n386892 , 
 n66078 , n386894 , n66080 , n66081 , n386897 , n66083 , n386899 , n386900 , n386901 , n386902 , 
 n386903 , n66089 , n66090 , n386906 , n66092 , n386908 , n66094 , n66095 , n386911 , n66097 , 
 n386913 , n66099 , n386915 , n386916 , n66102 , n386918 , n386919 , n386920 , n386921 , n66107 , 
 n386923 , n386924 , n66110 , n386926 , n386927 , n66113 , n66114 , n66115 , n386931 , n66117 , 
 n386933 , n386934 , n386935 , n386936 , n386937 , n66123 , n66124 , n386940 , n386941 , n386942 , 
 n386943 , n386944 , n66130 , n386946 , n386947 , n386948 , n386949 , n386950 , n66136 , n66137 , 
 n386953 , n386954 , n66140 , n386956 , n386957 , n66143 , n386959 , n66145 , n386961 , n386962 , 
 n386963 , n66149 , n386965 , n386966 , n66152 , n66153 , n386969 , n66155 , n386971 , n66157 , 
 n66158 , n386974 , n386975 , n66161 , n386977 , n386978 , n66164 , n386980 , n66166 , n66167 , 
 n66168 , n66169 , n386985 , n66171 , n66172 , n66173 , n386989 , n66175 , n386991 , n66177 , 
 n386993 , n66179 , n66180 , n386996 , n386997 , n66183 , n386999 , n387000 , n66186 , n387002 , 
 n387003 , n66189 , n387005 , n387006 , n66192 , n387008 , n387009 , n66195 , n387011 , n387012 , 
 n66198 , n387014 , n387015 , n387016 , n66202 , n387018 , n66204 , n387020 , n66206 , n387022 , 
 n387023 , n387024 , n387025 , n387026 , n387027 , n387028 , n387029 , n387030 , n387031 , n387032 , 
 n66218 , n387034 , n387035 , n66221 , n66222 , n387038 , n66224 , n387040 , n387041 , n66227 , 
 n387043 , n66229 , n387045 , n66231 , n66232 , n387048 , n387049 , n66235 , n387051 , n387052 , 
 n66238 , n387054 , n387055 , n66241 , n387057 , n66243 , n66244 , n387060 , n387061 , n66247 , 
 n66248 , n387064 , n66250 , n387066 , n66252 , n387068 , n66254 , n387070 , n387071 , n66257 , 
 n387073 , n387074 , n387075 , n387076 , n387077 , n66263 , n387079 , n387080 , n66266 , n387082 , 
 n387083 , n66269 , n66270 , n387086 , n66272 , n387088 , n387089 , n387090 , n387091 , n387092 , 
 n387093 , n387094 , n387095 , n66281 , n387097 , n387098 , n387099 , n387100 , n66286 , n387102 , 
 n387103 , n66289 , n387105 , n387106 , n66292 , n387108 , n387109 , n387110 , n387111 , n387112 , 
 n387113 , n387114 , n387115 , n387116 , n66302 , n387118 , n387119 , n387120 , n387121 , n387122 , 
 n66308 , n66309 , n387125 , n387126 , n66312 , n387128 , n66314 , n387130 , n387131 , n387132 , 
 n387133 , n387134 , n387135 , n66321 , n387137 , n66323 , n387139 , n387140 , n387141 , n387142 , 
 n66328 , n387144 , n387145 , n387146 , n387147 , n387148 , n387149 , n387150 , n387151 , n387152 , 
 n387153 , n387154 , n66340 , n387156 , n387157 , n66343 , n387159 , n387160 , n66346 , n387162 , 
 n387163 , n66349 , n387165 , n387166 , n387167 , n387168 , n387169 , n66355 , n387171 , n387172 , 
 n387173 , n66359 , n387175 , n387176 , n387177 , n387178 , n387179 , n387180 , n387181 , n387182 , 
 n387183 , n387184 , n387185 , n387186 , n387187 , n387188 , n387189 , n387190 , n387191 , n387192 , 
 n387193 , n66379 , n387195 , n66381 , n387197 , n387198 , n66384 , n387200 , n66386 , n387202 , 
 n387203 , n387204 , n66390 , n387206 , n387207 , n66393 , n387209 , n387210 , n387211 , n66397 , 
 n387213 , n387214 , n387215 , n387216 , n66402 , n66403 , n387219 , n66405 , n387221 , n387222 , 
 n66408 , n387224 , n387225 , n66411 , n387227 , n387228 , n66414 , n387230 , n387231 , n66417 , 
 n387233 , n387234 , n66420 , n66421 , n387237 , n66423 , n387239 , n387240 , n387241 , n387242 , 
 n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n387249 , n387250 , n387251 , n387252 , 
 n387253 , n66439 , n66440 , n66441 , n387257 , n387258 , n387259 , n387260 , n387261 , n387262 , 
 n387263 , n66449 , n387265 , n387266 , n387267 , n387268 , n66454 , n387270 , n66456 , n387272 , 
 n387273 , n66459 , n387275 , n387276 , n387277 , n66463 , n387279 , n387280 , n387281 , n387282 , 
 n387283 , n66469 , n66470 , n387286 , n66472 , n66473 , n387289 , n66475 , n387291 , n387292 , 
 n66478 , n387294 , n387295 , n387296 , n387297 , n387298 , n66484 , n387300 , n387301 , n387302 , 
 n66488 , n387304 , n387305 , n387306 , n387307 , n66493 , n387309 , n387310 , n66496 , n387312 , 
 n387313 , n387314 , n387315 , n66501 , n387317 , n387318 , n66504 , n66505 , n387321 , n387322 , 
 n387323 , n66509 , n387325 , n66511 , n387327 , n387328 , n387329 , n387330 , n66516 , n387332 , 
 n387333 , n387334 , n66520 , n66521 , n387337 , n387338 , n387339 , n387340 , n387341 , n66527 , 
 n66528 , n387344 , n66530 , n66531 , n387347 , n387348 , n387349 , n66535 , n387351 , n387352 , 
 n66538 , n387354 , n387355 , n387356 , n387357 , n387358 , n387359 , n66545 , n66546 , n387362 , 
 n387363 , n66549 , n387365 , n387366 , n66552 , n387368 , n387369 , n387370 , n387371 , n387372 , 
 n66558 , n387374 , n387375 , n66561 , n387377 , n387378 , n387379 , n387380 , n66566 , n387382 , 
 n387383 , n387384 , n387385 , n387386 , n387387 , n66573 , n387389 , n387390 , n66576 , n387392 , 
 n387393 , n387394 , n387395 , n387396 , n387397 , n66583 , n387399 , n387400 , n387401 , n66587 , 
 n387403 , n387404 , n387405 , n66591 , n387407 , n387408 , n387409 , n66595 , n387411 , n66597 , 
 n66598 , n387414 , n66600 , n387416 , n387417 , n66603 , n387419 , n387420 , n387421 , n387422 , 
 n387423 , n66609 , n66610 , n66611 , n387427 , n387428 , n387429 , n387430 , n387431 , n387432 , 
 n387433 , n66619 , n387435 , n387436 , n66622 , n387438 , n387439 , n387440 , n66626 , n387442 , 
 n387443 , n66629 , n387445 , n387446 , n66632 , n66633 , n387449 , n387450 , n66636 , n66637 , 
 n387453 , n387454 , n66640 , n66641 , n66642 , n387458 , n387459 , n66645 , n66646 , n66647 , 
 n387463 , n387464 , n66650 , n387466 , n387467 , n387468 , n66654 , n387470 , n387471 , n387472 , 
 n66658 , n387474 , n66660 , n66661 , n66662 , n387478 , n66664 , n387480 , n387481 , n66667 , 
 n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n387490 , n66676 , n387492 , 
 n66678 , n66679 , n387495 , n66681 , n387497 , n66683 , n66684 , n387500 , n387501 , n66687 , 
 n387503 , n387504 , n66690 , n387506 , n387507 , n387508 , n387509 , n387510 , n387511 , n387512 , 
 n387513 , n387514 , n387515 , n387516 , n387517 , n387518 , n387519 , n387520 , n387521 , n387522 , 
 n66708 , n66709 , n387525 , n387526 , n387527 , n387528 , n66714 , n387530 , n387531 , n387532 , 
 n387533 , n387534 , n387535 , n387536 , n387537 , n387538 , n387539 , n66725 , n387541 , n387542 , 
 n387543 , n66729 , n387545 , n387546 , n387547 , n66733 , n387549 , n387550 , n387551 , n66737 , 
 n66738 , n387554 , n66740 , n387556 , n387557 , n387558 , n66744 , n387560 , n387561 , n66747 , 
 n387563 , n387564 , n387565 , n387566 , n387567 , n387568 , n387569 , n387570 , n387571 , n66757 , 
 n66758 , n66759 , n387575 , n66761 , n387577 , n387578 , n387579 , n387580 , n387581 , n387582 , 
 n66768 , n387584 , n387585 , n387586 , n66772 , n387588 , n387589 , n66775 , n387591 , n387592 , 
 n387593 , n387594 , n387595 , n66781 , n387597 , n387598 , n66784 , n66785 , n387601 , n387602 , 
 n387603 , n387604 , n387605 , n387606 , n387607 , n66793 , n387609 , n387610 , n66796 , n387612 , 
 n66798 , n387614 , n387615 , n66801 , n387617 , n387618 , n387619 , n66805 , n66806 , n387622 , 
 n66808 , n387624 , n387625 , n66811 , n66812 , n387628 , n387629 , n66815 , n66816 , n387632 , 
 n387633 , n387634 , n66820 , n66821 , n387637 , n66823 , n66824 , n66825 , n387641 , n66827 , 
 n387643 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n387651 , n387652 , 
 n66838 , n387654 , n387655 , n387656 , n387657 , n66843 , n387659 , n387660 , n66846 , n387662 , 
 n387663 , n387664 , n387665 , n387666 , n387667 , n387668 , n66854 , n66855 , n387671 , n387672 , 
 n387673 , n387674 , n387675 , n387676 , n387677 , n387678 , n66864 , n387680 , n387681 , n387682 , 
 n66868 , n387684 , n387685 , n66871 , n387687 , n387688 , n387689 , n387690 , n66876 , n387692 , 
 n387693 , n387694 , n66880 , n66881 , n387697 , n387698 , n66884 , n387700 , n387701 , n66887 , 
 n387703 , n387704 , n66890 , n66891 , n387707 , n66893 , n66894 , n387710 , n387711 , n66897 , 
 n66898 , n387714 , n66900 , n66901 , n387717 , n66903 , n387719 , n66905 , n66906 , n387722 , 
 n387723 , n66909 , n387725 , n66911 , n66912 , n66913 , n66914 , n66915 , n387731 , n387732 , 
 n66918 , n387734 , n387735 , n387736 , n387737 , n66923 , n387739 , n387740 , n66926 , n387742 , 
 n387743 , n387744 , n387745 , n387746 , n387747 , n387748 , n387749 , n387750 , n66936 , n66937 , 
 n387753 , n387754 , n66940 , n387756 , n66942 , n66943 , n387759 , n387760 , n66946 , n66947 , 
 n387763 , n66949 , n387765 , n387766 , n387767 , n387768 , n387769 , n66955 , n387771 , n66957 , 
 n387773 , n387774 , n387775 , n387776 , n387777 , n387778 , n387779 , n387780 , n387781 , n66967 , 
 n387783 , n66969 , n66970 , n66971 , n66972 , n66973 , n387789 , n387790 , n66976 , n66977 , 
 n387793 , n387794 , n66980 , n387796 , n387797 , n387798 , n66984 , n387800 , n387801 , n387802 , 
 n387803 , n387804 , n387805 , n387806 , n387807 , n387808 , n66994 , n66995 , n387811 , n66997 , 
 n387813 , n66999 , n387815 , n67001 , n67002 , n387818 , n387819 , n67005 , n387821 , n387822 , 
 n67008 , n387824 , n387825 , n67011 , n387827 , n387828 , n67014 , n387830 , n67016 , n67017 , 
 n67018 , n387834 , n67020 , n387836 , n387837 , n387838 , n387839 , n67025 , n387841 , n387842 , 
 n67028 , n67029 , n67030 , n387846 , n67032 , n67033 , n67034 , n387850 , n387851 , n67037 , 
 n387853 , n67039 , n387855 , n67041 , n387857 , n387858 , n387859 , n387860 , n67046 , n387862 , 
 n387863 , n67049 , n387865 , n387866 , n387867 , n387868 , n387869 , n387870 , n387871 , n387872 , 
 n67058 , n387874 , n387875 , n387876 , n387877 , n387878 , n67064 , n387880 , n387881 , n67067 , 
 n67068 , n387884 , n67070 , n67071 , n387887 , n387888 , n67074 , n67075 , n67076 , n67077 , 
 n387893 , n387894 , n67080 , n387896 , n387897 , n387898 , n387899 , n67085 , n67086 , n387902 , 
 n387903 , n387904 , n67090 , n387906 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , 
 n67098 , n387914 , n387915 , n67101 , n387917 , n67103 , n387919 , n387920 , n67106 , n387922 , 
 n67108 , n67109 , n67110 , n67111 , n387927 , n67113 , n387929 , n67115 , n387931 , n67117 , 
 n387933 , n387934 , n387935 , n387936 , n387937 , n387938 , n387939 , n387940 , n387941 , n387942 , 
 n387943 , n387944 , n387945 , n387946 , n387947 , n387948 , n387949 , n387950 , n67118 , n67119 , 
 n387953 , n387954 , n387955 , n387956 , n387957 , n67125 , n387959 , n387960 , n387961 , n67129 , 
 n67130 , n387964 , n67132 , n387966 , n387967 , n67135 , n387969 , n387970 , n387971 , n387972 , 
 n387973 , n67141 , n387975 , n387976 , n67144 , n387978 , n387979 , n387980 , n67148 , n387982 , 
 n67150 , n387984 , n67152 , n387986 , n387987 , n387988 , n387989 , n387990 , n387991 , n387992 , 
 n387993 , n387994 , n387995 , n67163 , n387997 , n67165 , n67166 , n67167 , n388001 , n388002 , 
 n67170 , n388004 , n67172 , n67173 , n67174 , n388008 , n388009 , n67177 , n67178 , n388012 , 
 n388013 , n67181 , n67182 , n67183 , n388017 , n388018 , n67186 , n388020 , n67188 , n388022 , 
 n388023 , n388024 , n67192 , n67193 , n388027 , n67195 , n67196 , n67197 , n388031 , n388032 , 
 n388033 , n388034 , n67202 , n67203 , n388037 , n67205 , n388039 , n388040 , n67208 , n388042 , 
 n388043 , n67211 , n388045 , n388046 , n67214 , n388048 , n388049 , n388050 , n388051 , n388052 , 
 n388053 , n67221 , n388055 , n388056 , n388057 , n67225 , n388059 , n388060 , n388061 , n67229 , 
 n388063 , n388064 , n388065 , n67233 , n388067 , n388068 , n67236 , n388070 , n67237 , n67238 , 
 n67239 , n388074 , n67241 , n388076 , n67243 , n67244 , n388079 , n388080 , n67247 , n388082 , 
 n388083 , n67250 , n388085 , n388086 , n388087 , n388088 , n388089 , n388090 , n388091 , n388092 , 
 n388093 , n67260 , n388095 , n388096 , n388097 , n67264 , n388099 , n67266 , n67267 , n388102 , 
 n388103 , n388104 , n388105 , n388106 , n388107 , n67274 , n388109 , n67276 , n67277 , n388112 , 
 n67279 , n388114 , n388115 , n67282 , n388117 , n388118 , n388119 , n388120 , n388121 , n67288 , 
 n388123 , n388124 , n388125 , n388126 , n388127 , n388128 , n388129 , n67296 , n67297 , n388132 , 
 n388133 , n67300 , n388135 , n388136 , n67303 , n67304 , n388139 , n67306 , n388141 , n67308 , 
 n67309 , n388144 , n67311 , n67312 , n388147 , n388148 , n388149 , n388150 , n67317 , n388152 , 
 n388153 , n67320 , n67321 , n388156 , n67323 , n388158 , n388159 , n67326 , n388161 , n388162 , 
 n388163 , n67330 , n388165 , n67332 , n388167 , n67334 , n67335 , n388170 , n67337 , n388172 , 
 n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n388181 , n67348 , 
 n388183 , n388184 , n67351 , n388186 , n388187 , n67354 , n388189 , n388190 , n388191 , n388192 , 
 n388193 , n388194 , n388195 , n388196 , n67363 , n388198 , n67365 , n388200 , n67367 , n388202 , 
 n67369 , n388204 , n388205 , n388206 , n388207 , n388208 , n388209 , n388210 , n388211 , n67378 , 
 n388213 , n388214 , n388215 , n67382 , n67383 , n67384 , n67385 , n388220 , n67387 , n388222 , 
 n67389 , n388224 , n388225 , n388226 , n388227 , n388228 , n67395 , n388230 , n388231 , n67398 , 
 n67399 , n388234 , n67401 , n388236 , n388237 , n67404 , n388239 , n67406 , n388241 , n388242 , 
 n67409 , n388244 , n388245 , n67412 , n388247 , n388248 , n388249 , n388250 , n67417 , n67418 , 
 n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , 
 n388263 , n67430 , n67431 , n67432 , n67433 , n388268 , n67435 , n388270 , n388271 , n67438 , 
 n388273 , n388274 , n67441 , n67442 , n388277 , n67444 , n67445 , n388280 , n388281 , n67448 , 
 n67449 , n388284 , n67451 , n67452 , n67453 , n67454 , n388289 , n388290 , n388291 , n388292 , 
 n67459 , n67460 , n388295 , n388296 , n67463 , n388298 , n67465 , n67466 , n388301 , n388302 , 
 n67469 , n388304 , n388305 , n388306 , n388307 , n388308 , n67475 , n388310 , n67477 , n67478 , 
 n67479 , n67480 , n388315 , n388316 , n388317 , n388318 , n388319 , n67486 , n388321 , n388322 , 
 n67489 , n388324 , n388325 , n67492 , n67493 , n388328 , n388329 , n388330 , n388331 , n67498 , 
 n67499 , n388334 , n388335 , n388336 , n388337 , n388338 , n388339 , n388340 , n67507 , n388342 , 
 n67509 , n388344 , n67511 , n388346 , n388347 , n388348 , n67515 , n388350 , n388351 , n388352 , 
 n388353 , n388354 , n388355 , n67522 , n388357 , n388358 , n388359 , n67526 , n67527 , n67528 , 
 n67529 , n67530 , n67531 , n67532 , n388367 , n388368 , n388369 , n67536 , n388371 , n388372 , 
 n67539 , n388374 , n388375 , n67542 , n388377 , n388378 , n67545 , n67546 , n67547 , n388382 , 
 n388383 , n67550 , n67551 , n67552 , n388387 , n388388 , n388389 , n388390 , n388391 , n388392 , 
 n388393 , n67560 , n388395 , n388396 , n67563 , n388398 , n67565 , n67566 , n388401 , n67568 , 
 n388403 , n67570 , n388405 , n388406 , n388407 , n388408 , n388409 , n67576 , n388411 , n388412 , 
 n388413 , n388414 , n388415 , n388416 , n388417 , n388418 , n388419 , n388420 , n388421 , n388422 , 
 n388423 , n388424 , n388425 , n388426 , n388427 , n388428 , n67581 , n388430 , n388431 , n67584 , 
 n67585 , n67586 , n388435 , n67588 , n388437 , n67590 , n388439 , n388440 , n388441 , n388442 , 
 n388443 , n388444 , n388445 , n388446 , n388447 , n388448 , n388449 , n388450 , n67603 , n388452 , 
 n388453 , n67606 , n388455 , n67608 , n67609 , n388458 , n388459 , n67612 , n388461 , n388462 , 
 n388463 , n388464 , n388465 , n388466 , n67619 , n388468 , n388469 , n67622 , n388471 , n67624 , 
 n67625 , n67626 , n388475 , n388476 , n388477 , n388478 , n67631 , n388480 , n388481 , n388482 , 
 n67635 , n388484 , n388485 , n67638 , n388487 , n388488 , n67641 , n388490 , n67643 , n67644 , 
 n388493 , n67646 , n388495 , n388496 , n67649 , n67650 , n388499 , n388500 , n388501 , n388502 , 
 n388503 , n67656 , n67657 , n67658 , n67659 , n388508 , n388509 , n67662 , n388511 , n388512 , 
 n67665 , n388514 , n388515 , n67668 , n67669 , n388518 , n67671 , n388520 , n388521 , n67674 , 
 n67675 , n388524 , n67677 , n388526 , n388527 , n388528 , n388529 , n388530 , n388531 , n388532 , 
 n388533 , n67686 , n388535 , n388536 , n67689 , n388538 , n67691 , n67692 , n388541 , n388542 , 
 n388543 , n388544 , n388545 , n67698 , n388547 , n67700 , n67701 , n67702 , n388551 , n67704 , 
 n388553 , n67706 , n388555 , n388556 , n388557 , n388558 , n388559 , n388560 , n388561 , n388562 , 
 n388563 , n67716 , n67717 , n388566 , n67719 , n388568 , n67721 , n67722 , n67723 , n67724 , 
 n67725 , n388574 , n67727 , n388576 , n388577 , n388578 , n388579 , n67732 , n388581 , n388582 , 
 n388583 , n388584 , n388585 , n388586 , n388587 , n388588 , n388589 , n388590 , n388591 , n388592 , 
 n388593 , n67746 , n67747 , n388596 , n388597 , n67750 , n67751 , n388600 , n388601 , n67754 , 
 n388603 , n67756 , n388605 , n388606 , n388607 , n67759 , n388609 , n388610 , n67762 , n388612 , 
 n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n388621 , n388622 , 
 n67774 , n388624 , n388625 , n67777 , n67778 , n388628 , n67780 , n67781 , n67782 , n67783 , 
 n67784 , n67785 , n67786 , n67787 , n388637 , n388638 , n388639 , n388640 , n67792 , n388642 , 
 n67794 , n388644 , n388645 , n388646 , n388647 , n67799 , n388649 , n388650 , n67802 , n67803 , 
 n67804 , n388654 , n388655 , n388656 , n388657 , n388658 , n388659 , n388660 , n388661 , n388662 , 
 n388663 , n388664 , n388665 , n388666 , n388667 , n388668 , n388669 , n388670 , n388671 , n388672 , 
 n388673 , n388674 , n388675 , n388676 , n388677 , n388678 , n388679 , n388680 , n388681 , n67808 , 
 n388683 , n388684 , n388685 , n388686 , n67810 , n388688 , n388689 , n388690 , n388691 , n388692 , 
 n388693 , n388694 , n388695 , n388696 , n388697 , n388698 , n388699 , n388700 , n388701 , n388702 , 
 n388703 , n388704 , n388705 , n388706 , n388707 , n388708 , n388709 , n67814 , n388711 , n67816 , 
 n388713 , n67818 , n388715 , n67820 , n388717 , n67822 , n67823 , n388720 , n388721 , n388722 , 
 n388723 , n388724 , n67829 , n388726 , n388727 , n388728 , n388729 , n388730 , n388731 , n67836 , 
 n388733 , n388734 , n67839 , n388736 , n388737 , n67842 , n388739 , n67843 , n388741 , n67845 , 
 n67846 , n388744 , n67848 , n67849 , n67850 , n388748 , n67852 , n67853 , n67854 , n388752 , 
 n388753 , n67857 , n388755 , n388756 , n67860 , n388758 , n67862 , n388760 , n67864 , n388762 , 
 n67866 , n388764 , n67868 , n388766 , n388767 , n67871 , n67872 , n67873 , n67874 , n67875 , 
 n67876 , n388774 , n67878 , n388776 , n67880 , n388778 , n388779 , n388780 , n67884 , n388782 , 
 n67886 , n67887 , n67888 , n67889 , n388787 , n67891 , n388789 , n388790 , n67894 , n388792 , 
 n67896 , n388794 , n67898 , n388796 , n388797 , n388798 , n67902 , n388800 , n388801 , n388802 , 
 n67906 , n67907 , n388805 , n67909 , n388807 , n388808 , n67912 , n388810 , n388811 , n67915 , 
 n67916 , n67917 , n67918 , n67919 , n67920 , n388818 , n388819 , n388820 , n67924 , n388822 , 
 n388823 , n67927 , n388825 , n388826 , n388827 , n388828 , n67932 , n388830 , n67934 , n388832 , 
 n388833 , n67937 , n67938 , n67939 , n388837 , n67941 , n388839 , n388840 , n67944 , n67945 , 
 n67946 , n388844 , n388845 , n388846 , n67950 , n388848 , n388849 , n388850 , n388851 , n388852 , 
 n388853 , n388854 , n388855 , n388856 , n388857 , n388858 , n388859 , n388860 , n388861 , n388862 , 
 n388863 , n388864 , n388865 , n388866 , n388867 , n388868 , n388869 , n67954 , n388871 , n67956 , 
 n67957 , n388874 , n388875 , n388876 , n67961 , n388878 , n388879 , n67964 , n67965 , n67966 , 
 n67967 , n67968 , n388885 , n388886 , n67971 , n388888 , n67973 , n67974 , n67975 , n388892 , 
 n388893 , n388894 , n388895 , n67980 , n388897 , n388898 , n67983 , n388900 , n388901 , n67986 , 
 n67987 , n388904 , n388905 , n388906 , n67991 , n67992 , n67993 , n67994 , n67995 , n67996 , 
 n67997 , n67998 , n67999 , n68000 , n388917 , n68002 , n388919 , n388920 , n68005 , n388922 , 
 n388923 , n68008 , n388925 , n388926 , n68011 , n388928 , n388929 , n68014 , n388931 , n388932 , 
 n68017 , n388934 , n388935 , n68020 , n68021 , n388938 , n388939 , n388940 , n388941 , n68026 , 
 n388943 , n388944 , n388945 , n68030 , n388947 , n388948 , n388949 , n388950 , n388951 , n388952 , 
 n68037 , n388954 , n388955 , n388956 , n388957 , n388958 , n388959 , n388960 , n388961 , n388962 , 
 n388963 , n68048 , n388965 , n68050 , n388967 , n388968 , n68053 , n388970 , n388971 , n68056 , 
 n388973 , n68058 , n388975 , n68060 , n388977 , n68062 , n68063 , n388980 , n388981 , n68066 , 
 n388983 , n388984 , n68069 , n388986 , n388987 , n68072 , n388989 , n388990 , n388991 , n388992 , 
 n388993 , n388994 , n388995 , n388996 , n388997 , n388998 , n388999 , n389000 , n68085 , n389002 , 
 n389003 , n389004 , n68089 , n389006 , n389007 , n389008 , n389009 , n389010 , n389011 , n68096 , 
 n389013 , n389014 , n389015 , n389016 , n389017 , n389018 , n389019 , n389020 , n389021 , n389022 , 
 n389023 , n389024 , n389025 , n389026 , n389027 , n389028 , n389029 , n389030 , n389031 , n389032 , 
 n389033 , n389034 , n389035 , n68120 , n68121 , n68122 , n389039 , n68124 , n389041 , n68126 , 
 n389043 , n68128 , n389045 , n389046 , n68131 , n389048 , n68133 , n389050 , n389051 , n389052 , 
 n389053 , n389054 , n389055 , n389056 , n68141 , n389058 , n68143 , n68144 , n389061 , n389062 , 
 n68147 , n389064 , n68149 , n68150 , n389067 , n68152 , n389069 , n389070 , n389071 , n389072 , 
 n68157 , n389074 , n389075 , n389076 , n68161 , n389078 , n68163 , n389080 , n389081 , n68166 , 
 n389083 , n389084 , n389085 , n389086 , n389087 , n389088 , n68173 , n389090 , n389091 , n389092 , 
 n389093 , n389094 , n389095 , n389096 , n389097 , n389098 , n389099 , n389100 , n68185 , n68186 , 
 n389103 , n389104 , n68189 , n389106 , n389107 , n389108 , n389109 , n389110 , n389111 , n389112 , 
 n389113 , n389114 , n389115 , n68200 , n68201 , n389118 , n389119 , n389120 , n68205 , n68206 , 
 n68207 , n389124 , n68209 , n389126 , n68211 , n68212 , n68213 , n68214 , n68215 , n68216 , 
 n68217 , n389134 , n68219 , n389136 , n389137 , n389138 , n68223 , n389140 , n389141 , n389142 , 
 n68227 , n389144 , n389145 , n389146 , n68231 , n389148 , n389149 , n68234 , n68235 , n389152 , 
 n389153 , n389154 , n389155 , n389156 , n68241 , n389158 , n389159 , n389160 , n389161 , n68246 , 
 n389163 , n389164 , n68249 , n389166 , n389167 , n389168 , n389169 , n389170 , n68255 , n389172 , 
 n389173 , n389174 , n389175 , n389176 , n68261 , n389178 , n389179 , n68264 , n389181 , n389182 , 
 n389183 , n68268 , n389185 , n389186 , n389187 , n389188 , n68273 , n389190 , n389191 , n68276 , 
 n68277 , n389194 , n68279 , n68280 , n68281 , n68282 , n68283 , n389200 , n68285 , n389202 , 
 n68287 , n389204 , n389205 , n68290 , n68291 , n389208 , n389209 , n68294 , n389211 , n389212 , 
 n68297 , n389214 , n389215 , n389216 , n68301 , n389218 , n389219 , n389220 , n389221 , n389222 , 
 n389223 , n68308 , n68309 , n389226 , n389227 , n389228 , n389229 , n389230 , n389231 , n389232 , 
 n389233 , n389234 , n389235 , n389236 , n389237 , n68322 , n389239 , n389240 , n389241 , n68326 , 
 n389243 , n389244 , n68329 , n389246 , n389247 , n68332 , n389249 , n389250 , n68335 , n389252 , 
 n389253 , n389254 , n389255 , n389256 , n389257 , n389258 , n389259 , n68344 , n68345 , n389262 , 
 n389263 , n389264 , n68349 , n389266 , n389267 , n389268 , n68353 , n389270 , n389271 , n389272 , 
 n389273 , n389274 , n389275 , n389276 , n389277 , n389278 , n389279 , n389280 , n389281 , n389282 , 
 n68367 , n389284 , n389285 , n389286 , n389287 , n68372 , n389289 , n389290 , n68375 , n389292 , 
 n389293 , n68378 , n68379 , n389296 , n389297 , n68382 , n389299 , n389300 , n389301 , n68386 , 
 n68387 , n389304 , n389305 , n68390 , n68391 , n68392 , n389309 , n389310 , n68395 , n389312 , 
 n68397 , n389314 , n389315 , n68400 , n389317 , n68402 , n389319 , n389320 , n389321 , n68406 , 
 n389323 , n389324 , n68409 , n389326 , n389327 , n389328 , n68413 , n389330 , n389331 , n68416 , 
 n389333 , n389334 , n68419 , n389336 , n389337 , n389338 , n389339 , n68424 , n389341 , n389342 , 
 n68427 , n389344 , n389345 , n389346 , n389347 , n389348 , n389349 , n389350 , n389351 , n389352 , 
 n68437 , n389354 , n68439 , n68440 , n389357 , n389358 , n389359 , n389360 , n389361 , n68446 , 
 n389363 , n389364 , n389365 , n68450 , n389367 , n389368 , n389369 , n68454 , n389371 , n389372 , 
 n68457 , n389374 , n389375 , n389376 , n68461 , n389378 , n68463 , n389380 , n68465 , n68466 , 
 n389383 , n389384 , n389385 , n389386 , n68471 , n389388 , n389389 , n68474 , n68475 , n389392 , 
 n389393 , n389394 , n68479 , n389396 , n389397 , n68482 , n68483 , n389400 , n389401 , n68486 , 
 n389403 , n68488 , n389405 , n68490 , n68491 , n389408 , n389409 , n68494 , n389411 , n389412 , 
 n68497 , n68498 , n389415 , n389416 , n389417 , n68502 , n68503 , n389420 , n389421 , n68506 , 
 n68507 , n68508 , n389425 , n389426 , n68511 , n68512 , n68513 , n389430 , n389431 , n68516 , 
 n68517 , n68518 , n389435 , n389436 , n68521 , n389438 , n389439 , n389440 , n389441 , n389442 , 
 n68527 , n389444 , n389445 , n389446 , n68531 , n389448 , n68533 , n68534 , n389451 , n68536 , 
 n68537 , n68538 , n68539 , n68540 , n68541 , n68542 , n68543 , n389460 , n68545 , n68546 , 
 n389463 , n389464 , n68549 , n389466 , n68551 , n389468 , n68553 , n68554 , n68555 , n389472 , 
 n389473 , n389474 , n68559 , n389476 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , 
 n68567 , n68568 , n68569 , n68570 , n68571 , n68572 , n68573 , n68574 , n389491 , n68576 , 
 n68577 , n68578 , n68579 , n68580 , n68581 , n68582 , n68583 , n68584 , n389501 , n68586 , 
 n68587 , n68588 , n68589 , n68590 , n68591 , n389508 , n68593 , n389510 , n389511 , n389512 , 
 n389513 , n68598 , n389515 , n389516 , n389517 , n389518 , n389519 , n389520 , n389521 , n389522 , 
 n389523 , n68608 , n68609 , n68610 , n389527 , n68612 , n68613 , n389530 , n68615 , n389532 , 
 n68617 , n68618 , n68619 , n68620 , n389537 , n68622 , n389539 , n68624 , n389541 , n389542 , 
 n389543 , n68628 , n68629 , n389546 , n389547 , n68632 , n389549 , n389550 , n389551 , n389552 , 
 n68637 , n389554 , n68639 , n68640 , n389557 , n68642 , n68643 , n68644 , n68645 , n68646 , 
 n68647 , n68648 , n389565 , n68650 , n389567 , n389568 , n68653 , n389570 , n68655 , n389572 , 
 n389573 , n68658 , n389575 , n389576 , n389577 , n68662 , n389579 , n68664 , n68665 , n68666 , 
 n389583 , n389584 , n389585 , n389586 , n68671 , n389588 , n389589 , n389590 , n389591 , n68676 , 
 n389593 , n389594 , n389595 , n389596 , n389597 , n389598 , n68683 , n389600 , n389601 , n389602 , 
 n389603 , n68688 , n389605 , n68690 , n389607 , n68692 , n389609 , n389610 , n389611 , n389612 , 
 n389613 , n389614 , n389615 , n389616 , n389617 , n68702 , n389619 , n389620 , n68705 , n389622 , 
 n389623 , n68708 , n389625 , n389626 , n389627 , n389628 , n389629 , n389630 , n389631 , n389632 , 
 n68717 , n68718 , n68719 , n389636 , n389637 , n389638 , n389639 , n68724 , n68725 , n68726 , 
 n389643 , n68728 , n68729 , n389646 , n389647 , n389648 , n389649 , n389650 , n389651 , n389652 , 
 n68737 , n389654 , n68739 , n68740 , n389657 , n389658 , n389659 , n68744 , n389661 , n389662 , 
 n389663 , n389664 , n68745 , n389666 , n389667 , n389668 , n389669 , n389670 , n68750 , n389672 , 
 n389673 , n389674 , n389675 , n389676 , n389677 , n389678 , n68758 , n389680 , n389681 , n389682 , 
 n68762 , n389684 , n68764 , n68765 , n68766 , n68767 , n389689 , n68769 , n389691 , n389692 , 
 n68772 , n389694 , n389695 , n389696 , n389697 , n68777 , n68778 , n68779 , n68780 , n68781 , 
 n68782 , n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n389710 , n389711 , n68791 , 
 n389713 , n389714 , n68794 , n389716 , n389717 , n68797 , n389719 , n389720 , n68800 , n68801 , 
 n68802 , n389724 , n389725 , n389726 , n389727 , n389728 , n68808 , n389730 , n389731 , n68811 , 
 n389733 , n68813 , n389735 , n68815 , n389737 , n389738 , n389739 , n389740 , n389741 , n389742 , 
 n389743 , n68823 , n389745 , n389746 , n68826 , n68827 , n389749 , n389750 , n68830 , n389752 , 
 n68832 , n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , 
 n68842 , n68843 , n68844 , n389766 , n389767 , n389768 , n389769 , n389770 , n389771 , n389772 , 
 n68852 , n389774 , n389775 , n68855 , n389777 , n389778 , n389779 , n389780 , n389781 , n68861 , 
 n389783 , n68863 , n68864 , n68865 , n68866 , n389788 , n389789 , n68869 , n389791 , n389792 , 
 n68872 , n389794 , n389795 , n68875 , n389797 , n389798 , n68878 , n389800 , n68880 , n389802 , 
 n68882 , n389804 , n389805 , n68885 , n389807 , n389808 , n389809 , n389810 , n389811 , n389812 , 
 n389813 , n389814 , n389815 , n389816 , n68896 , n389818 , n389819 , n389820 , n389821 , n389822 , 
 n389823 , n68903 , n389825 , n389826 , n68906 , n389828 , n389829 , n68909 , n389831 , n68911 , 
 n68912 , n389834 , n389835 , n389836 , n389837 , n389838 , n68918 , n389840 , n389841 , n68921 , 
 n389843 , n389844 , n68924 , n389846 , n68926 , n68927 , n68928 , n68929 , n68930 , n389852 , 
 n389853 , n68933 , n389855 , n389856 , n68936 , n389858 , n68938 , n68939 , n68940 , n68941 , 
 n68942 , n68943 , n389865 , n68945 , n389867 , n68947 , n389869 , n68949 , n68950 , n68951 , 
 n68952 , n68953 , n68954 , n389876 , n389877 , n389878 , n68958 , n389880 , n389881 , n389882 , 
 n389883 , n389884 , n389885 , n389886 , n389887 , n389888 , n389889 , n68969 , n389891 , n389892 , 
 n68972 , n389894 , n389895 , n68975 , n389897 , n68977 , n389899 , n389900 , n389901 , n68981 , 
 n389903 , n389904 , n68984 , n68985 , n389907 , n68987 , n389909 , n389910 , n68990 , n389912 , 
 n389913 , n389914 , n68994 , n389916 , n389917 , n389918 , n68998 , n389920 , n389921 , n69001 , 
 n389923 , n69003 , n389925 , n69005 , n389927 , n389928 , n389929 , n389930 , n389931 , n69011 , 
 n69012 , n389934 , n389935 , n389936 , n389937 , n389938 , n389939 , n389940 , n389941 , n389942 , 
 n389943 , n389944 , n389945 , n389946 , n69026 , n69027 , n389949 , n389950 , n389951 , n69031 , 
 n389953 , n389954 , n389955 , n389956 , n69036 , n389958 , n389959 , n69039 , n389961 , n69041 , 
 n389963 , n389964 , n69044 , n69045 , n389967 , n69047 , n69048 , n389970 , n69050 , n389972 , 
 n389973 , n69053 , n389975 , n389976 , n69056 , n389978 , n69058 , n69059 , n389981 , n389982 , 
 n389983 , n389984 , n69064 , n389986 , n69066 , n389988 , n389989 , n69069 , n389991 , n69071 , 
 n389993 , n69073 , n389995 , n389996 , n69076 , n389998 , n389999 , n390000 , n69080 , n390002 , 
 n390003 , n390004 , n390005 , n390006 , n390007 , n69087 , n390009 , n390010 , n69090 , n69091 , 
 n390013 , n69093 , n390015 , n390016 , n69096 , n390018 , n69098 , n69099 , n390021 , n390022 , 
 n390023 , n69103 , n69104 , n390026 , n390027 , n69107 , n390029 , n390030 , n390031 , n390032 , 
 n69112 , n69113 , n69114 , n69115 , n69116 , n390038 , n390039 , n69119 , n390041 , n390042 , 
 n390043 , n390044 , n69124 , n390046 , n390047 , n390048 , n390049 , n69129 , n390051 , n69131 , 
 n69132 , n390054 , n390055 , n69135 , n390057 , n390058 , n390059 , n390060 , n390061 , n69141 , 
 n69142 , n390064 , n390065 , n69145 , n390067 , n390068 , n69148 , n390070 , n390071 , n69151 , 
 n390073 , n390074 , n69154 , n390076 , n390077 , n390078 , n390079 , n390080 , n390081 , n390082 , 
 n390083 , n69163 , n69164 , n69165 , n69166 , n69167 , n390089 , n69169 , n390091 , n69171 , 
 n390093 , n69173 , n390095 , n69175 , n390097 , n69177 , n69178 , n390100 , n390101 , n390102 , 
 n69182 , n390104 , n390105 , n390106 , n390107 , n390108 , n390109 , n390110 , n69190 , n390112 , 
 n390113 , n69193 , n69194 , n390116 , n69196 , n390118 , n69198 , n390120 , n69200 , n390122 , 
 n390123 , n69203 , n390125 , n390126 , n390127 , n390128 , n390129 , n69209 , n69210 , n390132 , 
 n390133 , n390134 , n69214 , n69215 , n69216 , n69217 , n69218 , n390140 , n390141 , n390142 , 
 n390143 , n390144 , n69224 , n390146 , n69226 , n390148 , n390149 , n390150 , n390151 , n390152 , 
 n69232 , n390154 , n390155 , n69235 , n390157 , n390158 , n69238 , n390160 , n390161 , n390162 , 
 n390163 , n390164 , n69244 , n390166 , n69246 , n390168 , n390169 , n69249 , n390171 , n69251 , 
 n390173 , n390174 , n69254 , n390176 , n390177 , n69257 , n390179 , n69259 , n390181 , n69261 , 
 n390183 , n69263 , n69264 , n390186 , n390187 , n390188 , n69268 , n390190 , n390191 , n390192 , 
 n69272 , n69273 , n390195 , n69275 , n390197 , n390198 , n390199 , n390200 , n69280 , n69281 , 
 n390203 , n390204 , n390205 , n390206 , n69286 , n390208 , n390209 , n69289 , n390211 , n390212 , 
 n69292 , n69293 , n69294 , n390216 , n390217 , n390218 , n69298 , n390220 , n390221 , n69301 , 
 n69302 , n390224 , n390225 , n390226 , n69306 , n390228 , n390229 , n69309 , n69310 , n390232 , 
 n390233 , n69313 , n69314 , n390236 , n69316 , n390238 , n390239 , n390240 , n390241 , n390242 , 
 n390243 , n390244 , n390245 , n390246 , n390247 , n390248 , n390249 , n390250 , n390251 , n69331 , 
 n390253 , n69333 , n390255 , n390256 , n390257 , n390258 , n390259 , n390260 , n69340 , n390262 , 
 n390263 , n390264 , n69344 , n69345 , n390267 , n390268 , n390269 , n69349 , n390271 , n390272 , 
 n69352 , n390274 , n390275 , n390276 , n390277 , n390278 , n390279 , n69359 , n390281 , n390282 , 
 n390283 , n390284 , n69364 , n390286 , n390287 , n390288 , n390289 , n69366 , n390291 , n69368 , 
 n390293 , n390294 , n390295 , n390296 , n390297 , n390298 , n390299 , n390300 , n390301 , n390302 , 
 n390303 , n390304 , n390305 , n390306 , n390307 , n390308 , n390309 , n390310 , n390311 , n390312 , 
 n390313 , n390314 , n390315 , n390316 , n390317 , n390318 , n390319 , n69373 , n390321 , n69375 , 
 n390323 , n390324 , n69378 , n390326 , n390327 , n69381 , n390329 , n390330 , n390331 , n390332 , 
 n390333 , n390334 , n390335 , n69389 , n390337 , n390338 , n390339 , n390340 , n390341 , n390342 , 
 n69396 , n69397 , n390345 , n390346 , n69400 , n390348 , n390349 , n69403 , n390351 , n390352 , 
 n69406 , n390354 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , 
 n69416 , n390364 , n69418 , n390366 , n390367 , n390368 , n390369 , n390370 , n390371 , n390372 , 
 n390373 , n390374 , n390375 , n390376 , n69430 , n390378 , n390379 , n69433 , n390381 , n390382 , 
 n69436 , n390384 , n390385 , n69439 , n390387 , n390388 , n390389 , n390390 , n390391 , n390392 , 
 n390393 , n69447 , n390395 , n390396 , n69450 , n390398 , n390399 , n69453 , n390401 , n69455 , 
 n390403 , n69457 , n69458 , n390406 , n390407 , n69461 , n69462 , n390410 , n69464 , n390412 , 
 n390413 , n390414 , n390415 , n390416 , n390417 , n69471 , n69472 , n390420 , n390421 , n69475 , 
 n390423 , n69477 , n390425 , n390426 , n69480 , n390428 , n69482 , n69483 , n69484 , n69485 , 
 n69486 , n69487 , n69488 , n69489 , n390437 , n390438 , n390439 , n390440 , n69494 , n390442 , 
 n390443 , n69497 , n390445 , n390446 , n69500 , n390448 , n390449 , n390450 , n390451 , n390452 , 
 n69506 , n69507 , n69508 , n69509 , n69510 , n390458 , n390459 , n390460 , n69514 , n390462 , 
 n390463 , n69517 , n390465 , n390466 , n390467 , n390468 , n390469 , n69523 , n390471 , n390472 , 
 n69526 , n390474 , n390475 , n69529 , n69530 , n390478 , n390479 , n390480 , n390481 , n390482 , 
 n390483 , n390484 , n390485 , n69538 , n390487 , n69540 , n390489 , n390490 , n69543 , n69544 , 
 n390493 , n69546 , n69547 , n390496 , n390497 , n69550 , n390499 , n390500 , n390501 , n390502 , 
 n390503 , n390504 , n390505 , n69558 , n390507 , n390508 , n69561 , n390510 , n69563 , n69564 , 
 n69565 , n69566 , n69567 , n69568 , n390517 , n390518 , n69571 , n390520 , n390521 , n390522 , 
 n390523 , n69576 , n390525 , n390526 , n69579 , n390528 , n390529 , n390530 , n390531 , n69584 , 
 n390533 , n69586 , n390535 , n390536 , n390537 , n390538 , n390539 , n390540 , n390541 , n69594 , 
 n390543 , n390544 , n69597 , n390546 , n390547 , n69600 , n390549 , n390550 , n390551 , n390552 , 
 n390553 , n390554 , n390555 , n69608 , n390557 , n390558 , n390559 , n390560 , n390561 , n69614 , 
 n390563 , n69616 , n390565 , n390566 , n69619 , n390568 , n390569 , n69622 , n390571 , n390572 , 
 n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n390579 , n69632 , n390581 , n69634 , 
 n69635 , n69636 , n390585 , n390586 , n390587 , n69640 , n69641 , n69642 , n69643 , n390592 , 
 n390593 , n390594 , n390595 , n390596 , n69649 , n390598 , n69651 , n390600 , n390601 , n69654 , 
 n390603 , n390604 , n390605 , n390606 , n69659 , n390608 , n69661 , n390610 , n69663 , n69664 , 
 n390613 , n390614 , n69667 , n390616 , n390617 , n69670 , n390619 , n390620 , n69673 , n390622 , 
 n69675 , n69676 , n390625 , n390626 , n69679 , n390628 , n390629 , n390630 , n390631 , n390632 , 
 n390633 , n69686 , n390635 , n390636 , n390637 , n390638 , n390639 , n390640 , n390641 , n390642 , 
 n390643 , n390644 , n390645 , n390646 , n390647 , n69700 , n390649 , n390650 , n390651 , n69704 , 
 n390653 , n390654 , n69707 , n390656 , n390657 , n69710 , n390659 , n390660 , n69713 , n390662 , 
 n390663 , n390664 , n390665 , n390666 , n69719 , n390668 , n390669 , n69722 , n390671 , n390672 , 
 n69725 , n390674 , n390675 , n69728 , n390677 , n69730 , n390679 , n390680 , n390681 , n69734 , 
 n390683 , n390684 , n69737 , n390686 , n390687 , n390688 , n390689 , n390690 , n390691 , n69744 , 
 n390693 , n390694 , n69747 , n390696 , n390697 , n69750 , n390699 , n390700 , n69753 , n390702 , 
 n69755 , n390704 , n390705 , n390706 , n390707 , n390708 , n390709 , n390710 , n390711 , n69764 , 
 n390713 , n69766 , n69767 , n390716 , n390717 , n69770 , n390719 , n390720 , n69773 , n390722 , 
 n69775 , n390724 , n69777 , n390726 , n390727 , n390728 , n390729 , n390730 , n69783 , n69784 , 
 n390733 , n390734 , n390735 , n390736 , n390737 , n390738 , n390739 , n390740 , n390741 , n390742 , 
 n69795 , n390744 , n390745 , n390746 , n390747 , n390748 , n69801 , n390750 , n69803 , n390752 , 
 n390753 , n390754 , n69807 , n390756 , n390757 , n69810 , n390759 , n390760 , n69813 , n390762 , 
 n390763 , n69816 , n390765 , n390766 , n69819 , n69820 , n390769 , n69822 , n390771 , n390772 , 
 n69825 , n390774 , n69827 , n390776 , n390777 , n69830 , n390779 , n390780 , n390781 , n390782 , 
 n69835 , n390784 , n390785 , n69838 , n390787 , n69840 , n69841 , n390790 , n390791 , n69844 , 
 n390793 , n69846 , n69847 , n390796 , n390797 , n69850 , n390799 , n390800 , n69853 , n390802 , 
 n390803 , n69856 , n390805 , n69858 , n69859 , n390808 , n390809 , n390810 , n390811 , n390812 , 
 n69865 , n390814 , n390815 , n390816 , n390817 , n390818 , n390819 , n390820 , n69873 , n390822 , 
 n390823 , n390824 , n390825 , n390826 , n69879 , n390828 , n390829 , n390830 , n390831 , n390832 , 
 n390833 , n390834 , n390835 , n390836 , n390837 , n390838 , n390839 , n390840 , n390841 , n69894 , 
 n69895 , n69896 , n390845 , n390846 , n69899 , n390848 , n390849 , n69902 , n390851 , n390852 , 
 n390853 , n390854 , n390855 , n69908 , n390857 , n390858 , n69911 , n69912 , n390861 , n69914 , 
 n69915 , n69916 , n390865 , n69918 , n69919 , n69920 , n390869 , n390870 , n69923 , n390872 , 
 n69925 , n69926 , n69927 , n390876 , n69929 , n69930 , n390879 , n390880 , n69933 , n69934 , 
 n390883 , n390884 , n69937 , n390886 , n390887 , n69940 , n69941 , n69942 , n390891 , n390892 , 
 n69945 , n69946 , n390895 , n69948 , n69949 , n390898 , n390899 , n69952 , n390901 , n390902 , 
 n390903 , n69956 , n390905 , n390906 , n390907 , n390908 , n69961 , n69962 , n390911 , n390912 , 
 n390913 , n69966 , n69967 , n69968 , n390917 , n390918 , n390919 , n390920 , n69973 , n390922 , 
 n390923 , n390924 , n69977 , n390926 , n390927 , n390928 , n390929 , n69982 , n390931 , n390932 , 
 n69985 , n390934 , n69987 , n390936 , n69989 , n69990 , n390939 , n390940 , n390941 , n390942 , 
 n390943 , n390944 , n390945 , n390946 , n390947 , n390948 , n390949 , n390950 , n390951 , n390952 , 
 n390953 , n390954 , n390955 , n390956 , n390957 , n390958 , n390959 , n390960 , n390961 , n390962 , 
 n390963 , n390964 , n390965 , n390966 , n390967 , n390968 , n390969 , n390970 , n390971 , n390972 , 
 n390973 , n390974 , n390975 , n390976 , n390977 , n390978 , n390979 , n69997 , n390981 , n69999 , 
 n70000 , n390984 , n390985 , n70003 , n70004 , n390988 , n70006 , n70007 , n390991 , n70009 , 
 n390993 , n70011 , n70012 , n390996 , n390997 , n70015 , n390999 , n391000 , n391001 , n391002 , 
 n391003 , n391004 , n391005 , n391006 , n391007 , n391008 , n391009 , n391010 , n391011 , n391012 , 
 n70030 , n391014 , n391015 , n70033 , n70034 , n391018 , n70036 , n70037 , n391021 , n391022 , 
 n391023 , n70041 , n391025 , n70043 , n391027 , n391028 , n391029 , n391030 , n391031 , n70049 , 
 n391033 , n391034 , n70052 , n391036 , n391037 , n391038 , n391039 , n391040 , n70058 , n391042 , 
 n391043 , n391044 , n70062 , n391046 , n391047 , n70065 , n391049 , n391050 , n70068 , n391052 , 
 n70070 , n391054 , n391055 , n391056 , n70074 , n391058 , n391059 , n70077 , n391061 , n391062 , 
 n70080 , n391064 , n70082 , n70083 , n391067 , n391068 , n70086 , n391070 , n391071 , n70089 , 
 n391073 , n391074 , n70092 , n391076 , n391077 , n70095 , n391079 , n391080 , n391081 , n391082 , 
 n391083 , n391084 , n391085 , n391086 , n391087 , n391088 , n391089 , n70107 , n391091 , n70109 , 
 n70110 , n70111 , n391095 , n70113 , n391097 , n391098 , n391099 , n70116 , n391101 , n391102 , 
 n391103 , n391104 , n391105 , n70121 , n391107 , n391108 , n391109 , n70125 , n391111 , n391112 , 
 n391113 , n391114 , n391115 , n391116 , n391117 , n391118 , n391119 , n391120 , n391121 , n391122 , 
 n391123 , n391124 , n391125 , n391126 , n391127 , n391128 , n391129 , n391130 , n391131 , n391132 , 
 n391133 , n391134 , n391135 , n391136 , n391137 , n391138 , n70131 , n70132 , n391141 , n391142 , 
 n70135 , n391144 , n70137 , n391146 , n391147 , n391148 , n391149 , n70142 , n391151 , n70144 , 
 n391153 , n391154 , n391155 , n70148 , n391157 , n391158 , n70151 , n391160 , n391161 , n70154 , 
 n391163 , n70156 , n391165 , n391166 , n391167 , n391168 , n391169 , n391170 , n70163 , n70164 , 
 n391173 , n70166 , n391175 , n391176 , n70169 , n391178 , n70171 , n391180 , n391181 , n391182 , 
 n391183 , n391184 , n70177 , n391186 , n391187 , n70180 , n70181 , n391190 , n70183 , n391192 , 
 n70185 , n70186 , n391195 , n70188 , n391197 , n70190 , n391199 , n391200 , n391201 , n391202 , 
 n391203 , n391204 , n391205 , n391206 , n391207 , n391208 , n70201 , n391210 , n391211 , n70204 , 
 n391213 , n391214 , n70207 , n391216 , n391217 , n391218 , n70211 , n391220 , n70213 , n391222 , 
 n391223 , n70216 , n70217 , n391226 , n391227 , n391228 , n70221 , n391230 , n70223 , n391232 , 
 n391233 , n70226 , n70227 , n70228 , n70229 , n391238 , n391239 , n70232 , n391241 , n391242 , 
 n391243 , n70236 , n391245 , n70238 , n391247 , n391248 , n70241 , n391250 , n391251 , n391252 , 
 n391253 , n70246 , n391255 , n391256 , n70249 , n391258 , n391259 , n391260 , n391261 , n70254 , 
 n391263 , n391264 , n70257 , n391266 , n391267 , n70260 , n391269 , n391270 , n70263 , n391272 , 
 n70265 , n391274 , n70267 , n391276 , n70269 , n70270 , n391279 , n391280 , n70273 , n391282 , 
 n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , 
 n391293 , n70286 , n70287 , n70288 , n70289 , n391298 , n391299 , n70292 , n391301 , n391302 , 
 n391303 , n391304 , n391305 , n391306 , n391307 , n70300 , n391309 , n391310 , n70303 , n391312 , 
 n391313 , n391314 , n391315 , n391316 , n70309 , n391318 , n391319 , n70312 , n70313 , n391322 , 
 n391323 , n70316 , n391325 , n391326 , n391327 , n391328 , n391329 , n391330 , n391331 , n70324 , 
 n391333 , n391334 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n391342 , 
 n70335 , n391344 , n391345 , n391346 , n391347 , n391348 , n391349 , n70342 , n70343 , n391352 , 
 n391353 , n391354 , n70347 , n70348 , n391357 , n391358 , n391359 , n391360 , n391361 , n70354 , 
 n391363 , n391364 , n391365 , n391366 , n391367 , n391368 , n391369 , n70362 , n391371 , n70364 , 
 n391373 , n391374 , n391375 , n391376 , n70369 , n391378 , n391379 , n70372 , n70373 , n391382 , 
 n391383 , n391384 , n391385 , n391386 , n391387 , n70380 , n391389 , n391390 , n70383 , n70384 , 
 n70385 , n391394 , n391395 , n70388 , n391397 , n391398 , n391399 , n391400 , n391401 , n391402 , 
 n391403 , n391404 , n70397 , n70398 , n70399 , n391408 , n391409 , n70402 , n70403 , n391412 , 
 n391413 , n70406 , n70407 , n391416 , n391417 , n70410 , n70411 , n70412 , n391421 , n70414 , 
 n70415 , n70416 , n391425 , n70418 , n391427 , n70420 , n391429 , n391430 , n391431 , n70424 , 
 n391433 , n391434 , n70427 , n391436 , n391437 , n391438 , n70431 , n391440 , n391441 , n391442 , 
 n391443 , n391444 , n391445 , n391446 , n70439 , n391448 , n70441 , n391450 , n391451 , n70444 , 
 n391453 , n391454 , n391455 , n391456 , n391457 , n70450 , n391459 , n391460 , n391461 , n391462 , 
 n391463 , n391464 , n391465 , n391466 , n70459 , n391468 , n391469 , n391470 , n391471 , n70464 , 
 n391473 , n391474 , n391475 , n391476 , n391477 , n391478 , n391479 , n70472 , n391481 , n391482 , 
 n391483 , n70476 , n391485 , n391486 , n70479 , n70480 , n391489 , n391490 , n391491 , n391492 , 
 n70485 , n391494 , n391495 , n70488 , n391497 , n391498 , n391499 , n391500 , n391501 , n391502 , 
 n391503 , n391504 , n391505 , n391506 , n70499 , n70500 , n391509 , n391510 , n391511 , n70504 , 
 n70505 , n391514 , n391515 , n391516 , n391517 , n391518 , n391519 , n391520 , n391521 , n391522 , 
 n391523 , n391524 , n391525 , n391526 , n70519 , n391528 , n391529 , n70522 , n391531 , n391532 , 
 n391533 , n70526 , n70527 , n391536 , n391537 , n391538 , n391539 , n391540 , n391541 , n391542 , 
 n391543 , n70536 , n70537 , n391546 , n391547 , n70540 , n391549 , n70542 , n391551 , n391552 , 
 n70545 , n391554 , n391555 , n70548 , n70549 , n391558 , n391559 , n70552 , n391561 , n391562 , 
 n391563 , n70556 , n391565 , n391566 , n70559 , n70560 , n391569 , n391570 , n70563 , n70564 , 
 n70565 , n391574 , n391575 , n391576 , n70569 , n391578 , n391579 , n391580 , n391581 , n391582 , 
 n70575 , n391584 , n70577 , n391586 , n391587 , n391588 , n391589 , n391590 , n70583 , n391592 , 
 n391593 , n70586 , n70587 , n391596 , n391597 , n391598 , n70591 , n391600 , n391601 , n70594 , 
 n391603 , n391604 , n391605 , n391606 , n391607 , n70600 , n391609 , n391610 , n391611 , n70604 , 
 n70605 , n391614 , n391615 , n391616 , n391617 , n391618 , n391619 , n70612 , n391621 , n70614 , 
 n70615 , n70616 , n70617 , n70618 , n391627 , n391628 , n391629 , n391630 , n391631 , n70624 , 
 n70625 , n391634 , n391635 , n391636 , n391637 , n391638 , n70631 , n391640 , n391641 , n391642 , 
 n391643 , n391644 , n391645 , n391646 , n391647 , n391648 , n391649 , n391650 , n391651 , n391652 , 
 n391653 , n391654 , n391655 , n391656 , n70649 , n70650 , n391659 , n391660 , n391661 , n391662 , 
 n391663 , n391664 , n391665 , n70658 , n391667 , n391668 , n391669 , n391670 , n70663 , n391672 , 
 n391673 , n391674 , n70667 , n391676 , n391677 , n391678 , n70671 , n391680 , n391681 , n70674 , 
 n391683 , n391684 , n70677 , n391686 , n391687 , n70680 , n391689 , n391690 , n391691 , n70684 , 
 n70685 , n391694 , n391695 , n391696 , n391697 , n391698 , n391699 , n70692 , n391701 , n391702 , 
 n70695 , n70696 , n391705 , n391706 , n70699 , n70700 , n70701 , n391710 , n391711 , n70704 , 
 n391713 , n70706 , n391715 , n70708 , n391717 , n70710 , n391719 , n391720 , n70713 , n391722 , 
 n391723 , n391724 , n391725 , n391726 , n70719 , n391728 , n391729 , n70722 , n391731 , n391732 , 
 n70725 , n391734 , n70727 , n391736 , n70729 , n391738 , n70731 , n70732 , n70733 , n391742 , 
 n70735 , n391744 , n391745 , n391746 , n70739 , n391748 , n70741 , n70742 , n391751 , n391752 , 
 n391753 , n391754 , n70747 , n391756 , n391757 , n70750 , n70751 , n391760 , n70753 , n70754 , 
 n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n391770 , n391771 , n70764 , 
 n391773 , n391774 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n391781 , n70774 , 
 n391783 , n391784 , n391785 , n391786 , n391787 , n70780 , n391789 , n70782 , n391791 , n391792 , 
 n391793 , n70786 , n391795 , n391796 , n391797 , n70790 , n391799 , n391800 , n70793 , n391802 , 
 n391803 , n70796 , n391805 , n391806 , n391807 , n391808 , n391809 , n391810 , n70803 , n391812 , 
 n391813 , n391814 , n391815 , n391816 , n391817 , n70810 , n391819 , n391820 , n70813 , n391822 , 
 n391823 , n70816 , n391825 , n391826 , n70819 , n391828 , n391829 , n70822 , n391831 , n391832 , 
 n391833 , n70826 , n391835 , n391836 , n391837 , n391838 , n391839 , n391840 , n70833 , n391842 , 
 n70835 , n70836 , n70837 , n70838 , n70839 , n391848 , n70841 , n391850 , n391851 , n70844 , 
 n391853 , n391854 , n391855 , n391856 , n70849 , n70850 , n391859 , n70852 , n391861 , n70854 , 
 n391863 , n391864 , n391865 , n391866 , n391867 , n391868 , n70861 , n391870 , n391871 , n391872 , 
 n391873 , n391874 , n391875 , n70868 , n70869 , n391878 , n70871 , n70872 , n391881 , n70874 , 
 n391883 , n70876 , n391885 , n391886 , n70879 , n391888 , n391889 , n70882 , n391891 , n391892 , 
 n70885 , n391894 , n391895 , n70888 , n391897 , n391898 , n70891 , n70892 , n391901 , n391902 , 
 n391903 , n391904 , n391905 , n391906 , n391907 , n391908 , n391909 , n391910 , n391911 , n391912 , 
 n391913 , n391914 , n70907 , n391916 , n391917 , n70910 , n391919 , n391920 , n391921 , n391922 , 
 n391923 , n70916 , n391925 , n391926 , n391927 , n391928 , n391929 , n391930 , n391931 , n70924 , 
 n391933 , n70926 , n70927 , n70928 , n391937 , n70930 , n391939 , n391940 , n391941 , n391942 , 
 n391943 , n391944 , n391945 , n391946 , n391947 , n391948 , n391949 , n391950 , n391951 , n391952 , 
 n391953 , n70946 , n391955 , n391956 , n70949 , n391958 , n391959 , n391960 , n391961 , n391962 , 
 n70955 , n391964 , n70957 , n391966 , n391967 , n391968 , n70961 , n391970 , n70963 , n70964 , 
 n70965 , n391974 , n391975 , n70968 , n391977 , n391978 , n70971 , n70972 , n391981 , n70974 , 
 n391983 , n70975 , n391985 , n391986 , n391987 , n70979 , n70980 , n391990 , n391991 , n70983 , 
 n70984 , n391994 , n391995 , n391996 , n391997 , n70989 , n391999 , n392000 , n392001 , n392002 , 
 n70994 , n392004 , n392005 , n392006 , n392007 , n392008 , n392009 , n71001 , n392011 , n392012 , 
 n392013 , n392014 , n392015 , n392016 , n392017 , n392018 , n392019 , n392020 , n392021 , n71013 , 
 n71014 , n392024 , n392025 , n71017 , n392027 , n71019 , n392029 , n71021 , n71022 , n71023 , 
 n71024 , n71025 , n71026 , n392036 , n71028 , n392038 , n392039 , n392040 , n71032 , n392042 , 
 n71034 , n392044 , n392045 , n392046 , n392047 , n392048 , n392049 , n392050 , n392051 , n392052 , 
 n392053 , n392054 , n392055 , n392056 , n392057 , n392058 , n71050 , n392060 , n392061 , n71053 , 
 n392063 , n392064 , n392065 , n392066 , n71058 , n392068 , n71060 , n392070 , n392071 , n71063 , 
 n392073 , n392074 , n392075 , n71067 , n392077 , n71069 , n392079 , n392080 , n71072 , n392082 , 
 n392083 , n71075 , n392085 , n71077 , n392087 , n71079 , n71080 , n71081 , n71082 , n71083 , 
 n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n392100 , n392101 , n392102 , 
 n392103 , n71095 , n392105 , n71097 , n392107 , n71099 , n71100 , n392110 , n392111 , n392112 , 
 n392113 , n392114 , n71106 , n392116 , n392117 , n392118 , n392119 , n392120 , n392121 , n392122 , 
 n392123 , n392124 , n392125 , n392126 , n392127 , n392128 , n392129 , n392130 , n392131 , n392132 , 
 n392133 , n392134 , n71126 , n392136 , n392137 , n71129 , n392139 , n392140 , n392141 , n71133 , 
 n392143 , n71135 , n392145 , n392146 , n71138 , n71139 , n392149 , n71141 , n392151 , n392152 , 
 n71144 , n392154 , n71146 , n392156 , n392157 , n71149 , n392159 , n392160 , n392161 , n71153 , 
 n392163 , n392164 , n392165 , n392166 , n392167 , n392168 , n392169 , n71161 , n392171 , n392172 , 
 n392173 , n392174 , n392175 , n392176 , n71168 , n71169 , n392179 , n392180 , n392181 , n392182 , 
 n71174 , n392184 , n392185 , n71177 , n71178 , n392188 , n392189 , n392190 , n392191 , n392192 , 
 n392193 , n71185 , n392195 , n392196 , n71188 , n71189 , n392199 , n392200 , n392201 , n71193 , 
 n71194 , n392204 , n392205 , n392206 , n392207 , n71199 , n392209 , n392210 , n71202 , n392212 , 
 n392213 , n392214 , n392215 , n71207 , n392217 , n392218 , n392219 , n392220 , n392221 , n392222 , 
 n71214 , n392224 , n392225 , n392226 , n392227 , n71219 , n392229 , n392230 , n392231 , n71223 , 
 n71224 , n392234 , n392235 , n71227 , n71228 , n392238 , n71230 , n392240 , n392241 , n392242 , 
 n392243 , n392244 , n392245 , n392246 , n71238 , n392248 , n392249 , n71241 , n71242 , n392252 , 
 n71244 , n392254 , n392255 , n71247 , n392257 , n392258 , n392259 , n71251 , n392261 , n392262 , 
 n71254 , n392264 , n392265 , n71257 , n71258 , n392268 , n392269 , n71261 , n392271 , n392272 , 
 n71264 , n71265 , n392275 , n392276 , n392277 , n71269 , n71270 , n392280 , n392281 , n71273 , 
 n71274 , n71275 , n392285 , n392286 , n71278 , n392288 , n392289 , n71281 , n392291 , n392292 , 
 n392293 , n71285 , n392295 , n392296 , n392297 , n392298 , n392299 , n392300 , n71292 , n392302 , 
 n392303 , n71295 , n71296 , n392306 , n392307 , n392308 , n71300 , n71301 , n392311 , n392312 , 
 n392313 , n71305 , n71306 , n392316 , n392317 , n392318 , n392319 , n392320 , n71312 , n392322 , 
 n392323 , n71315 , n392325 , n392326 , n392327 , n392328 , n71320 , n392330 , n71322 , n392332 , 
 n392333 , n392334 , n71326 , n392336 , n392337 , n71329 , n71330 , n392340 , n392341 , n71333 , 
 n71334 , n392344 , n392345 , n71337 , n392347 , n392348 , n392349 , n71341 , n392351 , n392352 , 
 n71344 , n392354 , n392355 , n392356 , n392357 , n392358 , n71350 , n71351 , n392361 , n392362 , 
 n392363 , n71355 , n71356 , n392366 , n71358 , n71359 , n392369 , n392370 , n71362 , n392372 , 
 n392373 , n392374 , n71366 , n71367 , n392377 , n392378 , n392379 , n392380 , n392381 , n71373 , 
 n392383 , n392384 , n71376 , n71377 , n392387 , n392388 , n392389 , n71381 , n392391 , n392392 , 
 n392393 , n392394 , n392395 , n71387 , n392397 , n392398 , n71390 , n71391 , n392401 , n392402 , 
 n392403 , n71395 , n392405 , n392406 , n392407 , n392408 , n392409 , n392410 , n392411 , n392412 , 
 n392413 , n392414 , n71406 , n392416 , n392417 , n392418 , n71410 , n392420 , n392421 , n71413 , 
 n392423 , n392424 , n71416 , n392426 , n392427 , n392428 , n392429 , n392430 , n71422 , n392432 , 
 n392433 , n392434 , n71426 , n392436 , n392437 , n392438 , n392439 , n392440 , n392441 , n392442 , 
 n71434 , n392444 , n392445 , n71437 , n71438 , n392448 , n392449 , n71441 , n392451 , n392452 , 
 n71444 , n392454 , n392455 , n71447 , n392457 , n392458 , n71450 , n71451 , n392461 , n392462 , 
 n392463 , n392464 , n71456 , n71457 , n392467 , n71459 , n392469 , n71461 , n71462 , n71463 , 
 n71464 , n71465 , n392475 , n71467 , n392477 , n71469 , n392479 , n392480 , n392481 , n392482 , 
 n392483 , n392484 , n71476 , n392486 , n392487 , n392488 , n392489 , n71481 , n392491 , n392492 , 
 n71484 , n392494 , n392495 , n392496 , n71488 , n392498 , n392499 , n392500 , n71492 , n71493 , 
 n392503 , n71495 , n71496 , n71497 , n392507 , n392508 , n71500 , n392510 , n71502 , n392512 , 
 n392513 , n392514 , n392515 , n392516 , n71508 , n392518 , n392519 , n392520 , n392521 , n392522 , 
 n392523 , n392524 , n392525 , n392526 , n392527 , n71519 , n71520 , n392530 , n392531 , n71523 , 
 n392533 , n392534 , n392535 , n392536 , n392537 , n392538 , n392539 , n71531 , n71532 , n71533 , 
 n71534 , n392544 , n392545 , n71537 , n392547 , n392548 , n392549 , n71541 , n71542 , n392552 , 
 n392553 , n71545 , n392555 , n392556 , n392557 , n392558 , n392559 , n392560 , n392561 , n392562 , 
 n392563 , n392564 , n71556 , n71557 , n392567 , n392568 , n392569 , n71561 , n392571 , n392572 , 
 n71564 , n392574 , n392575 , n71567 , n71568 , n71569 , n392579 , n392580 , n71572 , n392582 , 
 n392583 , n392584 , n392585 , n392586 , n392587 , n392588 , n392589 , n392590 , n71582 , n71583 , 
 n392593 , n392594 , n392595 , n71587 , n392597 , n392598 , n71590 , n392600 , n392601 , n71593 , 
 n392603 , n392604 , n71596 , n392606 , n392607 , n392608 , n392609 , n71601 , n392611 , n392612 , 
 n392613 , n71605 , n71606 , n392616 , n71608 , n392618 , n392619 , n392620 , n392621 , n71613 , 
 n392623 , n392624 , n71616 , n71617 , n392627 , n392628 , n392629 , n392630 , n71622 , n392632 , 
 n392633 , n71625 , n392635 , n392636 , n392637 , n71629 , n392639 , n392640 , n71632 , n392642 , 
 n392643 , n71635 , n71636 , n392646 , n392647 , n392648 , n392649 , n392650 , n71642 , n71643 , 
 n71644 , n392654 , n392655 , n71647 , n71648 , n392658 , n71650 , n392660 , n392661 , n71653 , 
 n392663 , n392664 , n392665 , n392666 , n392667 , n71659 , n71660 , n392670 , n392671 , n71663 , 
 n392673 , n392674 , n71666 , n392676 , n71668 , n71669 , n392679 , n71671 , n392681 , n71673 , 
 n71674 , n71675 , n71676 , n71677 , n392687 , n392688 , n71680 , n71681 , n71682 , n71683 , 
 n392693 , n392694 , n392695 , n392696 , n71688 , n392698 , n392699 , n71691 , n71692 , n392702 , 
 n392703 , n392704 , n71696 , n392706 , n392707 , n392708 , n392709 , n392710 , n392711 , n392712 , 
 n71704 , n392714 , n71706 , n392716 , n392717 , n71709 , n392719 , n392720 , n392721 , n392722 , 
 n392723 , n392724 , n71716 , n392726 , n392727 , n392728 , n71720 , n392730 , n392731 , n392732 , 
 n392733 , n71725 , n71726 , n392736 , n71728 , n71729 , n71730 , n392740 , n392741 , n71733 , 
 n71734 , n71735 , n71736 , n71737 , n392747 , n71739 , n71740 , n71741 , n392751 , n392752 , 
 n71744 , n392754 , n392755 , n71747 , n71748 , n392758 , n392759 , n392760 , n71752 , n392762 , 
 n392763 , n392764 , n71756 , n392766 , n71758 , n392768 , n392769 , n392770 , n71762 , n392772 , 
 n392773 , n71765 , n392775 , n392776 , n392777 , n392778 , n392779 , n392780 , n71772 , n392782 , 
 n392783 , n392784 , n392785 , n392786 , n392787 , n71779 , n392789 , n392790 , n71782 , n392792 , 
 n392793 , n392794 , n392795 , n392796 , n392797 , n392798 , n71790 , n71791 , n392801 , n71793 , 
 n71794 , n392804 , n71796 , n392806 , n71798 , n71799 , n71800 , n392810 , n392811 , n392812 , 
 n392813 , n392814 , n71806 , n392816 , n392817 , n71809 , n392819 , n392820 , n392821 , n392822 , 
 n392823 , n392824 , n71816 , n392826 , n71818 , n392828 , n71820 , n392830 , n392831 , n392832 , 
 n392833 , n392834 , n71826 , n71827 , n392837 , n392838 , n392839 , n392840 , n392841 , n71833 , 
 n392843 , n392844 , n71836 , n71837 , n392847 , n392848 , n71840 , n392850 , n392851 , n71843 , 
 n392853 , n392854 , n392855 , n392856 , n392857 , n71849 , n71850 , n71851 , n392861 , n71853 , 
 n71854 , n392864 , n392865 , n392866 , n71858 , n71859 , n392869 , n392870 , n392871 , n71863 , 
 n392873 , n392874 , n392875 , n392876 , n392877 , n392878 , n392879 , n392880 , n392881 , n392882 , 
 n392883 , n71875 , n71876 , n392886 , n392887 , n392888 , n392889 , n392890 , n392891 , n71883 , 
 n71884 , n392894 , n392895 , n392896 , n392897 , n71889 , n392899 , n392900 , n392901 , n392902 , 
 n71894 , n71895 , n71896 , n392906 , n71898 , n71899 , n71900 , n392910 , n392911 , n71903 , 
 n392913 , n71905 , n392915 , n71907 , n71908 , n71909 , n71910 , n71911 , n392921 , n71913 , 
 n392923 , n392924 , n71916 , n71917 , n392927 , n392928 , n71920 , n392930 , n392931 , n392932 , 
 n392933 , n392934 , n392935 , n392936 , n71928 , n392938 , n392939 , n392940 , n71932 , n392942 , 
 n392943 , n71935 , n392945 , n392946 , n392947 , n392948 , n392949 , n71941 , n71942 , n392952 , 
 n392953 , n392954 , n71946 , n392956 , n392957 , n71949 , n71950 , n392960 , n392961 , n392962 , 
 n392963 , n71955 , n392965 , n392966 , n71958 , n71959 , n392969 , n392970 , n71962 , n392972 , 
 n392973 , n392974 , n392975 , n392976 , n392977 , n392978 , n71970 , n71971 , n392981 , n71973 , 
 n392983 , n392984 , n71976 , n392986 , n392987 , n71979 , n392989 , n392990 , n392991 , n392992 , 
 n392993 , n392994 , n392995 , n71987 , n71988 , n392998 , n71990 , n71991 , n71992 , n393002 , 
 n71994 , n393004 , n71996 , n71997 , n393007 , n393008 , n393009 , n393010 , n393011 , n393012 , 
 n393013 , n393014 , n393015 , n393016 , n393017 , n72009 , n393019 , n72011 , n72012 , n393022 , 
 n72014 , n393024 , n393025 , n393026 , n393027 , n72019 , n393029 , n393030 , n72022 , n393032 , 
 n393033 , n393034 , n393035 , n393036 , n393037 , n72029 , n393039 , n393040 , n72032 , n72033 , 
 n393043 , n393044 , n393045 , n393046 , n393047 , n393048 , n393049 , n72041 , n393051 , n393052 , 
 n72044 , n393054 , n72046 , n393056 , n393057 , n393058 , n72050 , n393060 , n393061 , n393062 , 
 n393063 , n393064 , n393065 , n393066 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , 
 n393073 , n393074 , n72066 , n393076 , n393077 , n393078 , n72070 , n72071 , n393081 , n72073 , 
 n393083 , n393084 , n72076 , n393086 , n72078 , n393088 , n393089 , n72081 , n393091 , n393092 , 
 n72084 , n393094 , n72086 , n393096 , n72088 , n72089 , n72090 , n72091 , n393101 , n72093 , 
 n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , 
 n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n393122 , 
 n393123 , n72115 , n393125 , n393126 , n393127 , n393128 , n72120 , n393130 , n72122 , n393132 , 
 n393133 , n393134 , n393135 , n393136 , n393137 , n393138 , n393139 , n393140 , n393141 , n72133 , 
 n393143 , n393144 , n393145 , n72137 , n72138 , n393148 , n393149 , n393150 , n393151 , n393152 , 
 n393153 , n393154 , n393155 , n393156 , n72148 , n393158 , n393159 , n72151 , n393161 , n393162 , 
 n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n393171 , n72163 , 
 n393173 , n72165 , n72166 , n393176 , n72168 , n72169 , n393179 , n393180 , n393181 , n72173 , 
 n393183 , n393184 , n393185 , n72177 , n393187 , n393188 , n72180 , n393190 , n393191 , n72183 , 
 n393193 , n393194 , n72186 , n393196 , n393197 , n72189 , n393199 , n393200 , n393201 , n72193 , 
 n393203 , n393204 , n72196 , n72197 , n393207 , n393208 , n72200 , n393210 , n393211 , n393212 , 
 n393213 , n393214 , n393215 , n393216 , n72208 , n393218 , n72210 , n393220 , n393221 , n72213 , 
 n393223 , n393224 , n393225 , n393226 , n72218 , n72219 , n72220 , n393230 , n72222 , n72223 , 
 n393233 , n393234 , n72226 , n393236 , n393237 , n72229 , n393239 , n393240 , n72232 , n393242 , 
 n393243 , n393244 , n393245 , n72237 , n393247 , n393248 , n393249 , n393250 , n393251 , n393252 , 
 n393253 , n72245 , n393255 , n393256 , n72248 , n393258 , n393259 , n72251 , n393261 , n72253 , 
 n393263 , n393264 , n393265 , n393266 , n393267 , n393268 , n72260 , n393270 , n393271 , n72263 , 
 n393273 , n72265 , n393275 , n72267 , n393277 , n393278 , n393279 , n393280 , n72272 , n393282 , 
 n72274 , n72275 , n72276 , n72277 , n393287 , n72279 , n393289 , n72281 , n72282 , n393292 , 
 n393293 , n72285 , n393295 , n393296 , n72288 , n393298 , n72290 , n393300 , n393301 , n393302 , 
 n393303 , n393304 , n393305 , n72297 , n393307 , n72299 , n393309 , n72301 , n393311 , n393312 , 
 n393313 , n72305 , n72306 , n393316 , n393317 , n393318 , n393319 , n393320 , n72312 , n72313 , 
 n393323 , n393324 , n393325 , n393326 , n72318 , n393328 , n72320 , n72321 , n393331 , n393332 , 
 n72324 , n393334 , n393335 , n72327 , n393337 , n393338 , n393339 , n72331 , n393341 , n393342 , 
 n393343 , n72335 , n393345 , n393346 , n72338 , n72339 , n393349 , n393350 , n393351 , n72343 , 
 n393353 , n393354 , n72346 , n393356 , n393357 , n72349 , n72350 , n72351 , n393361 , n393362 , 
 n393363 , n72355 , n393365 , n393366 , n393367 , n393368 , n393369 , n393370 , n393371 , n393372 , 
 n393373 , n393374 , n393375 , n393376 , n72368 , n72369 , n393379 , n72371 , n72372 , n393382 , 
 n393383 , n72375 , n393385 , n393386 , n72378 , n72379 , n72380 , n393390 , n393391 , n393392 , 
 n393393 , n393394 , n393395 , n393396 , n72388 , n72389 , n393399 , n393400 , n393401 , n393402 , 
 n393403 , n393404 , n393405 , n393406 , n393407 , n393408 , n393409 , n393410 , n72402 , n393412 , 
 n393413 , n72405 , n393415 , n393416 , n393417 , n72409 , n393419 , n393420 , n393421 , n72413 , 
 n393423 , n393424 , n72416 , n393426 , n393427 , n72419 , n72420 , n393430 , n72422 , n72423 , 
 n393433 , n72425 , n72426 , n393436 , n393437 , n393438 , n72430 , n393440 , n393441 , n72433 , 
 n393443 , n393444 , n393445 , n393446 , n393447 , n393448 , n72440 , n393450 , n393451 , n393452 , 
 n393453 , n72445 , n393455 , n72447 , n393457 , n393458 , n72450 , n393460 , n393461 , n393462 , 
 n393463 , n393464 , n393465 , n393466 , n393467 , n393468 , n393469 , n72461 , n72462 , n393472 , 
 n393473 , n393474 , n72466 , n393476 , n393477 , n72469 , n72470 , n393480 , n393481 , n72473 , 
 n72474 , n393484 , n393485 , n72477 , n72478 , n72479 , n393489 , n393490 , n72482 , n72483 , 
 n72484 , n393494 , n393495 , n72487 , n393497 , n393498 , n393499 , n393500 , n72492 , n393502 , 
 n393503 , n72495 , n393505 , n393506 , n393507 , n72499 , n393509 , n393510 , n72502 , n72503 , 
 n393513 , n393514 , n72506 , n393516 , n393517 , n72509 , n72510 , n393520 , n393521 , n393522 , 
 n72514 , n393524 , n393525 , n393526 , n72518 , n72519 , n393529 , n393530 , n393531 , n393532 , 
 n393533 , n72525 , n393535 , n393536 , n72528 , n72529 , n393539 , n393540 , n393541 , n393542 , 
 n393543 , n393544 , n393545 , n72537 , n72538 , n393548 , n72540 , n72541 , n72542 , n393552 , 
 n393553 , n393554 , n72546 , n393556 , n393557 , n393558 , n393559 , n393560 , n393561 , n393562 , 
 n393563 , n393564 , n393565 , n393566 , n393567 , n393568 , n393569 , n393570 , n393571 , n393572 , 
 n393573 , n72565 , n393575 , n393576 , n72568 , n393578 , n393579 , n72571 , n393581 , n393582 , 
 n393583 , n72575 , n393585 , n393586 , n393587 , n72579 , n393589 , n393590 , n72582 , n393592 , 
 n393593 , n393594 , n72586 , n393596 , n72588 , n393598 , n393599 , n72591 , n72592 , n72593 , 
 n393603 , n393604 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , 
 n393613 , n72605 , n393615 , n393616 , n393617 , n72609 , n393619 , n393620 , n393621 , n72613 , 
 n72614 , n393624 , n393625 , n393626 , n393627 , n393628 , n393629 , n72621 , n72622 , n393632 , 
 n393633 , n393634 , n72626 , n393636 , n393637 , n72629 , n72630 , n393640 , n393641 , n393642 , 
 n393643 , n393644 , n393645 , n72637 , n393647 , n393648 , n393649 , n393650 , n393651 , n393652 , 
 n393653 , n393654 , n393655 , n72647 , n393657 , n393658 , n393659 , n72651 , n393661 , n72653 , 
 n72654 , n72655 , n72656 , n393666 , n393667 , n72659 , n72660 , n393670 , n393671 , n393672 , 
 n393673 , n393674 , n72666 , n393676 , n393677 , n393678 , n72670 , n393680 , n393681 , n393682 , 
 n72674 , n72675 , n393685 , n72677 , n393687 , n393688 , n393689 , n393690 , n72682 , n393692 , 
 n393693 , n72685 , n72686 , n393696 , n393697 , n393698 , n72690 , n393700 , n393701 , n393702 , 
 n72694 , n393704 , n393705 , n393706 , n72698 , n72699 , n393709 , n393710 , n393711 , n72703 , 
 n393713 , n393714 , n72706 , n393716 , n72708 , n393718 , n72710 , n72711 , n393721 , n393722 , 
 n72714 , n393724 , n393725 , n72717 , n393727 , n393728 , n393729 , n72721 , n393731 , n393732 , 
 n72724 , n72725 , n393735 , n393736 , n72728 , n393738 , n72730 , n72731 , n72732 , n393742 , 
 n393743 , n393744 , n72736 , n72737 , n393747 , n393748 , n72740 , n393750 , n393751 , n72743 , 
 n393753 , n393754 , n72746 , n393756 , n393757 , n72749 , n393759 , n72751 , n393761 , n72753 , 
 n393763 , n72755 , n393765 , n393766 , n72758 , n393768 , n393769 , n72761 , n393771 , n72763 , 
 n393773 , n393774 , n72766 , n393776 , n393777 , n72769 , n72770 , n393780 , n72772 , n393782 , 
 n72774 , n393784 , n393785 , n72777 , n393787 , n393788 , n393789 , n393790 , n393791 , n393792 , 
 n393793 , n393794 , n72786 , n393796 , n393797 , n72789 , n393799 , n393800 , n393801 , n72793 , 
 n393803 , n393804 , n393805 , n72797 , n393807 , n393808 , n72800 , n393810 , n393811 , n393812 , 
 n393813 , n393814 , n393815 , n72807 , n72808 , n393818 , n393819 , n393820 , n393821 , n393822 , 
 n393823 , n393824 , n72816 , n393826 , n393827 , n72819 , n393829 , n393830 , n393831 , n72823 , 
 n393833 , n393834 , n393835 , n393836 , n393837 , n72829 , n393839 , n393840 , n72832 , n72833 , 
 n72834 , n72835 , n393845 , n393846 , n72838 , n393848 , n393849 , n72841 , n393851 , n393852 , 
 n393853 , n393854 , n72846 , n72847 , n393857 , n72849 , n393859 , n393860 , n393861 , n72853 , 
 n393863 , n393864 , n72856 , n393866 , n393867 , n72859 , n393869 , n72861 , n393871 , n393872 , 
 n72864 , n393874 , n393875 , n72867 , n72868 , n393878 , n393879 , n393880 , n72872 , n393882 , 
 n393883 , n393884 , n393885 , n393886 , n393887 , n393888 , n72880 , n393890 , n393891 , n393892 , 
 n393893 , n393894 , n72886 , n393896 , n393897 , n393898 , n72890 , n393900 , n393901 , n393902 , 
 n393903 , n393904 , n393905 , n393906 , n393907 , n393908 , n393909 , n393910 , n393911 , n393912 , 
 n393913 , n72905 , n393915 , n393916 , n72908 , n72909 , n393919 , n72911 , n393921 , n393922 , 
 n393923 , n72915 , n393925 , n393926 , n72918 , n393928 , n393929 , n72921 , n393931 , n393932 , 
 n393933 , n393934 , n393935 , n393936 , n72928 , n72929 , n72930 , n393940 , n393941 , n72933 , 
 n393943 , n393944 , n393945 , n393946 , n393947 , n393948 , n393949 , n393950 , n393951 , n393952 , 
 n393953 , n393954 , n72946 , n393956 , n393957 , n72949 , n393959 , n393960 , n393961 , n393962 , 
 n393963 , n72955 , n393965 , n393966 , n393967 , n393968 , n393969 , n393970 , n72962 , n393972 , 
 n393973 , n393974 , n393975 , n393976 , n393977 , n393978 , n393979 , n393980 , n393981 , n393982 , 
 n393983 , n393984 , n393985 , n393986 , n393987 , n393988 , n72980 , n72981 , n393991 , n72983 , 
 n72984 , n393994 , n393995 , n393996 , n72988 , n393998 , n72990 , n394000 , n72992 , n394002 , 
 n394003 , n394004 , n394005 , n394006 , n72998 , n394008 , n394009 , n73001 , n394011 , n394012 , 
 n73004 , n394014 , n394015 , n73007 , n394017 , n394018 , n394019 , n394020 , n394021 , n73013 , 
 n394023 , n73015 , n394025 , n394026 , n394027 , n394028 , n394029 , n394030 , n73022 , n73023 , 
 n394033 , n73025 , n394035 , n73027 , n73028 , n394038 , n73030 , n394040 , n73032 , n394042 , 
 n394043 , n394044 , n394045 , n394046 , n394047 , n394048 , n73040 , n394050 , n394051 , n394052 , 
 n394053 , n394054 , n73046 , n394056 , n394057 , n394058 , n73050 , n394060 , n394061 , n394062 , 
 n73054 , n394064 , n394065 , n394066 , n73058 , n394068 , n394069 , n394070 , n394071 , n394072 , 
 n394073 , n394074 , n394075 , n394076 , n394077 , n394078 , n73070 , n394080 , n394081 , n73073 , 
 n394083 , n394084 , n394085 , n394086 , n394087 , n394088 , n394089 , n394090 , n394091 , n394092 , 
 n394093 , n394094 , n394095 , n394096 , n73088 , n394098 , n394099 , n394100 , n394101 , n394102 , 
 n73094 , n73095 , n394105 , n394106 , n73098 , n394108 , n73100 , n394110 , n73102 , n394112 , 
 n394113 , n73105 , n394115 , n394116 , n394117 , n394118 , n394119 , n394120 , n394121 , n394122 , 
 n73114 , n394124 , n394125 , n73117 , n73118 , n394128 , n73120 , n394130 , n394131 , n394132 , 
 n394133 , n394134 , n394135 , n394136 , n394137 , n394138 , n394139 , n73131 , n73132 , n73133 , 
 n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n394152 , 
 n73144 , n394154 , n394155 , n394156 , n394157 , n394158 , n73150 , n394160 , n394161 , n73153 , 
 n394163 , n394164 , n73156 , n394166 , n394167 , n73159 , n394169 , n394170 , n73162 , n394172 , 
 n394173 , n73165 , n394175 , n394176 , n73168 , n394178 , n73170 , n73171 , n73172 , n394182 , 
 n73174 , n394184 , n394185 , n73177 , n394187 , n394188 , n394189 , n394190 , n394191 , n394192 , 
 n73184 , n394194 , n394195 , n394196 , n73188 , n394198 , n394199 , n73191 , n394201 , n394202 , 
 n394203 , n394204 , n394205 , n73197 , n394207 , n394208 , n394209 , n394210 , n394211 , n394212 , 
 n73204 , n394214 , n394215 , n394216 , n394217 , n73209 , n394219 , n394220 , n394221 , n73213 , 
 n73214 , n394224 , n73216 , n394226 , n394227 , n73219 , n394229 , n73221 , n394231 , n394232 , 
 n394233 , n394234 , n394235 , n394236 , n73228 , n394238 , n394239 , n394240 , n394241 , n73233 , 
 n394243 , n73235 , n73236 , n394246 , n73238 , n394248 , n394249 , n73241 , n394251 , n394252 , 
 n394253 , n394254 , n394255 , n73247 , n394257 , n73249 , n73250 , n73251 , n73252 , n73253 , 
 n73254 , n73255 , n394265 , n394266 , n73258 , n394268 , n394269 , n394270 , n394271 , n394272 , 
 n394273 , n394274 , n394275 , n394276 , n394277 , n394278 , n394279 , n394280 , n394281 , n394282 , 
 n394283 , n394284 , n73276 , n394286 , n394287 , n73279 , n394289 , n394290 , n73282 , n73283 , 
 n394293 , n394294 , n73286 , n394296 , n394297 , n394298 , n394299 , n73291 , n394301 , n73293 , 
 n73294 , n73295 , n73296 , n73297 , n394307 , n73299 , n73300 , n73301 , n394311 , n394312 , 
 n73304 , n394314 , n73306 , n394316 , n394317 , n394318 , n394319 , n394320 , n394321 , n394322 , 
 n394323 , n394324 , n394325 , n394326 , n394327 , n394328 , n394329 , n394330 , n394331 , n394332 , 
 n394333 , n394334 , n394335 , n394336 , n394337 , n394338 , n394339 , n394340 , n394341 , n394342 , 
 n394343 , n394344 , n394345 , n394346 , n394347 , n394348 , n394349 , n73317 , n394351 , n394352 , 
 n394353 , n394354 , n394355 , n394356 , n394357 , n394358 , n394359 , n73327 , n73328 , n394362 , 
 n73330 , n394364 , n394365 , n394366 , n394367 , n394368 , n394369 , n394370 , n394371 , n394372 , 
 n394373 , n394374 , n73342 , n73343 , n73344 , n394378 , n394379 , n73347 , n394381 , n73349 , 
 n394383 , n73351 , n73352 , n394386 , n73354 , n394388 , n394389 , n73357 , n394391 , n394392 , 
 n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n394399 , n73367 , n394401 , n394402 , 
 n394403 , n394404 , n394405 , n394406 , n394407 , n394408 , n394409 , n394410 , n73378 , n394412 , 
 n73380 , n73381 , n73382 , n394416 , n73384 , n394418 , n394419 , n73387 , n73388 , n73389 , 
 n73390 , n73391 , n73392 , n73393 , n394427 , n394428 , n394429 , n394430 , n394431 , n394432 , 
 n394433 , n394434 , n394435 , n394436 , n394437 , n394438 , n394439 , n394440 , n73408 , n394442 , 
 n394443 , n73411 , n394445 , n394446 , n73414 , n394448 , n73416 , n73417 , n73418 , n394452 , 
 n73420 , n394454 , n394455 , n394456 , n394457 , n394458 , n394459 , n73427 , n394461 , n73429 , 
 n394463 , n394464 , n394465 , n394466 , n394467 , n394468 , n394469 , n394470 , n394471 , n394472 , 
 n394473 , n73441 , n394475 , n73443 , n394477 , n394478 , n73446 , n394480 , n394481 , n73449 , 
 n394483 , n394484 , n73452 , n394486 , n394487 , n73455 , n394489 , n394490 , n394491 , n73459 , 
 n394493 , n394494 , n394495 , n394496 , n394497 , n73465 , n394499 , n394500 , n394501 , n394502 , 
 n73470 , n394504 , n394505 , n73473 , n73474 , n394508 , n73476 , n73477 , n73478 , n73479 , 
 n73480 , n73481 , n394515 , n394516 , n394517 , n394518 , n394519 , n73487 , n394521 , n394522 , 
 n394523 , n73491 , n394525 , n394526 , n394527 , n394528 , n394529 , n394530 , n73498 , n394532 , 
 n394533 , n394534 , n394535 , n394536 , n394537 , n394538 , n394539 , n394540 , n73508 , n394542 , 
 n394543 , n73511 , n394545 , n73513 , n394547 , n73515 , n73516 , n394550 , n394551 , n73519 , 
 n394553 , n394554 , n394555 , n394556 , n394557 , n394558 , n73526 , n394560 , n394561 , n394562 , 
 n394563 , n394564 , n394565 , n394566 , n73534 , n73535 , n394569 , n394570 , n394571 , n394572 , 
 n394573 , n394574 , n73542 , n73543 , n394577 , n394578 , n394579 , n394580 , n73548 , n394582 , 
 n394583 , n394584 , n394585 , n73553 , n394587 , n394588 , n394589 , n73557 , n394591 , n394592 , 
 n73560 , n394594 , n394595 , n394596 , n394597 , n394598 , n394599 , n394600 , n73568 , n394602 , 
 n73570 , n73571 , n394605 , n394606 , n394607 , n394608 , n394609 , n73577 , n394611 , n394612 , 
 n73580 , n394614 , n394615 , n73583 , n394617 , n394618 , n73586 , n394620 , n394621 , n394622 , 
 n73590 , n73591 , n394625 , n394626 , n394627 , n394628 , n394629 , n73597 , n394631 , n394632 , 
 n394633 , n394634 , n394635 , n73603 , n394637 , n394638 , n394639 , n394640 , n394641 , n394642 , 
 n394643 , n73611 , n394645 , n394646 , n394647 , n73615 , n73616 , n394650 , n73618 , n394652 , 
 n394653 , n73621 , n394655 , n73623 , n394657 , n73625 , n394659 , n394660 , n73628 , n394662 , 
 n73630 , n73631 , n394665 , n394666 , n73634 , n394668 , n73636 , n394670 , n394671 , n394672 , 
 n394673 , n394674 , n394675 , n394676 , n394677 , n73645 , n394679 , n394680 , n394681 , n73649 , 
 n394683 , n394684 , n394685 , n394686 , n394687 , n394688 , n73656 , n73657 , n394691 , n394692 , 
 n394693 , n394694 , n73662 , n394696 , n394697 , n394698 , n73666 , n73667 , n394701 , n394702 , 
 n73670 , n394704 , n394705 , n73673 , n394707 , n394708 , n73676 , n394710 , n73678 , n394712 , 
 n73680 , n73681 , n394715 , n73683 , n394717 , n394718 , n394719 , n394720 , n394721 , n394722 , 
 n394723 , n394724 , n394725 , n394726 , n394727 , n394728 , n394729 , n394730 , n394731 , n73699 , 
 n394733 , n394734 , n394735 , n394736 , n394737 , n394738 , n394739 , n394740 , n394741 , n394742 , 
 n394743 , n73711 , n394745 , n394746 , n394747 , n73715 , n73716 , n394750 , n394751 , n73719 , 
 n394753 , n394754 , n73722 , n73723 , n394757 , n394758 , n73726 , n394760 , n73728 , n394762 , 
 n394763 , n73731 , n394765 , n394766 , n73734 , n394768 , n394769 , n394770 , n394771 , n73739 , 
 n394773 , n394774 , n394775 , n73743 , n73744 , n394778 , n394779 , n73747 , n394781 , n394782 , 
 n394783 , n73751 , n394785 , n394786 , n73754 , n394788 , n73756 , n73757 , n394791 , n394792 , 
 n394793 , n73761 , n394795 , n394796 , n394797 , n394798 , n394799 , n394800 , n394801 , n394802 , 
 n394803 , n394804 , n394805 , n73773 , n394807 , n394808 , n394809 , n73777 , n394811 , n394812 , 
 n73780 , n394814 , n394815 , n394816 , n394817 , n394818 , n73786 , n394820 , n394821 , n73789 , 
 n394823 , n73791 , n394825 , n394826 , n73794 , n394828 , n394829 , n394830 , n73798 , n394832 , 
 n394833 , n394834 , n394835 , n394836 , n394837 , n394838 , n394839 , n394840 , n394841 , n73809 , 
 n394843 , n394844 , n394845 , n394846 , n394847 , n394848 , n394849 , n394850 , n394851 , n394852 , 
 n394853 , n394854 , n73822 , n394856 , n394857 , n394858 , n394859 , n394860 , n394861 , n394862 , 
 n394863 , n394864 , n73832 , n394866 , n394867 , n394868 , n394869 , n394870 , n394871 , n394872 , 
 n394873 , n394874 , n73842 , n394876 , n394877 , n73845 , n394879 , n73847 , n394881 , n394882 , 
 n73850 , n73851 , n394885 , n73853 , n73854 , n394888 , n394889 , n394890 , n73858 , n394892 , 
 n394893 , n394894 , n394895 , n394896 , n73864 , n394898 , n394899 , n73867 , n394901 , n394902 , 
 n394903 , n73871 , n394905 , n394906 , n73874 , n73875 , n394909 , n394910 , n394911 , n394912 , 
 n394913 , n394914 , n73882 , n73883 , n394917 , n394918 , n394919 , n394920 , n394921 , n394922 , 
 n394923 , n394924 , n394925 , n394926 , n394927 , n394928 , n394929 , n394930 , n394931 , n394932 , 
 n73900 , n73901 , n394935 , n394936 , n73904 , n394938 , n394939 , n73907 , n73908 , n394942 , 
 n394943 , n394944 , n73912 , n394946 , n394947 , n73915 , n73916 , n394950 , n73918 , n394952 , 
 n394953 , n394954 , n73922 , n73923 , n394957 , n394958 , n73926 , n394960 , n394961 , n73929 , 
 n73930 , n394964 , n394965 , n394966 , n73934 , n73935 , n394969 , n394970 , n73938 , n394972 , 
 n394973 , n73941 , n394975 , n73943 , n73944 , n73945 , n394979 , n394980 , n73948 , n394982 , 
 n394983 , n73951 , n73952 , n73953 , n73954 , n73955 , n394989 , n73957 , n73958 , n394992 , 
 n394993 , n394994 , n394995 , n73963 , n394997 , n394998 , n73966 , n73967 , n395001 , n395002 , 
 n395003 , n395004 , n395005 , n395006 , n73974 , n73975 , n395009 , n395010 , n73978 , n395012 , 
 n395013 , n395014 , n395015 , n73983 , n73984 , n395018 , n73986 , n395020 , n395021 , n395022 , 
 n73990 , n395024 , n395025 , n73993 , n395027 , n395028 , n73996 , n73997 , n395031 , n395032 , 
 n395033 , n395034 , n74002 , n395036 , n395037 , n395038 , n395039 , n395040 , n395041 , n395042 , 
 n395043 , n395044 , n395045 , n395046 , n395047 , n395048 , n74016 , n395050 , n395051 , n395052 , 
 n395053 , n395054 , n395055 , n395056 , n74024 , n74025 , n395059 , n395060 , n395061 , n395062 , 
 n395063 , n395064 , n395065 , n395066 , n74034 , n395068 , n395069 , n395070 , n395071 , n395072 , 
 n395073 , n74041 , n395075 , n395076 , n395077 , n395078 , n395079 , n395080 , n395081 , n395082 , 
 n395083 , n395084 , n395085 , n395086 , n395087 , n395088 , n395089 , n395090 , n395091 , n74059 , 
 n74060 , n395094 , n395095 , n395096 , n395097 , n395098 , n395099 , n395100 , n395101 , n395102 , 
 n395103 , n395104 , n395105 , n395106 , n395107 , n395108 , n74076 , n74077 , n395111 , n395112 , 
 n74080 , n395114 , n395115 , n395116 , n395117 , n395118 , n395119 , n395120 , n74088 , n74089 , 
 n395123 , n395124 , n74092 , n395126 , n395127 , n395128 , n395129 , n395130 , n395131 , n395132 , 
 n395133 , n395134 , n395135 , n74103 , n395137 , n395138 , n395139 , n395140 , n74108 , n395142 , 
 n395143 , n74111 , n395145 , n395146 , n395147 , n395148 , n395149 , n74117 , n74118 , n395152 , 
 n74120 , n395154 , n395155 , n395156 , n395157 , n395158 , n395159 , n74127 , n395161 , n395162 , 
 n74130 , n395164 , n395165 , n395166 , n395167 , n395168 , n395169 , n74137 , n395171 , n395172 , 
 n395173 , n395174 , n395175 , n395176 , n395177 , n74145 , n395179 , n395180 , n74148 , n395182 , 
 n395183 , n395184 , n395185 , n74153 , n395187 , n395188 , n395189 , n74157 , n74158 , n395192 , 
 n74160 , n395194 , n395195 , n395196 , n395197 , n74165 , n395199 , n395200 , n395201 , n74169 , 
 n395203 , n395204 , n74172 , n395206 , n395207 , n74175 , n74176 , n74177 , n74178 , n74179 , 
 n395213 , n395214 , n395215 , n395216 , n395217 , n395218 , n395219 , n74187 , n74188 , n395222 , 
 n395223 , n395224 , n74192 , n395226 , n395227 , n74195 , n395229 , n395230 , n395231 , n395232 , 
 n395233 , n74201 , n395235 , n74203 , n395237 , n395238 , n74206 , n395240 , n395241 , n395242 , 
 n395243 , n74211 , n395245 , n395246 , n395247 , n395248 , n395249 , n395250 , n74218 , n395252 , 
 n395253 , n395254 , n395255 , n74223 , n74224 , n395258 , n395259 , n74227 , n395261 , n395262 , 
 n74230 , n395264 , n395265 , n74233 , n395267 , n395268 , n74236 , n395270 , n395271 , n74239 , 
 n395273 , n395274 , n395275 , n395276 , n74244 , n395278 , n395279 , n395280 , n74248 , n395282 , 
 n395283 , n395284 , n395285 , n395286 , n395287 , n395288 , n395289 , n395290 , n395291 , n395292 , 
 n395293 , n395294 , n395295 , n395296 , n74264 , n395298 , n395299 , n395300 , n395301 , n74269 , 
 n395303 , n395304 , n395305 , n395306 , n395307 , n395308 , n395309 , n74277 , n395311 , n74279 , 
 n74280 , n395314 , n395315 , n395316 , n395317 , n395318 , n395319 , n395320 , n395321 , n395322 , 
 n395323 , n74291 , n395325 , n395326 , n395327 , n395328 , n395329 , n395330 , n395331 , n395332 , 
 n395333 , n74301 , n395335 , n395336 , n395337 , n74305 , n74306 , n395340 , n74308 , n395342 , 
 n395343 , n74311 , n395345 , n395346 , n395347 , n74315 , n395349 , n395350 , n395351 , n395352 , 
 n395353 , n395354 , n395355 , n395356 , n395357 , n395358 , n395359 , n395360 , n74328 , n74329 , 
 n395363 , n74331 , n395365 , n395366 , n74334 , n395368 , n395369 , n395370 , n395371 , n74339 , 
 n74340 , n395374 , n395375 , n74343 , n395377 , n74345 , n395379 , n395380 , n74348 , n395382 , 
 n395383 , n74351 , n395385 , n395386 , n74354 , n74355 , n395389 , n395390 , n395391 , n395392 , 
 n395393 , n395394 , n395395 , n74363 , n395397 , n74365 , n395399 , n395400 , n74368 , n395402 , 
 n395403 , n395404 , n395405 , n395406 , n74374 , n395408 , n395409 , n395410 , n74378 , n395412 , 
 n395413 , n395414 , n395415 , n395416 , n74384 , n395418 , n74386 , n74387 , n395421 , n74389 , 
 n395423 , n74391 , n395425 , n395426 , n395427 , n74395 , n395429 , n74397 , n395431 , n395432 , 
 n395433 , n74401 , n74402 , n395436 , n395437 , n74405 , n74406 , n395440 , n74408 , n395442 , 
 n395443 , n395444 , n395445 , n74413 , n74414 , n395448 , n74416 , n74417 , n395451 , n74419 , 
 n395453 , n395454 , n74422 , n395456 , n74424 , n395458 , n395459 , n395460 , n74428 , n395462 , 
 n395463 , n74431 , n74432 , n395466 , n74434 , n395468 , n395469 , n395470 , n395471 , n395472 , 
 n395473 , n74441 , n395475 , n395476 , n395477 , n395478 , n74446 , n395480 , n395481 , n74449 , 
 n395483 , n395484 , n74452 , n395486 , n395487 , n74455 , n395489 , n395490 , n395491 , n395492 , 
 n395493 , n395494 , n395495 , n74463 , n395497 , n395498 , n74466 , n395500 , n395501 , n74469 , 
 n395503 , n395504 , n395505 , n395506 , n395507 , n395508 , n395509 , n395510 , n395511 , n74479 , 
 n74480 , n74481 , n74482 , n74483 , n74484 , n395518 , n395519 , n74487 , n395521 , n395522 , 
 n395523 , n395524 , n395525 , n395526 , n74494 , n395528 , n395529 , n74497 , n395531 , n395532 , 
 n395533 , n395534 , n74502 , n395536 , n395537 , n395538 , n395539 , n395540 , n395541 , n395542 , 
 n395543 , n395544 , n395545 , n395546 , n395547 , n395548 , n395549 , n74517 , n395551 , n395552 , 
 n74520 , n395554 , n74522 , n395556 , n395557 , n395558 , n395559 , n395560 , n395561 , n74529 , 
 n395563 , n395564 , n395565 , n74533 , n395567 , n395568 , n74536 , n395570 , n395571 , n395572 , 
 n395573 , n395574 , n395575 , n74543 , n395577 , n395578 , n395579 , n395580 , n74548 , n395582 , 
 n395583 , n74551 , n74552 , n395586 , n395587 , n395588 , n395589 , n395590 , n74558 , n395592 , 
 n74560 , n395594 , n395595 , n395596 , n395597 , n395598 , n395599 , n395600 , n74568 , n395602 , 
 n395603 , n74571 , n395605 , n395606 , n395607 , n395608 , n74576 , n395610 , n395611 , n74579 , 
 n395613 , n74581 , n395615 , n74583 , n395617 , n395618 , n395619 , n74587 , n395621 , n395622 , 
 n395623 , n395624 , n395625 , n395626 , n74594 , n74595 , n395629 , n395630 , n395631 , n395632 , 
 n395633 , n395634 , n395635 , n395636 , n395637 , n395638 , n395639 , n395640 , n395641 , n74609 , 
 n74610 , n74611 , n395645 , n395646 , n395647 , n74615 , n395649 , n395650 , n395651 , n395652 , 
 n395653 , n395654 , n395655 , n395656 , n395657 , n395658 , n74626 , n395660 , n395661 , n74629 , 
 n74630 , n395664 , n74632 , n74633 , n395667 , n395668 , n395669 , n395670 , n395671 , n395672 , 
 n395673 , n395674 , n395675 , n395676 , n74644 , n395678 , n395679 , n74647 , n395681 , n395682 , 
 n395683 , n395684 , n395685 , n395686 , n395687 , n395688 , n395689 , n395690 , n395691 , n395692 , 
 n395693 , n395694 , n395695 , n395696 , n395697 , n395698 , n395699 , n395700 , n395701 , n395702 , 
 n395703 , n395704 , n395705 , n395706 , n74674 , n395708 , n395709 , n74677 , n395711 , n395712 , 
 n395713 , n74681 , n74682 , n74683 , n395717 , n395718 , n74686 , n74687 , n74688 , n395722 , 
 n395723 , n74691 , n74692 , n395726 , n395727 , n395728 , n74696 , n395730 , n74698 , n395732 , 
 n74700 , n74701 , n395735 , n74703 , n395737 , n74705 , n395739 , n395740 , n74708 , n395742 , 
 n395743 , n74711 , n395745 , n395746 , n395747 , n395748 , n395749 , n395750 , n395751 , n395752 , 
 n395753 , n395754 , n395755 , n395756 , n395757 , n395758 , n395759 , n395760 , n395761 , n395762 , 
 n395763 , n74731 , n395765 , n395766 , n74734 , n395768 , n395769 , n74737 , n395771 , n395772 , 
 n74740 , n395774 , n395775 , n395776 , n395777 , n395778 , n74746 , n395780 , n395781 , n395782 , 
 n395783 , n395784 , n395785 , n74753 , n395787 , n395788 , n74756 , n395790 , n395791 , n395792 , 
 n74760 , n395794 , n395795 , n395796 , n74764 , n395798 , n395799 , n74767 , n395801 , n395802 , 
 n74770 , n395804 , n74772 , n74773 , n395807 , n74775 , n395809 , n395810 , n395811 , n395812 , 
 n74780 , n395814 , n395815 , n395816 , n395817 , n395818 , n74786 , n395820 , n74788 , n395822 , 
 n395823 , n74791 , n395825 , n74793 , n395827 , n395828 , n395829 , n395830 , n395831 , n395832 , 
 n395833 , n395834 , n395835 , n395836 , n395837 , n395838 , n395839 , n74807 , n395841 , n395842 , 
 n395843 , n395844 , n395845 , n74813 , n74814 , n74815 , n395849 , n74817 , n395851 , n74819 , 
 n395853 , n74821 , n74822 , n395856 , n74824 , n395858 , n395859 , n74827 , n395861 , n395862 , 
 n74830 , n395864 , n395865 , n74833 , n395867 , n395868 , n395869 , n395870 , n395871 , n395872 , 
 n395873 , n395874 , n395875 , n74843 , n395877 , n395878 , n395879 , n74847 , n74848 , n395882 , 
 n74850 , n395884 , n395885 , n74853 , n395887 , n395888 , n74856 , n395890 , n395891 , n74859 , 
 n395893 , n395894 , n395895 , n395896 , n395897 , n395898 , n74866 , n395900 , n395901 , n74869 , 
 n74870 , n395904 , n395905 , n395906 , n74874 , n74875 , n395909 , n395910 , n395911 , n395912 , 
 n395913 , n74881 , n74882 , n395916 , n395917 , n395918 , n395919 , n395920 , n395921 , n74889 , 
 n395923 , n395924 , n395925 , n395926 , n395927 , n74895 , n395929 , n395930 , n74898 , n395932 , 
 n395933 , n395934 , n395935 , n395936 , n395937 , n395938 , n395939 , n395940 , n395941 , n395942 , 
 n395943 , n74911 , n395945 , n74913 , n74914 , n74915 , n74916 , n395950 , n395951 , n395952 , 
 n74920 , n395954 , n395955 , n74923 , n74924 , n395958 , n395959 , n74927 , n395961 , n74929 , 
 n74930 , n395964 , n74932 , n395966 , n74934 , n74935 , n74936 , n395970 , n74938 , n395972 , 
 n395973 , n74941 , n395975 , n395976 , n395977 , n395978 , n395979 , n395980 , n74948 , n395982 , 
 n395983 , n395984 , n395985 , n395986 , n74954 , n395988 , n395989 , n74957 , n74958 , n395992 , 
 n395993 , n395994 , n395995 , n395996 , n395997 , n74965 , n395999 , n74967 , n74968 , n396002 , 
 n396003 , n396004 , n396005 , n396006 , n74974 , n396008 , n396009 , n396010 , n396011 , n396012 , 
 n396013 , n74975 , n74976 , n74977 , n396017 , n396018 , n396019 , n396020 , n396021 , n396022 , 
 n396023 , n396024 , n396025 , n396026 , n396027 , n396028 , n396029 , n396030 , n396031 , n74978 , 
 n74979 , n396034 , n396035 , n396036 , n396037 , n396038 , n396039 , n396040 , n396041 , n396042 , 
 n74989 , n74990 , n396045 , n396046 , n74993 , n396048 , n396049 , n396050 , n396051 , n396052 , 
 n396053 , n396054 , n396055 , n396056 , n396057 , n396058 , n396059 , n396060 , n396061 , n396062 , 
 n75009 , n75010 , n396065 , n396066 , n75013 , n396068 , n75015 , n396070 , n396071 , n396072 , 
 n396073 , n396074 , n396075 , n396076 , n396077 , n396078 , n396079 , n75026 , n75027 , n75028 , 
 n396083 , n396084 , n396085 , n396086 , n396087 , n396088 , n396089 , n396090 , n75037 , n75038 , 
 n396093 , n75040 , n396095 , n75042 , n396097 , n396098 , n396099 , n396100 , n75045 , n396102 , 
 n396103 , n396104 , n396105 , n396106 , n396107 , n396108 , n396109 , n396110 , n396111 , n396112 , 
 n396113 , n396114 , n396115 , n396116 , n396117 , n396118 , n75048 , n396120 , n396121 , n396122 , 
 n396123 , n396124 , n396125 , n396126 , n396127 , n396128 , n396129 , n396130 , n396131 , n396132 , 
 n396133 , n396134 , n396135 , n396136 , n396137 , n396138 , n396139 , n396140 , n396141 , n396142 , 
 n396143 , n396144 , n396145 , n396146 , n396147 , n396148 , n396149 , n396150 , n396151 , n396152 , 
 n396153 , n396154 , n396155 , n396156 , n396157 , n396158 , n396159 , n75063 , n396161 , n396162 , 
 n75066 , n396164 , n75068 , n396166 , n396167 , n396168 , n396169 , n396170 , n396171 , n396172 , 
 n396173 , n396174 , n396175 , n75076 , n396177 , n396178 , n75079 , n396180 , n396181 , n75082 , 
 n75083 , n396184 , n75085 , n396186 , n396187 , n396188 , n75089 , n75090 , n396191 , n75092 , 
 n396193 , n396194 , n396195 , n75096 , n396197 , n396198 , n75099 , n396200 , n396201 , n75102 , 
 n396203 , n396204 , n396205 , n396206 , n396207 , n396208 , n396209 , n396210 , n396211 , n396212 , 
 n396213 , n396214 , n396215 , n396216 , n396217 , n396218 , n396219 , n396220 , n396221 , n396222 , 
 n396223 , n396224 , n396225 , n396226 , n396227 , n75110 , n396229 , n75112 , n396231 , n396232 , 
 n396233 , n396234 , n396235 , n396236 , n75118 , n396238 , n396239 , n75121 , n396241 , n396242 , 
 n396243 , n75125 , n396245 , n75127 , n396247 , n396248 , n396249 , n396250 , n75132 , n396252 , 
 n396253 , n396254 , n396255 , n396256 , n396257 , n396258 , n396259 , n396260 , n396261 , n396262 , 
 n396263 , n396264 , n75146 , n396266 , n396267 , n75149 , n396269 , n75151 , n396271 , n396272 , 
 n75154 , n396274 , n75156 , n396276 , n396277 , n396278 , n396279 , n396280 , n396281 , n396282 , 
 n75164 , n396284 , n396285 , n396286 , n396287 , n396288 , n396289 , n396290 , n396291 , n396292 , 
 n396293 , n396294 , n396295 , n396296 , n396297 , n396298 , n396299 , n396300 , n396301 , n396302 , 
 n396303 , n396304 , n396305 , n396306 , n396307 , n396308 , n396309 , n396310 , n396311 , n75193 , 
 n396313 , n396314 , n75196 , n75197 , n75198 , n396318 , n75200 , n75201 , n396321 , n396322 , 
 n75204 , n396324 , n396325 , n396326 , n396327 , n396328 , n396329 , n396330 , n75212 , n396332 , 
 n396333 , n396334 , n396335 , n396336 , n396337 , n396338 , n396339 , n396340 , n75222 , n396342 , 
 n75224 , n396344 , n396345 , n396346 , n75228 , n75229 , n396349 , n75231 , n75232 , n396352 , 
 n396353 , n396354 , n396355 , n396356 , n75238 , n396358 , n396359 , n396360 , n75242 , n396362 , 
 n396363 , n396364 , n396365 , n396366 , n396367 , n396368 , n396369 , n396370 , n396371 , n396372 , 
 n75254 , n75255 , n396375 , n75257 , n396377 , n396378 , n75260 , n396380 , n75262 , n396382 , 
 n75264 , n396384 , n396385 , n396386 , n396387 , n396388 , n396389 , n396390 , n396391 , n396392 , 
 n396393 , n396394 , n75276 , n396396 , n396397 , n75279 , n396399 , n75281 , n396401 , n75283 , 
 n396403 , n75285 , n75286 , n75287 , n75288 , n396408 , n396409 , n396410 , n396411 , n396412 , 
 n396413 , n396414 , n396415 , n396416 , n75298 , n396418 , n75300 , n75301 , n75302 , n396422 , 
 n75304 , n396424 , n396425 , n75307 , n75308 , n396428 , n396429 , n396430 , n396431 , n396432 , 
 n75314 , n75315 , n396435 , n75317 , n75318 , n396438 , n396439 , n75321 , n396441 , n75323 , 
 n75324 , n396444 , n75326 , n75327 , n75328 , n75329 , n396449 , n75331 , n396451 , n396452 , 
 n396453 , n396454 , n396455 , n396456 , n75338 , n396458 , n396459 , n75341 , n396461 , n396462 , 
 n396463 , n396464 , n396465 , n396466 , n396467 , n75349 , n75350 , n396470 , n396471 , n75353 , 
 n396473 , n396474 , n75356 , n396476 , n396477 , n75359 , n75360 , n396480 , n396481 , n75363 , 
 n396483 , n75365 , n396485 , n396486 , n75368 , n396488 , n396489 , n396490 , n75372 , n396492 , 
 n396493 , n396494 , n75376 , n396496 , n396497 , n75379 , n396499 , n396500 , n396501 , n396502 , 
 n396503 , n396504 , n75386 , n396506 , n396507 , n396508 , n396509 , n396510 , n396511 , n396512 , 
 n75394 , n396514 , n396515 , n396516 , n396517 , n396518 , n396519 , n396520 , n396521 , n396522 , 
 n396523 , n396524 , n75406 , n396526 , n396527 , n396528 , n75410 , n75411 , n396531 , n396532 , 
 n75414 , n396534 , n396535 , n75417 , n75418 , n396538 , n396539 , n396540 , n396541 , n396542 , 
 n396543 , n396544 , n396545 , n396546 , n396547 , n396548 , n396549 , n396550 , n396551 , n396552 , 
 n396553 , n396554 , n396555 , n396556 , n396557 , n396558 , n396559 , n396560 , n396561 , n396562 , 
 n396563 , n396564 , n396565 , n396566 , n396567 , n396568 , n396569 , n396570 , n396571 , n75433 , 
 n396573 , n396574 , n75436 , n396576 , n75438 , n75439 , n396579 , n396580 , n396581 , n75443 , 
 n396583 , n396584 , n75446 , n396586 , n396587 , n75449 , n396589 , n75451 , n396591 , n396592 , 
 n396593 , n396594 , n75456 , n396596 , n396597 , n396598 , n396599 , n396600 , n75462 , n396602 , 
 n396603 , n396604 , n75466 , n75467 , n396607 , n396608 , n75470 , n396610 , n396611 , n75473 , 
 n396613 , n396614 , n396615 , n396616 , n396617 , n396618 , n396619 , n396620 , n396621 , n396622 , 
 n396623 , n396624 , n396625 , n75487 , n396627 , n396628 , n396629 , n396630 , n396631 , n75493 , 
 n396633 , n396634 , n396635 , n396636 , n396637 , n396638 , n396639 , n396640 , n396641 , n396642 , 
 n396643 , n75505 , n396645 , n396646 , n396647 , n75509 , n396649 , n396650 , n75512 , n75513 , 
 n75514 , n396654 , n396655 , n75517 , n396657 , n396658 , n396659 , n396660 , n396661 , n396662 , 
 n396663 , n396664 , n396665 , n396666 , n396667 , n75529 , n396669 , n396670 , n396671 , n396672 , 
 n396673 , n396674 , n396675 , n396676 , n75538 , n396678 , n396679 , n396680 , n396681 , n75543 , 
 n75544 , n396684 , n75546 , n75547 , n396687 , n396688 , n75550 , n396690 , n396691 , n396692 , 
 n75554 , n396694 , n396695 , n75557 , n396697 , n75559 , n396699 , n396700 , n396701 , n396702 , 
 n396703 , n396704 , n396705 , n396706 , n75568 , n75569 , n396709 , n396710 , n75572 , n396712 , 
 n396713 , n75575 , n396715 , n396716 , n75578 , n396718 , n75580 , n396720 , n396721 , n75583 , 
 n396723 , n396724 , n396725 , n396726 , n396727 , n396728 , n75590 , n396730 , n396731 , n396732 , 
 n75594 , n75595 , n396735 , n75597 , n396737 , n75599 , n396739 , n396740 , n396741 , n396742 , 
 n396743 , n75605 , n396745 , n396746 , n396747 , n396748 , n75610 , n396750 , n396751 , n75613 , 
 n396753 , n396754 , n396755 , n396756 , n396757 , n75619 , n75620 , n396760 , n75622 , n396762 , 
 n396763 , n396764 , n396765 , n396766 , n396767 , n396768 , n396769 , n396770 , n75632 , n75633 , 
 n396773 , n396774 , n75636 , n396776 , n396777 , n396778 , n396779 , n396780 , n396781 , n396782 , 
 n396783 , n396784 , n75646 , n75647 , n396787 , n396788 , n396789 , n75651 , n396791 , n396792 , 
 n75654 , n396794 , n396795 , n75657 , n396797 , n396798 , n396799 , n396800 , n396801 , n75663 , 
 n75664 , n396804 , n75666 , n75667 , n396807 , n396808 , n396809 , n396810 , n396811 , n396812 , 
 n75674 , n396814 , n396815 , n396816 , n396817 , n396818 , n396819 , n396820 , n75682 , n75683 , 
 n396823 , n396824 , n396825 , n75687 , n396827 , n396828 , n75690 , n396830 , n75692 , n396832 , 
 n396833 , n75695 , n396835 , n396836 , n396837 , n396838 , n75700 , n75701 , n396841 , n396842 , 
 n75704 , n396844 , n396845 , n75707 , n396847 , n396848 , n396849 , n396850 , n396851 , n75713 , 
 n396853 , n396854 , n75716 , n75717 , n396857 , n396858 , n75720 , n396860 , n75722 , n75723 , 
 n75724 , n75725 , n75726 , n396866 , n396867 , n75729 , n396869 , n396870 , n396871 , n75733 , 
 n396873 , n396874 , n396875 , n75737 , n396877 , n396878 , n75740 , n75741 , n396881 , n396882 , 
 n396883 , n75745 , n396885 , n75747 , n396887 , n396888 , n396889 , n396890 , n75752 , n396892 , 
 n396893 , n396894 , n75756 , n396896 , n396897 , n396898 , n75760 , n396900 , n396901 , n396902 , 
 n75764 , n396904 , n396905 , n75767 , n396907 , n75769 , n75770 , n75771 , n396911 , n75773 , 
 n396913 , n396914 , n396915 , n396916 , n396917 , n396918 , n396919 , n75781 , n75782 , n396922 , 
 n396923 , n396924 , n75786 , n396926 , n396927 , n396928 , n75790 , n75791 , n396931 , n396932 , 
 n396933 , n396934 , n396935 , n75797 , n396937 , n396938 , n75800 , n396940 , n396941 , n396942 , 
 n75804 , n396944 , n396945 , n396946 , n75808 , n396948 , n396949 , n75811 , n396951 , n396952 , 
 n396953 , n75815 , n396955 , n396956 , n396957 , n396958 , n396959 , n396960 , n396961 , n75823 , 
 n396963 , n396964 , n396965 , n396966 , n396967 , n396968 , n396969 , n396970 , n75832 , n75833 , 
 n396973 , n396974 , n396975 , n396976 , n396977 , n396978 , n396979 , n396980 , n396981 , n396982 , 
 n396983 , n396984 , n396985 , n75847 , n396987 , n396988 , n396989 , n396990 , n396991 , n396992 , 
 n396993 , n396994 , n75856 , n396996 , n396997 , n396998 , n396999 , n397000 , n397001 , n397002 , 
 n397003 , n397004 , n397005 , n75867 , n397007 , n397008 , n397009 , n75871 , n397011 , n397012 , 
 n397013 , n397014 , n397015 , n397016 , n75878 , n75879 , n397019 , n397020 , n397021 , n397022 , 
 n397023 , n397024 , n397025 , n397026 , n75888 , n397028 , n397029 , n75891 , n75892 , n397032 , 
 n397033 , n397034 , n75896 , n397036 , n397037 , n397038 , n75900 , n397040 , n397041 , n397042 , 
 n75904 , n397044 , n397045 , n397046 , n397047 , n75909 , n397049 , n397050 , n397051 , n397052 , 
 n397053 , n397054 , n397055 , n397056 , n397057 , n397058 , n397059 , n397060 , n397061 , n397062 , 
 n397063 , n397064 , n397065 , n397066 , n397067 , n397068 , n397069 , n397070 , n397071 , n397072 , 
 n397073 , n397074 , n397075 , n397076 , n397077 , n75939 , n75940 , n397080 , n397081 , n75943 , 
 n397083 , n397084 , n75946 , n75947 , n397087 , n397088 , n397089 , n397090 , n397091 , n397092 , 
 n75954 , n397094 , n397095 , n397096 , n397097 , n397098 , n75960 , n397100 , n397101 , n397102 , 
 n75964 , n397104 , n397105 , n397106 , n397107 , n397108 , n397109 , n75971 , n75972 , n75973 , 
 n75974 , n75975 , n75976 , n397116 , n397117 , n397118 , n75980 , n75981 , n397121 , n75983 , 
 n75984 , n75985 , n75986 , n75987 , n397127 , n397128 , n397129 , n397130 , n397131 , n397132 , 
 n397133 , n397134 , n397135 , n397136 , n75998 , n397138 , n397139 , n76001 , n397141 , n397142 , 
 n76004 , n397144 , n397145 , n76007 , n397147 , n76009 , n397149 , n76011 , n397151 , n76013 , 
 n397153 , n76015 , n397155 , n397156 , n397157 , n397158 , n397159 , n397160 , n76022 , n76023 , 
 n397163 , n397164 , n397165 , n397166 , n397167 , n76029 , n76030 , n397170 , n397171 , n76033 , 
 n76034 , n397174 , n397175 , n397176 , n397177 , n76039 , n76040 , n397180 , n76042 , n76043 , 
 n397183 , n397184 , n397185 , n397186 , n397187 , n397188 , n76050 , n397190 , n397191 , n76053 , 
 n397193 , n397194 , n397195 , n397196 , n397197 , n397198 , n76060 , n397200 , n397201 , n397202 , 
 n397203 , n76065 , n397205 , n397206 , n397207 , n397208 , n397209 , n76071 , n397211 , n397212 , 
 n76074 , n76075 , n397215 , n397216 , n76078 , n397218 , n397219 , n76081 , n76082 , n397222 , 
 n397223 , n76085 , n397225 , n397226 , n397227 , n76089 , n397229 , n397230 , n397231 , n397232 , 
 n76094 , n397234 , n397235 , n76097 , n76098 , n397238 , n397239 , n76101 , n397241 , n397242 , 
 n397243 , n397244 , n397245 , n76107 , n397247 , n397248 , n76110 , n397250 , n76112 , n397252 , 
 n397253 , n397254 , n397255 , n397256 , n397257 , n397258 , n397259 , n397260 , n397261 , n76123 , 
 n397263 , n397264 , n397265 , n76127 , n397267 , n397268 , n397269 , n397270 , n76132 , n397272 , 
 n397273 , n76135 , n397275 , n397276 , n397277 , n397278 , n397279 , n76141 , n397281 , n397282 , 
 n397283 , n397284 , n397285 , n397286 , n76148 , n397288 , n397289 , n76151 , n76152 , n397292 , 
 n76154 , n76155 , n397295 , n397296 , n76158 , n76159 , n397299 , n397300 , n76162 , n397302 , 
 n76164 , n397304 , n76166 , n76167 , n397307 , n397308 , n397309 , n397310 , n397311 , n397312 , 
 n397313 , n397314 , n397315 , n397316 , n397317 , n397318 , n397319 , n397320 , n397321 , n397322 , 
 n397323 , n397324 , n397325 , n397326 , n76188 , n397328 , n76190 , n397330 , n76192 , n397332 , 
 n76194 , n397334 , n397335 , n397336 , n397337 , n397338 , n397339 , n397340 , n397341 , n397342 , 
 n397343 , n397344 , n397345 , n397346 , n397347 , n76209 , n397349 , n76211 , n76212 , n76213 , 
 n397353 , n76215 , n397355 , n397356 , n397357 , n397358 , n397359 , n397360 , n397361 , n76223 , 
 n397363 , n397364 , n76226 , n397366 , n397367 , n397368 , n76230 , n397370 , n76232 , n397372 , 
 n397373 , n76235 , n397375 , n397376 , n76238 , n397378 , n397379 , n76241 , n76242 , n397382 , 
 n76244 , n397384 , n397385 , n397386 , n397387 , n397388 , n397389 , n397390 , n397391 , n397392 , 
 n397393 , n76255 , n76256 , n397396 , n397397 , n397398 , n397399 , n76261 , n397401 , n76263 , 
 n76264 , n397404 , n397405 , n76267 , n397407 , n397408 , n76270 , n397410 , n397411 , n397412 , 
 n397413 , n397414 , n397415 , n397416 , n397417 , n397418 , n397419 , n397420 , n397421 , n397422 , 
 n397423 , n397424 , n76273 , n397426 , n397427 , n397428 , n397429 , n397430 , n397431 , n397432 , 
 n397433 , n397434 , n397435 , n397436 , n397437 , n397438 , n397439 , n397440 , n397441 , n397442 , 
 n397443 , n397444 , n397445 , n397446 , n397447 , n397448 , n397449 , n397450 , n397451 , n397452 , 
 n397453 , n397454 , n397455 , n397456 , n397457 , n397458 , n397459 , n397460 , n397461 , n397462 , 
 n76290 , n76291 , n76292 , n397466 , n397467 , n397468 , n397469 , n76297 , n397471 , n397472 , 
 n397473 , n397474 , n397475 , n397476 , n76304 , n397478 , n397479 , n397480 , n397481 , n76309 , 
 n397483 , n397484 , n76312 , n397486 , n397487 , n397488 , n397489 , n397490 , n397491 , n397492 , 
 n397493 , n397494 , n397495 , n397496 , n397497 , n397498 , n76326 , n397500 , n397501 , n76329 , 
 n397503 , n397504 , n76332 , n397506 , n397507 , n76335 , n397509 , n397510 , n76338 , n397512 , 
 n397513 , n76341 , n397515 , n76343 , n397517 , n397518 , n76346 , n76347 , n397521 , n397522 , 
 n76350 , n397524 , n76352 , n397526 , n397527 , n397528 , n397529 , n397530 , n76358 , n76359 , 
 n397533 , n397534 , n76362 , n76363 , n397537 , n397538 , n397539 , n397540 , n397541 , n397542 , 
 n397543 , n397544 , n397545 , n76372 , n76373 , n397548 , n397549 , n397550 , n76377 , n76378 , 
 n397553 , n397554 , n76381 , n76382 , n397557 , n76384 , n397559 , n397560 , n397561 , n397562 , 
 n397563 , n76390 , n397565 , n397566 , n76393 , n397568 , n397569 , n76396 , n397571 , n397572 , 
 n397573 , n397574 , n397575 , n397576 , n397577 , n397578 , n397579 , n76406 , n397581 , n76408 , 
 n397583 , n397584 , n76411 , n397586 , n397587 , n397588 , n76415 , n397590 , n397591 , n397592 , 
 n397593 , n397594 , n397595 , n397596 , n397597 , n397598 , n397599 , n76426 , n397601 , n397602 , 
 n397603 , n76430 , n397605 , n397606 , n76433 , n76434 , n397609 , n76436 , n397611 , n397612 , 
 n397613 , n76440 , n397615 , n397616 , n397617 , n397618 , n397619 , n397620 , n76447 , n397622 , 
 n397623 , n397624 , n76451 , n397626 , n397627 , n397628 , n397629 , n397630 , n397631 , n76458 , 
 n397633 , n397634 , n397635 , n397636 , n397637 , n397638 , n397639 , n397640 , n397641 , n76468 , 
 n397643 , n76470 , n397645 , n76472 , n76473 , n397648 , n397649 , n76476 , n76477 , n397652 , 
 n76479 , n397654 , n397655 , n397656 , n397657 , n397658 , n397659 , n397660 , n397661 , n397662 , 
 n397663 , n397664 , n397665 , n397666 , n397667 , n397668 , n397669 , n397670 , n397671 , n397672 , 
 n397673 , n397674 , n397675 , n397676 , n397677 , n397678 , n397679 , n397680 , n397681 , n76482 , 
 n397683 , n397684 , n397685 , n397686 , n397687 , n76488 , n397689 , n397690 , n397691 , n397692 , 
 n76493 , n397694 , n397695 , n76496 , n76497 , n397698 , n76499 , n397700 , n397701 , n397702 , 
 n397703 , n397704 , n397705 , n76506 , n397707 , n76508 , n397709 , n397710 , n397711 , n397712 , 
 n397713 , n397714 , n397715 , n76516 , n76517 , n397718 , n76519 , n397720 , n397721 , n76522 , 
 n397723 , n397724 , n397725 , n397726 , n76527 , n397728 , n397729 , n397730 , n397731 , n397732 , 
 n397733 , n397734 , n76535 , n397736 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , 
 n76543 , n397744 , n397745 , n397746 , n397747 , n397748 , n397749 , n397750 , n397751 , n76552 , 
 n76553 , n76554 , n76555 , n397756 , n76557 , n397758 , n397759 , n397760 , n397761 , n397762 , 
 n397763 , n76564 , n397765 , n397766 , n397767 , n76568 , n397769 , n397770 , n397771 , n397772 , 
 n397773 , n76574 , n397775 , n397776 , n76577 , n397778 , n397779 , n76580 , n397781 , n397782 , 
 n76583 , n76584 , n397785 , n76586 , n397787 , n397788 , n397789 , n76590 , n397791 , n397792 , 
 n76593 , n397794 , n397795 , n76596 , n76597 , n397798 , n76599 , n397800 , n397801 , n397802 , 
 n397803 , n397804 , n397805 , n397806 , n397807 , n397808 , n397809 , n76610 , n397811 , n76612 , 
 n397813 , n76614 , n397815 , n397816 , n397817 , n397818 , n397819 , n397820 , n397821 , n397822 , 
 n397823 , n397824 , n397825 , n397826 , n397827 , n397828 , n397829 , n397830 , n397831 , n76632 , 
 n397833 , n397834 , n76635 , n397836 , n76637 , n397838 , n397839 , n397840 , n397841 , n397842 , 
 n397843 , n397844 , n397845 , n397846 , n397847 , n397848 , n397849 , n397850 , n76651 , n397852 , 
 n397853 , n397854 , n397855 , n76656 , n76657 , n397858 , n397859 , n397860 , n397861 , n397862 , 
 n397863 , n397864 , n397865 , n397866 , n397867 , n397868 , n397869 , n397870 , n397871 , n397872 , 
 n397873 , n397874 , n397875 , n397876 , n397877 , n397878 , n397879 , n76664 , n76665 , n397882 , 
 n76667 , n76668 , n76669 , n397886 , n397887 , n76672 , n397889 , n397890 , n76675 , n397892 , 
 n397893 , n397894 , n397895 , n397896 , n76681 , n397898 , n397899 , n76684 , n397901 , n397902 , 
 n397903 , n397904 , n397905 , n397906 , n397907 , n76692 , n397909 , n397910 , n397911 , n397912 , 
 n397913 , n397914 , n397915 , n397916 , n397917 , n397918 , n76696 , n76697 , n76698 , n397922 , 
 n76700 , n397924 , n397925 , n397926 , n397927 , n397928 , n397929 , n397930 , n76708 , n76709 , 
 n397933 , n397934 , n397935 , n397936 , n397937 , n397938 , n76716 , n76717 , n397941 , n76719 , 
 n397943 , n76721 , n397945 , n397946 , n76724 , n76725 , n76726 , n397950 , n397951 , n397952 , 
 n397953 , n397954 , n76732 , n76733 , n397957 , n76735 , n76736 , n397960 , n397961 , n397962 , 
 n76740 , n397964 , n76742 , n397966 , n397967 , n397968 , n397969 , n397970 , n397971 , n397972 , 
 n76750 , n397974 , n76752 , n397976 , n76754 , n397978 , n397979 , n397980 , n397981 , n397982 , 
 n397983 , n397984 , n397985 , n397986 , n397987 , n76765 , n397989 , n397990 , n397991 , n76769 , 
 n397993 , n397994 , n397995 , n397996 , n397997 , n397998 , n397999 , n398000 , n398001 , n398002 , 
 n398003 , n398004 , n398005 , n398006 , n398007 , n398008 , n398009 , n398010 , n398011 , n398012 , 
 n76790 , n398014 , n398015 , n398016 , n398017 , n398018 , n398019 , n398020 , n398021 , n76799 , 
 n76800 , n398024 , n398025 , n76803 , n398027 , n398028 , n398029 , n398030 , n398031 , n76809 , 
 n76810 , n398034 , n398035 , n76813 , n398037 , n398038 , n398039 , n76817 , n76818 , n398042 , 
 n398043 , n398044 , n398045 , n76823 , n398047 , n398048 , n398049 , n76827 , n398051 , n398052 , 
 n76830 , n76831 , n398055 , n398056 , n76834 , n76835 , n398059 , n398060 , n398061 , n398062 , 
 n76840 , n398064 , n398065 , n398066 , n76842 , n398068 , n398069 , n76845 , n398071 , n398072 , 
 n76848 , n398074 , n398075 , n76851 , n398077 , n398078 , n76854 , n398080 , n76856 , n398082 , 
 n398083 , n76859 , n398085 , n398086 , n398087 , n398088 , n76864 , n398090 , n398091 , n398092 , 
 n398093 , n398094 , n398095 , n398096 , n398097 , n76873 , n398099 , n76875 , n398101 , n76877 , 
 n398103 , n398104 , n76880 , n76881 , n398107 , n398108 , n76884 , n76885 , n398111 , n76887 , 
 n76888 , n398114 , n76890 , n76891 , n398117 , n76893 , n398119 , n76895 , n398121 , n76897 , 
 n398123 , n398124 , n76900 , n398126 , n398127 , n76903 , n398129 , n398130 , n76906 , n398132 , 
 n398133 , n76909 , n398135 , n398136 , n76912 , n398138 , n398139 , n398140 , n398141 , n398142 , 
 n76918 , n398144 , n398145 , n398146 , n398147 , n398148 , n398149 , n76925 , n398151 , n76927 , 
 n398153 , n398154 , n398155 , n398156 , n398157 , n398158 , n398159 , n398160 , n398161 , n398162 , 
 n398163 , n398164 , n398165 , n398166 , n398167 , n398168 , n398169 , n398170 , n398171 , n398172 , 
 n398173 , n398174 , n398175 , n398176 , n398177 , n398178 , n398179 , n398180 , n76930 , n76931 , 
 n398183 , n398184 , n398185 , n398186 , n398187 , n76936 , n398189 , n398190 , n398191 , n76940 , 
 n398193 , n398194 , n76943 , n398196 , n398197 , n76946 , n76947 , n398200 , n76949 , n398202 , 
 n398203 , n398204 , n398205 , n76954 , n398207 , n76956 , n398209 , n76958 , n76959 , n76960 , 
 n398213 , n398214 , n398215 , n398216 , n398217 , n398218 , n398219 , n398220 , n398221 , n76970 , 
 n398223 , n398224 , n76973 , n398226 , n398227 , n76976 , n398229 , n398230 , n76979 , n398232 , 
 n76981 , n398234 , n398235 , n398236 , n398237 , n398238 , n398239 , n76988 , n76989 , n398242 , 
 n398243 , n398244 , n398245 , n398246 , n398247 , n76996 , n398249 , n398250 , n398251 , n398252 , 
 n398253 , n77002 , n398255 , n77004 , n77005 , n398258 , n398259 , n77008 , n77009 , n398262 , 
 n398263 , n398264 , n398265 , n398266 , n77015 , n398268 , n398269 , n77018 , n77019 , n398272 , 
 n77021 , n398274 , n398275 , n398276 , n77025 , n77026 , n77027 , n77028 , n77029 , n398282 , 
 n77031 , n398284 , n398285 , n398286 , n398287 , n398288 , n77037 , n77038 , n77039 , n398292 , 
 n398293 , n398294 , n77043 , n77044 , n398297 , n398298 , n398299 , n398300 , n398301 , n398302 , 
 n77051 , n398304 , n398305 , n77054 , n77055 , n398308 , n77057 , n398310 , n398311 , n398312 , 
 n398313 , n77062 , n77063 , n398316 , n398317 , n77066 , n398319 , n398320 , n398321 , n398322 , 
 n398323 , n398324 , n398325 , n77074 , n398327 , n77076 , n398329 , n398330 , n398331 , n398332 , 
 n398333 , n77082 , n398335 , n77084 , n398337 , n398338 , n77087 , n398340 , n398341 , n77090 , 
 n398343 , n398344 , n77093 , n398346 , n398347 , n77096 , n77097 , n398350 , n398351 , n398352 , 
 n398353 , n398354 , n77103 , n398356 , n398357 , n398358 , n77107 , n398360 , n77109 , n77110 , 
 n398363 , n398364 , n398365 , n398366 , n77115 , n398368 , n398369 , n398370 , n398371 , n398372 , 
 n398373 , n398374 , n398375 , n398376 , n398377 , n77126 , n398379 , n398380 , n77129 , n398382 , 
 n398383 , n398384 , n398385 , n77134 , n398387 , n398388 , n398389 , n398390 , n398391 , n398392 , 
 n398393 , n398394 , n398395 , n77144 , n398397 , n77146 , n398399 , n398400 , n398401 , n398402 , 
 n398403 , n77152 , n398405 , n398406 , n398407 , n398408 , n398409 , n398410 , n398411 , n398412 , 
 n398413 , n398414 , n398415 , n77164 , n398417 , n398418 , n398419 , n398420 , n398421 , n398422 , 
 n398423 , n398424 , n398425 , n398426 , n398427 , n398428 , n77177 , n398430 , n77179 , n398432 , 
 n77181 , n398434 , n398435 , n398436 , n398437 , n398438 , n398439 , n398440 , n398441 , n398442 , 
 n398443 , n398444 , n398445 , n398446 , n398447 , n398448 , n398449 , n398450 , n77190 , n77191 , 
 n398453 , n398454 , n77194 , n398456 , n77196 , n77197 , n398459 , n398460 , n398461 , n77201 , 
 n398463 , n398464 , n77204 , n398466 , n398467 , n398468 , n398469 , n398470 , n398471 , n398472 , 
 n398473 , n398474 , n398475 , n398476 , n398477 , n398478 , n398479 , n398480 , n398481 , n398482 , 
 n398483 , n398484 , n398485 , n398486 , n398487 , n398488 , n398489 , n398490 , n398491 , n398492 , 
 n398493 , n398494 , n398495 , n398496 , n398497 , n398498 , n398499 , n398500 , n398501 , n77213 , 
 n398503 , n398504 , n77216 , n398506 , n398507 , n398508 , n77220 , n77221 , n398511 , n77223 , 
 n398513 , n398514 , n398515 , n398516 , n77228 , n398518 , n398519 , n398520 , n77232 , n398522 , 
 n77234 , n398524 , n398525 , n77237 , n398527 , n398528 , n398529 , n398530 , n398531 , n398532 , 
 n398533 , n398534 , n77246 , n398536 , n77248 , n398538 , n398539 , n398540 , n398541 , n77253 , 
 n398543 , n398544 , n398545 , n77257 , n77258 , n398548 , n77260 , n398550 , n398551 , n398552 , 
 n398553 , n398554 , n77266 , n398556 , n398557 , n398558 , n77270 , n398560 , n398561 , n398562 , 
 n398563 , n77275 , n398565 , n398566 , n77278 , n398568 , n398569 , n398570 , n398571 , n77283 , 
 n398573 , n398574 , n77286 , n398576 , n398577 , n77289 , n77290 , n398580 , n398581 , n398582 , 
 n398583 , n398584 , n398585 , n398586 , n398587 , n398588 , n77300 , n398590 , n398591 , n398592 , 
 n398593 , n398594 , n398595 , n398596 , n398597 , n398598 , n398599 , n398600 , n77312 , n398602 , 
 n398603 , n398604 , n398605 , n398606 , n77318 , n398608 , n398609 , n77321 , n398611 , n398612 , 
 n398613 , n77325 , n77326 , n77327 , n398617 , n398618 , n398619 , n398620 , n77332 , n398622 , 
 n398623 , n398624 , n398625 , n398626 , n398627 , n398628 , n398629 , n398630 , n77342 , n398632 , 
 n398633 , n398634 , n77346 , n398636 , n398637 , n77349 , n398639 , n398640 , n398641 , n398642 , 
 n398643 , n398644 , n398645 , n398646 , n398647 , n398648 , n398649 , n398650 , n398651 , n398652 , 
 n398653 , n77365 , n398655 , n398656 , n398657 , n77369 , n398659 , n398660 , n398661 , n398662 , 
 n398663 , n398664 , n77376 , n398666 , n398667 , n77379 , n398669 , n398670 , n398671 , n398672 , 
 n77384 , n398674 , n398675 , n398676 , n77388 , n77389 , n398679 , n77391 , n398681 , n398682 , 
 n77394 , n398684 , n398685 , n398686 , n398687 , n398688 , n398689 , n398690 , n398691 , n398692 , 
 n398693 , n398694 , n77406 , n398696 , n398697 , n398698 , n77410 , n398700 , n77412 , n398702 , 
 n398703 , n398704 , n398705 , n398706 , n398707 , n398708 , n77420 , n398710 , n398711 , n77423 , 
 n398713 , n398714 , n398715 , n398716 , n398717 , n398718 , n398719 , n398720 , n398721 , n398722 , 
 n77434 , n77435 , n398725 , n398726 , n77438 , n398728 , n77440 , n398730 , n77442 , n77443 , 
 n398733 , n77445 , n398735 , n398736 , n398737 , n398738 , n398739 , n77451 , n398741 , n398742 , 
 n77454 , n398744 , n398745 , n398746 , n398747 , n398748 , n398749 , n77461 , n398751 , n398752 , 
 n398753 , n398754 , n398755 , n398756 , n77468 , n398758 , n398759 , n398760 , n77472 , n398762 , 
 n77474 , n398764 , n77476 , n398766 , n398767 , n398768 , n398769 , n398770 , n398771 , n398772 , 
 n398773 , n398774 , n398775 , n398776 , n77488 , n398778 , n398779 , n398780 , n398781 , n398782 , 
 n77494 , n398784 , n398785 , n398786 , n398787 , n77499 , n398789 , n77501 , n398791 , n398792 , 
 n398793 , n398794 , n77506 , n398796 , n398797 , n77509 , n398799 , n398800 , n77512 , n398802 , 
 n398803 , n398804 , n77516 , n398806 , n398807 , n77519 , n398809 , n398810 , n398811 , n398812 , 
 n398813 , n398814 , n398815 , n398816 , n77528 , n77529 , n398819 , n77531 , n398821 , n398822 , 
 n77534 , n77535 , n77536 , n398826 , n77538 , n77539 , n398829 , n398830 , n77542 , n398832 , 
 n398833 , n77545 , n77546 , n398836 , n398837 , n398838 , n77550 , n398840 , n398841 , n77553 , 
 n77554 , n398844 , n398845 , n398846 , n398847 , n398848 , n398849 , n398850 , n77562 , n77563 , 
 n398853 , n398854 , n398855 , n398856 , n398857 , n398858 , n398859 , n77571 , n398861 , n398862 , 
 n398863 , n77575 , n398865 , n398866 , n398867 , n398868 , n398869 , n77581 , n398871 , n398872 , 
 n77584 , n398874 , n77586 , n398876 , n398877 , n77589 , n398879 , n398880 , n398881 , n77593 , 
 n398883 , n398884 , n398885 , n77597 , n398887 , n398888 , n398889 , n77601 , n77602 , n77603 , 
 n77604 , n398894 , n77606 , n398896 , n398897 , n398898 , n398899 , n398900 , n398901 , n398902 , 
 n398903 , n77615 , n398905 , n398906 , n77618 , n398908 , n398909 , n77621 , n77622 , n398912 , 
 n77624 , n398914 , n398915 , n398916 , n398917 , n398918 , n398919 , n398920 , n398921 , n398922 , 
 n398923 , n398924 , n398925 , n398926 , n398927 , n398928 , n398929 , n77641 , n398931 , n398932 , 
 n398933 , n398934 , n398935 , n398936 , n398937 , n398938 , n398939 , n398940 , n398941 , n77653 , 
 n398943 , n77655 , n398945 , n77657 , n398947 , n77659 , n398949 , n77661 , n398951 , n398952 , 
 n398953 , n77665 , n398955 , n398956 , n77668 , n398958 , n398959 , n398960 , n398961 , n77673 , 
 n398963 , n398964 , n77676 , n398966 , n398967 , n77679 , n398969 , n398970 , n398971 , n398972 , 
 n398973 , n398974 , n398975 , n398976 , n398977 , n398978 , n398979 , n398980 , n398981 , n398982 , 
 n398983 , n398984 , n398985 , n398986 , n398987 , n398988 , n77700 , n77701 , n398991 , n398992 , 
 n77704 , n77705 , n77706 , n77707 , n77708 , n398998 , n77710 , n77711 , n399001 , n399002 , 
 n77714 , n399004 , n77716 , n77717 , n399007 , n77719 , n77720 , n399010 , n399011 , n77723 , 
 n399013 , n399014 , n77726 , n77727 , n399017 , n399018 , n77730 , n399020 , n77732 , n399022 , 
 n77734 , n399024 , n399025 , n399026 , n399027 , n399028 , n399029 , n77741 , n77742 , n399032 , 
 n77744 , n399034 , n77746 , n77747 , n399037 , n399038 , n77750 , n77751 , n77752 , n399042 , 
 n399043 , n77755 , n399045 , n399046 , n399047 , n399048 , n399049 , n399050 , n399051 , n399052 , 
 n399053 , n399054 , n77766 , n399056 , n77768 , n399058 , n399059 , n399060 , n399061 , n399062 , 
 n399063 , n399064 , n399065 , n77777 , n399067 , n399068 , n77780 , n399070 , n399071 , n77783 , 
 n399073 , n399074 , n77786 , n399076 , n399077 , n77789 , n399079 , n399080 , n399081 , n77793 , 
 n77794 , n399084 , n399085 , n77797 , n399087 , n399088 , n77800 , n399090 , n399091 , n77803 , 
 n399093 , n399094 , n399095 , n399096 , n399097 , n399098 , n399099 , n77811 , n399101 , n77813 , 
 n399103 , n399104 , n399105 , n399106 , n399107 , n399108 , n77819 , n399110 , n399111 , n77822 , 
 n77823 , n399114 , n399115 , n77826 , n399117 , n399118 , n399119 , n399120 , n399121 , n77832 , 
 n399123 , n399124 , n399125 , n399126 , n399127 , n399128 , n77839 , n399130 , n399131 , n399132 , 
 n399133 , n77844 , n77845 , n77846 , n399137 , n77848 , n77849 , n399140 , n77851 , n399142 , 
 n399143 , n77854 , n399145 , n77856 , n399147 , n77858 , n77859 , n399150 , n399151 , n399152 , 
 n399153 , n77864 , n77865 , n77866 , n77867 , n399158 , n399159 , n399160 , n399161 , n399162 , 
 n399163 , n77874 , n399165 , n399166 , n77877 , n399168 , n399169 , n77880 , n399171 , n399172 , 
 n77883 , n399174 , n399175 , n399176 , n399177 , n77888 , n399179 , n77890 , n399181 , n77892 , 
 n77893 , n77894 , n399185 , n399186 , n399187 , n399188 , n399189 , n399190 , n399191 , n399192 , 
 n399193 , n399194 , n399195 , n399196 , n399197 , n399198 , n399199 , n399200 , n399201 , n399202 , 
 n399203 , n399204 , n77901 , n399206 , n77903 , n399208 , n399209 , n399210 , n399211 , n399212 , 
 n399213 , n77909 , n399215 , n399216 , n77912 , n399218 , n77914 , n399220 , n399221 , n399222 , 
 n399223 , n399224 , n399225 , n399226 , n399227 , n399228 , n399229 , n399230 , n399231 , n399232 , 
 n399233 , n399234 , n399235 , n399236 , n399237 , n399238 , n399239 , n77935 , n399241 , n399242 , 
 n77938 , n399244 , n77940 , n399246 , n399247 , n399248 , n399249 , n399250 , n399251 , n399252 , 
 n399253 , n399254 , n399255 , n399256 , n399257 , n77953 , n399259 , n399260 , n77956 , n77957 , 
 n399263 , n77959 , n399265 , n77961 , n399267 , n399268 , n399269 , n77965 , n399271 , n399272 , 
 n399273 , n399274 , n399275 , n399276 , n399277 , n77973 , n399279 , n399280 , n399281 , n77977 , 
 n399283 , n399284 , n399285 , n77981 , n399287 , n399288 , n77984 , n399290 , n399291 , n399292 , 
 n77988 , n399294 , n399295 , n399296 , n399297 , n399298 , n77994 , n399300 , n399301 , n399302 , 
 n399303 , n399304 , n399305 , n399306 , n399307 , n399308 , n399309 , n399310 , n399311 , n78007 , 
 n399313 , n399314 , n78010 , n78011 , n399317 , n78013 , n78014 , n399320 , n399321 , n399322 , 
 n399323 , n399324 , n399325 , n399326 , n399327 , n399328 , n399329 , n399330 , n399331 , n78027 , 
 n399333 , n399334 , n78030 , n399336 , n399337 , n78033 , n399339 , n399340 , n399341 , n78037 , 
 n78038 , n399344 , n399345 , n78041 , n399347 , n399348 , n78044 , n399350 , n399351 , n399352 , 
 n399353 , n78049 , n399355 , n399356 , n78052 , n399358 , n399359 , n399360 , n399361 , n78057 , 
 n399363 , n399364 , n78060 , n399366 , n399367 , n399368 , n78064 , n78065 , n399371 , n399372 , 
 n399373 , n78069 , n399375 , n78071 , n399377 , n399378 , n399379 , n399380 , n399381 , n399382 , 
 n399383 , n399384 , n399385 , n399386 , n78082 , n78083 , n399389 , n399390 , n399391 , n399392 , 
 n399393 , n78089 , n399395 , n399396 , n399397 , n399398 , n78094 , n399400 , n399401 , n399402 , 
 n399403 , n399404 , n399405 , n78101 , n399407 , n399408 , n399409 , n78105 , n399411 , n399412 , 
 n399413 , n78109 , n399415 , n399416 , n399417 , n78113 , n78114 , n78115 , n399421 , n399422 , 
 n78118 , n399424 , n399425 , n399426 , n78122 , n399428 , n399429 , n399430 , n78126 , n399432 , 
 n78128 , n399434 , n399435 , n399436 , n399437 , n78133 , n399439 , n399440 , n78136 , n399442 , 
 n399443 , n78139 , n78140 , n78141 , n399447 , n399448 , n78144 , n78145 , n78146 , n399452 , 
 n78148 , n78149 , n399455 , n399456 , n399457 , n399458 , n399459 , n399460 , n399461 , n399462 , 
 n399463 , n78159 , n78160 , n399466 , n399467 , n399468 , n399469 , n399470 , n399471 , n78167 , 
 n78168 , n399474 , n399475 , n399476 , n399477 , n399478 , n399479 , n399480 , n399481 , n399482 , 
 n399483 , n399484 , n399485 , n399486 , n399487 , n399488 , n399489 , n399490 , n399491 , n399492 , 
 n399493 , n78189 , n399495 , n399496 , n78192 , n399498 , n78194 , n399500 , n399501 , n399502 , 
 n78198 , n399504 , n78200 , n399506 , n399507 , n399508 , n399509 , n399510 , n399511 , n399512 , 
 n78208 , n399514 , n399515 , n399516 , n399517 , n399518 , n78214 , n78215 , n399521 , n399522 , 
 n78218 , n78219 , n399525 , n399526 , n399527 , n399528 , n78224 , n78225 , n78226 , n399532 , 
 n399533 , n78229 , n399535 , n399536 , n78232 , n399538 , n399539 , n399540 , n399541 , n399542 , 
 n399543 , n399544 , n399545 , n399546 , n399547 , n399548 , n399549 , n78245 , n399551 , n399552 , 
 n399553 , n399554 , n78250 , n399556 , n78252 , n399558 , n399559 , n78255 , n399561 , n399562 , 
 n399563 , n399564 , n78260 , n78261 , n399567 , n399568 , n399569 , n78265 , n399571 , n399572 , 
 n399573 , n78269 , n78270 , n399576 , n78272 , n78273 , n399579 , n399580 , n78276 , n399582 , 
 n399583 , n78279 , n78280 , n399586 , n399587 , n78283 , n399589 , n399590 , n78286 , n399592 , 
 n399593 , n399594 , n399595 , n399596 , n399597 , n78293 , n399599 , n399600 , n78296 , n399602 , 
 n399603 , n78299 , n399605 , n399606 , n78302 , n399608 , n399609 , n78305 , n399611 , n399612 , 
 n399613 , n78309 , n399615 , n399616 , n399617 , n399618 , n399619 , n399620 , n78316 , n399622 , 
 n399623 , n399624 , n399625 , n399626 , n399627 , n399628 , n399629 , n399630 , n78326 , n399632 , 
 n399633 , n78329 , n399635 , n399636 , n78332 , n399638 , n399639 , n399640 , n399641 , n399642 , 
 n399643 , n399644 , n78340 , n78341 , n399647 , n399648 , n78344 , n399650 , n399651 , n399652 , 
 n399653 , n399654 , n78350 , n399656 , n78352 , n399658 , n78354 , n399660 , n399661 , n399662 , 
 n399663 , n78359 , n78360 , n78361 , n399667 , n399668 , n399669 , n399670 , n399671 , n78367 , 
 n399673 , n78369 , n399675 , n78371 , n399677 , n399678 , n78374 , n399680 , n399681 , n399682 , 
 n399683 , n399684 , n78380 , n399686 , n399687 , n78383 , n399689 , n78385 , n78386 , n399692 , 
 n399693 , n78389 , n399695 , n399696 , n399697 , n399698 , n399699 , n399700 , n78396 , n78397 , 
 n399703 , n78399 , n78400 , n399706 , n399707 , n399708 , n399709 , n399710 , n399711 , n399712 , 
 n78408 , n399714 , n399715 , n399716 , n399717 , n399718 , n399719 , n399720 , n399721 , n399722 , 
 n399723 , n399724 , n399725 , n399726 , n78422 , n78423 , n399729 , n399730 , n399731 , n399732 , 
 n399733 , n399734 , n399735 , n78431 , n399737 , n399738 , n399739 , n399740 , n399741 , n399742 , 
 n399743 , n399744 , n399745 , n399746 , n399747 , n399748 , n399749 , n78445 , n78446 , n78447 , 
 n399753 , n399754 , n78450 , n78451 , n399757 , n399758 , n78454 , n78455 , n399761 , n399762 , 
 n399763 , n78459 , n399765 , n399766 , n399767 , n399768 , n78464 , n399770 , n399771 , n399772 , 
 n399773 , n399774 , n399775 , n399776 , n399777 , n399778 , n399779 , n78475 , n399781 , n399782 , 
 n399783 , n399784 , n399785 , n399786 , n78482 , n78483 , n399789 , n78485 , n399791 , n399792 , 
 n399793 , n399794 , n399795 , n399796 , n399797 , n78493 , n399799 , n78495 , n399801 , n399802 , 
 n78498 , n399804 , n78500 , n78501 , n78502 , n399808 , n399809 , n399810 , n78506 , n399812 , 
 n399813 , n78509 , n399815 , n78511 , n399817 , n78513 , n399819 , n399820 , n78516 , n399822 , 
 n399823 , n78519 , n399825 , n78521 , n78522 , n399828 , n399829 , n399830 , n78526 , n399832 , 
 n399833 , n78529 , n399835 , n399836 , n399837 , n78533 , n399839 , n399840 , n78536 , n78537 , 
 n399843 , n399844 , n78540 , n78541 , n78542 , n399848 , n399849 , n78545 , n399851 , n399852 , 
 n399853 , n399854 , n399855 , n78551 , n399857 , n399858 , n78554 , n399860 , n399861 , n78557 , 
 n399863 , n399864 , n78560 , n78561 , n78562 , n78563 , n78564 , n78565 , n399871 , n399872 , 
 n399873 , n78569 , n399875 , n399876 , n78572 , n399878 , n399879 , n78575 , n399881 , n399882 , 
 n78578 , n78579 , n399885 , n399886 , n399887 , n399888 , n399889 , n399890 , n78586 , n399892 , 
 n399893 , n399894 , n399895 , n78591 , n399897 , n399898 , n78594 , n399900 , n78596 , n78597 , 
 n78598 , n78599 , n399905 , n78601 , n399907 , n399908 , n399909 , n399910 , n399911 , n399912 , 
 n399913 , n78609 , n399915 , n78611 , n399917 , n78613 , n399919 , n78615 , n399921 , n399922 , 
 n399923 , n399924 , n399925 , n78621 , n399927 , n78623 , n78624 , n399930 , n399931 , n78627 , 
 n78628 , n399934 , n78630 , n399936 , n399937 , n399938 , n399939 , n399940 , n78636 , n399942 , 
 n399943 , n399944 , n399945 , n78641 , n399947 , n399948 , n399949 , n78645 , n399951 , n78647 , 
 n78648 , n78649 , n399955 , n399956 , n78652 , n399958 , n399959 , n78655 , n399961 , n399962 , 
 n399963 , n399964 , n399965 , n399966 , n399967 , n78663 , n399969 , n399970 , n78666 , n399972 , 
 n399973 , n78669 , n78670 , n399976 , n78672 , n399978 , n399979 , n78675 , n399981 , n399982 , 
 n399983 , n399984 , n399985 , n399986 , n399987 , n399988 , n399989 , n78685 , n78686 , n399992 , 
 n399993 , n78689 , n399995 , n78691 , n399997 , n399998 , n78694 , n400000 , n400001 , n400002 , 
 n400003 , n400004 , n400005 , n400006 , n400007 , n400008 , n400009 , n78705 , n400011 , n400012 , 
 n400013 , n400014 , n400015 , n78711 , n400017 , n400018 , n400019 , n400020 , n400021 , n78717 , 
 n400023 , n78719 , n400025 , n400026 , n78722 , n400028 , n78724 , n400030 , n400031 , n78727 , 
 n400033 , n78729 , n78730 , n400036 , n400037 , n400038 , n400039 , n400040 , n400041 , n78737 , 
 n78738 , n78739 , n78740 , n78741 , n78742 , n400048 , n400049 , n400050 , n400051 , n78747 , 
 n400053 , n400054 , n400055 , n400056 , n400057 , n400058 , n400059 , n400060 , n78756 , n78757 , 
 n78758 , n400064 , n78760 , n78761 , n400067 , n78763 , n400069 , n400070 , n78766 , n400072 , 
 n400073 , n78769 , n400075 , n400076 , n78772 , n400078 , n400079 , n78775 , n400081 , n78777 , 
 n78778 , n400084 , n400085 , n400086 , n400087 , n400088 , n400089 , n78785 , n400091 , n400092 , 
 n78788 , n400094 , n78790 , n400096 , n400097 , n400098 , n78794 , n400100 , n400101 , n78797 , 
 n400103 , n400104 , n400105 , n400106 , n400107 , n400108 , n78804 , n400110 , n400111 , n400112 , 
 n400113 , n400114 , n400115 , n400116 , n400117 , n400118 , n400119 , n78815 , n400121 , n400122 , 
 n400123 , n400124 , n400125 , n78821 , n400127 , n78823 , n400129 , n400130 , n78826 , n400132 , 
 n400133 , n400134 , n400135 , n400136 , n400137 , n400138 , n400139 , n400140 , n400141 , n78837 , 
 n400143 , n400144 , n400145 , n78841 , n400147 , n400148 , n400149 , n400150 , n400151 , n78847 , 
 n400153 , n78849 , n400155 , n78851 , n78852 , n78853 , n78854 , n78855 , n400161 , n400162 , 
 n400163 , n400164 , n400165 , n400166 , n400167 , n400168 , n400169 , n400170 , n400171 , n400172 , 
 n400173 , n400174 , n400175 , n400176 , n400177 , n400178 , n400179 , n400180 , n400181 , n400182 , 
 n400183 , n400184 , n400185 , n78858 , n400187 , n400188 , n78861 , n400190 , n400191 , n400192 , 
 n400193 , n400194 , n400195 , n400196 , n400197 , n78870 , n400199 , n400200 , n400201 , n78874 , 
 n78875 , n400204 , n400205 , n400206 , n400207 , n78880 , n400209 , n400210 , n78883 , n400212 , 
 n400213 , n78886 , n400215 , n400216 , n400217 , n400218 , n400219 , n78892 , n400221 , n400222 , 
 n400223 , n78896 , n400225 , n400226 , n400227 , n400228 , n78901 , n400230 , n400231 , n400232 , 
 n400233 , n400234 , n78907 , n400236 , n78909 , n400238 , n400239 , n400240 , n400241 , n400242 , 
 n78915 , n400244 , n400245 , n78918 , n400247 , n400248 , n78921 , n400250 , n400251 , n78924 , 
 n400253 , n400254 , n400255 , n400256 , n400257 , n400258 , n400259 , n400260 , n400261 , n400262 , 
 n400263 , n400264 , n400265 , n400266 , n400267 , n400268 , n400269 , n400270 , n400271 , n400272 , 
 n400273 , n400274 , n400275 , n400276 , n400277 , n400278 , n400279 , n400280 , n78936 , n400282 , 
 n400283 , n400284 , n78940 , n400286 , n400287 , n400288 , n400289 , n400290 , n400291 , n400292 , 
 n400293 , n400294 , n400295 , n400296 , n400297 , n400298 , n400299 , n400300 , n400301 , n400302 , 
 n400303 , n400304 , n400305 , n400306 , n400307 , n400308 , n400309 , n400310 , n400311 , n400312 , 
 n400313 , n400314 , n400315 , n400316 , n78950 , n400318 , n400319 , n400320 , n400321 , n400322 , 
 n400323 , n400324 , n400325 , n400326 , n78960 , n400328 , n78962 , n400330 , n78964 , n400332 , 
 n400333 , n78967 , n400335 , n400336 , n400337 , n400338 , n400339 , n400340 , n400341 , n400342 , 
 n400343 , n400344 , n400345 , n400346 , n400347 , n400348 , n78982 , n78983 , n78984 , n78985 , 
 n78986 , n78987 , n400355 , n400356 , n400357 , n400358 , n400359 , n78993 , n400361 , n78995 , 
 n78996 , n78997 , n400365 , n78999 , n79000 , n400368 , n79002 , n400370 , n79004 , n400372 , 
 n400373 , n79007 , n400375 , n79009 , n79010 , n400378 , n400379 , n400380 , n400381 , n400382 , 
 n79016 , n400384 , n79018 , n79019 , n79020 , n79021 , n79022 , n79023 , n79024 , n400392 , 
 n79026 , n400394 , n79028 , n400396 , n400397 , n400398 , n400399 , n400400 , n400401 , n400402 , 
 n400403 , n400404 , n400405 , n400406 , n79040 , n400408 , n400409 , n400410 , n400411 , n400412 , 
 n79046 , n400414 , n400415 , n79049 , n400417 , n400418 , n79052 , n400420 , n400421 , n79055 , 
 n400423 , n400424 , n400425 , n400426 , n400427 , n79061 , n400429 , n400430 , n400431 , n400432 , 
 n400433 , n400434 , n79068 , n400436 , n400437 , n79071 , n400439 , n400440 , n400441 , n79075 , 
 n400443 , n400444 , n79078 , n400446 , n400447 , n79081 , n400449 , n400450 , n79084 , n79085 , 
 n400453 , n400454 , n400455 , n79089 , n400457 , n400458 , n400459 , n400460 , n400461 , n400462 , 
 n400463 , n400464 , n79098 , n400466 , n400467 , n400468 , n79102 , n400470 , n400471 , n400472 , 
 n400473 , n400474 , n400475 , n400476 , n400477 , n400478 , n400479 , n400480 , n79114 , n400482 , 
 n400483 , n79117 , n400485 , n400486 , n400487 , n400488 , n400489 , n79123 , n400491 , n400492 , 
 n400493 , n400494 , n400495 , n79129 , n79130 , n79131 , n400499 , n400500 , n79134 , n400502 , 
 n400503 , n400504 , n400505 , n79139 , n400507 , n400508 , n400509 , n400510 , n400511 , n400512 , 
 n400513 , n400514 , n400515 , n400516 , n400517 , n400518 , n400519 , n400520 , n79154 , n400522 , 
 n400523 , n400524 , n79158 , n400526 , n400527 , n400528 , n400529 , n400530 , n79164 , n400532 , 
 n400533 , n400534 , n400535 , n79169 , n400537 , n400538 , n79172 , n400540 , n400541 , n400542 , 
 n79176 , n79177 , n400545 , n79179 , n79180 , n400548 , n400549 , n400550 , n400551 , n400552 , 
 n400553 , n79187 , n400555 , n400556 , n400557 , n400558 , n400559 , n400560 , n79194 , n79195 , 
 n400563 , n400564 , n400565 , n400566 , n79199 , n400568 , n400569 , n79202 , n400571 , n400572 , 
 n400573 , n400574 , n400575 , n79205 , n400577 , n400578 , n79208 , n79209 , n400581 , n400582 , 
 n400583 , n79213 , n79214 , n79215 , n400587 , n79217 , n79218 , n400590 , n400591 , n79221 , 
 n79222 , n400594 , n79224 , n79225 , n400597 , n400598 , n400599 , n79229 , n400601 , n400602 , 
 n79232 , n79233 , n400605 , n400606 , n400607 , n79237 , n400609 , n400610 , n400611 , n79241 , 
 n79242 , n400614 , n400615 , n79245 , n400617 , n400618 , n79248 , n400620 , n400621 , n79251 , 
 n400623 , n400624 , n400625 , n400626 , n400627 , n400628 , n400629 , n400630 , n400631 , n400632 , 
 n400633 , n400634 , n400635 , n79265 , n400637 , n400638 , n79268 , n79269 , n400641 , n400642 , 
 n400643 , n400644 , n400645 , n400646 , n79276 , n79277 , n400649 , n400650 , n400651 , n79281 , 
 n400653 , n400654 , n400655 , n79285 , n400657 , n400658 , n79288 , n79289 , n400661 , n400662 , 
 n400663 , n400664 , n400665 , n400666 , n400667 , n400668 , n400669 , n400670 , n400671 , n400672 , 
 n400673 , n400674 , n400675 , n400676 , n400677 , n400678 , n400679 , n400680 , n400681 , n400682 , 
 n400683 , n79299 , n79300 , n400686 , n400687 , n400688 , n79304 , n400690 , n400691 , n79307 , 
 n79308 , n400694 , n79310 , n400696 , n79312 , n400698 , n400699 , n400700 , n400701 , n79317 , 
 n79318 , n400704 , n400705 , n400706 , n400707 , n79323 , n79324 , n400710 , n79326 , n400712 , 
 n400713 , n79329 , n400715 , n400716 , n79332 , n79333 , n400719 , n400720 , n400721 , n79337 , 
 n400723 , n400724 , n79340 , n79341 , n400727 , n400728 , n400729 , n400730 , n79346 , n400732 , 
 n400733 , n79349 , n79350 , n400736 , n400737 , n79353 , n79354 , n400740 , n400741 , n400742 , 
 n79358 , n400744 , n79360 , n400746 , n400747 , n400748 , n400749 , n400750 , n400751 , n400752 , 
 n400753 , n400754 , n400755 , n400756 , n79372 , n400758 , n400759 , n400760 , n79376 , n79377 , 
 n400763 , n400764 , n400765 , n400766 , n400767 , n400768 , n79384 , n400770 , n400771 , n400772 , 
 n79388 , n400774 , n79390 , n400776 , n400777 , n400778 , n79394 , n400780 , n400781 , n400782 , 
 n400783 , n400784 , n79400 , n400786 , n400787 , n79403 , n400789 , n400790 , n400791 , n400792 , 
 n400793 , n400794 , n400795 , n400796 , n79412 , n400798 , n400799 , n79415 , n400801 , n400802 , 
 n400803 , n400804 , n400805 , n79421 , n79422 , n400808 , n400809 , n400810 , n400811 , n79427 , 
 n400813 , n400814 , n400815 , n400816 , n400817 , n79433 , n79434 , n400820 , n400821 , n400822 , 
 n400823 , n400824 , n79440 , n400826 , n400827 , n79443 , n400829 , n79445 , n400831 , n79447 , 
 n79448 , n400834 , n400835 , n400836 , n79452 , n400838 , n400839 , n400840 , n79456 , n79457 , 
 n400843 , n400844 , n400845 , n400846 , n400847 , n79463 , n400849 , n400850 , n400851 , n400852 , 
 n400853 , n79469 , n400855 , n400856 , n400857 , n400858 , n400859 , n400860 , n400861 , n79477 , 
 n400863 , n400864 , n400865 , n79481 , n79482 , n400868 , n79484 , n400870 , n400871 , n400872 , 
 n400873 , n79489 , n79490 , n400876 , n400877 , n400878 , n400879 , n400880 , n400881 , n400882 , 
 n400883 , n79499 , n79500 , n400886 , n400887 , n400888 , n79504 , n79505 , n400891 , n400892 , 
 n400893 , n400894 , n79510 , n79511 , n400897 , n400898 , n400899 , n79515 , n400901 , n79517 , 
 n79518 , n400904 , n400905 , n79521 , n400907 , n400908 , n79524 , n400910 , n400911 , n400912 , 
 n400913 , n400914 , n79530 , n400916 , n400917 , n400918 , n79534 , n400920 , n400921 , n79537 , 
 n79538 , n400924 , n79540 , n400926 , n400927 , n400928 , n400929 , n400930 , n79546 , n79547 , 
 n400933 , n400934 , n79550 , n400936 , n400937 , n400938 , n400939 , n400940 , n400941 , n400942 , 
 n400943 , n400944 , n400945 , n400946 , n400947 , n400948 , n400949 , n400950 , n400951 , n400952 , 
 n400953 , n400954 , n400955 , n400956 , n400957 , n400958 , n400959 , n400960 , n400961 , n400962 , 
 n400963 , n400964 , n400965 , n400966 , n400967 , n79558 , n400969 , n400970 , n79561 , n400972 , 
 n79563 , n400974 , n400975 , n400976 , n400977 , n400978 , n400979 , n79570 , n79571 , n79572 , 
 n400983 , n79574 , n79575 , n400986 , n400987 , n400988 , n400989 , n400990 , n400991 , n400992 , 
 n400993 , n400994 , n400995 , n400996 , n400997 , n400998 , n400999 , n401000 , n401001 , n401002 , 
 n401003 , n401004 , n401005 , n401006 , n401007 , n401008 , n401009 , n79581 , n401011 , n401012 , 
 n401013 , n79585 , n401015 , n401016 , n401017 , n401018 , n79590 , n401020 , n401021 , n401022 , 
 n401023 , n401024 , n79596 , n401026 , n401027 , n79599 , n401029 , n401030 , n401031 , n401032 , 
 n401033 , n401034 , n401035 , n401036 , n401037 , n401038 , n401039 , n401040 , n401041 , n79613 , 
 n79614 , n401044 , n401045 , n79617 , n79618 , n79619 , n401049 , n401050 , n79622 , n79623 , 
 n79624 , n401054 , n401055 , n401056 , n401057 , n79629 , n401059 , n401060 , n401061 , n401062 , 
 n401063 , n401064 , n401065 , n401066 , n79638 , n79639 , n401069 , n401070 , n79642 , n401072 , 
 n401073 , n401074 , n79646 , n401076 , n401077 , n401078 , n401079 , n401080 , n401081 , n401082 , 
 n401083 , n401084 , n401085 , n79657 , n401087 , n401088 , n401089 , n401090 , n401091 , n79663 , 
 n401093 , n401094 , n401095 , n79667 , n79668 , n401098 , n79670 , n401100 , n401101 , n79673 , 
 n401103 , n401104 , n401105 , n79677 , n401107 , n79679 , n79680 , n401110 , n79682 , n401112 , 
 n79684 , n79685 , n401115 , n401116 , n401117 , n79689 , n401119 , n79691 , n79692 , n401122 , 
 n401123 , n401124 , n401125 , n401126 , n401127 , n401128 , n401129 , n401130 , n401131 , n401132 , 
 n401133 , n401134 , n401135 , n401136 , n401137 , n401138 , n401139 , n401140 , n401141 , n79713 , 
 n401143 , n79715 , n401145 , n401146 , n401147 , n401148 , n79720 , n401150 , n401151 , n79723 , 
 n401153 , n401154 , n401155 , n401156 , n401157 , n401158 , n401159 , n401160 , n79732 , n401162 , 
 n401163 , n401164 , n401165 , n401166 , n401167 , n401168 , n401169 , n79741 , n79742 , n401172 , 
 n401173 , n79745 , n401175 , n401176 , n79748 , n401178 , n401179 , n401180 , n79752 , n401182 , 
 n401183 , n401184 , n401185 , n401186 , n401187 , n401188 , n401189 , n401190 , n79762 , n401192 , 
 n79764 , n79765 , n401195 , n401196 , n79768 , n401198 , n401199 , n401200 , n401201 , n401202 , 
 n401203 , n79775 , n401205 , n401206 , n401207 , n401208 , n79780 , n401210 , n401211 , n79783 , 
 n401213 , n401214 , n401215 , n401216 , n401217 , n79789 , n401219 , n401220 , n79792 , n401222 , 
 n79794 , n401224 , n401225 , n401226 , n79798 , n401228 , n401229 , n79801 , n401231 , n401232 , 
 n401233 , n401234 , n401235 , n401236 , n401237 , n401238 , n79810 , n401240 , n79812 , n79813 , 
 n401243 , n401244 , n79816 , n401246 , n401247 , n401248 , n401249 , n401250 , n401251 , n79823 , 
 n401253 , n401254 , n401255 , n401256 , n401257 , n401258 , n401259 , n79831 , n401261 , n401262 , 
 n79834 , n79835 , n79836 , n401266 , n401267 , n79839 , n79840 , n79841 , n401271 , n401272 , 
 n401273 , n401274 , n79846 , n79847 , n401277 , n79849 , n401279 , n401280 , n401281 , n401282 , 
 n401283 , n401284 , n79856 , n401286 , n401287 , n401288 , n401289 , n401290 , n79862 , n401292 , 
 n401293 , n79865 , n401295 , n401296 , n79868 , n401298 , n79870 , n401300 , n401301 , n401302 , 
 n401303 , n401304 , n79876 , n401306 , n401307 , n401308 , n401309 , n401310 , n401311 , n401312 , 
 n79884 , n401314 , n401315 , n401316 , n79888 , n401318 , n401319 , n401320 , n401321 , n401322 , 
 n79894 , n401324 , n401325 , n401326 , n79898 , n401328 , n401329 , n401330 , n79902 , n79903 , 
 n401333 , n401334 , n79906 , n79907 , n401337 , n401338 , n401339 , n401340 , n401341 , n401342 , 
 n401343 , n401344 , n401345 , n401346 , n79918 , n401348 , n401349 , n79921 , n401351 , n401352 , 
 n401353 , n401354 , n79926 , n401356 , n401357 , n401358 , n401359 , n401360 , n401361 , n79933 , 
 n401363 , n401364 , n79936 , n401366 , n401367 , n79939 , n401369 , n401370 , n401371 , n401372 , 
 n79944 , n79945 , n401375 , n79947 , n401377 , n401378 , n401379 , n401380 , n79952 , n401382 , 
 n401383 , n79955 , n401385 , n401386 , n401387 , n79959 , n79960 , n401390 , n79962 , n79963 , 
 n401393 , n401394 , n401395 , n401396 , n401397 , n401398 , n401399 , n401400 , n401401 , n401402 , 
 n401403 , n401404 , n401405 , n401406 , n401407 , n401408 , n401409 , n401410 , n401411 , n401412 , 
 n79984 , n401414 , n401415 , n79987 , n401417 , n401418 , n401419 , n401420 , n401421 , n401422 , 
 n401423 , n79995 , n401425 , n401426 , n401427 , n79999 , n401429 , n80001 , n401431 , n401432 , 
 n401433 , n401434 , n401435 , n401436 , n401437 , n401438 , n401439 , n80011 , n80012 , n401442 , 
 n401443 , n401444 , n80016 , n401446 , n401447 , n401448 , n401449 , n401450 , n401451 , n401452 , 
 n401453 , n401454 , n401455 , n401456 , n401457 , n401458 , n401459 , n401460 , n401461 , n401462 , 
 n401463 , n401464 , n401465 , n401466 , n401467 , n401468 , n401469 , n401470 , n401471 , n80022 , 
 n401473 , n401474 , n401475 , n80026 , n401477 , n401478 , n80029 , n80030 , n80031 , n401482 , 
 n401483 , n80034 , n401485 , n401486 , n401487 , n80038 , n80039 , n401490 , n80041 , n80042 , 
 n401493 , n401494 , n80045 , n401496 , n401497 , n80048 , n80049 , n401500 , n401501 , n401502 , 
 n80053 , n401504 , n401505 , n80056 , n401507 , n401508 , n401509 , n401510 , n401511 , n401512 , 
 n401513 , n80064 , n401515 , n401516 , n80067 , n401518 , n401519 , n401520 , n401521 , n401522 , 
 n401523 , n80074 , n401525 , n401526 , n80077 , n401528 , n401529 , n401530 , n80081 , n401532 , 
 n401533 , n401534 , n80085 , n401536 , n401537 , n401538 , n401539 , n401540 , n401541 , n401542 , 
 n80093 , n401544 , n401545 , n80096 , n401547 , n401548 , n80099 , n401550 , n401551 , n401552 , 
 n401553 , n401554 , n401555 , n401556 , n80107 , n401558 , n401559 , n401560 , n401561 , n401562 , 
 n401563 , n401564 , n401565 , n401566 , n401567 , n401568 , n401569 , n401570 , n401571 , n401572 , 
 n401573 , n401574 , n401575 , n80126 , n401577 , n401578 , n401579 , n401580 , n401581 , n80132 , 
 n401583 , n401584 , n80135 , n401586 , n401587 , n401588 , n80139 , n401590 , n401591 , n401592 , 
 n80143 , n401594 , n401595 , n80146 , n401597 , n401598 , n401599 , n80150 , n401601 , n401602 , 
 n401603 , n401604 , n401605 , n80156 , n401607 , n80158 , n80159 , n80160 , n401611 , n401612 , 
 n401613 , n80164 , n401615 , n80166 , n401617 , n80168 , n401619 , n401620 , n401621 , n401622 , 
 n401623 , n80174 , n80175 , n401626 , n401627 , n401628 , n401629 , n401630 , n80181 , n80182 , 
 n401633 , n80184 , n401635 , n401636 , n80187 , n401638 , n401639 , n401640 , n401641 , n401642 , 
 n80193 , n401644 , n401645 , n401646 , n401647 , n401648 , n80199 , n401650 , n401651 , n80202 , 
 n401653 , n401654 , n401655 , n401656 , n401657 , n401658 , n401659 , n401660 , n401661 , n401662 , 
 n401663 , n401664 , n401665 , n80216 , n401667 , n401668 , n80219 , n401670 , n401671 , n401672 , 
 n401673 , n401674 , n80225 , n401676 , n401677 , n401678 , n401679 , n401680 , n401681 , n401682 , 
 n401683 , n401684 , n401685 , n401686 , n401687 , n80238 , n401689 , n401690 , n401691 , n401692 , 
 n401693 , n80244 , n401695 , n401696 , n80247 , n401698 , n401699 , n80250 , n401701 , n401702 , 
 n401703 , n401704 , n401705 , n401706 , n401707 , n401708 , n401709 , n401710 , n401711 , n401712 , 
 n80263 , n401714 , n80265 , n80266 , n80267 , n401718 , n401719 , n401720 , n401721 , n80272 , 
 n401723 , n80274 , n401725 , n401726 , n80277 , n401728 , n80279 , n80280 , n401731 , n401732 , 
 n80283 , n401734 , n401735 , n80286 , n401737 , n401738 , n401739 , n80290 , n401741 , n401742 , 
 n80293 , n401744 , n401745 , n401746 , n80297 , n80298 , n80299 , n401750 , n401751 , n401752 , 
 n401753 , n401754 , n80305 , n401756 , n401757 , n80308 , n401759 , n401760 , n401761 , n401762 , 
 n401763 , n401764 , n401765 , n80316 , n401767 , n401768 , n401769 , n80320 , n401771 , n401772 , 
 n401773 , n401774 , n401775 , n80326 , n401777 , n401778 , n401779 , n80330 , n401781 , n80332 , 
 n401783 , n401784 , n401785 , n401786 , n401787 , n401788 , n401789 , n401790 , n401791 , n401792 , 
 n401793 , n401794 , n401795 , n80346 , n401797 , n401798 , n80349 , n80350 , n401801 , n80352 , 
 n401803 , n401804 , n401805 , n401806 , n401807 , n401808 , n80359 , n401810 , n401811 , n401812 , 
 n80363 , n401814 , n401815 , n401816 , n80367 , n401818 , n401819 , n80370 , n401821 , n401822 , 
 n401823 , n401824 , n401825 , n80376 , n401827 , n401828 , n401829 , n401830 , n80381 , n401832 , 
 n401833 , n401834 , n401835 , n401836 , n401837 , n401838 , n401839 , n401840 , n401841 , n401842 , 
 n401843 , n401844 , n80395 , n401846 , n401847 , n401848 , n80399 , n401850 , n401851 , n401852 , 
 n80403 , n401854 , n401855 , n80406 , n401857 , n401858 , n401859 , n401860 , n80411 , n401862 , 
 n401863 , n401864 , n80415 , n401866 , n401867 , n401868 , n401869 , n401870 , n80421 , n401872 , 
 n401873 , n80424 , n401875 , n401876 , n80427 , n80428 , n401879 , n401880 , n401881 , n401882 , 
 n401883 , n80434 , n401885 , n401886 , n401887 , n80438 , n401889 , n401890 , n401891 , n401892 , 
 n401893 , n401894 , n80445 , n401896 , n401897 , n401898 , n401899 , n401900 , n401901 , n401902 , 
 n401903 , n401904 , n401905 , n401906 , n401907 , n401908 , n401909 , n401910 , n401911 , n80462 , 
 n80463 , n401914 , n80465 , n80466 , n80467 , n80468 , n401919 , n401920 , n401921 , n401922 , 
 n401923 , n401924 , n401925 , n401926 , n401927 , n401928 , n401929 , n401930 , n401931 , n401932 , 
 n80483 , n401934 , n401935 , n80486 , n401937 , n401938 , n401939 , n401940 , n401941 , n401942 , 
 n80493 , n80494 , n401945 , n401946 , n401947 , n401948 , n401949 , n401950 , n80501 , n401952 , 
 n401953 , n401954 , n401955 , n401956 , n401957 , n401958 , n401959 , n401960 , n401961 , n401962 , 
 n401963 , n80514 , n80515 , n80516 , n80517 , n80518 , n80519 , n80520 , n80521 , n401972 , 
 n401973 , n401974 , n401975 , n401976 , n401977 , n80528 , n401979 , n401980 , n401981 , n401982 , 
 n80533 , n401984 , n401985 , n80536 , n401987 , n401988 , n80539 , n80540 , n401991 , n401992 , 
 n401993 , n80544 , n80545 , n401996 , n401997 , n80548 , n80549 , n402000 , n402001 , n402002 , 
 n80553 , n402004 , n402005 , n402006 , n402007 , n402008 , n402009 , n402010 , n402011 , n402012 , 
 n402013 , n80564 , n80565 , n402016 , n402017 , n80568 , n402019 , n402020 , n402021 , n402022 , 
 n402023 , n80574 , n402025 , n402026 , n402027 , n402028 , n80579 , n402030 , n402031 , n402032 , 
 n402033 , n402034 , n80585 , n80586 , n402037 , n402038 , n402039 , n402040 , n402041 , n402042 , 
 n402043 , n402044 , n80595 , n402046 , n402047 , n402048 , n402049 , n402050 , n80601 , n402052 , 
 n402053 , n402054 , n402055 , n80606 , n402057 , n402058 , n80609 , n402060 , n402061 , n402062 , 
 n80613 , n402064 , n402065 , n80616 , n80617 , n80618 , n402069 , n402070 , n80621 , n402072 , 
 n402073 , n402074 , n402075 , n402076 , n80627 , n402078 , n402079 , n402080 , n402081 , n402082 , 
 n402083 , n80634 , n402085 , n80636 , n80637 , n402088 , n402089 , n80640 , n402091 , n402092 , 
 n80643 , n402094 , n402095 , n402096 , n402097 , n80648 , n80649 , n402100 , n402101 , n80652 , 
 n402103 , n402104 , n402105 , n402106 , n402107 , n402108 , n80659 , n80660 , n402111 , n402112 , 
 n402113 , n80664 , n402115 , n402116 , n402117 , n80668 , n402119 , n402120 , n402121 , n402122 , 
 n402123 , n402124 , n80675 , n402126 , n402127 , n402128 , n402129 , n80680 , n402131 , n402132 , 
 n80683 , n80684 , n402135 , n402136 , n402137 , n80688 , n402139 , n80690 , n402141 , n402142 , 
 n402143 , n80694 , n80695 , n402146 , n80697 , n80698 , n80699 , n80700 , n402151 , n402152 , 
 n402153 , n80704 , n80705 , n402156 , n402157 , n80708 , n80709 , n402160 , n80711 , n80712 , 
 n80713 , n402164 , n80715 , n80716 , n80717 , n80718 , n80719 , n80720 , n80721 , n80722 , 
 n80723 , n80724 , n80725 , n80726 , n80727 , n402178 , n80729 , n402180 , n80731 , n80732 , 
 n402183 , n80734 , n402185 , n402186 , n402187 , n402188 , n402189 , n402190 , n402191 , n402192 , 
 n402193 , n402194 , n402195 , n402196 , n402197 , n402198 , n402199 , n402200 , n402201 , n402202 , 
 n402203 , n402204 , n402205 , n402206 , n80742 , n402208 , n402209 , n402210 , n402211 , n402212 , 
 n402213 , n402214 , n402215 , n402216 , n402217 , n402218 , n80754 , n402220 , n402221 , n402222 , 
 n402223 , n402224 , n402225 , n80761 , n402227 , n402228 , n402229 , n80765 , n402231 , n402232 , 
 n402233 , n402234 , n402235 , n402236 , n402237 , n80773 , n402239 , n402240 , n402241 , n402242 , 
 n402243 , n402244 , n80780 , n402246 , n402247 , n80783 , n402249 , n80785 , n80786 , n402252 , 
 n402253 , n80789 , n402255 , n402256 , n402257 , n402258 , n402259 , n80795 , n402261 , n402262 , 
 n402263 , n402264 , n80800 , n402266 , n402267 , n402268 , n402269 , n80805 , n402271 , n402272 , 
 n80808 , n80809 , n402275 , n80811 , n402277 , n402278 , n402279 , n402280 , n402281 , n402282 , 
 n80818 , n402284 , n402285 , n402286 , n80822 , n402288 , n402289 , n402290 , n402291 , n402292 , 
 n80828 , n402294 , n80830 , n402296 , n402297 , n402298 , n80834 , n80835 , n80836 , n80837 , 
 n80838 , n402304 , n80840 , n402306 , n402307 , n80843 , n402309 , n402310 , n402311 , n402312 , 
 n402313 , n402314 , n402315 , n402316 , n402317 , n402318 , n402319 , n80855 , n402321 , n402322 , 
 n80858 , n402324 , n402325 , n80861 , n402327 , n402328 , n402329 , n402330 , n402331 , n402332 , 
 n402333 , n402334 , n402335 , n80871 , n80872 , n402338 , n402339 , n402340 , n402341 , n402342 , 
 n402343 , n80879 , n80880 , n402346 , n402347 , n80883 , n402349 , n80885 , n402351 , n402352 , 
 n402353 , n80889 , n402355 , n402356 , n402357 , n402358 , n402359 , n80895 , n402361 , n402362 , 
 n80898 , n80899 , n402365 , n80901 , n402367 , n402368 , n402369 , n402370 , n402371 , n402372 , 
 n402373 , n402374 , n402375 , n402376 , n80912 , n80913 , n402379 , n402380 , n80916 , n80917 , 
 n80918 , n402384 , n402385 , n80921 , n80922 , n402388 , n402389 , n402390 , n80926 , n402392 , 
 n402393 , n402394 , n402395 , n402396 , n402397 , n402398 , n402399 , n402400 , n402401 , n402402 , 
 n402403 , n402404 , n402405 , n402406 , n402407 , n402408 , n402409 , n402410 , n402411 , n402412 , 
 n402413 , n402414 , n402415 , n402416 , n402417 , n402418 , n402419 , n402420 , n402421 , n80932 , 
 n80933 , n402424 , n402425 , n402426 , n402427 , n80937 , n402429 , n402430 , n402431 , n402432 , 
 n402433 , n402434 , n402435 , n402436 , n80946 , n402438 , n402439 , n402440 , n402441 , n80951 , 
 n402443 , n402444 , n80954 , n402446 , n402447 , n402448 , n80958 , n80959 , n402451 , n402452 , 
 n402453 , n402454 , n402455 , n80965 , n402457 , n402458 , n80968 , n402460 , n80970 , n402462 , 
 n402463 , n402464 , n402465 , n402466 , n402467 , n402468 , n402469 , n402470 , n402471 , n402472 , 
 n402473 , n402474 , n402475 , n402476 , n402477 , n402478 , n402479 , n402480 , n80990 , n402482 , 
 n80992 , n402484 , n402485 , n402486 , n402487 , n402488 , n402489 , n402490 , n402491 , n402492 , 
 n402493 , n402494 , n402495 , n402496 , n402497 , n81007 , n81008 , n81009 , n81010 , n81011 , 
 n402503 , n402504 , n402505 , n402506 , n81016 , n402508 , n402509 , n402510 , n402511 , n402512 , 
 n402513 , n402514 , n402515 , n402516 , n81026 , n402518 , n402519 , n81029 , n402521 , n402522 , 
 n81032 , n402524 , n402525 , n402526 , n402527 , n402528 , n402529 , n402530 , n81040 , n402532 , 
 n81042 , n402534 , n402535 , n402536 , n81046 , n402538 , n402539 , n402540 , n402541 , n402542 , 
 n402543 , n402544 , n402545 , n402546 , n402547 , n402548 , n81058 , n402550 , n402551 , n402552 , 
 n402553 , n402554 , n402555 , n81065 , n402557 , n402558 , n81068 , n81069 , n402561 , n402562 , 
 n402563 , n81073 , n402565 , n81075 , n402567 , n402568 , n81078 , n81079 , n81080 , n402572 , 
 n402573 , n81083 , n81084 , n402576 , n81086 , n402578 , n402579 , n402580 , n402581 , n402582 , 
 n402583 , n402584 , n402585 , n402586 , n402587 , n402588 , n402589 , n402590 , n402591 , n402592 , 
 n402593 , n402594 , n81090 , n402596 , n81092 , n402598 , n81094 , n402600 , n402601 , n402602 , 
 n402603 , n402604 , n402605 , n402606 , n402607 , n402608 , n402609 , n402610 , n402611 , n402612 , 
 n402613 , n402614 , n402615 , n81099 , n402617 , n402618 , n402619 , n81103 , n402621 , n402622 , 
 n402623 , n81107 , n81108 , n402626 , n402627 , n402628 , n402629 , n402630 , n81114 , n402632 , 
 n402633 , n81117 , n402635 , n402636 , n402637 , n402638 , n402639 , n402640 , n402641 , n402642 , 
 n402643 , n402644 , n402645 , n402646 , n402647 , n402648 , n402649 , n402650 , n402651 , n402652 , 
 n402653 , n81125 , n402655 , n402656 , n81128 , n402658 , n402659 , n402660 , n402661 , n402662 , 
 n81134 , n402664 , n402665 , n402666 , n402667 , n402668 , n402669 , n402670 , n402671 , n402672 , 
 n402673 , n402674 , n402675 , n81147 , n402677 , n402678 , n402679 , n81151 , n81152 , n402682 , 
 n402683 , n81155 , n402685 , n81157 , n402687 , n402688 , n81160 , n402690 , n81162 , n81163 , 
 n402693 , n402694 , n402695 , n402696 , n402697 , n81169 , n402699 , n402700 , n402701 , n402702 , 
 n402703 , n402704 , n402705 , n402706 , n81178 , n402708 , n402709 , n402710 , n402711 , n402712 , 
 n81184 , n402714 , n81186 , n81187 , n402717 , n402718 , n402719 , n402720 , n402721 , n402722 , 
 n402723 , n81195 , n402725 , n402726 , n81198 , n402728 , n402729 , n81201 , n402731 , n81203 , 
 n402733 , n81205 , n81206 , n81207 , n81208 , n81209 , n81210 , n81211 , n402741 , n81213 , 
 n402743 , n402744 , n402745 , n402746 , n402747 , n402748 , n402749 , n402750 , n402751 , n402752 , 
 n402753 , n81225 , n402755 , n402756 , n402757 , n402758 , n402759 , n81231 , n402761 , n81233 , 
 n402763 , n402764 , n402765 , n402766 , n402767 , n81239 , n402769 , n402770 , n81242 , n402772 , 
 n402773 , n402774 , n402775 , n402776 , n81248 , n402778 , n402779 , n402780 , n81252 , n402782 , 
 n402783 , n402784 , n402785 , n402786 , n402787 , n402788 , n81260 , n402790 , n402791 , n402792 , 
 n402793 , n402794 , n402795 , n81267 , n81268 , n402798 , n81270 , n402800 , n402801 , n402802 , 
 n402803 , n81275 , n402805 , n402806 , n402807 , n81279 , n402809 , n81281 , n402811 , n402812 , 
 n402813 , n402814 , n81286 , n81287 , n81288 , n402818 , n81290 , n81291 , n81292 , n81293 , 
 n81294 , n81295 , n81296 , n402826 , n81298 , n81299 , n81300 , n81301 , n81302 , n81303 , 
 n81304 , n81305 , n81306 , n402836 , n402837 , n402838 , n402839 , n402840 , n402841 , n402842 , 
 n81314 , n81315 , n402845 , n402846 , n402847 , n402848 , n402849 , n402850 , n402851 , n402852 , 
 n402853 , n402854 , n402855 , n402856 , n402857 , n402858 , n402859 , n402860 , n81332 , n402862 , 
 n402863 , n81335 , n402865 , n402866 , n81338 , n402868 , n402869 , n81341 , n402871 , n402872 , 
 n402873 , n402874 , n402875 , n402876 , n402877 , n81349 , n402879 , n402880 , n81352 , n81353 , 
 n81354 , n81355 , n81356 , n402886 , n402887 , n402888 , n81360 , n402890 , n402891 , n402892 , 
 n402893 , n402894 , n402895 , n402896 , n402897 , n81369 , n402899 , n402900 , n81372 , n402902 , 
 n81374 , n81375 , n402905 , n402906 , n402907 , n402908 , n402909 , n402910 , n402911 , n402912 , 
 n81384 , n402914 , n402915 , n402916 , n402917 , n402918 , n81390 , n81391 , n402921 , n402922 , 
 n81394 , n81395 , n402925 , n81397 , n81398 , n402928 , n81400 , n402930 , n402931 , n402932 , 
 n402933 , n402934 , n402935 , n402936 , n402937 , n402938 , n402939 , n81408 , n402941 , n402942 , 
 n402943 , n402944 , n402945 , n402946 , n402947 , n402948 , n402949 , n402950 , n402951 , n402952 , 
 n402953 , n402954 , n402955 , n402956 , n402957 , n402958 , n402959 , n402960 , n402961 , n402962 , 
 n402963 , n402964 , n402965 , n402966 , n402967 , n402968 , n402969 , n402970 , n402971 , n402972 , 
 n402973 , n81422 , n402975 , n81424 , n81425 , n402978 , n402979 , n402980 , n402981 , n81430 , 
 n402983 , n402984 , n402985 , n402986 , n81435 , n402988 , n402989 , n402990 , n402991 , n81440 , 
 n402993 , n402994 , n402995 , n402996 , n81445 , n402998 , n402999 , n403000 , n403001 , n403002 , 
 n403003 , n403004 , n403005 , n403006 , n403007 , n403008 , n403009 , n403010 , n403011 , n403012 , 
 n403013 , n403014 , n403015 , n403016 , n403017 , n403018 , n403019 , n403020 , n403021 , n403022 , 
 n403023 , n403024 , n403025 , n403026 , n403027 , n403028 , n403029 , n403030 , n81451 , n403032 , 
 n403033 , n403034 , n403035 , n403036 , n403037 , n403038 , n403039 , n403040 , n403041 , n403042 , 
 n403043 , n81461 , n403045 , n403046 , n403047 , n81465 , n403049 , n403050 , n403051 , n403052 , 
 n403053 , n403054 , n403055 , n403056 , n403057 , n403058 , n403059 , n403060 , n403061 , n81479 , 
 n403063 , n403064 , n403065 , n403066 , n403067 , n403068 , n403069 , n403070 , n403071 , n81489 , 
 n403073 , n403074 , n81492 , n81493 , n403077 , n81495 , n403079 , n403080 , n403081 , n403082 , 
 n403083 , n403084 , n403085 , n81503 , n403087 , n81505 , n81506 , n403090 , n403091 , n81509 , 
 n403093 , n403094 , n403095 , n403096 , n403097 , n403098 , n403099 , n403100 , n81518 , n403102 , 
 n403103 , n403104 , n403105 , n403106 , n403107 , n403108 , n403109 , n403110 , n403111 , n81529 , 
 n403113 , n403114 , n403115 , n403116 , n403117 , n403118 , n403119 , n403120 , n403121 , n403122 , 
 n81540 , n403124 , n403125 , n403126 , n403127 , n403128 , n403129 , n403130 , n403131 , n403132 , 
 n403133 , n403134 , n81549 , n403136 , n403137 , n403138 , n403139 , n403140 , n81555 , n403142 , 
 n403143 , n81558 , n403145 , n403146 , n403147 , n81562 , n403149 , n403150 , n81565 , n403152 , 
 n403153 , n403154 , n403155 , n403156 , n403157 , n403158 , n403159 , n81574 , n403161 , n403162 , 
 n403163 , n403164 , n403165 , n403166 , n403167 , n403168 , n403169 , n403170 , n403171 , n403172 , 
 n403173 , n403174 , n403175 , n403176 , n403177 , n403178 , n403179 , n403180 , n403181 , n403182 , 
 n403183 , n403184 , n403185 , n81579 , n81580 , n403188 , n81582 , n403190 , n403191 , n403192 , 
 n403193 , n403194 , n403195 , n403196 , n403197 , n403198 , n403199 , n403200 , n403201 , n403202 , 
 n403203 , n403204 , n403205 , n403206 , n403207 , n403208 , n403209 , n403210 , n403211 , n403212 , 
 n403213 , n403214 , n403215 , n403216 , n403217 , n403218 , n403219 , n81586 , n403221 , n403222 , 
 n81587 , n403224 , n403225 , n403226 , n81591 , n81592 , n403229 , n403230 , n81595 , n403232 , 
 n403233 , n403234 , n403235 , n403236 , n403237 , n403238 , n81603 , n403240 , n403241 , n81606 , 
 n81607 , n403244 , n81609 , n403246 , n403247 , n403248 , n403249 , n403250 , n403251 , n403252 , 
 n81617 , n81618 , n403255 , n403256 , n403257 , n403258 , n403259 , n403260 , n81625 , n403262 , 
 n403263 , n403264 , n81629 , n403266 , n403267 , n403268 , n403269 , n403270 , n403271 , n403272 , 
 n81637 , n81638 , n403275 , n403276 , n81641 , n403278 , n403279 , n403280 , n81645 , n403282 , 
 n403283 , n403284 , n403285 , n81650 , n403287 , n403288 , n81653 , n403290 , n403291 , n403292 , 
 n403293 , n403294 , n403295 , n403296 , n403297 , n81662 , n403299 , n403300 , n403301 , n81666 , 
 n403303 , n403304 , n403305 , n81670 , n81671 , n403308 , n81673 , n403310 , n403311 , n81676 , 
 n403313 , n403314 , n403315 , n403316 , n81681 , n403318 , n403319 , n403320 , n403321 , n403322 , 
 n403323 , n81688 , n403325 , n403326 , n403327 , n403328 , n403329 , n403330 , n81695 , n403332 , 
 n403333 , n403334 , n81699 , n403336 , n403337 , n81702 , n403339 , n403340 , n403341 , n403342 , 
 n403343 , n81708 , n403345 , n403346 , n403347 , n403348 , n81713 , n403350 , n403351 , n403352 , 
 n81717 , n403354 , n403355 , n403356 , n403357 , n403358 , n403359 , n403360 , n81725 , n403362 , 
 n403363 , n81728 , n403365 , n81730 , n81731 , n403368 , n403369 , n81734 , n403371 , n403372 , 
 n403373 , n81738 , n403375 , n403376 , n403377 , n403378 , n81743 , n403380 , n403381 , n81746 , 
 n81747 , n403384 , n403385 , n403386 , n81751 , n403388 , n81753 , n403390 , n403391 , n403392 , 
 n81757 , n403394 , n403395 , n81760 , n403397 , n81762 , n403399 , n81764 , n403401 , n403402 , 
 n403403 , n81768 , n403405 , n403406 , n81771 , n403408 , n403409 , n403410 , n403411 , n81776 , 
 n403413 , n403414 , n403415 , n81780 , n81781 , n403418 , n403419 , n403420 , n403421 , n403422 , 
 n403423 , n403424 , n403425 , n403426 , n403427 , n403428 , n403429 , n403430 , n403431 , n403432 , 
 n81797 , n81798 , n81799 , n403436 , n403437 , n403438 , n81803 , n81804 , n403441 , n403442 , 
 n81807 , n403444 , n403445 , n403446 , n403447 , n403448 , n403449 , n403450 , n81815 , n403452 , 
 n403453 , n81818 , n403455 , n403456 , n403457 , n403458 , n81823 , n403460 , n403461 , n403462 , 
 n403463 , n403464 , n81829 , n81830 , n403467 , n403468 , n81833 , n403470 , n403471 , n403472 , 
 n403473 , n403474 , n81839 , n403476 , n403477 , n81842 , n81843 , n403480 , n403481 , n403482 , 
 n81847 , n81848 , n81849 , n403486 , n81851 , n81852 , n403489 , n403490 , n81855 , n403492 , 
 n403493 , n81858 , n403495 , n403496 , n81861 , n81862 , n81863 , n81864 , n403501 , n403502 , 
 n81867 , n403504 , n403505 , n403506 , n81871 , n403508 , n81873 , n403510 , n403511 , n403512 , 
 n403513 , n403514 , n81879 , n403516 , n403517 , n403518 , n403519 , n403520 , n403521 , n403522 , 
 n403523 , n403524 , n403525 , n403526 , n81891 , n403528 , n403529 , n403530 , n403531 , n403532 , 
 n403533 , n403534 , n403535 , n403536 , n403537 , n403538 , n81903 , n403540 , n403541 , n403542 , 
 n403543 , n403544 , n403545 , n403546 , n81911 , n81912 , n403549 , n403550 , n403551 , n403552 , 
 n403553 , n403554 , n403555 , n403556 , n81921 , n81922 , n403559 , n403560 , n403561 , n403562 , 
 n403563 , n403564 , n81929 , n403566 , n403567 , n403568 , n403569 , n81934 , n403571 , n403572 , 
 n403573 , n81938 , n81939 , n403576 , n403577 , n81942 , n403579 , n403580 , n403581 , n81946 , 
 n403583 , n403584 , n81949 , n81950 , n403587 , n81952 , n403589 , n403590 , n403591 , n403592 , 
 n403593 , n403594 , n81959 , n403596 , n403597 , n403598 , n403599 , n403600 , n403601 , n403602 , 
 n403603 , n403604 , n403605 , n403606 , n403607 , n403608 , n403609 , n403610 , n403611 , n403612 , 
 n403613 , n81967 , n403615 , n403616 , n403617 , n403618 , n403619 , n81973 , n403621 , n403622 , 
 n403623 , n403624 , n403625 , n403626 , n403627 , n403628 , n403629 , n81983 , n403631 , n403632 , 
 n403633 , n81987 , n403635 , n403636 , n403637 , n81991 , n403639 , n403640 , n403641 , n81995 , 
 n403643 , n81997 , n403645 , n403646 , n403647 , n82001 , n403649 , n403650 , n403651 , n403652 , 
 n403653 , n403654 , n403655 , n403656 , n403657 , n403658 , n403659 , n403660 , n403661 , n403662 , 
 n403663 , n403664 , n403665 , n82005 , n403667 , n403668 , n403669 , n403670 , n403671 , n403672 , 
 n82012 , n403674 , n403675 , n82015 , n403677 , n403678 , n403679 , n403680 , n82020 , n82021 , 
 n403683 , n403684 , n403685 , n82025 , n403687 , n403688 , n403689 , n403690 , n403691 , n403692 , 
 n403693 , n403694 , n82034 , n403696 , n403697 , n403698 , n403699 , n403700 , n403701 , n403702 , 
 n403703 , n403704 , n403705 , n82045 , n403707 , n82047 , n82048 , n403710 , n403711 , n403712 , 
 n403713 , n403714 , n403715 , n403716 , n403717 , n403718 , n403719 , n403720 , n82060 , n403722 , 
 n403723 , n82063 , n403725 , n403726 , n82066 , n403728 , n403729 , n82069 , n403731 , n403732 , 
 n82072 , n403734 , n403735 , n403736 , n82076 , n82077 , n403739 , n403740 , n82080 , n82081 , 
 n403743 , n403744 , n82084 , n403746 , n403747 , n82087 , n403749 , n403750 , n403751 , n403752 , 
 n403753 , n403754 , n403755 , n82095 , n403757 , n403758 , n403759 , n403760 , n403761 , n403762 , 
 n403763 , n403764 , n403765 , n82105 , n403767 , n403768 , n403769 , n82109 , n403771 , n403772 , 
 n403773 , n403774 , n403775 , n403776 , n403777 , n403778 , n403779 , n403780 , n403781 , n403782 , 
 n82122 , n403784 , n403785 , n82125 , n403787 , n403788 , n403789 , n82129 , n403791 , n403792 , 
 n403793 , n82133 , n403795 , n403796 , n82136 , n403798 , n403799 , n403800 , n403801 , n403802 , 
 n403803 , n403804 , n82144 , n82145 , n82146 , n403808 , n403809 , n403810 , n403811 , n403812 , 
 n403813 , n403814 , n403815 , n403816 , n403817 , n82157 , n403819 , n403820 , n82160 , n82161 , 
 n403823 , n403824 , n82164 , n403826 , n403827 , n82167 , n82168 , n403830 , n403831 , n403832 , 
 n403833 , n403834 , n403835 , n403836 , n403837 , n82177 , n82178 , n403840 , n403841 , n403842 , 
 n82182 , n403844 , n403845 , n403846 , n82186 , n403848 , n403849 , n403850 , n82190 , n403852 , 
 n403853 , n82193 , n403855 , n82195 , n403857 , n403858 , n403859 , n403860 , n403861 , n82201 , 
 n403863 , n403864 , n82204 , n82205 , n403867 , n403868 , n82208 , n403870 , n403871 , n82211 , 
 n403873 , n403874 , n82214 , n403876 , n403877 , n82217 , n403879 , n403880 , n403881 , n403882 , 
 n403883 , n403884 , n403885 , n403886 , n403887 , n403888 , n82228 , n82229 , n403891 , n403892 , 
 n82232 , n82233 , n403895 , n403896 , n403897 , n403898 , n403899 , n403900 , n82240 , n82241 , 
 n403903 , n403904 , n403905 , n82245 , n403907 , n403908 , n403909 , n82249 , n82250 , n403912 , 
 n82252 , n403914 , n403915 , n403916 , n403917 , n403918 , n403919 , n82259 , n403921 , n403922 , 
 n82262 , n403924 , n403925 , n82265 , n403927 , n403928 , n82268 , n82269 , n82270 , n403932 , 
 n403933 , n403934 , n403935 , n82275 , n403937 , n403938 , n403939 , n82279 , n82280 , n403942 , 
 n403943 , n82283 , n403945 , n403946 , n82286 , n403948 , n403949 , n403950 , n403951 , n403952 , 
 n403953 , n403954 , n403955 , n82295 , n82296 , n403958 , n403959 , n403960 , n82300 , n403962 , 
 n403963 , n82303 , n403965 , n403966 , n403967 , n403968 , n403969 , n403970 , n82310 , n403972 , 
 n403973 , n82313 , n403975 , n403976 , n403977 , n403978 , n403979 , n403980 , n403981 , n403982 , 
 n82322 , n403984 , n403985 , n403986 , n403987 , n403988 , n403989 , n403990 , n403991 , n82331 , 
 n82332 , n403994 , n403995 , n403996 , n403997 , n403998 , n403999 , n404000 , n404001 , n404002 , 
 n82342 , n404004 , n82344 , n404006 , n82346 , n82347 , n82348 , n82349 , n82350 , n404012 , 
 n82352 , n82353 , n82354 , n404016 , n404017 , n404018 , n404019 , n404020 , n404021 , n404022 , 
 n404023 , n404024 , n82364 , n82365 , n404027 , n404028 , n404029 , n404030 , n404031 , n82371 , 
 n82372 , n404034 , n404035 , n82375 , n82376 , n82377 , n404039 , n404040 , n404041 , n404042 , 
 n82382 , n404044 , n404045 , n82385 , n82386 , n404048 , n404049 , n404050 , n404051 , n404052 , 
 n404053 , n82393 , n82394 , n404056 , n404057 , n404058 , n404059 , n404060 , n82398 , n82399 , 
 n404063 , n404064 , n404065 , n82403 , n404067 , n82405 , n404069 , n404070 , n404071 , n404072 , 
 n82410 , n404074 , n82412 , n404076 , n82414 , n404078 , n82416 , n404080 , n404081 , n82419 , 
 n404083 , n82421 , n82422 , n404086 , n404087 , n82425 , n404089 , n404090 , n404091 , n82429 , 
 n404093 , n404094 , n404095 , n82433 , n404097 , n82435 , n404099 , n404100 , n404101 , n404102 , 
 n82440 , n404104 , n404105 , n82443 , n404107 , n404108 , n404109 , n82447 , n404111 , n404112 , 
 n404113 , n404114 , n404115 , n404116 , n82454 , n404118 , n404119 , n404120 , n404121 , n404122 , 
 n404123 , n404124 , n404125 , n404126 , n404127 , n404128 , n404129 , n404130 , n404131 , n404132 , 
 n404133 , n404134 , n404135 , n82461 , n404137 , n404138 , n82464 , n404140 , n404141 , n404142 , 
 n404143 , n82469 , n404145 , n82470 , n404147 , n404148 , n404149 , n82473 , n404151 , n82475 , 
 n404153 , n82477 , n82478 , n404156 , n404157 , n82481 , n404159 , n404160 , n404161 , n404162 , 
 n404163 , n404164 , n404165 , n404166 , n404167 , n404168 , n404169 , n404170 , n404171 , n404172 , 
 n404173 , n404174 , n404175 , n82486 , n404177 , n404178 , n404179 , n82490 , n404181 , n404182 , 
 n82493 , n404184 , n404185 , n404186 , n82497 , n82498 , n82499 , n404190 , n404191 , n82502 , 
 n82503 , n404194 , n404195 , n404196 , n404197 , n404198 , n404199 , n404200 , n404201 , n404202 , 
 n404203 , n404204 , n404205 , n404206 , n404207 , n404208 , n404209 , n404210 , n404211 , n404212 , 
 n404213 , n404214 , n404215 , n404216 , n404217 , n404218 , n404219 , n404220 , n404221 , n404222 , 
 n82510 , n404224 , n404225 , n404226 , n82514 , n82515 , n404229 , n404230 , n404231 , n404232 , 
 n82520 , n82521 , n404235 , n404236 , n404237 , n404238 , n404239 , n404240 , n404241 , n404242 , 
 n404243 , n404244 , n404245 , n82533 , n404247 , n404248 , n82536 , n404250 , n82538 , n404252 , 
 n82540 , n404254 , n404255 , n82543 , n404257 , n404258 , n82546 , n404260 , n404261 , n82549 , 
 n404263 , n404264 , n404265 , n404266 , n404267 , n404268 , n404269 , n404270 , n404271 , n404272 , 
 n404273 , n404274 , n404275 , n404276 , n404277 , n404278 , n404279 , n404280 , n404281 , n404282 , 
 n404283 , n404284 , n404285 , n404286 , n404287 , n404288 , n404289 , n404290 , n404291 , n404292 , 
 n404293 , n404294 , n404295 , n404296 , n404297 , n404298 , n82561 , n82562 , n404301 , n404302 , 
 n82565 , n404304 , n82566 , n404306 , n404307 , n82569 , n82570 , n404310 , n404311 , n404312 , 
 n404313 , n404314 , n404315 , n404316 , n404317 , n404318 , n404319 , n404320 , n404321 , n404322 , 
 n404323 , n404324 , n404325 , n404326 , n404327 , n404328 , n404329 , n404330 , n82573 , n404332 , 
 n404333 , n82575 , n82576 , n404336 , n404337 , n404338 , n404339 , n82581 , n404341 , n404342 , 
 n404343 , n82585 , n404345 , n404346 , n404347 , n404348 , n82590 , n404350 , n404351 , n82593 , 
 n82594 , n404354 , n82596 , n82597 , n82598 , n404358 , n404359 , n404360 , n404361 , n82603 , 
 n404363 , n404364 , n404365 , n404366 , n404367 , n404368 , n404369 , n404370 , n404371 , n404372 , 
 n404373 , n404374 , n404375 , n404376 , n82618 , n404378 , n404379 , n404380 , n82622 , n82623 , 
 n404383 , n404384 , n404385 , n404386 , n82628 , n404388 , n404389 , n82631 , n82632 , n82633 , 
 n82634 , n82635 , n82636 , n404396 , n404397 , n82639 , n404399 , n404400 , n404401 , n404402 , 
 n404403 , n404404 , n404405 , n404406 , n404407 , n82649 , n404409 , n404410 , n82652 , n404412 , 
 n404413 , n404414 , n404415 , n404416 , n404417 , n404418 , n404419 , n404420 , n404421 , n404422 , 
 n404423 , n404424 , n404425 , n404426 , n404427 , n404428 , n404429 , n404430 , n82672 , n404432 , 
 n404433 , n82675 , n404435 , n404436 , n82678 , n404438 , n404439 , n404440 , n404441 , n82683 , 
 n404443 , n82685 , n82686 , n404446 , n404447 , n404448 , n82690 , n404450 , n404451 , n404452 , 
 n404453 , n404454 , n82696 , n404456 , n404457 , n82699 , n82700 , n82701 , n404461 , n404462 , 
 n82704 , n404464 , n404465 , n404466 , n82708 , n404468 , n82710 , n82711 , n404471 , n404472 , 
 n82714 , n404474 , n404475 , n82717 , n82718 , n404478 , n404479 , n82721 , n82722 , n82723 , 
 n404483 , n404484 , n82726 , n82727 , n82728 , n404488 , n82730 , n404490 , n404491 , n82733 , 
 n404493 , n404494 , n82736 , n82737 , n404497 , n404498 , n82740 , n404500 , n404501 , n404502 , 
 n82744 , n404504 , n82746 , n404506 , n82748 , n82749 , n404509 , n82751 , n82752 , n404512 , 
 n404513 , n82755 , n82756 , n404516 , n82758 , n82759 , n404519 , n82761 , n404521 , n404522 , 
 n404523 , n404524 , n404525 , n404526 , n404527 , n404528 , n404529 , n404530 , n82772 , n82773 , 
 n404533 , n404534 , n404535 , n82777 , n404537 , n404538 , n404539 , n404540 , n404541 , n404542 , 
 n404543 , n404544 , n404545 , n404546 , n404547 , n404548 , n404549 , n404550 , n404551 , n404552 , 
 n404553 , n404554 , n404555 , n404556 , n404557 , n82780 , n82781 , n82782 , n82783 , n82784 , 
 n82785 , n82786 , n82787 , n82788 , n82789 , n82790 , n404569 , n404570 , n404571 , n404572 , 
 n404573 , n404574 , n404575 , n404576 , n404577 , n404578 , n82801 , n404580 , n404581 , n404582 , 
 n404583 , n404584 , n404585 , n404586 , n404587 , n404588 , n404589 , n404590 , n82813 , n404592 , 
 n82815 , n404594 , n82817 , n404596 , n404597 , n404598 , n404599 , n404600 , n404601 , n404602 , 
 n82824 , n404604 , n404605 , n404606 , n404607 , n82829 , n82830 , n82831 , n82832 , n404612 , 
 n82834 , n404614 , n404615 , n404616 , n404617 , n404618 , n404619 , n404620 , n404621 , n404622 , 
 n404623 , n404624 , n404625 , n404626 , n404627 , n404628 , n404629 , n404630 , n404631 , n404632 , 
 n404633 , n82855 , n404635 , n404636 , n82858 , n404638 , n404639 , n404640 , n404641 , n82863 , 
 n404643 , n404644 , n404645 , n404646 , n404647 , n82869 , n404649 , n404650 , n82872 , n404652 , 
 n404653 , n404654 , n404655 , n82877 , n404657 , n404658 , n82880 , n404660 , n404661 , n404662 , 
 n404663 , n82885 , n404665 , n82887 , n82888 , n404668 , n404669 , n404670 , n404671 , n404672 , 
 n404673 , n404674 , n404675 , n404676 , n404677 , n404678 , n404679 , n404680 , n404681 , n404682 , 
 n404683 , n404684 , n82906 , n404686 , n404687 , n404688 , n82910 , n404690 , n404691 , n404692 , 
 n404693 , n404694 , n404695 , n82917 , n404697 , n404698 , n404699 , n404700 , n82922 , n82923 , 
 n82924 , n82925 , n404705 , n82927 , n82928 , n404708 , n82930 , n82931 , n82932 , n404712 , 
 n404713 , n404714 , n82936 , n404716 , n404717 , n404718 , n82940 , n404720 , n404721 , n404722 , 
 n404723 , n404724 , n404725 , n404726 , n404727 , n404728 , n404729 , n404730 , n404731 , n404732 , 
 n404733 , n404734 , n404735 , n404736 , n404737 , n404738 , n404739 , n404740 , n82950 , n404742 , 
 n82952 , n404744 , n82954 , n404746 , n404747 , n404748 , n404749 , n404750 , n404751 , n404752 , 
 n404753 , n404754 , n82964 , n404756 , n404757 , n82967 , n404759 , n404760 , n404761 , n404762 , 
 n404763 , n404764 , n404765 , n404766 , n404767 , n404768 , n404769 , n404770 , n404771 , n404772 , 
 n404773 , n404774 , n404775 , n404776 , n404777 , n404778 , n404779 , n404780 , n404781 , n404782 , 
 n404783 , n404784 , n404785 , n404786 , n404787 , n404788 , n404789 , n404790 , n404791 , n404792 , 
 n404793 , n404794 , n404795 , n82982 , n404797 , n404798 , n82985 , n404800 , n404801 , n82988 , 
 n404803 , n404804 , n404805 , n404806 , n82993 , n82994 , n82995 , n82996 , n404811 , n82998 , 
 n404813 , n404814 , n83001 , n404816 , n404817 , n404818 , n404819 , n404820 , n83007 , n404822 , 
 n404823 , n83010 , n404825 , n404826 , n83013 , n404828 , n404829 , n404830 , n404831 , n404832 , 
 n404833 , n404834 , n404835 , n404836 , n404837 , n83023 , n404839 , n404840 , n404841 , n404842 , 
 n404843 , n404844 , n404845 , n83031 , n404847 , n404848 , n83034 , n404850 , n404851 , n404852 , 
 n404853 , n404854 , n83040 , n404856 , n404857 , n404858 , n404859 , n404860 , n404861 , n404862 , 
 n404863 , n404864 , n83050 , n404866 , n404867 , n404868 , n404869 , n404870 , n83056 , n404872 , 
 n404873 , n404874 , n404875 , n404876 , n404877 , n404878 , n404879 , n404880 , n404881 , n404882 , 
 n83068 , n83069 , n83070 , n83071 , n83072 , n83073 , n83074 , n83075 , n83076 , n404892 , 
 n83078 , n404894 , n404895 , n83081 , n404897 , n404898 , n83084 , n404900 , n404901 , n404902 , 
 n404903 , n83089 , n83090 , n404906 , n404907 , n83093 , n404909 , n404910 , n404911 , n83097 , 
 n404913 , n404914 , n404915 , n404916 , n404917 , n404918 , n404919 , n404920 , n404921 , n404922 , 
 n404923 , n404924 , n404925 , n404926 , n404927 , n404928 , n404929 , n404930 , n404931 , n83104 , 
 n404933 , n404934 , n83107 , n404936 , n404937 , n404938 , n83111 , n404940 , n404941 , n404942 , 
 n404943 , n404944 , n404945 , n404946 , n404947 , n404948 , n404949 , n404950 , n404951 , n404952 , 
 n404953 , n404954 , n83113 , n404956 , n404957 , n83116 , n404959 , n404960 , n404961 , n404962 , 
 n404963 , n83122 , n404965 , n404966 , n83125 , n404968 , n404969 , n404970 , n404971 , n404972 , 
 n404973 , n404974 , n404975 , n83134 , n404977 , n404978 , n404979 , n404980 , n404981 , n404982 , 
 n83141 , n83142 , n404985 , n404986 , n404987 , n404988 , n404989 , n83148 , n404991 , n404992 , 
 n404993 , n83152 , n83153 , n404996 , n404997 , n404998 , n404999 , n405000 , n405001 , n405002 , 
 n405003 , n405004 , n405005 , n405006 , n405007 , n405008 , n405009 , n405010 , n405011 , n405012 , 
 n405013 , n405014 , n405015 , n83160 , n83161 , n405018 , n405019 , n405020 , n83165 , n405022 , 
 n405023 , n83168 , n405025 , n405026 , n83171 , n405028 , n405029 , n83174 , n405031 , n405032 , 
 n83177 , n405034 , n405035 , n405036 , n83181 , n83182 , n83183 , n405040 , n405041 , n405042 , 
 n405043 , n83188 , n405045 , n405046 , n405047 , n405048 , n83193 , n83194 , n83195 , n405052 , 
 n83197 , n405054 , n405055 , n405056 , n405057 , n83202 , n405059 , n405060 , n405061 , n83206 , 
 n405063 , n405064 , n405065 , n83210 , n405067 , n405068 , n83213 , n83214 , n405071 , n405072 , 
 n405073 , n405074 , n405075 , n405076 , n405077 , n405078 , n405079 , n405080 , n83225 , n83226 , 
 n405083 , n405084 , n405085 , n405086 , n83231 , n83232 , n405089 , n405090 , n83235 , n83236 , 
 n83237 , n405094 , n83239 , n405096 , n405097 , n405098 , n405099 , n405100 , n405101 , n405102 , 
 n405103 , n405104 , n405105 , n405106 , n83251 , n405108 , n405109 , n405110 , n405111 , n405112 , 
 n405113 , n405114 , n405115 , n405116 , n405117 , n405118 , n83263 , n405120 , n405121 , n405122 , 
 n405123 , n83268 , n83269 , n405126 , n83271 , n405128 , n405129 , n405130 , n83275 , n83276 , 
 n405133 , n405134 , n83279 , n405136 , n83281 , n405138 , n83283 , n405140 , n83285 , n83286 , 
 n83287 , n83288 , n405145 , n405146 , n83291 , n405148 , n405149 , n83294 , n405151 , n83296 , 
 n405153 , n405154 , n405155 , n405156 , n83301 , n405158 , n83303 , n405160 , n405161 , n405162 , 
 n83307 , n405164 , n405165 , n405166 , n405167 , n405168 , n83313 , n405170 , n405171 , n83316 , 
 n405173 , n405174 , n405175 , n405176 , n405177 , n405178 , n405179 , n83324 , n405181 , n83326 , 
 n405183 , n83328 , n405185 , n405186 , n83331 , n405188 , n405189 , n405190 , n405191 , n83336 , 
 n405193 , n405194 , n405195 , n83340 , n405197 , n405198 , n405199 , n83344 , n405201 , n405202 , 
 n405203 , n405204 , n405205 , n405206 , n405207 , n405208 , n405209 , n405210 , n405211 , n405212 , 
 n405213 , n405214 , n405215 , n83360 , n405217 , n405218 , n405219 , n83364 , n405221 , n405222 , 
 n405223 , n405224 , n405225 , n405226 , n83371 , n405228 , n405229 , n83374 , n405231 , n405232 , 
 n405233 , n83378 , n405235 , n405236 , n83381 , n405238 , n405239 , n83384 , n405241 , n405242 , 
 n83387 , n405244 , n405245 , n405246 , n405247 , n405248 , n405249 , n405250 , n405251 , n405252 , 
 n405253 , n405254 , n405255 , n405256 , n405257 , n405258 , n405259 , n405260 , n405261 , n405262 , 
 n405263 , n405264 , n405265 , n405266 , n405267 , n405268 , n405269 , n405270 , n405271 , n405272 , 
 n405273 , n405274 , n83391 , n405276 , n405277 , n83392 , n405279 , n405280 , n83395 , n405282 , 
 n83397 , n405284 , n83399 , n405286 , n83401 , n83402 , n83403 , n405290 , n83405 , n405292 , 
 n405293 , n83408 , n405295 , n405296 , n405297 , n405298 , n405299 , n405300 , n405301 , n405302 , 
 n405303 , n405304 , n405305 , n405306 , n405307 , n405308 , n405309 , n405310 , n405311 , n405312 , 
 n405313 , n405314 , n405315 , n405316 , n405317 , n405318 , n405319 , n405320 , n83414 , n405322 , 
 n405323 , n405324 , n405325 , n405326 , n83420 , n405328 , n405329 , n405330 , n405331 , n405332 , 
 n405333 , n405334 , n405335 , n83429 , n83430 , n83431 , n405339 , n405340 , n83434 , n405342 , 
 n405343 , n83437 , n405345 , n405346 , n83440 , n405348 , n405349 , n405350 , n405351 , n405352 , 
 n405353 , n405354 , n405355 , n405356 , n405357 , n83451 , n83452 , n405360 , n405361 , n405362 , 
 n405363 , n405364 , n405365 , n83459 , n405367 , n405368 , n405369 , n405370 , n405371 , n405372 , 
 n405373 , n405374 , n83468 , n405376 , n405377 , n405378 , n405379 , n405380 , n405381 , n405382 , 
 n405383 , n405384 , n405385 , n405386 , n83480 , n405388 , n405389 , n405390 , n405391 , n405392 , 
 n405393 , n405394 , n405395 , n405396 , n405397 , n405398 , n405399 , n405400 , n405401 , n405402 , 
 n405403 , n405404 , n405405 , n405406 , n405407 , n405408 , n405409 , n405410 , n405411 , n405412 , 
 n405413 , n405414 , n405415 , n405416 , n405417 , n405418 , n405419 , n405420 , n405421 , n405422 , 
 n405423 , n83486 , n405425 , n83488 , n405427 , n405428 , n405429 , n83492 , n405431 , n405432 , 
 n405433 , n405434 , n405435 , n405436 , n405437 , n405438 , n405439 , n405440 , n83503 , n405442 , 
 n405443 , n405444 , n405445 , n405446 , n83509 , n405448 , n405449 , n83512 , n405451 , n405452 , 
 n83515 , n405454 , n405455 , n405456 , n83519 , n405458 , n83521 , n405460 , n83523 , n405462 , 
 n405463 , n405464 , n405465 , n405466 , n405467 , n405468 , n405469 , n83532 , n405471 , n83534 , 
 n83535 , n405474 , n405475 , n405476 , n405477 , n83540 , n405479 , n405480 , n405481 , n405482 , 
 n405483 , n405484 , n405485 , n405486 , n405487 , n405488 , n405489 , n405490 , n405491 , n405492 , 
 n405493 , n405494 , n405495 , n83555 , n405497 , n405498 , n405499 , n405500 , n405501 , n405502 , 
 n405503 , n405504 , n83564 , n405506 , n405507 , n405508 , n405509 , n83569 , n405511 , n405512 , 
 n83572 , n83573 , n405515 , n83575 , n83576 , n405518 , n405519 , n405520 , n405521 , n405522 , 
 n83582 , n405524 , n405525 , n405526 , n405527 , n405528 , n405529 , n405530 , n83590 , n405532 , 
 n405533 , n405534 , n405535 , n405536 , n83596 , n405538 , n405539 , n405540 , n405541 , n405542 , 
 n83602 , n405544 , n405545 , n405546 , n405547 , n405548 , n405549 , n405550 , n405551 , n83611 , 
 n405553 , n405554 , n405555 , n405556 , n405557 , n83617 , n405559 , n405560 , n83620 , n405562 , 
 n405563 , n83623 , n405565 , n405566 , n83626 , n83627 , n83628 , n405570 , n405571 , n83631 , 
 n405573 , n83633 , n405575 , n405576 , n83636 , n405578 , n405579 , n83639 , n405581 , n405582 , 
 n83642 , n83643 , n405585 , n83645 , n405587 , n405588 , n405589 , n405590 , n405591 , n405592 , 
 n405593 , n405594 , n405595 , n405596 , n405597 , n83657 , n405599 , n83659 , n405601 , n405602 , 
 n83662 , n405604 , n405605 , n83665 , n405607 , n405608 , n83668 , n405610 , n405611 , n405612 , 
 n83672 , n405614 , n405615 , n405616 , n405617 , n405618 , n405619 , n405620 , n405621 , n405622 , 
 n405623 , n405624 , n405625 , n405626 , n405627 , n405628 , n405629 , n405630 , n405631 , n405632 , 
 n405633 , n405634 , n405635 , n405636 , n405637 , n405638 , n405639 , n405640 , n83678 , n405642 , 
 n405643 , n83681 , n405645 , n405646 , n83684 , n83685 , n405649 , n83687 , n83688 , n83689 , 
 n405653 , n405654 , n83692 , n405656 , n83694 , n405658 , n405659 , n405660 , n405661 , n405662 , 
 n405663 , n405664 , n405665 , n405666 , n405667 , n405668 , n405669 , n405670 , n83706 , n405672 , 
 n83708 , n83709 , n405675 , n405676 , n405677 , n405678 , n405679 , n405680 , n405681 , n405682 , 
 n405683 , n405684 , n405685 , n405686 , n405687 , n405688 , n405689 , n405690 , n405691 , n83727 , 
 n405693 , n405694 , n405695 , n83731 , n405697 , n405698 , n83732 , n405700 , n405701 , n405702 , 
 n405703 , n405704 , n405705 , n405706 , n405707 , n405708 , n405709 , n405710 , n405711 , n405712 , 
 n405713 , n405714 , n405715 , n405716 , n405717 , n405718 , n405719 , n405720 , n405721 , n405722 , 
 n405723 , n405724 , n405725 , n405726 , n405727 , n405728 , n405729 , n405730 , n405731 , n405732 , 
 n83744 , n405734 , n405735 , n405736 , n405737 , n405738 , n405739 , n405740 , n405741 , n405742 , 
 n405743 , n405744 , n405745 , n405746 , n405747 , n405748 , n405749 , n405750 , n405751 , n405752 , 
 n405753 , n405754 , n405755 , n405756 , n83750 , n405758 , n405759 , n405760 , n405761 , n83753 , 
 n405763 , n405764 , n83756 , n405766 , n405767 , n83759 , n405769 , n405770 , n405771 , n405772 , 
 n405773 , n405774 , n405775 , n405776 , n405777 , n405778 , n83766 , n405780 , n405781 , n405782 , 
 n83770 , n83771 , n405785 , n83773 , n405787 , n405788 , n405789 , n405790 , n405791 , n405792 , 
 n405793 , n405794 , n405795 , n405796 , n405797 , n405798 , n405799 , n83787 , n405801 , n405802 , 
 n405803 , n405804 , n405805 , n405806 , n405807 , n405808 , n405809 , n405810 , n405811 , n405812 , 
 n405813 , n405814 , n405815 , n405816 , n405817 , n405818 , n405819 , n405820 , n405821 , n405822 , 
 n83794 , n405824 , n405825 , n405826 , n405827 , n83799 , n405829 , n405830 , n405831 , n405832 , 
 n405833 , n405834 , n405835 , n405836 , n405837 , n405838 , n405839 , n405840 , n405841 , n83808 , 
 n405843 , n405844 , n83810 , n83811 , n405847 , n405848 , n405849 , n83813 , n405851 , n405852 , 
 n405853 , n83816 , n83817 , n83818 , n405857 , n405858 , n405859 , n405860 , n405861 , n405862 , 
 n405863 , n405864 , n405865 , n405866 , n405867 , n405868 , n405869 , n405870 , n405871 , n405872 , 
 n405873 , n405874 , n405875 , n405876 , n405877 , n405878 , n405879 , n405880 , n405881 , n405882 , 
 n405883 , n83827 , n83828 , n405886 , n405887 , n83831 , n405889 , n405890 , n83834 , n83835 , 
 n405893 , n405894 , n405895 , n405896 , n405897 , n83840 , n405899 , n405900 , n405901 , n405902 , 
 n83845 , n83846 , n405905 , n405906 , n83849 , n83850 , n83851 , n405910 , n405911 , n405912 , 
 n405913 , n405914 , n405915 , n405916 , n405917 , n405918 , n405919 , n405920 , n405921 , n405922 , 
 n405923 , n405924 , n405925 , n405926 , n405927 , n405928 , n405929 , n405930 , n405931 , n405932 , 
 n405933 , n405934 , n83858 , n83859 , n405937 , n405938 , n405939 , n405940 , n405941 , n405942 , 
 n405943 , n405944 , n405945 , n405946 , n405947 , n405948 , n83872 , n405950 , n405951 , n405952 , 
 n405953 , n405954 , n405955 , n405956 , n405957 , n405958 , n405959 , n405960 , n405961 , n405962 , 
 n405963 , n405964 , n405965 , n405966 , n405967 , n405968 , n405969 , n405970 , n405971 , n405972 , 
 n405973 , n405974 , n405975 , n405976 , n405977 , n405978 , n405979 , n83892 , n405981 , n405982 , 
 n405983 , n405984 , n405985 , n83896 , n405987 , n405988 , n83899 , n83900 , n83901 , n83902 , 
 n83903 , n83904 , n405995 , n405996 , n83907 , n405998 , n405999 , n406000 , n83908 , n83909 , 
 n406003 , n406004 , n406005 , n406006 , n406007 , n406008 , n406009 , n406010 , n406011 , n406012 , 
 n406013 , n406014 , n406015 , n406016 , n406017 , n406018 , n406019 , n406020 , n406021 , n406022 , 
 n83913 , n83914 , n406025 , n406026 , n83917 , n406028 , n83919 , n406030 , n406031 , n83922 , 
 n406033 , n406034 , n406035 , n406036 , n406037 , n406038 , n406039 , n406040 , n406041 , n406042 , 
 n83932 , n83933 , n406045 , n406046 , n83936 , n406048 , n406049 , n406050 , n406051 , n406052 , 
 n406053 , n406054 , n83940 , n83941 , n83942 , n406058 , n406059 , n406060 , n406061 , n406062 , 
 n83948 , n406064 , n406065 , n406066 , n406067 , n406068 , n83954 , n406070 , n83956 , n83957 , 
 n406073 , n83958 , n83959 , n406076 , n406077 , n406078 , n406079 , n406080 , n406081 , n406082 , 
 n406083 , n406084 , n406085 , n406086 , n406087 , n406088 , n406089 , n406090 , n406091 , n406092 , 
 n406093 , n406094 , n406095 , n406096 , n406097 , n406098 , n406099 , n406100 , n406101 , n406102 , 
 n406103 , n406104 , n406105 , n406106 , n406107 , n406108 , n406109 , n406110 , n406111 , n406112 , 
 n406113 , n406114 , n406115 , n406116 , n406117 , n406118 , n83965 , n83966 , n406121 , n406122 , 
 n406123 , n406124 , n406125 , n83972 , n406127 , n406128 , n406129 , n406130 , n406131 , n406132 , 
 n406133 , n406134 , n406135 , n406136 , n406137 , n406138 , n406139 , n406140 , n406141 , n406142 , 
 n406143 , n406144 , n406145 , n406146 , n406147 , n406148 , n406149 , n406150 , n406151 , n406152 , 
 n406153 , n406154 , n406155 , n406156 , n406157 , n406158 , n406159 , n406160 , n406161 , n406162 , 
 n406163 , n406164 , n406165 , n406166 , n406167 , n406168 , n406169 , n406170 , n406171 , n406172 , 
 n406173 , n406174 , n406175 , n406176 , n406177 , n406178 , n406179 , n406180 , n406181 , n406182 , 
 n406183 , n406184 , n406185 , n406186 , n406187 , n406188 , n406189 , n406190 , n406191 , n406192 , 
 n406193 , n406194 , n406195 , n406196 , n406197 , n406198 , n406199 , n406200 , n406201 , n406202 , 
 n406203 , n406204 , n406205 , n406206 , n406207 , n406208 , n83992 , n406210 , n406211 , n406212 , 
 n406213 , n406214 , n406215 , n406216 , n406217 , n406218 , n406219 , n406220 , n406221 , n406222 , 
 n406223 , n406224 , n406225 , n406226 , n406227 , n406228 , n406229 , n406230 , n406231 , n406232 , 
 n406233 , n406234 , n406235 , n406236 , n406237 , n406238 , n406239 , n406240 , n406241 , n406242 , 
 n406243 , n406244 , n406245 , n406246 , n406247 , n406248 , n406249 , n406250 , n406251 , n406252 , 
 n406253 , n406254 , n84018 , n406256 , n406257 , n406258 , n84022 , n406260 , n406261 , n84025 , 
 n406263 , n406264 , n406265 , n406266 , n406267 , n406268 , n406269 , n406270 , n84034 , n84035 , 
 n406273 , n84037 , n84038 , n406276 , n406277 , n84041 , n84042 , n406280 , n406281 , n406282 , 
 n406283 , n84047 , n406285 , n406286 , n406287 , n406288 , n406289 , n84053 , n406291 , n406292 , 
 n406293 , n406294 , n406295 , n406296 , n406297 , n406298 , n406299 , n406300 , n406301 , n406302 , 
 n406303 , n406304 , n406305 , n406306 , n406307 , n406308 , n406309 , n406310 , n406311 , n406312 , 
 n406313 , n406314 , n406315 , n406316 , n406317 , n406318 , n406319 , n406320 , n406321 , n406322 , 
 n406323 , n406324 , n84071 , n406326 , n84073 , n406328 , n84075 , n406330 , n406331 , n406332 , 
 n406333 , n406334 , n406335 , n406336 , n406337 , n84084 , n406339 , n406340 , n84087 , n406342 , 
 n406343 , n84090 , n406345 , n406346 , n406347 , n406348 , n84095 , n406350 , n406351 , n406352 , 
 n406353 , n406354 , n84101 , n406356 , n406357 , n406358 , n406359 , n84106 , n406361 , n406362 , 
 n406363 , n406364 , n406365 , n406366 , n406367 , n406368 , n406369 , n84116 , n406371 , n406372 , 
 n406373 , n406374 , n84121 , n406376 , n84123 , n406378 , n406379 , n84126 , n406381 , n406382 , 
 n406383 , n406384 , n406385 , n406386 , n84129 , n406388 , n84131 , n84132 , n84133 , n84134 , 
 n406393 , n84136 , n84137 , n406396 , n84139 , n406398 , n406399 , n406400 , n84143 , n406402 , 
 n406403 , n406404 , n406405 , n84148 , n406407 , n406408 , n406409 , n406410 , n406411 , n406412 , 
 n406413 , n406414 , n406415 , n406416 , n406417 , n406418 , n406419 , n406420 , n406421 , n406422 , 
 n406423 , n406424 , n406425 , n406426 , n406427 , n406428 , n406429 , n84154 , n406431 , n406432 , 
 n406433 , n406434 , n84159 , n406436 , n406437 , n84162 , n406439 , n406440 , n84165 , n84166 , 
 n406443 , n406444 , n406445 , n406446 , n406447 , n406448 , n406449 , n84174 , n406451 , n406452 , 
 n406453 , n406454 , n406455 , n406456 , n406457 , n406458 , n84182 , n84183 , n406461 , n84185 , 
 n406463 , n406464 , n406465 , n406466 , n406467 , n406468 , n406469 , n84193 , n84194 , n406472 , 
 n406473 , n406474 , n84198 , n406476 , n406477 , n84201 , n406479 , n406480 , n406481 , n406482 , 
 n406483 , n406484 , n406485 , n406486 , n84210 , n84211 , n406489 , n406490 , n406491 , n406492 , 
 n84216 , n406494 , n406495 , n406496 , n406497 , n406498 , n406499 , n406500 , n406501 , n406502 , 
 n406503 , n406504 , n84226 , n406506 , n406507 , n406508 , n84230 , n406510 , n406511 , n406512 , 
 n406513 , n406514 , n406515 , n406516 , n406517 , n84239 , n406519 , n406520 , n406521 , n406522 , 
 n406523 , n406524 , n406525 , n406526 , n406527 , n84249 , n406529 , n406530 , n84252 , n406532 , 
 n406533 , n84255 , n406535 , n406536 , n84258 , n84259 , n406539 , n406540 , n406541 , n84263 , 
 n406543 , n406544 , n406545 , n406546 , n406547 , n84269 , n406549 , n406550 , n406551 , n406552 , 
 n406553 , n406554 , n84276 , n406556 , n406557 , n84279 , n406559 , n406560 , n406561 , n84283 , 
 n406563 , n406564 , n84286 , n84287 , n406567 , n406568 , n406569 , n406570 , n406571 , n406572 , 
 n406573 , n84295 , n406575 , n406576 , n84298 , n406578 , n84300 , n406580 , n84302 , n406582 , 
 n406583 , n406584 , n84306 , n406586 , n406587 , n406588 , n406589 , n84311 , n406591 , n406592 , 
 n406593 , n84315 , n406595 , n406596 , n406597 , n406598 , n406599 , n406600 , n84322 , n406602 , 
 n406603 , n84325 , n406605 , n406606 , n406607 , n406608 , n406609 , n84331 , n84332 , n406612 , 
 n406613 , n406614 , n84336 , n406616 , n406617 , n84339 , n84340 , n406620 , n84342 , n84343 , 
 n406623 , n406624 , n84346 , n84347 , n84348 , n406628 , n406629 , n406630 , n84352 , n406632 , 
 n406633 , n406634 , n406635 , n406636 , n84358 , n406638 , n406639 , n406640 , n406641 , n84363 , 
 n406643 , n406644 , n406645 , n84367 , n406647 , n406648 , n406649 , n84371 , n406651 , n406652 , 
 n84374 , n84375 , n406655 , n406656 , n406657 , n406658 , n406659 , n406660 , n406661 , n406662 , 
 n406663 , n406664 , n406665 , n406666 , n406667 , n84389 , n84390 , n406670 , n84392 , n84393 , 
 n84394 , n84395 , n406675 , n406676 , n84398 , n406678 , n84400 , n406680 , n84402 , n84403 , 
 n406683 , n406684 , n406685 , n84407 , n406687 , n84409 , n406689 , n406690 , n406691 , n406692 , 
 n406693 , n406694 , n406695 , n406696 , n84418 , n406698 , n84420 , n406700 , n406701 , n84423 , 
 n84424 , n406704 , n406705 , n406706 , n406707 , n84429 , n406709 , n406710 , n84432 , n84433 , 
 n406713 , n406714 , n406715 , n84437 , n406717 , n406718 , n406719 , n84440 , n406721 , n406722 , 
 n406723 , n84444 , n406725 , n406726 , n84447 , n406728 , n406729 , n406730 , n84451 , n406732 , 
 n406733 , n84454 , n406735 , n406736 , n406737 , n84458 , n406739 , n406740 , n84461 , n406742 , 
 n406743 , n406744 , n406745 , n406746 , n406747 , n406748 , n406749 , n406750 , n406751 , n406752 , 
 n406753 , n406754 , n406755 , n84476 , n84477 , n406758 , n84479 , n406760 , n406761 , n406762 , 
 n84483 , n406764 , n406765 , n84486 , n406767 , n406768 , n406769 , n84490 , n406771 , n406772 , 
 n84493 , n406774 , n406775 , n406776 , n406777 , n406778 , n84499 , n406780 , n406781 , n406782 , 
 n406783 , n406784 , n406785 , n406786 , n406787 , n406788 , n406789 , n406790 , n406791 , n406792 , 
 n406793 , n406794 , n406795 , n406796 , n406797 , n406798 , n406799 , n406800 , n406801 , n406802 , 
 n406803 , n406804 , n406805 , n406806 , n406807 , n406808 , n406809 , n84507 , n406811 , n406812 , 
 n406813 , n406814 , n406815 , n406816 , n406817 , n406818 , n406819 , n406820 , n406821 , n406822 , 
 n84514 , n406824 , n406825 , n406826 , n84518 , n84519 , n84520 , n406830 , n406831 , n406832 , 
 n84524 , n406834 , n406835 , n406836 , n406837 , n84529 , n406839 , n406840 , n84532 , n406842 , 
 n406843 , n84535 , n84536 , n406846 , n84537 , n406848 , n84539 , n84540 , n84541 , n84542 , 
 n84543 , n84544 , n84545 , n84546 , n84547 , n84548 , n406859 , n84550 , n406861 , n84552 , 
 n406863 , n84554 , n84555 , n406866 , n406867 , n406868 , n406869 , n406870 , n84561 , n406872 , 
 n406873 , n84564 , n406875 , n406876 , n406877 , n406878 , n406879 , n406880 , n406881 , n406882 , 
 n84573 , n406884 , n84575 , n84576 , n406887 , n406888 , n84579 , n84580 , n84581 , n406892 , 
 n84583 , n406894 , n406895 , n84586 , n406897 , n84588 , n406899 , n406900 , n84591 , n406902 , 
 n84593 , n406904 , n406905 , n406906 , n84597 , n406908 , n406909 , n84600 , n406911 , n406912 , 
 n406913 , n406914 , n406915 , n406916 , n406917 , n406918 , n84609 , n84610 , n84611 , n84612 , 
 n84613 , n84614 , n84615 , n406926 , n406927 , n406928 , n84619 , n406930 , n406931 , n84622 , 
 n406933 , n406934 , n84625 , n84626 , n406937 , n406938 , n84629 , n406940 , n406941 , n84632 , 
 n84633 , n84634 , n84635 , n406946 , n406947 , n406948 , n84639 , n406950 , n406951 , n406952 , 
 n406953 , n406954 , n84645 , n406956 , n406957 , n406958 , n406959 , n406960 , n406961 , n406962 , 
 n406963 , n406964 , n406965 , n406966 , n406967 , n84658 , n84659 , n84660 , n84661 , n84662 , 
 n84663 , n84664 , n84665 , n406976 , n84667 , n406978 , n406979 , n84670 , n406981 , n84672 , 
 n84673 , n406984 , n406985 , n406986 , n84677 , n84678 , n406989 , n406990 , n406991 , n406992 , 
 n406993 , n84684 , n406995 , n84686 , n406997 , n406998 , n406999 , n84690 , n407001 , n84692 , 
 n407003 , n407004 , n407005 , n407006 , n407007 , n407008 , n407009 , n84700 , n84701 , n407012 , 
 n407013 , n84704 , n407015 , n407016 , n407017 , n407018 , n407019 , n407020 , n407021 , n407022 , 
 n407023 , n407024 , n407025 , n407026 , n407027 , n407028 , n84719 , n407030 , n407031 , n407032 , 
 n84723 , n407034 , n84725 , n407036 , n407037 , n407038 , n407039 , n407040 , n407041 , n84732 , 
 n407043 , n407044 , n407045 , n84736 , n407047 , n407048 , n407049 , n407050 , n407051 , n407052 , 
 n84743 , n84744 , n407055 , n407056 , n407057 , n407058 , n407059 , n407060 , n407061 , n407062 , 
 n84753 , n84754 , n84755 , n407066 , n407067 , n84758 , n84759 , n84760 , n407071 , n407072 , 
 n84763 , n84764 , n84765 , n407076 , n407077 , n84768 , n407079 , n407080 , n84771 , n407082 , 
 n407083 , n84774 , n407085 , n407086 , n407087 , n84778 , n407089 , n407090 , n407091 , n407092 , 
 n407093 , n407094 , n407095 , n407096 , n407097 , n407098 , n407099 , n407100 , n407101 , n407102 , 
 n407103 , n407104 , n407105 , n407106 , n84781 , n84782 , n84783 , n84784 , n84785 , n84786 , 
 n84787 , n84788 , n407115 , n84790 , n407117 , n407118 , n84793 , n407120 , n407121 , n84796 , 
 n407123 , n407124 , n84799 , n407126 , n407127 , n407128 , n407129 , n407130 , n407131 , n407132 , 
 n407133 , n407134 , n407135 , n407136 , n84811 , n407138 , n407139 , n407140 , n84815 , n84816 , 
 n407143 , n407144 , n407145 , n407146 , n407147 , n84822 , n407149 , n407150 , n407151 , n84826 , 
 n407153 , n407154 , n407155 , n407156 , n407157 , n407158 , n407159 , n407160 , n407161 , n84836 , 
 n84837 , n407164 , n407165 , n407166 , n84841 , n84842 , n407169 , n407170 , n84845 , n407172 , 
 n407173 , n84848 , n407175 , n407176 , n407177 , n84852 , n407179 , n407180 , n407181 , n407182 , 
 n407183 , n407184 , n407185 , n407186 , n84861 , n407188 , n84863 , n407190 , n84865 , n407192 , 
 n407193 , n84868 , n407195 , n407196 , n84871 , n407198 , n407199 , n407200 , n407201 , n407202 , 
 n407203 , n407204 , n84879 , n407206 , n407207 , n407208 , n84883 , n407210 , n84885 , n84886 , 
 n84887 , n84888 , n84889 , n84890 , n84891 , n407218 , n84893 , n407220 , n407221 , n407222 , 
 n84897 , n407224 , n407225 , n407226 , n407227 , n407228 , n407229 , n407230 , n407231 , n407232 , 
 n407233 , n407234 , n84909 , n407236 , n84911 , n407238 , n407239 , n407240 , n407241 , n407242 , 
 n407243 , n407244 , n407245 , n84914 , n407247 , n84916 , n84917 , n407250 , n407251 , n407252 , 
 n84921 , n407254 , n407255 , n84924 , n407257 , n84926 , n407259 , n407260 , n84929 , n407262 , 
 n407263 , n407264 , n407265 , n84934 , n407267 , n84936 , n84937 , n84938 , n84939 , n84940 , 
 n84941 , n407274 , n84943 , n407276 , n407277 , n407278 , n407279 , n407280 , n407281 , n407282 , 
 n84951 , n407284 , n84953 , n84954 , n407287 , n407288 , n407289 , n407290 , n84959 , n407292 , 
 n407293 , n407294 , n84963 , n407296 , n84965 , n407298 , n407299 , n407300 , n407301 , n84970 , 
 n84971 , n407304 , n407305 , n407306 , n407307 , n407308 , n407309 , n407310 , n407311 , n407312 , 
 n84981 , n407314 , n407315 , n407316 , n407317 , n407318 , n407319 , n407320 , n84989 , n407322 , 
 n84991 , n407324 , n407325 , n407326 , n407327 , n407328 , n407329 , n407330 , n407331 , n407332 , 
 n407333 , n407334 , n407335 , n407336 , n407337 , n85004 , n407339 , n407340 , n407341 , n407342 , 
 n407343 , n407344 , n407345 , n85009 , n407347 , n85011 , n407349 , n407350 , n407351 , n407352 , 
 n407353 , n407354 , n407355 , n407356 , n407357 , n407358 , n407359 , n407360 , n407361 , n407362 , 
 n407363 , n85022 , n407365 , n85024 , n85025 , n407368 , n407369 , n407370 , n407371 , n85030 , 
 n407373 , n85032 , n85033 , n407376 , n407377 , n407378 , n407379 , n407380 , n85039 , n407382 , 
 n407383 , n85042 , n407385 , n407386 , n407387 , n407388 , n407389 , n407390 , n407391 , n407392 , 
 n407393 , n407394 , n407395 , n407396 , n407397 , n407398 , n407399 , n85058 , n407401 , n407402 , 
 n407403 , n407404 , n407405 , n407406 , n85065 , n407408 , n407409 , n407410 , n407411 , n407412 , 
 n407413 , n407414 , n407415 , n407416 , n407417 , n407418 , n85077 , n407420 , n407421 , n407422 , 
 n407423 , n85082 , n407425 , n85084 , n407427 , n85086 , n85087 , n407430 , n407431 , n407432 , 
 n407433 , n407434 , n407435 , n407436 , n407437 , n407438 , n407439 , n407440 , n407441 , n407442 , 
 n407443 , n407444 , n407445 , n407446 , n85105 , n85106 , n407449 , n85108 , n407451 , n407452 , 
 n85111 , n407454 , n407455 , n85114 , n407457 , n407458 , n407459 , n407460 , n407461 , n407462 , 
 n407463 , n407464 , n407465 , n407466 , n407467 , n407468 , n407469 , n407470 , n407471 , n407472 , 
 n407473 , n407474 , n407475 , n407476 , n407477 , n407478 , n407479 , n407480 , n407481 , n407482 , 
 n407483 , n407484 , n85120 , n85121 , n85122 , n407488 , n85124 , n407490 , n407491 , n85127 , 
 n407493 , n407494 , n407495 , n85131 , n407497 , n407498 , n407499 , n85135 , n407501 , n407502 , 
 n407503 , n407504 , n407505 , n85141 , n407507 , n407508 , n407509 , n407510 , n85146 , n407512 , 
 n85148 , n85149 , n407515 , n407516 , n407517 , n407518 , n407519 , n407520 , n407521 , n407522 , 
 n407523 , n407524 , n407525 , n407526 , n407527 , n407528 , n407529 , n407530 , n407531 , n407532 , 
 n407533 , n407534 , n407535 , n407536 , n407537 , n85163 , n407539 , n407540 , n407541 , n407542 , 
 n85168 , n407544 , n407545 , n407546 , n407547 , n407548 , n407549 , n407550 , n407551 , n407552 , 
 n407553 , n85179 , n407555 , n407556 , n407557 , n407558 , n85184 , n407560 , n407561 , n85187 , 
 n407563 , n407564 , n85190 , n407566 , n407567 , n407568 , n407569 , n407570 , n85196 , n407572 , 
 n407573 , n407574 , n85200 , n407576 , n407577 , n407578 , n85204 , n407580 , n407581 , n85207 , 
 n407583 , n407584 , n85210 , n85211 , n407587 , n85213 , n407589 , n85215 , n85216 , n407592 , 
 n407593 , n85219 , n407595 , n407596 , n407597 , n407598 , n407599 , n407600 , n85226 , n407602 , 
 n407603 , n85229 , n407605 , n407606 , n85232 , n407608 , n85234 , n407610 , n407611 , n407612 , 
 n407613 , n407614 , n85240 , n407616 , n407617 , n85243 , n85244 , n407620 , n407621 , n407622 , 
 n407623 , n407624 , n407625 , n407626 , n85252 , n407628 , n407629 , n407630 , n407631 , n407632 , 
 n407633 , n85259 , n407635 , n407636 , n85262 , n85263 , n85264 , n85265 , n85266 , n85267 , 
 n85268 , n85269 , n85270 , n85271 , n85272 , n85273 , n85274 , n407650 , n407651 , n85277 , 
 n407653 , n407654 , n85280 , n85281 , n407657 , n85283 , n407659 , n85285 , n407661 , n85287 , 
 n407663 , n407664 , n407665 , n407666 , n407667 , n407668 , n407669 , n407670 , n407671 , n407672 , 
 n407673 , n85299 , n85300 , n407676 , n85302 , n85303 , n407679 , n407680 , n85306 , n407682 , 
 n407683 , n407684 , n85310 , n407686 , n407687 , n407688 , n85314 , n85315 , n407691 , n407692 , 
 n407693 , n407694 , n407695 , n407696 , n85322 , n407698 , n407699 , n85325 , n407701 , n407702 , 
 n85328 , n407704 , n407705 , n85331 , n407707 , n407708 , n85334 , n407710 , n407711 , n407712 , 
 n407713 , n407714 , n407715 , n407716 , n407717 , n407718 , n407719 , n407720 , n407721 , n85347 , 
 n407723 , n407724 , n407725 , n85351 , n85352 , n407728 , n407729 , n85355 , n407731 , n407732 , 
 n407733 , n407734 , n407735 , n407736 , n85362 , n407738 , n407739 , n407740 , n85366 , n85367 , 
 n407743 , n407744 , n85370 , n85371 , n407747 , n85373 , n407749 , n407750 , n407751 , n407752 , 
 n407753 , n407754 , n407755 , n407756 , n407757 , n407758 , n407759 , n407760 , n85386 , n407762 , 
 n407763 , n85389 , n407765 , n407766 , n85392 , n407768 , n407769 , n85395 , n407771 , n85397 , 
 n407773 , n407774 , n85400 , n407776 , n407777 , n85403 , n85404 , n407780 , n407781 , n407782 , 
 n85408 , n407784 , n407785 , n407786 , n85412 , n407788 , n85414 , n85415 , n85416 , n407792 , 
 n407793 , n85419 , n407795 , n407796 , n407797 , n85423 , n407799 , n407800 , n407801 , n85427 , 
 n407803 , n407804 , n407805 , n85431 , n407807 , n407808 , n407809 , n85435 , n407811 , n85437 , 
 n85438 , n407814 , n407815 , n407816 , n407817 , n407818 , n85444 , n407820 , n407821 , n85447 , 
 n85448 , n407824 , n407825 , n407826 , n85452 , n407828 , n407829 , n85455 , n85456 , n407832 , 
 n85458 , n407834 , n407835 , n85461 , n407837 , n407838 , n407839 , n407840 , n407841 , n407842 , 
 n407843 , n407844 , n407845 , n407846 , n407847 , n407848 , n407849 , n407850 , n407851 , n407852 , 
 n407853 , n407854 , n407855 , n407856 , n407857 , n407858 , n407859 , n407860 , n85464 , n407862 , 
 n407863 , n85467 , n407865 , n407866 , n85470 , n85471 , n407869 , n407870 , n407871 , n407872 , 
 n407873 , n85477 , n407875 , n407876 , n407877 , n85481 , n407879 , n407880 , n85484 , n407882 , 
 n407883 , n407884 , n85488 , n85489 , n407887 , n85491 , n407889 , n407890 , n407891 , n407892 , 
 n407893 , n407894 , n85498 , n85499 , n407897 , n407898 , n407899 , n407900 , n407901 , n407902 , 
 n407903 , n407904 , n407905 , n85509 , n407907 , n407908 , n407909 , n85513 , n407911 , n407912 , 
 n85516 , n407914 , n407915 , n407916 , n85520 , n85521 , n407919 , n85523 , n85524 , n407922 , 
 n85526 , n407924 , n85528 , n407926 , n407927 , n407928 , n407929 , n85533 , n407931 , n407932 , 
 n407933 , n85537 , n407935 , n407936 , n85540 , n407938 , n407939 , n85543 , n407941 , n407942 , 
 n407943 , n407944 , n85548 , n407946 , n407947 , n85551 , n407949 , n407950 , n407951 , n407952 , 
 n407953 , n407954 , n407955 , n407956 , n407957 , n407958 , n407959 , n407960 , n85564 , n407962 , 
 n407963 , n407964 , n407965 , n407966 , n407967 , n85571 , n407969 , n407970 , n85574 , n407972 , 
 n407973 , n407974 , n407975 , n407976 , n407977 , n85581 , n407979 , n407980 , n407981 , n407982 , 
 n407983 , n407984 , n407985 , n85589 , n85590 , n407988 , n85592 , n407990 , n85594 , n407992 , 
 n407993 , n407994 , n407995 , n407996 , n407997 , n407998 , n407999 , n408000 , n408001 , n408002 , 
 n408003 , n408004 , n408005 , n408006 , n408007 , n408008 , n408009 , n408010 , n408011 , n85597 , 
 n408013 , n408014 , n408015 , n408016 , n408017 , n408018 , n85602 , n408020 , n408021 , n85605 , 
 n85606 , n85607 , n85608 , n408026 , n85610 , n85611 , n85612 , n408030 , n408031 , n85615 , 
 n85616 , n85617 , n408035 , n85619 , n408037 , n85621 , n408039 , n85623 , n85624 , n85625 , 
 n408043 , n408044 , n85628 , n408046 , n408047 , n408048 , n85632 , n408050 , n408051 , n408052 , 
 n85636 , n408054 , n408055 , n408056 , n408057 , n408058 , n408059 , n85642 , n85643 , n408062 , 
 n408063 , n408064 , n408065 , n408066 , n408067 , n408068 , n85651 , n85652 , n408071 , n408072 , 
 n408073 , n408074 , n408075 , n408076 , n408077 , n85660 , n85661 , n408080 , n85663 , n85664 , 
 n408083 , n408084 , n408085 , n408086 , n85669 , n85670 , n408089 , n408090 , n408091 , n408092 , 
 n85675 , n408094 , n408095 , n85678 , n85679 , n408098 , n408099 , n408100 , n408101 , n408102 , 
 n85685 , n85686 , n408105 , n408106 , n408107 , n408108 , n408109 , n408110 , n85693 , n408112 , 
 n408113 , n408114 , n408115 , n408116 , n408117 , n408118 , n408119 , n408120 , n85703 , n408122 , 
 n408123 , n408124 , n408125 , n85708 , n85709 , n408128 , n85711 , n85712 , n85713 , n408132 , 
 n85715 , n408134 , n408135 , n408136 , n85719 , n408138 , n408139 , n85722 , n85723 , n408142 , 
 n408143 , n408144 , n85727 , n408146 , n408147 , n85730 , n408149 , n408150 , n408151 , n408152 , 
 n408153 , n85736 , n408155 , n408156 , n408157 , n408158 , n85741 , n408160 , n408161 , n85744 , 
 n85745 , n85746 , n85747 , n85748 , n408167 , n85750 , n85751 , n408170 , n408171 , n408172 , 
 n408173 , n408174 , n408175 , n408176 , n408177 , n408178 , n408179 , n408180 , n408181 , n408182 , 
 n408183 , n408184 , n408185 , n408186 , n408187 , n408188 , n408189 , n408190 , n408191 , n408192 , 
 n408193 , n408194 , n408195 , n85755 , n85756 , n408198 , n85758 , n85759 , n408201 , n408202 , 
 n408203 , n408204 , n408205 , n408206 , n408207 , n408208 , n408209 , n408210 , n408211 , n408212 , 
 n408213 , n408214 , n408215 , n408216 , n408217 , n408218 , n408219 , n408220 , n408221 , n85778 , 
 n408223 , n408224 , n408225 , n408226 , n408227 , n85784 , n408229 , n408230 , n85787 , n408232 , 
 n408233 , n408234 , n408235 , n408236 , n408237 , n408238 , n85795 , n408240 , n408241 , n85798 , 
 n85799 , n408244 , n85801 , n408246 , n408247 , n408248 , n408249 , n408250 , n408251 , n85808 , 
 n408253 , n408254 , n408255 , n408256 , n408257 , n408258 , n85815 , n408260 , n408261 , n85818 , 
 n408263 , n408264 , n408265 , n408266 , n408267 , n408268 , n408269 , n408270 , n85827 , n408272 , 
 n408273 , n408274 , n408275 , n408276 , n85833 , n408278 , n408279 , n408280 , n408281 , n408282 , 
 n85839 , n408284 , n85841 , n408286 , n408287 , n408288 , n408289 , n408290 , n408291 , n408292 , 
 n408293 , n408294 , n408295 , n408296 , n408297 , n408298 , n408299 , n408300 , n85846 , n408302 , 
 n408303 , n408304 , n408305 , n408306 , n408307 , n85853 , n85854 , n408310 , n408311 , n408312 , 
 n85858 , n408314 , n408315 , n408316 , n408317 , n408318 , n85864 , n408320 , n408321 , n408322 , 
 n408323 , n408324 , n408325 , n85871 , n408327 , n408328 , n408329 , n85875 , n408331 , n408332 , 
 n408333 , n408334 , n408335 , n408336 , n85882 , n408338 , n408339 , n85885 , n408341 , n85887 , 
 n85888 , n408344 , n408345 , n85891 , n408347 , n408348 , n85894 , n408350 , n408351 , n85897 , 
 n408353 , n85899 , n408355 , n408356 , n408357 , n408358 , n408359 , n408360 , n408361 , n408362 , 
 n408363 , n408364 , n408365 , n408366 , n408367 , n408368 , n408369 , n408370 , n408371 , n408372 , 
 n408373 , n408374 , n408375 , n408376 , n408377 , n408378 , n408379 , n408380 , n408381 , n408382 , 
 n408383 , n408384 , n408385 , n408386 , n408387 , n408388 , n408389 , n408390 , n408391 , n408392 , 
 n408393 , n408394 , n408395 , n408396 , n85917 , n408398 , n408399 , n85920 , n85921 , n408402 , 
 n408403 , n408404 , n408405 , n408406 , n408407 , n408408 , n408409 , n408410 , n408411 , n408412 , 
 n408413 , n408414 , n85933 , n408416 , n408417 , n408418 , n85936 , n408420 , n85938 , n85939 , 
 n408423 , n408424 , n408425 , n408426 , n85944 , n85945 , n408429 , n408430 , n85948 , n408432 , 
 n408433 , n85951 , n408435 , n408436 , n85954 , n85955 , n408439 , n408440 , n408441 , n408442 , 
 n408443 , n85961 , n85962 , n85963 , n85964 , n85965 , n85966 , n408450 , n408451 , n85969 , 
 n408453 , n408454 , n408455 , n408456 , n408457 , n408458 , n408459 , n408460 , n85978 , n85979 , 
 n408463 , n408464 , n85982 , n408466 , n408467 , n408468 , n85986 , n85987 , n85988 , n85989 , 
 n408473 , n85991 , n408475 , n408476 , n408477 , n85995 , n85996 , n408480 , n408481 , n85999 , 
 n408483 , n408484 , n86002 , n408486 , n86004 , n86005 , n408489 , n408490 , n408491 , n86009 , 
 n408493 , n86011 , n86012 , n408496 , n86014 , n408498 , n408499 , n86017 , n408501 , n408502 , 
 n86020 , n408504 , n408505 , n408506 , n408507 , n408508 , n408509 , n408510 , n408511 , n408512 , 
 n86027 , n86028 , n408515 , n408516 , n408517 , n86031 , n86032 , n408520 , n408521 , n86035 , 
 n408523 , n408524 , n86038 , n408526 , n408527 , n408528 , n408529 , n408530 , n408531 , n408532 , 
 n408533 , n408534 , n86048 , n408536 , n86050 , n408538 , n408539 , n86053 , n408541 , n408542 , 
 n408543 , n408544 , n86058 , n408546 , n86060 , n408548 , n408549 , n86063 , n408551 , n408552 , 
 n86066 , n408554 , n408555 , n408556 , n408557 , n408558 , n408559 , n408560 , n408561 , n408562 , 
 n408563 , n408564 , n408565 , n86079 , n408567 , n86081 , n408569 , n408570 , n86084 , n408572 , 
 n408573 , n408574 , n86088 , n86089 , n408577 , n86091 , n86092 , n408580 , n408581 , n408582 , 
 n408583 , n408584 , n408585 , n408586 , n408587 , n408588 , n408589 , n86099 , n408591 , n408592 , 
 n408593 , n408594 , n408595 , n408596 , n408597 , n408598 , n408599 , n408600 , n408601 , n408602 , 
 n408603 , n408604 , n408605 , n408606 , n86102 , n408608 , n408609 , n408610 , n408611 , n408612 , 
 n408613 , n408614 , n408615 , n408616 , n86112 , n408618 , n408619 , n408620 , n408621 , n408622 , 
 n408623 , n86119 , n408625 , n408626 , n408627 , n86123 , n408629 , n408630 , n408631 , n408632 , 
 n86128 , n408634 , n408635 , n86131 , n408637 , n408638 , n408639 , n408640 , n408641 , n408642 , 
 n408643 , n408644 , n408645 , n408646 , n408647 , n86137 , n408649 , n408650 , n86140 , n408652 , 
 n408653 , n86143 , n408655 , n408656 , n408657 , n86147 , n408659 , n408660 , n408661 , n408662 , 
 n408663 , n408664 , n408665 , n408666 , n86156 , n86157 , n408669 , n408670 , n86160 , n86161 , 
 n408673 , n408674 , n408675 , n408676 , n408677 , n408678 , n408679 , n408680 , n408681 , n408682 , 
 n408683 , n408684 , n86172 , n408686 , n408687 , n408688 , n408689 , n86177 , n408691 , n86179 , 
 n408693 , n408694 , n408695 , n86183 , n408697 , n408698 , n86186 , n408700 , n408701 , n408702 , 
 n408703 , n86191 , n86192 , n408706 , n408707 , n408708 , n408709 , n408710 , n408711 , n408712 , 
 n408713 , n408714 , n86202 , n408716 , n408717 , n86205 , n408719 , n408720 , n408721 , n408722 , 
 n408723 , n408724 , n408725 , n408726 , n408727 , n408728 , n408729 , n86217 , n408731 , n408732 , 
 n408733 , n408734 , n408735 , n86223 , n408737 , n408738 , n86226 , n408740 , n408741 , n408742 , 
 n408743 , n408744 , n408745 , n86233 , n408747 , n408748 , n86236 , n408750 , n408751 , n86239 , 
 n408753 , n408754 , n408755 , n408756 , n86244 , n408758 , n408759 , n408760 , n408761 , n408762 , 
 n408763 , n408764 , n408765 , n408766 , n86254 , n408768 , n86256 , n86257 , n408771 , n86259 , 
 n408773 , n86261 , n86262 , n86263 , n86264 , n86265 , n408779 , n86267 , n408781 , n408782 , 
 n408783 , n86271 , n408785 , n86273 , n408787 , n408788 , n408789 , n86277 , n408791 , n408792 , 
 n408793 , n408794 , n408795 , n408796 , n408797 , n408798 , n408799 , n86287 , n86288 , n86289 , 
 n86290 , n408804 , n408805 , n86293 , n408807 , n408808 , n86296 , n408810 , n86298 , n408812 , 
 n408813 , n408814 , n86302 , n408816 , n408817 , n408818 , n408819 , n408820 , n408821 , n408822 , 
 n408823 , n408824 , n408825 , n408826 , n408827 , n408828 , n86316 , n408830 , n408831 , n408832 , 
 n86320 , n408834 , n408835 , n408836 , n86324 , n408838 , n86326 , n86327 , n86328 , n408842 , 
 n86330 , n408844 , n408845 , n408846 , n408847 , n408848 , n408849 , n408850 , n408851 , n408852 , 
 n86340 , n86341 , n86342 , n86343 , n408857 , n86345 , n408859 , n408860 , n408861 , n86349 , 
 n408863 , n86351 , n408865 , n408866 , n86354 , n408868 , n86356 , n408870 , n408871 , n408872 , 
 n408873 , n408874 , n86362 , n408876 , n408877 , n86365 , n408879 , n408880 , n408881 , n408882 , 
 n408883 , n408884 , n408885 , n408886 , n408887 , n408888 , n408889 , n408890 , n408891 , n408892 , 
 n86380 , n408894 , n408895 , n86383 , n86384 , n86385 , n86386 , n86387 , n408901 , n408902 , 
 n86390 , n408904 , n86392 , n408906 , n408907 , n86395 , n408909 , n408910 , n86398 , n408912 , 
 n408913 , n408914 , n408915 , n408916 , n86404 , n408918 , n408919 , n408920 , n408921 , n408922 , 
 n408923 , n408924 , n86412 , n408926 , n408927 , n408928 , n408929 , n408930 , n86418 , n86419 , 
 n408933 , n408934 , n408935 , n86423 , n408937 , n86425 , n408939 , n408940 , n408941 , n408942 , 
 n86430 , n408944 , n408945 , n408946 , n86434 , n408948 , n408949 , n86437 , n408951 , n86439 , 
 n408953 , n408954 , n86442 , n408956 , n408957 , n86445 , n408959 , n408960 , n86448 , n408962 , 
 n86450 , n86451 , n408965 , n408966 , n86454 , n408968 , n408969 , n86457 , n408971 , n408972 , 
 n408973 , n86461 , n86462 , n408976 , n408977 , n408978 , n86466 , n408980 , n408981 , n408982 , 
 n408983 , n408984 , n408985 , n408986 , n408987 , n408988 , n408989 , n408990 , n408991 , n408992 , 
 n86480 , n86481 , n408995 , n408996 , n86484 , n408998 , n408999 , n86487 , n409001 , n409002 , 
 n409003 , n409004 , n409005 , n409006 , n409007 , n409008 , n409009 , n409010 , n409011 , n409012 , 
 n409013 , n86501 , n409015 , n409016 , n86504 , n409018 , n409019 , n409020 , n409021 , n409022 , 
 n409023 , n86511 , n86512 , n409026 , n86514 , n409028 , n409029 , n409030 , n409031 , n409032 , 
 n86520 , n409034 , n409035 , n409036 , n86524 , n409038 , n409039 , n86527 , n409041 , n409042 , 
 n409043 , n409044 , n409045 , n409046 , n86534 , n409048 , n409049 , n409050 , n409051 , n409052 , 
 n409053 , n409054 , n409055 , n409056 , n86544 , n86545 , n409059 , n86547 , n409061 , n409062 , 
 n86550 , n409064 , n409065 , n86553 , n409067 , n409068 , n86556 , n86557 , n409071 , n86559 , 
 n86560 , n409074 , n409075 , n86563 , n409077 , n409078 , n409079 , n409080 , n409081 , n409082 , 
 n409083 , n409084 , n409085 , n409086 , n409087 , n409088 , n86576 , n409090 , n86578 , n409092 , 
 n409093 , n409094 , n409095 , n86583 , n409097 , n86585 , n86586 , n409100 , n86588 , n409102 , 
 n86590 , n86591 , n409105 , n409106 , n86594 , n409108 , n409109 , n409110 , n409111 , n409112 , 
 n409113 , n86601 , n409115 , n409116 , n86604 , n86605 , n409119 , n86607 , n409121 , n409122 , 
 n409123 , n409124 , n409125 , n86613 , n409127 , n409128 , n409129 , n86617 , n409131 , n86619 , 
 n86620 , n409134 , n409135 , n409136 , n409137 , n409138 , n86626 , n409140 , n409141 , n86629 , 
 n409143 , n86631 , n409145 , n409146 , n409147 , n409148 , n86636 , n409150 , n409151 , n409152 , 
 n409153 , n86641 , n409155 , n409156 , n86644 , n409158 , n409159 , n409160 , n86648 , n409162 , 
 n86650 , n409164 , n409165 , n409166 , n86654 , n409168 , n409169 , n409170 , n409171 , n409172 , 
 n409173 , n409174 , n86662 , n409176 , n409177 , n409178 , n409179 , n409180 , n409181 , n409182 , 
 n409183 , n409184 , n409185 , n86673 , n409187 , n409188 , n86676 , n86677 , n86678 , n409192 , 
 n409193 , n409194 , n86682 , n409196 , n86684 , n409198 , n86686 , n86687 , n409201 , n409202 , 
 n86690 , n409204 , n409205 , n86693 , n409207 , n409208 , n86696 , n409210 , n409211 , n409212 , 
 n409213 , n409214 , n409215 , n409216 , n409217 , n409218 , n409219 , n409220 , n409221 , n409222 , 
 n86710 , n86711 , n86712 , n86713 , n86714 , n409228 , n409229 , n409230 , n409231 , n409232 , 
 n86720 , n409234 , n409235 , n409236 , n409237 , n409238 , n409239 , n409240 , n86728 , n86729 , 
 n409243 , n86731 , n409245 , n409246 , n409247 , n409248 , n409249 , n409250 , n409251 , n409252 , 
 n409253 , n409254 , n409255 , n409256 , n409257 , n409258 , n86746 , n409260 , n409261 , n409262 , 
 n86750 , n86751 , n409265 , n86753 , n409267 , n409268 , n409269 , n409270 , n409271 , n409272 , 
 n409273 , n409274 , n86762 , n409276 , n409277 , n409278 , n409279 , n409280 , n409281 , n409282 , 
 n409283 , n409284 , n409285 , n409286 , n86774 , n86775 , n409289 , n409290 , n409291 , n409292 , 
 n409293 , n86781 , n409295 , n409296 , n86784 , n409298 , n86786 , n86787 , n409301 , n409302 , 
 n409303 , n409304 , n86792 , n409306 , n86794 , n409308 , n86796 , n86797 , n409311 , n86799 , 
 n409313 , n86801 , n409315 , n409316 , n409317 , n86805 , n86806 , n409320 , n409321 , n409322 , 
 n409323 , n86811 , n409325 , n409326 , n86814 , n409328 , n86816 , n86817 , n86818 , n409332 , 
 n409333 , n86821 , n86822 , n409336 , n409337 , n86825 , n409339 , n409340 , n86828 , n409342 , 
 n409343 , n409344 , n86832 , n409346 , n86834 , n86835 , n409349 , n409350 , n86838 , n409352 , 
 n409353 , n409354 , n409355 , n409356 , n86844 , n409358 , n409359 , n86847 , n409361 , n409362 , 
 n409363 , n409364 , n409365 , n409366 , n409367 , n409368 , n86856 , n409370 , n409371 , n409372 , 
 n409373 , n409374 , n409375 , n409376 , n409377 , n409378 , n409379 , n409380 , n409381 , n409382 , 
 n409383 , n409384 , n409385 , n86873 , n409387 , n86875 , n409389 , n409390 , n409391 , n86879 , 
 n409393 , n409394 , n409395 , n409396 , n409397 , n86885 , n409399 , n86887 , n409401 , n409402 , 
 n409403 , n86891 , n409405 , n409406 , n409407 , n409408 , n409409 , n409410 , n409411 , n409412 , 
 n409413 , n86901 , n409415 , n409416 , n86904 , n409418 , n409419 , n86907 , n409421 , n409422 , 
 n86910 , n409424 , n409425 , n86913 , n86914 , n409428 , n409429 , n86917 , n409431 , n409432 , 
 n409433 , n409434 , n86922 , n409436 , n86924 , n409438 , n409439 , n86927 , n86928 , n409442 , 
 n409443 , n409444 , n409445 , n86933 , n409447 , n409448 , n86936 , n409450 , n409451 , n86939 , 
 n86940 , n409454 , n86942 , n409456 , n409457 , n86945 , n86946 , n409460 , n409461 , n409462 , 
 n86950 , n86951 , n409465 , n409466 , n409467 , n409468 , n409469 , n409470 , n409471 , n409472 , 
 n409473 , n409474 , n86962 , n86963 , n409477 , n86965 , n409479 , n409480 , n409481 , n86969 , 
 n86970 , n409484 , n409485 , n86973 , n86974 , n409488 , n409489 , n409490 , n86978 , n409492 , 
 n409493 , n409494 , n409495 , n409496 , n86984 , n86985 , n409499 , n409500 , n86988 , n409502 , 
 n409503 , n409504 , n409505 , n409506 , n409507 , n409508 , n409509 , n409510 , n409511 , n409512 , 
 n409513 , n409514 , n409515 , n409516 , n409517 , n87005 , n409519 , n409520 , n409521 , n409522 , 
 n409523 , n409524 , n409525 , n409526 , n409527 , n409528 , n409529 , n409530 , n409531 , n409532 , 
 n409533 , n87021 , n409535 , n409536 , n409537 , n409538 , n87026 , n409540 , n87028 , n87029 , 
 n409543 , n409544 , n409545 , n87033 , n409547 , n409548 , n87036 , n87037 , n87038 , n87039 , 
 n87040 , n87041 , n409555 , n409556 , n409557 , n409558 , n409559 , n87047 , n409561 , n409562 , 
 n409563 , n409564 , n87052 , n409566 , n409567 , n409568 , n87056 , n409570 , n409571 , n409572 , 
 n409573 , n409574 , n87062 , n409576 , n409577 , n409578 , n409579 , n87067 , n87068 , n87069 , 
 n87070 , n87071 , n87072 , n87073 , n87074 , n87075 , n87076 , n409590 , n409591 , n409592 , 
 n409593 , n409594 , n409595 , n409596 , n87084 , n409598 , n409599 , n87087 , n409601 , n409602 , 
 n409603 , n409604 , n87092 , n409606 , n409607 , n409608 , n409609 , n409610 , n87098 , n409612 , 
 n409613 , n409614 , n87102 , n409616 , n409617 , n409618 , n409619 , n409620 , n409621 , n409622 , 
 n409623 , n409624 , n409625 , n409626 , n409627 , n87115 , n409629 , n409630 , n87118 , n409632 , 
 n409633 , n409634 , n409635 , n409636 , n87124 , n409638 , n409639 , n409640 , n409641 , n409642 , 
 n409643 , n409644 , n87132 , n87133 , n87134 , n87135 , n87136 , n87137 , n409651 , n409652 , 
 n409653 , n409654 , n409655 , n409656 , n409657 , n87145 , n409659 , n409660 , n87148 , n409662 , 
 n409663 , n409664 , n87152 , n409666 , n409667 , n87155 , n409669 , n409670 , n87158 , n409672 , 
 n409673 , n409674 , n409675 , n409676 , n409677 , n409678 , n409679 , n409680 , n409681 , n409682 , 
 n409683 , n87171 , n87172 , n409686 , n87174 , n409688 , n409689 , n87177 , n409691 , n87179 , 
 n87180 , n87181 , n409695 , n409696 , n409697 , n87185 , n409699 , n87187 , n409701 , n409702 , 
 n87190 , n87191 , n409705 , n87193 , n87194 , n409708 , n409709 , n409710 , n409711 , n87199 , 
 n409713 , n409714 , n409715 , n409716 , n409717 , n409718 , n87203 , n87204 , n409721 , n409722 , 
 n87207 , n409724 , n409725 , n409726 , n87211 , n409728 , n409729 , n87214 , n409731 , n409732 , 
 n409733 , n87218 , n409735 , n87220 , n409737 , n87222 , n87223 , n409740 , n409741 , n87226 , 
 n409743 , n409744 , n87229 , n409746 , n409747 , n87232 , n409749 , n409750 , n409751 , n409752 , 
 n87237 , n409754 , n87239 , n87240 , n409757 , n409758 , n409759 , n409760 , n409761 , n409762 , 
 n409763 , n87248 , n87249 , n409766 , n87251 , n409768 , n409769 , n87254 , n409771 , n409772 , 
 n409773 , n409774 , n409775 , n409776 , n409777 , n409778 , n87263 , n409780 , n409781 , n409782 , 
 n409783 , n409784 , n409785 , n409786 , n87271 , n409788 , n409789 , n409790 , n87275 , n409792 , 
 n409793 , n409794 , n409795 , n409796 , n409797 , n409798 , n87283 , n87284 , n409801 , n409802 , 
 n409803 , n87288 , n409805 , n409806 , n409807 , n87292 , n87293 , n87294 , n409811 , n409812 , 
 n87297 , n409814 , n409815 , n87300 , n409817 , n409818 , n409819 , n409820 , n409821 , n409822 , 
 n409823 , n409824 , n409825 , n409826 , n87311 , n409828 , n87313 , n409830 , n409831 , n409832 , 
 n87317 , n409834 , n87319 , n409836 , n409837 , n409838 , n409839 , n409840 , n409841 , n409842 , 
 n87327 , n87328 , n409845 , n409846 , n409847 , n409848 , n409849 , n409850 , n87335 , n87336 , 
 n409853 , n87338 , n409855 , n409856 , n409857 , n409858 , n409859 , n409860 , n409861 , n409862 , 
 n409863 , n409864 , n409865 , n409866 , n87351 , n409868 , n409869 , n87354 , n409871 , n409872 , 
 n409873 , n409874 , n409875 , n409876 , n409877 , n87362 , n409879 , n409880 , n409881 , n87366 , 
 n409883 , n409884 , n87369 , n409886 , n409887 , n409888 , n87373 , n87374 , n409891 , n409892 , 
 n409893 , n87378 , n409895 , n409896 , n87381 , n409898 , n87383 , n409900 , n409901 , n409902 , 
 n409903 , n409904 , n409905 , n87390 , n409907 , n409908 , n87393 , n87394 , n409911 , n409912 , 
 n87397 , n409914 , n409915 , n87400 , n409917 , n409918 , n87403 , n409920 , n87405 , n409922 , 
 n409923 , n409924 , n409925 , n409926 , n409927 , n409928 , n87413 , n87414 , n409931 , n409932 , 
 n409933 , n409934 , n409935 , n87420 , n409937 , n409938 , n409939 , n409940 , n409941 , n409942 , 
 n409943 , n409944 , n409945 , n409946 , n409947 , n409948 , n409949 , n409950 , n409951 , n87436 , 
 n409953 , n409954 , n409955 , n409956 , n409957 , n409958 , n409959 , n409960 , n409961 , n409962 , 
 n409963 , n87448 , n409965 , n409966 , n409967 , n409968 , n409969 , n409970 , n409971 , n87456 , 
 n409973 , n409974 , n87459 , n409976 , n409977 , n409978 , n409979 , n409980 , n409981 , n409982 , 
 n409983 , n409984 , n87469 , n409986 , n87471 , n87472 , n87473 , n409990 , n409991 , n409992 , 
 n87477 , n409994 , n409995 , n87480 , n87481 , n409998 , n409999 , n87484 , n410001 , n410002 , 
 n87487 , n410004 , n410005 , n87490 , n87491 , n410008 , n410009 , n87494 , n410011 , n87496 , 
 n87497 , n87498 , n410015 , n410016 , n87501 , n87502 , n410019 , n410020 , n410021 , n410022 , 
 n87507 , n410024 , n87509 , n410026 , n87511 , n410028 , n410029 , n410030 , n410031 , n410032 , 
 n410033 , n410034 , n410035 , n410036 , n410037 , n410038 , n87523 , n410040 , n410041 , n410042 , 
 n87527 , n87528 , n410045 , n87530 , n410047 , n410048 , n410049 , n410050 , n410051 , n87536 , 
 n87537 , n410054 , n87539 , n410056 , n87541 , n87542 , n410059 , n410060 , n87545 , n410062 , 
 n410063 , n410064 , n410065 , n410066 , n410067 , n410068 , n410069 , n410070 , n87555 , n410072 , 
 n410073 , n87558 , n87559 , n87560 , n87561 , n87562 , n410079 , n410080 , n87565 , n87566 , 
 n87567 , n410084 , n410085 , n87570 , n410087 , n410088 , n410089 , n87574 , n410091 , n410092 , 
 n410093 , n87578 , n410095 , n410096 , n87581 , n410098 , n410099 , n410100 , n410101 , n410102 , 
 n410103 , n410104 , n410105 , n410106 , n410107 , n410108 , n410109 , n410110 , n410111 , n410112 , 
 n410113 , n410114 , n87599 , n410116 , n410117 , n410118 , n410119 , n410120 , n410121 , n410122 , 
 n410123 , n410124 , n410125 , n87610 , n87611 , n410128 , n87613 , n410130 , n410131 , n87616 , 
 n87617 , n410134 , n410135 , n87620 , n410137 , n410138 , n87623 , n410140 , n410141 , n410142 , 
 n410143 , n87628 , n87629 , n87630 , n410147 , n410148 , n87633 , n410150 , n87635 , n410152 , 
 n410153 , n410154 , n410155 , n410156 , n410157 , n410158 , n410159 , n410160 , n410161 , n410162 , 
 n87647 , n410164 , n410165 , n410166 , n87651 , n87652 , n410169 , n87654 , n410171 , n410172 , 
 n410173 , n410174 , n410175 , n410176 , n87658 , n410178 , n87660 , n87661 , n410181 , n410182 , 
 n410183 , n410184 , n87666 , n410186 , n410187 , n410188 , n410189 , n410190 , n410191 , n410192 , 
 n410193 , n410194 , n410195 , n410196 , n410197 , n410198 , n87680 , n410200 , n410201 , n410202 , 
 n410203 , n410204 , n410205 , n410206 , n410207 , n410208 , n410209 , n410210 , n410211 , n410212 , 
 n410213 , n410214 , n87696 , n410216 , n410217 , n87699 , n410219 , n410220 , n410221 , n410222 , 
 n410223 , n410224 , n410225 , n410226 , n410227 , n87709 , n410229 , n410230 , n410231 , n410232 , 
 n410233 , n410234 , n410235 , n410236 , n87718 , n410238 , n87720 , n87721 , n410241 , n410242 , 
 n410243 , n410244 , n87726 , n410246 , n410247 , n410248 , n410249 , n410250 , n410251 , n410252 , 
 n410253 , n410254 , n410255 , n87737 , n87738 , n410258 , n87740 , n410260 , n87742 , n410262 , 
 n410263 , n410264 , n410265 , n87747 , n410267 , n410268 , n87750 , n410270 , n410271 , n87753 , 
 n87754 , n87755 , n87756 , n410276 , n410277 , n87759 , n87760 , n410280 , n87762 , n87763 , 
 n410283 , n410284 , n410285 , n410286 , n410287 , n410288 , n87770 , n410290 , n87772 , n87773 , 
 n410293 , n410294 , n87776 , n410296 , n410297 , n410298 , n410299 , n410300 , n87782 , n410302 , 
 n87784 , n87785 , n410305 , n87787 , n410307 , n87789 , n87790 , n410310 , n410311 , n87793 , 
 n410313 , n410314 , n87796 , n87797 , n87798 , n410318 , n410319 , n87801 , n410321 , n410322 , 
 n410323 , n87805 , n410325 , n410326 , n410327 , n87809 , n410329 , n410330 , n87812 , n410332 , 
 n410333 , n410334 , n410335 , n410336 , n410337 , n410338 , n410339 , n87821 , n87822 , n410342 , 
 n410343 , n410344 , n87826 , n410346 , n410347 , n87829 , n410349 , n410350 , n410351 , n87833 , 
 n410353 , n410354 , n87836 , n410356 , n410357 , n410358 , n87840 , n410360 , n410361 , n87843 , 
 n87844 , n410364 , n410365 , n87847 , n410367 , n410368 , n410369 , n87851 , n410371 , n410372 , 
 n410373 , n410374 , n87856 , n410376 , n410377 , n87859 , n410379 , n410380 , n410381 , n410382 , 
 n410383 , n87865 , n410385 , n410386 , n410387 , n410388 , n410389 , n410390 , n87872 , n410392 , 
 n410393 , n87875 , n410395 , n410396 , n410397 , n410398 , n87880 , n410400 , n410401 , n410402 , 
 n410403 , n410404 , n410405 , n410406 , n87888 , n410408 , n410409 , n87891 , n410411 , n410412 , 
 n410413 , n410414 , n87896 , n410416 , n87898 , n410418 , n410419 , n410420 , n87902 , n410422 , 
 n410423 , n87905 , n410425 , n410426 , n87908 , n410428 , n410429 , n87911 , n410431 , n410432 , 
 n87914 , n410434 , n410435 , n87917 , n410437 , n410438 , n87920 , n410440 , n87922 , n87923 , 
 n410443 , n410444 , n87926 , n410446 , n410447 , n87929 , n87930 , n410450 , n410451 , n87933 , 
 n410453 , n87935 , n410455 , n410456 , n87938 , n410458 , n410459 , n410460 , n410461 , n410462 , 
 n410463 , n410464 , n410465 , n87947 , n410467 , n410468 , n410469 , n410470 , n410471 , n410472 , 
 n410473 , n410474 , n410475 , n410476 , n87958 , n410478 , n410479 , n410480 , n410481 , n410482 , 
 n410483 , n410484 , n410485 , n87967 , n87968 , n410488 , n410489 , n410490 , n410491 , n87973 , 
 n87974 , n410494 , n410495 , n410496 , n410497 , n410498 , n87980 , n410500 , n87982 , n87983 , 
 n410503 , n410504 , n87986 , n410506 , n410507 , n87989 , n87990 , n410510 , n87992 , n410512 , 
 n87994 , n87995 , n410515 , n410516 , n87998 , n410518 , n410519 , n410520 , n410521 , n410522 , 
 n88004 , n88005 , n88006 , n410526 , n410527 , n88009 , n410529 , n410530 , n88012 , n410532 , 
 n410533 , n88015 , n410535 , n88017 , n88018 , n410538 , n410539 , n88021 , n410541 , n410542 , 
 n88024 , n410544 , n410545 , n88027 , n410547 , n410548 , n88030 , n410550 , n88032 , n410552 , 
 n410553 , n88035 , n410555 , n88037 , n88038 , n410558 , n410559 , n410560 , n88042 , n88043 , 
 n410563 , n410564 , n88046 , n410566 , n88048 , n410568 , n88050 , n410570 , n410571 , n88053 , 
 n410573 , n88055 , n88056 , n410576 , n88058 , n410578 , n410579 , n410580 , n410581 , n410582 , 
 n410583 , n410584 , n410585 , n410586 , n410587 , n410588 , n410589 , n410590 , n410591 , n410592 , 
 n410593 , n410594 , n410595 , n410596 , n410597 , n410598 , n410599 , n410600 , n410601 , n410602 , 
 n410603 , n410604 , n88086 , n410606 , n88088 , n410608 , n410609 , n88091 , n410611 , n88093 , 
 n88094 , n410614 , n410615 , n410616 , n410617 , n410618 , n410619 , n410620 , n410621 , n410622 , 
 n88104 , n410624 , n410625 , n88107 , n410627 , n410628 , n88110 , n410630 , n410631 , n88113 , 
 n88114 , n410634 , n410635 , n88117 , n410637 , n410638 , n88120 , n410640 , n410641 , n410642 , 
 n410643 , n410644 , n410645 , n88127 , n410647 , n410648 , n410649 , n410650 , n410651 , n410652 , 
 n88134 , n410654 , n410655 , n410656 , n88138 , n410658 , n410659 , n88141 , n410661 , n410662 , 
 n410663 , n410664 , n410665 , n88147 , n410667 , n410668 , n410669 , n410670 , n410671 , n410672 , 
 n410673 , n410674 , n410675 , n410676 , n88158 , n410678 , n410679 , n88161 , n88162 , n88163 , 
 n88164 , n88165 , n88166 , n88167 , n410687 , n410688 , n410689 , n410690 , n88172 , n410692 , 
 n410693 , n410694 , n88176 , n410696 , n410697 , n88179 , n410699 , n410700 , n410701 , n410702 , 
 n410703 , n410704 , n410705 , n410706 , n88188 , n410708 , n410709 , n88191 , n410711 , n410712 , 
 n88194 , n410714 , n410715 , n88197 , n88198 , n410718 , n88200 , n410720 , n88202 , n410722 , 
 n410723 , n410724 , n410725 , n410726 , n410727 , n88209 , n88210 , n410730 , n88212 , n410732 , 
 n88214 , n410734 , n410735 , n88217 , n410737 , n88219 , n88220 , n88221 , n88222 , n410742 , 
 n88224 , n410744 , n410745 , n410746 , n88228 , n88229 , n410749 , n410750 , n88232 , n88233 , 
 n88234 , n410754 , n410755 , n410756 , n88238 , n410758 , n410759 , n410760 , n88242 , n410762 , 
 n410763 , n410764 , n410765 , n410766 , n410767 , n410768 , n410769 , n410770 , n88247 , n88248 , 
 n410773 , n410774 , n410775 , n410776 , n410777 , n88254 , n410779 , n410780 , n88257 , n410782 , 
 n410783 , n410784 , n410785 , n88262 , n410787 , n88264 , n88265 , n410790 , n410791 , n88268 , 
 n88269 , n410794 , n410795 , n88272 , n88273 , n410798 , n410799 , n88276 , n88277 , n88278 , 
 n410803 , n410804 , n88281 , n88282 , n410807 , n410808 , n88285 , n88286 , n88287 , n410812 , 
 n410813 , n410814 , n88291 , n410816 , n410817 , n410818 , n88295 , n88296 , n88297 , n410822 , 
 n410823 , n88300 , n410825 , n88302 , n410827 , n88304 , n88305 , n88306 , n410831 , n410832 , 
 n88309 , n410834 , n410835 , n88312 , n410837 , n410838 , n410839 , n410840 , n410841 , n88318 , 
 n410843 , n410844 , n88321 , n410846 , n410847 , n410848 , n410849 , n410850 , n410851 , n410852 , 
 n410853 , n410854 , n88331 , n410856 , n410857 , n88334 , n410859 , n410860 , n410861 , n410862 , 
 n410863 , n410864 , n410865 , n410866 , n88343 , n410868 , n410869 , n410870 , n410871 , n88348 , 
 n410873 , n410874 , n88351 , n410876 , n88353 , n88354 , n410879 , n410880 , n410881 , n410882 , 
 n410883 , n410884 , n410885 , n410886 , n410887 , n88364 , n410889 , n88366 , n410891 , n88368 , 
 n410893 , n410894 , n410895 , n410896 , n88373 , n410898 , n410899 , n410900 , n410901 , n410902 , 
 n410903 , n88380 , n410905 , n410906 , n410907 , n410908 , n410909 , n410910 , n410911 , n410912 , 
 n410913 , n410914 , n88391 , n88392 , n410917 , n410918 , n88395 , n410920 , n410921 , n410922 , 
 n410923 , n410924 , n88401 , n410926 , n410927 , n410928 , n410929 , n410930 , n410931 , n410932 , 
 n410933 , n410934 , n410935 , n410936 , n410937 , n410938 , n88415 , n410940 , n410941 , n88418 , 
 n410943 , n410944 , n410945 , n410946 , n410947 , n410948 , n410949 , n410950 , n410951 , n410952 , 
 n410953 , n410954 , n410955 , n410956 , n410957 , n88434 , n410959 , n88436 , n410961 , n88438 , 
 n410963 , n410964 , n410965 , n410966 , n410967 , n410968 , n410969 , n410970 , n88447 , n410972 , 
 n410973 , n410974 , n88451 , n410976 , n410977 , n410978 , n410979 , n410980 , n410981 , n410982 , 
 n410983 , n88460 , n410985 , n88462 , n88463 , n410988 , n410989 , n88466 , n410991 , n410992 , 
 n88469 , n410994 , n410995 , n410996 , n88473 , n88474 , n410999 , n411000 , n411001 , n88478 , 
 n88479 , n411004 , n411005 , n411006 , n88483 , n411008 , n411009 , n88486 , n411011 , n411012 , 
 n411013 , n411014 , n411015 , n411016 , n411017 , n88494 , n88495 , n411020 , n411021 , n411022 , 
 n411023 , n88500 , n411025 , n411026 , n411027 , n411028 , n411029 , n411030 , n411031 , n411032 , 
 n411033 , n411034 , n411035 , n411036 , n88513 , n411038 , n411039 , n88516 , n411041 , n411042 , 
 n411043 , n411044 , n88521 , n411046 , n411047 , n88524 , n411049 , n411050 , n88527 , n411052 , 
 n411053 , n88530 , n411055 , n411056 , n88533 , n411058 , n411059 , n411060 , n411061 , n411062 , 
 n411063 , n411064 , n411065 , n411066 , n88543 , n411068 , n88545 , n411070 , n411071 , n88548 , 
 n411073 , n88550 , n88551 , n411076 , n411077 , n88554 , n411079 , n411080 , n88557 , n411082 , 
 n411083 , n411084 , n88561 , n411086 , n411087 , n88564 , n411089 , n411090 , n88567 , n88568 , 
 n88569 , n88570 , n88571 , n88572 , n411097 , n411098 , n411099 , n411100 , n411101 , n411102 , 
 n88579 , n88580 , n411105 , n88582 , n411107 , n88584 , n88585 , n411110 , n411111 , n88588 , 
 n411113 , n411114 , n88591 , n411116 , n411117 , n411118 , n88595 , n411120 , n411121 , n411122 , 
 n411123 , n411124 , n88601 , n411126 , n411127 , n88604 , n411129 , n411130 , n411131 , n88608 , 
 n411133 , n88610 , n88611 , n411136 , n88613 , n88614 , n88615 , n411140 , n411141 , n88618 , 
 n88619 , n88620 , n411145 , n411146 , n88623 , n88624 , n411149 , n411150 , n88627 , n411152 , 
 n88629 , n411154 , n88631 , n411156 , n411157 , n411158 , n411159 , n411160 , n88637 , n411162 , 
 n411163 , n88640 , n411165 , n411166 , n88643 , n411168 , n411169 , n411170 , n411171 , n88648 , 
 n411173 , n411174 , n411175 , n411176 , n411177 , n88654 , n411179 , n88656 , n411181 , n411182 , 
 n88659 , n411184 , n88661 , n411186 , n411187 , n411188 , n88665 , n411190 , n411191 , n411192 , 
 n411193 , n88670 , n88671 , n88672 , n88673 , n88674 , n88675 , n88676 , n411201 , n88678 , 
 n411203 , n411204 , n88681 , n88682 , n88683 , n411208 , n411209 , n411210 , n411211 , n411212 , 
 n411213 , n411214 , n88691 , n411216 , n411217 , n411218 , n88695 , n88696 , n411221 , n411222 , 
 n88699 , n88700 , n411225 , n411226 , n411227 , n411228 , n411229 , n411230 , n411231 , n411232 , 
 n411233 , n88706 , n411235 , n411236 , n88709 , n411238 , n411239 , n411240 , n88713 , n88714 , 
 n88715 , n411244 , n88717 , n411246 , n411247 , n88720 , n411249 , n411250 , n411251 , n411252 , 
 n411253 , n411254 , n88727 , n88728 , n411257 , n88730 , n411259 , n88732 , n411261 , n411262 , 
 n88735 , n411264 , n88737 , n411266 , n411267 , n88740 , n411269 , n411270 , n88743 , n411272 , 
 n411273 , n411274 , n411275 , n411276 , n411277 , n411278 , n411279 , n411280 , n411281 , n411282 , 
 n411283 , n411284 , n411285 , n411286 , n88759 , n411288 , n411289 , n411290 , n411291 , n88764 , 
 n411293 , n411294 , n88767 , n411296 , n411297 , n411298 , n411299 , n411300 , n88773 , n411302 , 
 n411303 , n411304 , n411305 , n411306 , n411307 , n88780 , n411309 , n411310 , n411311 , n411312 , 
 n411313 , n411314 , n411315 , n411316 , n411317 , n88790 , n411319 , n411320 , n411321 , n411322 , 
 n411323 , n411324 , n411325 , n88798 , n88799 , n411328 , n411329 , n88802 , n411331 , n411332 , 
 n411333 , n411334 , n411335 , n411336 , n88809 , n88810 , n88811 , n411340 , n411341 , n411342 , 
 n411343 , n88816 , n411345 , n411346 , n411347 , n411348 , n411349 , n88822 , n411351 , n411352 , 
 n88825 , n411354 , n411355 , n411356 , n411357 , n411358 , n88831 , n411360 , n411361 , n88834 , 
 n88835 , n411364 , n411365 , n88838 , n88839 , n411368 , n88841 , n411370 , n411371 , n411372 , 
 n411373 , n411374 , n88847 , n411376 , n411377 , n88850 , n411379 , n411380 , n411381 , n411382 , 
 n411383 , n88856 , n411385 , n411386 , n411387 , n88860 , n411389 , n411390 , n411391 , n411392 , 
 n411393 , n411394 , n411395 , n411396 , n411397 , n411398 , n411399 , n411400 , n411401 , n411402 , 
 n411403 , n88876 , n88877 , n411406 , n411407 , n88880 , n411409 , n88882 , n411411 , n411412 , 
 n411413 , n411414 , n411415 , n411416 , n88889 , n411418 , n411419 , n411420 , n411421 , n411422 , 
 n411423 , n411424 , n411425 , n411426 , n411427 , n88900 , n88901 , n88902 , n411431 , n88904 , 
 n411433 , n411434 , n411435 , n411436 , n411437 , n411438 , n411439 , n411440 , n411441 , n88914 , 
 n411443 , n411444 , n411445 , n411446 , n411447 , n411448 , n411449 , n88922 , n411451 , n411452 , 
 n88925 , n411454 , n411455 , n88928 , n411457 , n411458 , n411459 , n411460 , n411461 , n411462 , 
 n411463 , n411464 , n411465 , n411466 , n411467 , n88940 , n411469 , n411470 , n88943 , n411472 , 
 n411473 , n88946 , n88947 , n88948 , n411477 , n411478 , n88951 , n411480 , n88953 , n411482 , 
 n88955 , n88956 , n411485 , n88958 , n411487 , n88960 , n411489 , n411490 , n411491 , n411492 , 
 n411493 , n411494 , n411495 , n411496 , n411497 , n411498 , n88971 , n411500 , n411501 , n88974 , 
 n411503 , n411504 , n88977 , n411506 , n411507 , n411508 , n411509 , n411510 , n411511 , n411512 , 
 n411513 , n411514 , n88987 , n411516 , n88989 , n88990 , n88991 , n88992 , n411521 , n411522 , 
 n88995 , n411524 , n411525 , n411526 , n411527 , n411528 , n89001 , n89002 , n411531 , n411532 , 
 n411533 , n89006 , n89007 , n89008 , n411537 , n411538 , n89011 , n411540 , n411541 , n411542 , 
 n411543 , n411544 , n411545 , n411546 , n89019 , n411548 , n89021 , n411550 , n411551 , n89024 , 
 n411553 , n411554 , n411555 , n411556 , n411557 , n89030 , n411559 , n411560 , n89033 , n411562 , 
 n411563 , n411564 , n411565 , n89038 , n411567 , n411568 , n89041 , n411570 , n411571 , n411572 , 
 n411573 , n89046 , n411575 , n411576 , n89049 , n411578 , n411579 , n411580 , n411581 , n411582 , 
 n411583 , n411584 , n411585 , n411586 , n411587 , n411588 , n411589 , n89062 , n89063 , n89064 , 
 n411593 , n411594 , n411595 , n411596 , n411597 , n411598 , n411599 , n411600 , n411601 , n411602 , 
 n89074 , n411604 , n411605 , n411606 , n411607 , n411608 , n411609 , n411610 , n411611 , n411612 , 
 n411613 , n89085 , n411615 , n411616 , n89088 , n411618 , n411619 , n89091 , n411621 , n411622 , 
 n89094 , n411624 , n411625 , n411626 , n411627 , n411628 , n411629 , n411630 , n411631 , n411632 , 
 n411633 , n411634 , n411635 , n411636 , n411637 , n411638 , n89110 , n411640 , n411641 , n411642 , 
 n411643 , n411644 , n411645 , n411646 , n89118 , n411648 , n411649 , n89121 , n411651 , n411652 , 
 n411653 , n411654 , n411655 , n411656 , n411657 , n411658 , n89130 , n411660 , n411661 , n89133 , 
 n411663 , n89135 , n89136 , n411666 , n411667 , n89139 , n89140 , n411670 , n411671 , n89143 , 
 n89144 , n89145 , n89146 , n411676 , n411677 , n89149 , n411679 , n411680 , n411681 , n89153 , 
 n411683 , n89155 , n411685 , n411686 , n89158 , n411688 , n411689 , n411690 , n411691 , n411692 , 
 n89164 , n89165 , n89166 , n411696 , n411697 , n89169 , n411699 , n89171 , n411701 , n411702 , 
 n411703 , n89175 , n411705 , n411706 , n411707 , n89179 , n89180 , n411710 , n411711 , n411712 , 
 n411713 , n411714 , n89186 , n411716 , n411717 , n411718 , n411719 , n89191 , n89192 , n411722 , 
 n411723 , n411724 , n89196 , n411726 , n411727 , n89199 , n411729 , n411730 , n411731 , n411732 , 
 n411733 , n411734 , n411735 , n411736 , n89208 , n411738 , n411739 , n89211 , n411741 , n411742 , 
 n89214 , n411744 , n411745 , n89217 , n89218 , n411748 , n89220 , n411750 , n411751 , n411752 , 
 n411753 , n411754 , n411755 , n411756 , n411757 , n89229 , n411759 , n411760 , n411761 , n89233 , 
 n411763 , n411764 , n89236 , n411766 , n411767 , n89239 , n411769 , n411770 , n89242 , n89243 , 
 n411773 , n89245 , n411775 , n411776 , n89248 , n411778 , n411779 , n411780 , n89252 , n411782 , 
 n411783 , n411784 , n411785 , n411786 , n411787 , n89259 , n411789 , n411790 , n411791 , n411792 , 
 n411793 , n411794 , n89266 , n89267 , n411797 , n89269 , n411799 , n411800 , n411801 , n411802 , 
 n89274 , n411804 , n411805 , n411806 , n411807 , n411808 , n411809 , n411810 , n411811 , n411812 , 
 n411813 , n411814 , n89286 , n411816 , n89288 , n89289 , n411819 , n411820 , n411821 , n411822 , 
 n89294 , n411824 , n411825 , n411826 , n89298 , n89299 , n411829 , n411830 , n89302 , n411832 , 
 n411833 , n89305 , n411835 , n411836 , n411837 , n89309 , n411839 , n411840 , n89312 , n411842 , 
 n411843 , n89315 , n411845 , n89317 , n411847 , n411848 , n411849 , n411850 , n411851 , n89323 , 
 n411853 , n411854 , n89326 , n411856 , n411857 , n411858 , n411859 , n411860 , n411861 , n89333 , 
 n411863 , n411864 , n411865 , n411866 , n89338 , n89339 , n411869 , n89341 , n411871 , n411872 , 
 n89344 , n411874 , n411875 , n89347 , n411877 , n411878 , n89350 , n89351 , n411881 , n89353 , 
 n411883 , n411884 , n89356 , n411886 , n411887 , n411888 , n411889 , n89361 , n89362 , n411892 , 
 n411893 , n411894 , n411895 , n411896 , n89368 , n411898 , n89370 , n89371 , n411901 , n411902 , 
 n411903 , n411904 , n411905 , n89377 , n411907 , n411908 , n411909 , n89381 , n411911 , n411912 , 
 n411913 , n411914 , n411915 , n89387 , n411917 , n411918 , n89390 , n411920 , n411921 , n411922 , 
 n89394 , n411924 , n411925 , n411926 , n89398 , n411928 , n411929 , n89401 , n89402 , n411932 , 
 n411933 , n411934 , n411935 , n411936 , n411937 , n411938 , n411939 , n89411 , n411941 , n411942 , 
 n89414 , n411944 , n411945 , n89417 , n411947 , n411948 , n411949 , n411950 , n411951 , n411952 , 
 n89424 , n411954 , n411955 , n89427 , n411957 , n411958 , n89430 , n411960 , n411961 , n89433 , 
 n411963 , n411964 , n411965 , n411966 , n411967 , n411968 , n89440 , n411970 , n411971 , n411972 , 
 n89444 , n411974 , n411975 , n411976 , n89448 , n411978 , n411979 , n89451 , n89452 , n89453 , 
 n89454 , n89455 , n89456 , n411986 , n89458 , n89459 , n89460 , n89461 , n411991 , n89463 , 
 n89464 , n411994 , n411995 , n411996 , n411997 , n89469 , n411999 , n412000 , n89472 , n89473 , 
 n412003 , n412004 , n412005 , n412006 , n412007 , n412008 , n89480 , n412010 , n412011 , n412012 , 
 n412013 , n412014 , n412015 , n412016 , n412017 , n412018 , n412019 , n412020 , n89492 , n412022 , 
 n412023 , n89495 , n89496 , n412026 , n89498 , n412028 , n412029 , n412030 , n89502 , n412032 , 
 n89504 , n412034 , n412035 , n412036 , n89505 , n89506 , n412039 , n412040 , n89509 , n412042 , 
 n412043 , n412044 , n412045 , n89514 , n412047 , n412048 , n89517 , n412050 , n412051 , n412052 , 
 n412053 , n412054 , n89523 , n89524 , n412057 , n412058 , n412059 , n412060 , n412061 , n89530 , 
 n412063 , n412064 , n89533 , n412066 , n412067 , n412068 , n412069 , n412070 , n412071 , n412072 , 
 n412073 , n89542 , n412075 , n412076 , n89545 , n412078 , n89547 , n412080 , n412081 , n412082 , 
 n412083 , n89552 , n412085 , n412086 , n412087 , n412088 , n412089 , n412090 , n412091 , n89560 , 
 n412093 , n412094 , n412095 , n89564 , n412097 , n412098 , n412099 , n412100 , n412101 , n412102 , 
 n412103 , n412104 , n412105 , n412106 , n412107 , n412108 , n412109 , n89578 , n412111 , n412112 , 
 n412113 , n412114 , n412115 , n412116 , n89585 , n412118 , n412119 , n89588 , n89589 , n412122 , 
 n412123 , n412124 , n412125 , n412126 , n412127 , n412128 , n412129 , n412130 , n412131 , n412132 , 
 n412133 , n412134 , n89603 , n89604 , n89605 , n412138 , n89607 , n412140 , n412141 , n412142 , 
 n89611 , n89612 , n89613 , n412146 , n412147 , n412148 , n89617 , n89618 , n412151 , n89620 , 
 n412153 , n412154 , n89623 , n89624 , n412157 , n412158 , n412159 , n412160 , n412161 , n412162 , 
 n412163 , n412164 , n89633 , n89634 , n412167 , n412168 , n89637 , n412170 , n412171 , n412172 , 
 n412173 , n412174 , n412175 , n89644 , n89645 , n89646 , n412179 , n412180 , n412181 , n89650 , 
 n89651 , n412184 , n412185 , n412186 , n89655 , n89656 , n412189 , n412190 , n89659 , n89660 , 
 n89661 , n412194 , n412195 , n412196 , n412197 , n89666 , n412199 , n412200 , n89669 , n412202 , 
 n412203 , n412204 , n412205 , n89674 , n412207 , n412208 , n412209 , n412210 , n89679 , n412212 , 
 n412213 , n412214 , n412215 , n412216 , n89685 , n412218 , n412219 , n89688 , n412221 , n412222 , 
 n412223 , n412224 , n412225 , n412226 , n89695 , n89696 , n412229 , n412230 , n89699 , n412232 , 
 n412233 , n89702 , n412235 , n412236 , n412237 , n412238 , n412239 , n412240 , n89709 , n412242 , 
 n412243 , n412244 , n412245 , n412246 , n89715 , n89716 , n412249 , n412250 , n412251 , n89720 , 
 n89721 , n412254 , n412255 , n412256 , n412257 , n412258 , n89727 , n412260 , n89729 , n412262 , 
 n89731 , n412264 , n412265 , n89734 , n412267 , n412268 , n412269 , n89738 , n89739 , n412272 , 
 n89741 , n412274 , n412275 , n89744 , n412277 , n89746 , n412279 , n412280 , n412281 , n89750 , 
 n412283 , n412284 , n89753 , n412286 , n412287 , n412288 , n89757 , n412290 , n412291 , n412292 , 
 n412293 , n412294 , n412295 , n89764 , n89765 , n412298 , n412299 , n89768 , n412301 , n412302 , 
 n412303 , n89772 , n412305 , n412306 , n412307 , n412308 , n412309 , n412310 , n412311 , n412312 , 
 n412313 , n89782 , n412315 , n89784 , n89785 , n412318 , n412319 , n412320 , n412321 , n412322 , 
 n89791 , n412324 , n412325 , n412326 , n412327 , n412328 , n89797 , n89798 , n412331 , n412332 , 
 n89801 , n89802 , n89803 , n412336 , n412337 , n89806 , n412339 , n412340 , n412341 , n412342 , 
 n412343 , n89812 , n89813 , n412346 , n412347 , n89816 , n412349 , n412350 , n412351 , n412352 , 
 n412353 , n412354 , n89823 , n412356 , n89825 , n89826 , n412359 , n412360 , n89829 , n412362 , 
 n412363 , n412364 , n89833 , n412366 , n412367 , n89836 , n89837 , n412370 , n412371 , n412372 , 
 n89841 , n412374 , n412375 , n412376 , n89845 , n412378 , n89847 , n412380 , n412381 , n89850 , 
 n412383 , n412384 , n89853 , n412386 , n412387 , n89856 , n412389 , n412390 , n89859 , n89860 , 
 n89861 , n412394 , n412395 , n89864 , n89865 , n412398 , n412399 , n412400 , n412401 , n89870 , 
 n412403 , n412404 , n89873 , n89874 , n89875 , n412408 , n412409 , n412410 , n89879 , n412412 , 
 n412413 , n412414 , n89883 , n412416 , n89885 , n412418 , n412419 , n89888 , n89889 , n89890 , 
 n412423 , n412424 , n412425 , n89894 , n412427 , n412428 , n412429 , n412430 , n412431 , n412432 , 
 n89901 , n412434 , n412435 , n89904 , n412437 , n412438 , n89907 , n412440 , n89909 , n412442 , 
 n89911 , n412444 , n89913 , n412446 , n89915 , n89916 , n412449 , n412450 , n89919 , n412452 , 
 n412453 , n412454 , n412455 , n412456 , n412457 , n89926 , n412459 , n412460 , n89929 , n412462 , 
 n412463 , n89932 , n412465 , n412466 , n412467 , n89936 , n412469 , n89938 , n89939 , n412472 , 
 n412473 , n412474 , n412475 , n412476 , n412477 , n412478 , n412479 , n412480 , n89943 , n89944 , 
 n412483 , n412484 , n89947 , n412486 , n412487 , n412488 , n89951 , n412490 , n412491 , n412492 , 
 n412493 , n412494 , n412495 , n89958 , n412497 , n412498 , n412499 , n89962 , n412501 , n412502 , 
 n89965 , n412504 , n412505 , n412506 , n89969 , n412508 , n412509 , n412510 , n412511 , n412512 , 
 n412513 , n412514 , n412515 , n412516 , n412517 , n89980 , n89981 , n412520 , n89983 , n412522 , 
 n412523 , n412524 , n89987 , n89988 , n412527 , n89990 , n412529 , n412530 , n412531 , n89994 , 
 n89995 , n412534 , n412535 , n89998 , n412537 , n412538 , n90001 , n412540 , n412541 , n90004 , 
 n412543 , n412544 , n412545 , n412546 , n90009 , n412548 , n412549 , n90012 , n412551 , n412552 , 
 n412553 , n412554 , n412555 , n412556 , n412557 , n412558 , n412559 , n412560 , n90023 , n412562 , 
 n412563 , n412564 , n412565 , n412566 , n412567 , n412568 , n412569 , n412570 , n412571 , n412572 , 
 n412573 , n412574 , n412575 , n90038 , n412577 , n412578 , n412579 , n412580 , n412581 , n412582 , 
 n412583 , n90046 , n412585 , n412586 , n412587 , n412588 , n412589 , n412590 , n412591 , n412592 , 
 n412593 , n412594 , n90057 , n412596 , n90059 , n90060 , n412599 , n412600 , n90063 , n412602 , 
 n412603 , n412604 , n412605 , n412606 , n90069 , n412608 , n412609 , n90072 , n412611 , n412612 , 
 n90075 , n412614 , n412615 , n412616 , n412617 , n412618 , n90081 , n412620 , n90083 , n412622 , 
 n412623 , n412624 , n412625 , n90088 , n412627 , n412628 , n90091 , n90092 , n412631 , n90094 , 
 n412633 , n412634 , n90097 , n412636 , n412637 , n412638 , n412639 , n412640 , n412641 , n412642 , 
 n412643 , n90106 , n412645 , n90108 , n90109 , n412648 , n412649 , n90112 , n90113 , n412652 , 
 n90115 , n412654 , n412655 , n90118 , n90119 , n412658 , n412659 , n412660 , n412661 , n90124 , 
 n412663 , n412664 , n412665 , n412666 , n412667 , n412668 , n412669 , n412670 , n412671 , n412672 , 
 n412673 , n412674 , n90137 , n412676 , n412677 , n90140 , n412679 , n412680 , n412681 , n412682 , 
 n412683 , n412684 , n90147 , n412686 , n412687 , n412688 , n412689 , n412690 , n412691 , n412692 , 
 n90155 , n412694 , n90157 , n412696 , n412697 , n412698 , n90161 , n412700 , n90163 , n412702 , 
 n412703 , n412704 , n412705 , n412706 , n412707 , n90170 , n412709 , n412710 , n90173 , n412712 , 
 n412713 , n90176 , n412715 , n412716 , n90179 , n412718 , n412719 , n412720 , n412721 , n412722 , 
 n412723 , n412724 , n90187 , n412726 , n412727 , n90190 , n412729 , n412730 , n412731 , n90194 , 
 n90195 , n412734 , n412735 , n412736 , n412737 , n412738 , n412739 , n412740 , n412741 , n412742 , 
 n412743 , n412744 , n412745 , n412746 , n412747 , n412748 , n412749 , n412750 , n412751 , n412752 , 
 n412753 , n90216 , n412755 , n412756 , n90219 , n412758 , n412759 , n412760 , n90223 , n412762 , 
 n412763 , n412764 , n412765 , n412766 , n412767 , n412768 , n412769 , n412770 , n412771 , n90234 , 
 n412773 , n412774 , n90237 , n412776 , n412777 , n412778 , n412779 , n412780 , n412781 , n412782 , 
 n412783 , n412784 , n412785 , n90245 , n412787 , n412788 , n412789 , n90249 , n412791 , n412792 , 
 n412793 , n90253 , n412795 , n412796 , n90256 , n412798 , n412799 , n412800 , n412801 , n90261 , 
 n412803 , n412804 , n412805 , n90265 , n412807 , n412808 , n90268 , n412810 , n90270 , n412812 , 
 n412813 , n412814 , n412815 , n90275 , n412817 , n412818 , n90278 , n412820 , n412821 , n90281 , 
 n412823 , n412824 , n90284 , n90285 , n412827 , n412828 , n412829 , n412830 , n412831 , n412832 , 
 n412833 , n412834 , n90294 , n412836 , n412837 , n412838 , n412839 , n412840 , n412841 , n412842 , 
 n412843 , n412844 , n412845 , n412846 , n90306 , n412848 , n412849 , n90309 , n412851 , n412852 , 
 n412853 , n90313 , n412855 , n412856 , n412857 , n90317 , n412859 , n412860 , n90320 , n90321 , 
 n90322 , n412864 , n412865 , n412866 , n412867 , n90327 , n412869 , n412870 , n90330 , n90331 , 
 n412873 , n412874 , n412875 , n412876 , n412877 , n412878 , n90338 , n412880 , n412881 , n412882 , 
 n412883 , n412884 , n412885 , n412886 , n90346 , n412888 , n412889 , n90349 , n412891 , n412892 , 
 n412893 , n90353 , n412895 , n412896 , n90356 , n90357 , n412899 , n412900 , n90360 , n412902 , 
 n90362 , n90363 , n412905 , n412906 , n412907 , n90367 , n90368 , n412910 , n90370 , n90371 , 
 n412913 , n412914 , n90374 , n412916 , n412917 , n412918 , n90378 , n412920 , n412921 , n90381 , 
 n412923 , n412924 , n412925 , n90385 , n412927 , n412928 , n412929 , n412930 , n412931 , n412932 , 
 n90392 , n90393 , n90394 , n90395 , n90396 , n412938 , n412939 , n412940 , n412941 , n412942 , 
 n412943 , n412944 , n412945 , n412946 , n412947 , n412948 , n90408 , n412950 , n90410 , n412952 , 
 n412953 , n90413 , n412955 , n412956 , n412957 , n412958 , n90418 , n412960 , n412961 , n412962 , 
 n90422 , n90423 , n412965 , n412966 , n90426 , n412968 , n412969 , n90429 , n412971 , n412972 , 
 n90432 , n90433 , n90434 , n90435 , n90436 , n90437 , n90438 , n90439 , n412981 , n90441 , 
 n412983 , n90443 , n90444 , n412986 , n412987 , n412988 , n412989 , n412990 , n90450 , n412992 , 
 n90452 , n90453 , n90454 , n412996 , n412997 , n412998 , n412999 , n413000 , n90460 , n413002 , 
 n90462 , n413004 , n413005 , n413006 , n413007 , n413008 , n413009 , n413010 , n413011 , n413012 , 
 n413013 , n413014 , n413015 , n413016 , n413017 , n413018 , n413019 , n413020 , n413021 , n413022 , 
 n413023 , n90483 , n413025 , n413026 , n90486 , n413028 , n90488 , n413030 , n413031 , n90491 , 
 n413033 , n413034 , n413035 , n413036 , n413037 , n90497 , n90498 , n413040 , n413041 , n413042 , 
 n413043 , n413044 , n90504 , n413046 , n413047 , n90507 , n413049 , n413050 , n90510 , n413052 , 
 n413053 , n413054 , n413055 , n90515 , n90516 , n90517 , n413059 , n413060 , n413061 , n413062 , 
 n90522 , n413064 , n413065 , n90525 , n90526 , n90527 , n413069 , n413070 , n413071 , n90531 , 
 n90532 , n413074 , n413075 , n90535 , n413077 , n413078 , n413079 , n90539 , n413081 , n90541 , 
 n413083 , n413084 , n90544 , n90545 , n413087 , n90547 , n413089 , n90549 , n90550 , n413092 , 
 n413093 , n90553 , n90554 , n413096 , n413097 , n90557 , n413099 , n90559 , n413101 , n90561 , 
 n413103 , n90563 , n90564 , n413106 , n90566 , n413108 , n413109 , n90569 , n413111 , n413112 , 
 n413113 , n413114 , n413115 , n413116 , n413117 , n413118 , n413119 , n413120 , n413121 , n413122 , 
 n413123 , n413124 , n413125 , n90585 , n413127 , n413128 , n413129 , n413130 , n413131 , n413132 , 
 n413133 , n90593 , n413135 , n413136 , n413137 , n413138 , n413139 , n413140 , n413141 , n90601 , 
 n413143 , n90603 , n413145 , n413146 , n90606 , n413148 , n413149 , n90609 , n413151 , n413152 , 
 n90612 , n413154 , n413155 , n90615 , n413157 , n413158 , n90618 , n413160 , n413161 , n413162 , 
 n413163 , n413164 , n90624 , n413166 , n413167 , n90627 , n413169 , n90629 , n90630 , n90631 , 
 n90632 , n90633 , n90634 , n90635 , n90636 , n90637 , n90638 , n90639 , n90640 , n413182 , 
 n413183 , n413184 , n413185 , n413186 , n413187 , n413188 , n413189 , n90649 , n413191 , n90651 , 
 n413193 , n413194 , n413195 , n90655 , n413197 , n413198 , n90658 , n90659 , n90660 , n90661 , 
 n90662 , n90663 , n90664 , n90665 , n90666 , n90667 , n413209 , n90669 , n413211 , n413212 , 
 n90672 , n90673 , n90674 , n90675 , n413217 , n90677 , n90678 , n413220 , n413221 , n413222 , 
 n90682 , n413224 , n413225 , n90685 , n413227 , n413228 , n90688 , n413230 , n413231 , n90691 , 
 n413233 , n90693 , n413235 , n413236 , n90696 , n413238 , n413239 , n413240 , n90700 , n90701 , 
 n413243 , n413244 , n90704 , n413246 , n413247 , n90707 , n413249 , n413250 , n413251 , n413252 , 
 n413253 , n413254 , n413255 , n413256 , n413257 , n90717 , n413259 , n413260 , n413261 , n413262 , 
 n413263 , n413264 , n413265 , n413266 , n413267 , n413268 , n413269 , n413270 , n90730 , n90731 , 
 n413273 , n413274 , n90734 , n413276 , n413277 , n413278 , n413279 , n413280 , n90740 , n413282 , 
 n90742 , n90743 , n90744 , n90745 , n90746 , n413288 , n90748 , n413290 , n413291 , n413292 , 
 n90752 , n413294 , n90754 , n413296 , n413297 , n413298 , n413299 , n413300 , n413301 , n413302 , 
 n413303 , n413304 , n413305 , n413306 , n413307 , n413308 , n413309 , n90769 , n413311 , n90771 , 
 n413313 , n90773 , n90774 , n413316 , n413317 , n90777 , n90778 , n90779 , n413321 , n413322 , 
 n413323 , n90783 , n413325 , n413326 , n413327 , n90787 , n90788 , n413330 , n413331 , n90791 , 
 n413333 , n413334 , n413335 , n413336 , n90796 , n413338 , n413339 , n413340 , n413341 , n413342 , 
 n413343 , n90803 , n413345 , n413346 , n90806 , n90807 , n90808 , n90809 , n90810 , n413352 , 
 n90812 , n413354 , n413355 , n90815 , n413357 , n90817 , n413359 , n413360 , n413361 , n413362 , 
 n413363 , n413364 , n413365 , n413366 , n90826 , n413368 , n413369 , n413370 , n90830 , n413372 , 
 n413373 , n90833 , n413375 , n90835 , n90836 , n413378 , n413379 , n90839 , n413381 , n90841 , 
 n90842 , n413384 , n413385 , n90845 , n413387 , n413388 , n413389 , n413390 , n413391 , n413392 , 
 n413393 , n413394 , n413395 , n413396 , n90856 , n413398 , n413399 , n413400 , n413401 , n90861 , 
 n413403 , n413404 , n90864 , n413406 , n413407 , n90867 , n413409 , n413410 , n413411 , n413412 , 
 n413413 , n413414 , n413415 , n90875 , n413417 , n413418 , n413419 , n413420 , n413421 , n413422 , 
 n90882 , n413424 , n413425 , n413426 , n90886 , n413428 , n413429 , n413430 , n413431 , n413432 , 
 n413433 , n413434 , n413435 , n90895 , n413437 , n413438 , n90898 , n413440 , n90900 , n90901 , 
 n90902 , n413444 , n90904 , n413446 , n90906 , n413448 , n413449 , n413450 , n413451 , n413452 , 
 n413453 , n413454 , n413455 , n90915 , n413457 , n413458 , n90918 , n413460 , n90920 , n90921 , 
 n413463 , n413464 , n90924 , n413466 , n413467 , n90927 , n413469 , n90929 , n413471 , n90931 , 
 n413473 , n90933 , n413475 , n90935 , n413477 , n413478 , n413479 , n90939 , n90940 , n413482 , 
 n90942 , n413484 , n413485 , n413486 , n90946 , n413488 , n413489 , n90949 , n90950 , n413492 , 
 n413493 , n413494 , n413495 , n413496 , n90956 , n413498 , n90958 , n413500 , n413501 , n90961 , 
 n413503 , n413504 , n413505 , n413506 , n413507 , n90967 , n413509 , n413510 , n90970 , n413512 , 
 n413513 , n413514 , n413515 , n413516 , n413517 , n413518 , n413519 , n413520 , n413521 , n413522 , 
 n413523 , n413524 , n413525 , n413526 , n413527 , n413528 , n413529 , n413530 , n413531 , n413532 , 
 n413533 , n90985 , n413535 , n413536 , n413537 , n413538 , n413539 , n413540 , n413541 , n413542 , 
 n413543 , n413544 , n413545 , n413546 , n413547 , n413548 , n413549 , n413550 , n413551 , n91003 , 
 n413553 , n91005 , n91006 , n413556 , n413557 , n91009 , n413559 , n413560 , n91012 , n413562 , 
 n91014 , n91015 , n91016 , n413566 , n91018 , n413568 , n413569 , n413570 , n413571 , n91023 , 
 n413573 , n413574 , n91026 , n91027 , n413577 , n413578 , n91030 , n91031 , n413581 , n413582 , 
 n413583 , n413584 , n413585 , n413586 , n413587 , n413588 , n413589 , n91041 , n413591 , n413592 , 
 n413593 , n413594 , n91046 , n413596 , n413597 , n91049 , n413599 , n91051 , n413601 , n413602 , 
 n91054 , n413604 , n413605 , n413606 , n413607 , n91059 , n413609 , n413610 , n413611 , n413612 , 
 n413613 , n413614 , n91066 , n413616 , n91068 , n413618 , n413619 , n91071 , n413621 , n91073 , 
 n413623 , n91075 , n413625 , n413626 , n91078 , n91079 , n91080 , n91081 , n413631 , n413632 , 
 n413633 , n413634 , n413635 , n413636 , n413637 , n413638 , n413639 , n413640 , n413641 , n413642 , 
 n91094 , n413644 , n413645 , n413646 , n413647 , n91099 , n413649 , n413650 , n91102 , n413652 , 
 n413653 , n91105 , n413655 , n413656 , n413657 , n413658 , n413659 , n413660 , n413661 , n413662 , 
 n413663 , n413664 , n91116 , n413666 , n413667 , n413668 , n91120 , n91121 , n91122 , n413672 , 
 n91124 , n91125 , n413675 , n91127 , n413677 , n91129 , n91130 , n413680 , n413681 , n413682 , 
 n413683 , n413684 , n91136 , n413686 , n91138 , n413688 , n413689 , n413690 , n91142 , n413692 , 
 n413693 , n413694 , n413695 , n413696 , n413697 , n413698 , n413699 , n91151 , n91152 , n413702 , 
 n91154 , n413704 , n91156 , n91157 , n91158 , n413708 , n91160 , n91161 , n91162 , n91163 , 
 n91164 , n91165 , n413715 , n413716 , n413717 , n413718 , n413719 , n413720 , n413721 , n91173 , 
 n91174 , n413724 , n91176 , n413726 , n413727 , n91179 , n413729 , n413730 , n413731 , n413732 , 
 n413733 , n413734 , n413735 , n413736 , n413737 , n91189 , n413739 , n413740 , n413741 , n413742 , 
 n413743 , n91195 , n413745 , n413746 , n413747 , n413748 , n413749 , n413750 , n413751 , n91203 , 
 n413753 , n91205 , n413755 , n413756 , n413757 , n413758 , n413759 , n413760 , n413761 , n413762 , 
 n413763 , n413764 , n413765 , n413766 , n413767 , n413768 , n413769 , n413770 , n413771 , n413772 , 
 n413773 , n413774 , n91226 , n413776 , n413777 , n91229 , n413779 , n413780 , n91232 , n413782 , 
 n413783 , n91235 , n413785 , n413786 , n413787 , n91239 , n91240 , n91241 , n413791 , n413792 , 
 n413793 , n413794 , n413795 , n413796 , n413797 , n413798 , n413799 , n91251 , n91252 , n91253 , 
 n413803 , n91255 , n91256 , n413806 , n91258 , n413808 , n413809 , n413810 , n91262 , n91263 , 
 n413813 , n91265 , n413815 , n413816 , n413817 , n413818 , n91270 , n413820 , n91272 , n91273 , 
 n413823 , n91275 , n413825 , n91277 , n413827 , n413828 , n413829 , n413830 , n413831 , n413832 , 
 n413833 , n413834 , n413835 , n413836 , n413837 , n413838 , n413839 , n91291 , n413841 , n413842 , 
 n413843 , n91295 , n91296 , n413846 , n413847 , n91299 , n91300 , n413850 , n91302 , n413852 , 
 n91304 , n413854 , n91306 , n413856 , n91308 , n91309 , n91310 , n413860 , n91312 , n413862 , 
 n91314 , n413864 , n413865 , n91317 , n413867 , n413868 , n91320 , n413870 , n91322 , n413872 , 
 n413873 , n413874 , n413875 , n413876 , n91328 , n413878 , n91330 , n413880 , n413881 , n413882 , 
 n413883 , n413884 , n413885 , n91337 , n91338 , n413888 , n91340 , n413890 , n91342 , n91343 , 
 n413893 , n91345 , n413895 , n413896 , n413897 , n413898 , n413899 , n413900 , n91352 , n91353 , 
 n91354 , n413904 , n413905 , n413906 , n413907 , n413908 , n91360 , n413910 , n91362 , n413912 , 
 n91364 , n91365 , n413915 , n413916 , n413917 , n413918 , n413919 , n413920 , n413921 , n413922 , 
 n413923 , n413924 , n413925 , n413926 , n413927 , n413928 , n91380 , n413930 , n413931 , n413932 , 
 n413933 , n413934 , n413935 , n413936 , n413937 , n413938 , n413939 , n413940 , n91392 , n413942 , 
 n413943 , n413944 , n413945 , n91397 , n413947 , n413948 , n413949 , n91401 , n413951 , n413952 , 
 n91404 , n413954 , n413955 , n413956 , n413957 , n413958 , n413959 , n413960 , n413961 , n413962 , 
 n413963 , n413964 , n413965 , n91417 , n413967 , n413968 , n91420 , n413970 , n413971 , n91423 , 
 n91424 , n91425 , n91426 , n91427 , n413977 , n91429 , n91430 , n413980 , n413981 , n91433 , 
 n413983 , n413984 , n413985 , n413986 , n413987 , n413988 , n413989 , n91441 , n413991 , n91443 , 
 n91444 , n413994 , n413995 , n91447 , n413997 , n413998 , n91450 , n414000 , n414001 , n414002 , 
 n91454 , n414004 , n91456 , n414006 , n414007 , n414008 , n414009 , n414010 , n414011 , n91463 , 
 n414013 , n414014 , n414015 , n414016 , n414017 , n91469 , n414019 , n414020 , n414021 , n91473 , 
 n414023 , n414024 , n414025 , n414026 , n414027 , n414028 , n414029 , n414030 , n414031 , n414032 , 
 n414033 , n414034 , n414035 , n414036 , n414037 , n414038 , n414039 , n91491 , n91492 , n414042 , 
 n91494 , n414044 , n414045 , n91497 , n414047 , n414048 , n414049 , n91501 , n91502 , n91503 , 
 n91504 , n414054 , n91506 , n414056 , n414057 , n414058 , n414059 , n414060 , n91512 , n414062 , 
 n414063 , n91515 , n414065 , n414066 , n91518 , n91519 , n91520 , n414070 , n414071 , n91523 , 
 n414073 , n414074 , n414075 , n91527 , n91528 , n414078 , n414079 , n414080 , n414081 , n414082 , 
 n414083 , n414084 , n414085 , n414086 , n414087 , n91539 , n414089 , n91541 , n91542 , n91543 , 
 n91544 , n91545 , n91546 , n91547 , n414097 , n414098 , n91550 , n414100 , n414101 , n91553 , 
 n414103 , n414104 , n414105 , n91557 , n414107 , n414108 , n414109 , n414110 , n414111 , n414112 , 
 n414113 , n414114 , n414115 , n414116 , n91566 , n414118 , n414119 , n414120 , n414121 , n414122 , 
 n414123 , n414124 , n414125 , n91575 , n414127 , n91577 , n414129 , n414130 , n414131 , n414132 , 
 n414133 , n414134 , n414135 , n414136 , n414137 , n414138 , n414139 , n414140 , n414141 , n91591 , 
 n414143 , n414144 , n414145 , n414146 , n414147 , n91597 , n414149 , n414150 , n414151 , n91601 , 
 n414153 , n414154 , n91604 , n414156 , n414157 , n91607 , n91608 , n414160 , n91610 , n414162 , 
 n91612 , n414164 , n414165 , n91615 , n414167 , n91617 , n91618 , n414170 , n414171 , n91621 , 
 n91622 , n414174 , n414175 , n414176 , n414177 , n91627 , n414179 , n91629 , n91630 , n414182 , 
 n91632 , n91633 , n91634 , n414186 , n414187 , n91637 , n91638 , n91639 , n91640 , n414192 , 
 n91642 , n414194 , n91644 , n414196 , n414197 , n414198 , n91648 , n414200 , n414201 , n91651 , 
 n414203 , n91653 , n91654 , n91655 , n414207 , n414208 , n91658 , n414210 , n414211 , n91661 , 
 n414213 , n414214 , n91664 , n91665 , n91666 , n414218 , n414219 , n414220 , n414221 , n414222 , 
 n414223 , n91673 , n414225 , n414226 , n91676 , n414228 , n414229 , n414230 , n414231 , n91681 , 
 n91682 , n91683 , n414235 , n91685 , n91686 , n414238 , n91688 , n414240 , n91690 , n91691 , 
 n91692 , n91693 , n414245 , n414246 , n91696 , n414248 , n91698 , n91699 , n91700 , n91701 , 
 n414253 , n414254 , n414255 , n414256 , n414257 , n91707 , n414259 , n414260 , n414261 , n414262 , 
 n414263 , n91713 , n414265 , n414266 , n91716 , n414268 , n414269 , n91719 , n414271 , n414272 , 
 n91722 , n414274 , n414275 , n91725 , n414277 , n91727 , n414279 , n414280 , n414281 , n414282 , 
 n414283 , n414284 , n414285 , n414286 , n414287 , n414288 , n91738 , n414290 , n91740 , n414292 , 
 n414293 , n414294 , n414295 , n414296 , n414297 , n414298 , n414299 , n414300 , n414301 , n91751 , 
 n414303 , n414304 , n414305 , n91755 , n414307 , n414308 , n414309 , n414310 , n414311 , n414312 , 
 n91762 , n414314 , n414315 , n91765 , n414317 , n414318 , n414319 , n91769 , n414321 , n91771 , 
 n414323 , n414324 , n91774 , n414326 , n414327 , n91777 , n414329 , n91779 , n414331 , n414332 , 
 n91782 , n414334 , n414335 , n91785 , n414337 , n414338 , n91788 , n414340 , n414341 , n414342 , 
 n91792 , n414344 , n91794 , n414346 , n414347 , n91797 , n414349 , n91799 , n91800 , n91801 , 
 n91802 , n91803 , n414355 , n414356 , n414357 , n91807 , n414359 , n414360 , n91810 , n414362 , 
 n414363 , n414364 , n414365 , n91815 , n414367 , n414368 , n91818 , n91819 , n414371 , n91821 , 
 n414373 , n91823 , n91824 , n414376 , n414377 , n414378 , n414379 , n414380 , n414381 , n414382 , 
 n414383 , n414384 , n414385 , n414386 , n414387 , n414388 , n414389 , n414390 , n414391 , n91841 , 
 n414393 , n414394 , n414395 , n91845 , n414397 , n414398 , n91848 , n414400 , n414401 , n414402 , 
 n414403 , n414404 , n91854 , n414406 , n91856 , n414408 , n414409 , n414410 , n91860 , n414412 , 
 n414413 , n91863 , n414415 , n414416 , n414417 , n91867 , n414419 , n414420 , n91870 , n414422 , 
 n414423 , n91873 , n414425 , n414426 , n414427 , n414428 , n414429 , n414430 , n91880 , n414432 , 
 n414433 , n414434 , n414435 , n91885 , n414437 , n414438 , n91888 , n414440 , n414441 , n414442 , 
 n414443 , n414444 , n414445 , n414446 , n91891 , n414448 , n414449 , n91894 , n414451 , n414452 , 
 n414453 , n414454 , n91899 , n414456 , n414457 , n414458 , n414459 , n414460 , n414461 , n414462 , 
 n414463 , n414464 , n414465 , n414466 , n91911 , n414468 , n414469 , n414470 , n414471 , n414472 , 
 n414473 , n91918 , n414475 , n414476 , n414477 , n414478 , n91923 , n91924 , n91925 , n414482 , 
 n91927 , n91928 , n414485 , n91930 , n91931 , n414488 , n91933 , n91934 , n91935 , n414492 , 
 n414493 , n91938 , n91939 , n91940 , n414497 , n91942 , n91943 , n414500 , n414501 , n91946 , 
 n414503 , n91948 , n414505 , n414506 , n414507 , n414508 , n414509 , n414510 , n414511 , n414512 , 
 n414513 , n414514 , n414515 , n91960 , n414517 , n414518 , n414519 , n91964 , n91965 , n414522 , 
 n414523 , n414524 , n414525 , n414526 , n414527 , n414528 , n91973 , n414530 , n91975 , n91976 , 
 n91977 , n91978 , n414535 , n414536 , n414537 , n414538 , n414539 , n414540 , n91985 , n414542 , 
 n414543 , n414544 , n414545 , n414546 , n414547 , n91992 , n414549 , n414550 , n414551 , n414552 , 
 n414553 , n414554 , n414555 , n414556 , n414557 , n414558 , n92003 , n414560 , n414561 , n92006 , 
 n414563 , n414564 , n92009 , n414566 , n414567 , n414568 , n414569 , n414570 , n92015 , n92016 , 
 n414573 , n92018 , n414575 , n92020 , n414577 , n414578 , n92023 , n414580 , n414581 , n414582 , 
 n414583 , n92028 , n414585 , n92030 , n414587 , n92032 , n92033 , n414590 , n414591 , n92036 , 
 n414593 , n414594 , n92039 , n414596 , n414597 , n92042 , n92043 , n92044 , n414601 , n92046 , 
 n414603 , n414604 , n92049 , n414606 , n414607 , n92052 , n414609 , n414610 , n414611 , n414612 , 
 n414613 , n92058 , n414615 , n414616 , n92061 , n414618 , n414619 , n414620 , n414621 , n414622 , 
 n92067 , n414624 , n414625 , n414626 , n414627 , n414628 , n414629 , n414630 , n414631 , n92076 , 
 n414633 , n92078 , n414635 , n414636 , n92081 , n414638 , n414639 , n414640 , n92085 , n414642 , 
 n414643 , n414644 , n414645 , n414646 , n414647 , n414648 , n414649 , n92094 , n92095 , n414652 , 
 n414653 , n414654 , n414655 , n414656 , n414657 , n414658 , n92103 , n414660 , n414661 , n92106 , 
 n414663 , n414664 , n92109 , n414666 , n414667 , n92112 , n414669 , n414670 , n414671 , n414672 , 
 n414673 , n414674 , n92119 , n92120 , n414677 , n414678 , n414679 , n414680 , n414681 , n92126 , 
 n414683 , n414684 , n414685 , n414686 , n414687 , n92132 , n92133 , n414690 , n414691 , n414692 , 
 n414693 , n92138 , n414695 , n414696 , n414697 , n414698 , n92143 , n414700 , n414701 , n92146 , 
 n92147 , n414704 , n414705 , n414706 , n92151 , n414708 , n414709 , n92154 , n414711 , n414712 , 
 n414713 , n414714 , n92159 , n92160 , n414717 , n414718 , n414719 , n92164 , n92165 , n414722 , 
 n414723 , n414724 , n92169 , n414726 , n414727 , n92172 , n414729 , n92174 , n414731 , n92176 , 
 n414733 , n92178 , n92179 , n92180 , n414737 , n414738 , n414739 , n414740 , n92185 , n414742 , 
 n414743 , n414744 , n414745 , n414746 , n414747 , n414748 , n414749 , n414750 , n414751 , n414752 , 
 n92197 , n414754 , n92199 , n92200 , n414757 , n414758 , n414759 , n414760 , n414761 , n414762 , 
 n414763 , n414764 , n92209 , n414766 , n414767 , n92212 , n414769 , n414770 , n92215 , n414772 , 
 n414773 , n414774 , n414775 , n414776 , n414777 , n414778 , n414779 , n414780 , n414781 , n92226 , 
 n92227 , n414784 , n414785 , n414786 , n414787 , n414788 , n92233 , n414790 , n414791 , n92236 , 
 n414793 , n92238 , n414795 , n92240 , n92241 , n414798 , n414799 , n414800 , n414801 , n414802 , 
 n414803 , n414804 , n414805 , n92250 , n414807 , n414808 , n92253 , n414810 , n414811 , n414812 , 
 n414813 , n414814 , n92259 , n414816 , n414817 , n414818 , n92263 , n414820 , n414821 , n414822 , 
 n414823 , n92268 , n414825 , n414826 , n92271 , n92272 , n92273 , n414830 , n414831 , n414832 , 
 n414833 , n92278 , n414835 , n92280 , n414837 , n92282 , n414839 , n92284 , n414841 , n414842 , 
 n414843 , n414844 , n414845 , n414846 , n414847 , n92292 , n414849 , n92294 , n92295 , n92296 , 
 n92297 , n92298 , n92299 , n414856 , n92301 , n414858 , n414859 , n414860 , n92305 , n414862 , 
 n92307 , n414864 , n414865 , n414866 , n92311 , n92312 , n414869 , n92314 , n414871 , n414872 , 
 n92317 , n414874 , n414875 , n414876 , n414877 , n92322 , n414879 , n414880 , n414881 , n414882 , 
 n414883 , n414884 , n414885 , n414886 , n414887 , n414888 , n414889 , n414890 , n92335 , n414892 , 
 n414893 , n92338 , n414895 , n414896 , n414897 , n414898 , n414899 , n414900 , n414901 , n414902 , 
 n414903 , n414904 , n414905 , n414906 , n92351 , n414908 , n414909 , n414910 , n92355 , n414912 , 
 n414913 , n414914 , n92359 , n414916 , n414917 , n92362 , n92363 , n414920 , n414921 , n414922 , 
 n414923 , n414924 , n414925 , n92370 , n414927 , n92372 , n414929 , n92374 , n92375 , n414932 , 
 n414933 , n414934 , n92379 , n414936 , n414937 , n92382 , n414939 , n414940 , n92385 , n414942 , 
 n414943 , n92388 , n414945 , n92390 , n414947 , n92392 , n92393 , n414950 , n92395 , n414952 , 
 n414953 , n414954 , n92399 , n414956 , n414957 , n414958 , n414959 , n414960 , n414961 , n414962 , 
 n414963 , n92408 , n414965 , n92410 , n92411 , n414968 , n414969 , n414970 , n414971 , n414972 , 
 n92417 , n92418 , n414975 , n92420 , n414977 , n414978 , n414979 , n414980 , n414981 , n414982 , 
 n414983 , n414984 , n414985 , n414986 , n92431 , n414988 , n414989 , n92434 , n414991 , n92436 , 
 n414993 , n414994 , n414995 , n414996 , n414997 , n414998 , n92443 , n415000 , n92445 , n92446 , 
 n92447 , n415004 , n92449 , n92450 , n415007 , n92452 , n415009 , n415010 , n92455 , n415012 , 
 n92457 , n92458 , n415015 , n92460 , n415017 , n415018 , n415019 , n415020 , n415021 , n415022 , 
 n415023 , n415024 , n92469 , n415026 , n415027 , n415028 , n415029 , n415030 , n92475 , n415032 , 
 n415033 , n92478 , n92479 , n415036 , n415037 , n415038 , n92483 , n415040 , n92485 , n415042 , 
 n415043 , n92488 , n415045 , n92490 , n92491 , n92492 , n415049 , n415050 , n92495 , n415052 , 
 n92497 , n415054 , n415055 , n415056 , n415057 , n92502 , n92503 , n415060 , n92505 , n415062 , 
 n415063 , n415064 , n415065 , n415066 , n415067 , n92512 , n415069 , n415070 , n92515 , n415072 , 
 n415073 , n92518 , n415075 , n92520 , n415077 , n92522 , n415079 , n415080 , n92525 , n92526 , 
 n415083 , n415084 , n415085 , n415086 , n415087 , n415088 , n92533 , n415090 , n415091 , n415092 , 
 n415093 , n415094 , n415095 , n415096 , n415097 , n415098 , n92543 , n92544 , n415101 , n415102 , 
 n92547 , n415104 , n415105 , n415106 , n92551 , n415108 , n415109 , n92554 , n415111 , n415112 , 
 n415113 , n92558 , n415115 , n415116 , n92561 , n415118 , n415119 , n92564 , n415121 , n415122 , 
 n415123 , n92568 , n415125 , n415126 , n92571 , n415128 , n415129 , n92574 , n415131 , n415132 , 
 n92577 , n415134 , n415135 , n92580 , n92581 , n415138 , n92583 , n415140 , n92585 , n415142 , 
 n415143 , n92588 , n415145 , n415146 , n92591 , n415148 , n415149 , n415150 , n415151 , n415152 , 
 n92597 , n415154 , n415155 , n415156 , n415157 , n415158 , n415159 , n415160 , n92605 , n415162 , 
 n415163 , n92608 , n415165 , n415166 , n415167 , n415168 , n92613 , n415170 , n415171 , n415172 , 
 n92617 , n92618 , n92619 , n92620 , n415177 , n415178 , n92623 , n92624 , n92625 , n92626 , 
 n92627 , n415184 , n415185 , n92630 , n415187 , n415188 , n415189 , n415190 , n415191 , n415192 , 
 n415193 , n92638 , n415195 , n415196 , n415197 , n415198 , n415199 , n415200 , n415201 , n415202 , 
 n415203 , n415204 , n92649 , n415206 , n415207 , n92652 , n415209 , n415210 , n92655 , n92656 , 
 n415213 , n92658 , n415215 , n92660 , n415217 , n415218 , n415219 , n415220 , n415221 , n415222 , 
 n92667 , n415224 , n92669 , n415226 , n415227 , n415228 , n415229 , n415230 , n415231 , n92676 , 
 n415233 , n92678 , n415235 , n415236 , n92681 , n415238 , n415239 , n92684 , n415241 , n415242 , 
 n92687 , n415244 , n415245 , n415246 , n415247 , n415248 , n415249 , n92694 , n415251 , n415252 , 
 n92697 , n92698 , n415255 , n92700 , n92701 , n415258 , n415259 , n415260 , n415261 , n415262 , 
 n415263 , n415264 , n92709 , n415266 , n92711 , n415268 , n415269 , n415270 , n92715 , n92716 , 
 n415273 , n92718 , n415275 , n415276 , n92721 , n415278 , n415279 , n92724 , n415281 , n415282 , 
 n92727 , n415284 , n415285 , n415286 , n415287 , n92732 , n415289 , n92734 , n92735 , n415292 , 
 n415293 , n92738 , n415295 , n415296 , n415297 , n92742 , n415299 , n92744 , n92745 , n415302 , 
 n415303 , n415304 , n92749 , n92750 , n415307 , n92752 , n92753 , n415310 , n415311 , n92756 , 
 n415313 , n415314 , n415315 , n92760 , n415317 , n415318 , n415319 , n415320 , n415321 , n92766 , 
 n92767 , n415324 , n92769 , n92770 , n415327 , n415328 , n415329 , n415330 , n415331 , n415332 , 
 n415333 , n415334 , n92779 , n92780 , n415337 , n92782 , n415339 , n415340 , n92785 , n415342 , 
 n415343 , n92788 , n415345 , n92790 , n415347 , n92792 , n92793 , n415350 , n415351 , n92796 , 
 n92797 , n415354 , n92799 , n92800 , n415357 , n415358 , n415359 , n415360 , n415361 , n415362 , 
 n92807 , n415364 , n415365 , n92810 , n415367 , n415368 , n415369 , n415370 , n415371 , n92816 , 
 n415373 , n415374 , n92819 , n415376 , n415377 , n92822 , n415379 , n415380 , n92825 , n415382 , 
 n92827 , n92828 , n415385 , n92830 , n415387 , n92832 , n92833 , n92834 , n415391 , n415392 , 
 n415393 , n415394 , n415395 , n415396 , n415397 , n92842 , n415399 , n92844 , n92845 , n415402 , 
 n92847 , n415404 , n92849 , n415406 , n415407 , n92852 , n415409 , n415410 , n415411 , n415412 , 
 n415413 , n92858 , n415415 , n415416 , n92861 , n415418 , n415419 , n415420 , n415421 , n92866 , 
 n415423 , n415424 , n415425 , n415426 , n92871 , n92872 , n415429 , n415430 , n415431 , n415432 , 
 n415433 , n415434 , n415435 , n92880 , n92881 , n415438 , n415439 , n415440 , n92885 , n415442 , 
 n92887 , n415444 , n415445 , n415446 , n92891 , n415448 , n415449 , n92894 , n92895 , n415452 , 
 n415453 , n415454 , n415455 , n415456 , n415457 , n92902 , n415459 , n415460 , n92905 , n92906 , 
 n415463 , n415464 , n415465 , n92910 , n92911 , n415468 , n92913 , n92914 , n415471 , n92916 , 
 n415473 , n415474 , n92919 , n415476 , n92921 , n415478 , n415479 , n415480 , n415481 , n415482 , 
 n92927 , n92928 , n415485 , n415486 , n415487 , n415488 , n92933 , n415490 , n415491 , n92936 , 
 n92937 , n415494 , n415495 , n415496 , n415497 , n415498 , n92943 , n415500 , n415501 , n415502 , 
 n92947 , n92948 , n92949 , n415506 , n415507 , n415508 , n415509 , n415510 , n415511 , n415512 , 
 n415513 , n415514 , n415515 , n415516 , n415517 , n92962 , n415519 , n415520 , n415521 , n415522 , 
 n92967 , n92968 , n92969 , n415526 , n415527 , n92972 , n415529 , n92974 , n415531 , n415532 , 
 n92977 , n415534 , n92979 , n415536 , n415537 , n92982 , n92983 , n415540 , n415541 , n415542 , 
 n415543 , n415544 , n415545 , n92990 , n415547 , n92992 , n92993 , n92994 , n92995 , n92996 , 
 n92997 , n415554 , n92999 , n415556 , n415557 , n415558 , n93003 , n415560 , n415561 , n93006 , 
 n93007 , n415564 , n93009 , n415566 , n415567 , n415568 , n415569 , n415570 , n415571 , n415572 , 
 n93017 , n415574 , n415575 , n93020 , n93021 , n93022 , n415579 , n415580 , n93025 , n415582 , 
 n415583 , n415584 , n415585 , n415586 , n93031 , n415588 , n415589 , n415590 , n93035 , n415592 , 
 n415593 , n415594 , n415595 , n415596 , n93041 , n415598 , n415599 , n93044 , n93045 , n415602 , 
 n415603 , n93048 , n415605 , n415606 , n93051 , n415608 , n415609 , n93054 , n93055 , n415612 , 
 n415613 , n415614 , n93059 , n415616 , n415617 , n415618 , n415619 , n415620 , n415621 , n415622 , 
 n415623 , n415624 , n93069 , n415626 , n415627 , n93072 , n415629 , n415630 , n93075 , n93076 , 
 n415633 , n93078 , n415635 , n415636 , n93081 , n415638 , n415639 , n415640 , n93085 , n415642 , 
 n415643 , n415644 , n415645 , n415646 , n415647 , n415648 , n415649 , n415650 , n415651 , n415652 , 
 n415653 , n93098 , n93099 , n415656 , n93101 , n415658 , n415659 , n415660 , n415661 , n415662 , 
 n93107 , n415664 , n415665 , n415666 , n415667 , n415668 , n93113 , n415670 , n415671 , n415672 , 
 n93117 , n415674 , n415675 , n415676 , n415677 , n415678 , n415679 , n415680 , n415681 , n415682 , 
 n415683 , n415684 , n93129 , n415686 , n415687 , n415688 , n415689 , n415690 , n93135 , n415692 , 
 n415693 , n93138 , n93139 , n415696 , n415697 , n415698 , n93143 , n415700 , n415701 , n415702 , 
 n415703 , n415704 , n415705 , n415706 , n415707 , n415708 , n415709 , n415710 , n415711 , n415712 , 
 n415713 , n415714 , n415715 , n93160 , n415717 , n415718 , n93163 , n415720 , n415721 , n93166 , 
 n415723 , n415724 , n93169 , n415726 , n415727 , n93172 , n93173 , n415730 , n93175 , n415732 , 
 n415733 , n415734 , n415735 , n415736 , n93181 , n93182 , n415739 , n415740 , n93185 , n93186 , 
 n93187 , n415744 , n415745 , n93190 , n415747 , n93192 , n93193 , n415750 , n93195 , n415752 , 
 n415753 , n415754 , n415755 , n415756 , n415757 , n415758 , n415759 , n415760 , n415761 , n93206 , 
 n415763 , n415764 , n415765 , n415766 , n93211 , n415768 , n415769 , n415770 , n415771 , n415772 , 
 n415773 , n93218 , n415775 , n415776 , n93221 , n93222 , n415779 , n415780 , n415781 , n415782 , 
 n93227 , n415784 , n415785 , n415786 , n415787 , n93232 , n93233 , n415790 , n415791 , n93236 , 
 n415793 , n415794 , n415795 , n415796 , n415797 , n415798 , n415799 , n93244 , n415801 , n415802 , 
 n415803 , n415804 , n415805 , n93250 , n415807 , n415808 , n93253 , n415810 , n415811 , n415812 , 
 n415813 , n415814 , n415815 , n415816 , n415817 , n415818 , n93263 , n93264 , n415821 , n415822 , 
 n415823 , n415824 , n415825 , n415826 , n93271 , n415828 , n415829 , n415830 , n415831 , n415832 , 
 n415833 , n415834 , n415835 , n415836 , n415837 , n93282 , n415839 , n415840 , n415841 , n415842 , 
 n415843 , n415844 , n415845 , n93290 , n415847 , n93292 , n93293 , n93294 , n415851 , n415852 , 
 n93297 , n415854 , n415855 , n415856 , n93301 , n415858 , n93303 , n415860 , n93305 , n93306 , 
 n93307 , n93308 , n415865 , n415866 , n93311 , n415868 , n415869 , n93314 , n93315 , n415872 , 
 n415873 , n415874 , n415875 , n415876 , n415877 , n93322 , n415879 , n93324 , n415881 , n415882 , 
 n93327 , n415884 , n415885 , n93330 , n415887 , n415888 , n93333 , n415890 , n93335 , n93336 , 
 n93337 , n93338 , n93339 , n93340 , n93341 , n93342 , n93343 , n415900 , n415901 , n415902 , 
 n415903 , n415904 , n93349 , n415906 , n93351 , n415908 , n415909 , n415910 , n93355 , n415912 , 
 n415913 , n93358 , n93359 , n415916 , n415917 , n93362 , n93363 , n93364 , n93365 , n415922 , 
 n415923 , n415924 , n415925 , n415926 , n93371 , n93372 , n415929 , n415930 , n415931 , n415932 , 
 n415933 , n93378 , n415935 , n93380 , n93381 , n415938 , n415939 , n415940 , n93385 , n415942 , 
 n93387 , n415944 , n415945 , n93390 , n93391 , n93392 , n415949 , n415950 , n415951 , n93396 , 
 n415953 , n415954 , n93399 , n415956 , n415957 , n415958 , n415959 , n93404 , n415961 , n415962 , 
 n93407 , n415964 , n415965 , n415966 , n93411 , n415968 , n415969 , n415970 , n415971 , n415972 , 
 n415973 , n415974 , n415975 , n415976 , n415977 , n93422 , n415979 , n93424 , n415981 , n415982 , 
 n93427 , n415984 , n415985 , n93430 , n415987 , n93432 , n415989 , n415990 , n415991 , n415992 , 
 n415993 , n415994 , n415995 , n415996 , n415997 , n415998 , n415999 , n416000 , n416001 , n416002 , 
 n416003 , n416004 , n416005 , n93450 , n93451 , n93452 , n416009 , n416010 , n416011 , n416012 , 
 n93457 , n416014 , n416015 , n416016 , n93461 , n93462 , n416019 , n416020 , n93465 , n416022 , 
 n416023 , n416024 , n416025 , n416026 , n416027 , n416028 , n93473 , n416030 , n416031 , n416032 , 
 n416033 , n93478 , n416035 , n93480 , n416037 , n416038 , n416039 , n416040 , n416041 , n416042 , 
 n416043 , n416044 , n416045 , n416046 , n416047 , n93492 , n93493 , n416050 , n416051 , n416052 , 
 n416053 , n416054 , n416055 , n416056 , n93501 , n93502 , n416059 , n416060 , n416061 , n93506 , 
 n416063 , n416064 , n416065 , n416066 , n416067 , n416068 , n416069 , n416070 , n416071 , n416072 , 
 n93517 , n416074 , n416075 , n93520 , n93521 , n416078 , n416079 , n93524 , n416081 , n416082 , 
 n416083 , n93528 , n416085 , n416086 , n416087 , n93532 , n93533 , n93534 , n93535 , n416092 , 
 n416093 , n416094 , n416095 , n416096 , n93541 , n416098 , n416099 , n416100 , n416101 , n416102 , 
 n416103 , n93548 , n416105 , n93550 , n416107 , n93552 , n93553 , n93554 , n93555 , n416112 , 
 n416113 , n416114 , n416115 , n93560 , n416117 , n416118 , n416119 , n93564 , n416121 , n416122 , 
 n93567 , n416124 , n416125 , n93570 , n93571 , n416128 , n93573 , n416130 , n416131 , n93576 , 
 n416133 , n416134 , n416135 , n416136 , n416137 , n416138 , n93583 , n93584 , n416141 , n416142 , 
 n93587 , n416144 , n416145 , n416146 , n93591 , n416148 , n416149 , n416150 , n93595 , n416152 , 
 n93597 , n416154 , n93599 , n416156 , n93601 , n416158 , n416159 , n93604 , n416161 , n416162 , 
 n416163 , n416164 , n416165 , n416166 , n93611 , n416168 , n416169 , n416170 , n93615 , n416172 , 
 n416173 , n416174 , n93619 , n416176 , n93621 , n416178 , n416179 , n93624 , n416181 , n93626 , 
 n416183 , n416184 , n416185 , n416186 , n416187 , n416188 , n416189 , n416190 , n416191 , n416192 , 
 n416193 , n416194 , n416195 , n416196 , n416197 , n416198 , n416199 , n93644 , n416201 , n416202 , 
 n416203 , n416204 , n416205 , n416206 , n93651 , n93652 , n416209 , n416210 , n416211 , n416212 , 
 n416213 , n93658 , n93659 , n416216 , n416217 , n416218 , n416219 , n416220 , n93665 , n416222 , 
 n416223 , n416224 , n416225 , n93670 , n93671 , n416228 , n416229 , n416230 , n416231 , n416232 , 
 n93677 , n93678 , n416235 , n93680 , n416237 , n416238 , n93683 , n416240 , n416241 , n93686 , 
 n416243 , n416244 , n416245 , n416246 , n416247 , n416248 , n93693 , n416250 , n416251 , n416252 , 
 n416253 , n416254 , n93699 , n93700 , n416257 , n416258 , n416259 , n416260 , n416261 , n416262 , 
 n93707 , n416264 , n416265 , n416266 , n416267 , n416268 , n416269 , n416270 , n93715 , n416272 , 
 n416273 , n93718 , n416275 , n93720 , n416277 , n416278 , n416279 , n93724 , n416281 , n416282 , 
 n416283 , n416284 , n416285 , n93730 , n93731 , n93732 , n416289 , n93734 , n416291 , n93736 , 
 n416293 , n416294 , n416295 , n416296 , n416297 , n416298 , n416299 , n416300 , n416301 , n416302 , 
 n416303 , n416304 , n416305 , n93750 , n416307 , n416308 , n416309 , n416310 , n416311 , n416312 , 
 n416313 , n416314 , n93759 , n416316 , n416317 , n416318 , n416319 , n416320 , n93765 , n93766 , 
 n416323 , n416324 , n416325 , n93770 , n416327 , n416328 , n416329 , n93774 , n93775 , n416332 , 
 n416333 , n416334 , n416335 , n416336 , n93781 , n93782 , n416339 , n93784 , n416341 , n93786 , 
 n93787 , n93788 , n416345 , n416346 , n93791 , n416348 , n416349 , n93794 , n416351 , n416352 , 
 n416353 , n416354 , n93799 , n416356 , n416357 , n416358 , n93803 , n416360 , n416361 , n416362 , 
 n93807 , n416364 , n416365 , n93810 , n416367 , n416368 , n416369 , n416370 , n416371 , n416372 , 
 n93817 , n416374 , n416375 , n416376 , n93821 , n93822 , n416379 , n93824 , n416381 , n93826 , 
 n416383 , n416384 , n93829 , n93830 , n416387 , n416388 , n93833 , n93834 , n93835 , n416392 , 
 n93837 , n93838 , n93839 , n416396 , n93841 , n416398 , n93843 , n93844 , n93845 , n416402 , 
 n93847 , n416404 , n416405 , n93850 , n416407 , n416408 , n93853 , n416410 , n416411 , n416412 , 
 n416413 , n93858 , n416415 , n416416 , n416417 , n93862 , n416419 , n93864 , n416421 , n93866 , 
 n93867 , n416424 , n93869 , n416426 , n416427 , n416428 , n416429 , n416430 , n416431 , n416432 , 
 n416433 , n93878 , n416435 , n416436 , n416437 , n416438 , n416439 , n93884 , n93885 , n416442 , 
 n416443 , n416444 , n93889 , n416446 , n416447 , n93892 , n416449 , n416450 , n416451 , n416452 , 
 n416453 , n416454 , n416455 , n416456 , n416457 , n416458 , n416459 , n93904 , n416461 , n93906 , 
 n416463 , n416464 , n93909 , n416466 , n416467 , n416468 , n416469 , n416470 , n416471 , n416472 , 
 n416473 , n93918 , n93919 , n416476 , n416477 , n416478 , n416479 , n416480 , n93925 , n93926 , 
 n416483 , n416484 , n93929 , n93930 , n416487 , n416488 , n93933 , n416490 , n416491 , n416492 , 
 n416493 , n416494 , n93939 , n93940 , n416497 , n416498 , n416499 , n93944 , n416501 , n416502 , 
 n416503 , n93948 , n416505 , n416506 , n416507 , n416508 , n416509 , n416510 , n416511 , n416512 , 
 n416513 , n416514 , n93959 , n416516 , n416517 , n416518 , n416519 , n416520 , n416521 , n416522 , 
 n93967 , n416524 , n416525 , n416526 , n416527 , n93972 , n416529 , n416530 , n416531 , n416532 , 
 n93977 , n416534 , n416535 , n416536 , n93981 , n93982 , n93983 , n93984 , n93985 , n416542 , 
 n93987 , n416544 , n93989 , n416546 , n416547 , n416548 , n93993 , n416550 , n416551 , n416552 , 
 n93997 , n416554 , n93999 , n94000 , n416557 , n416558 , n416559 , n416560 , n416561 , n416562 , 
 n416563 , n416564 , n416565 , n416566 , n416567 , n416568 , n416569 , n416570 , n416571 , n416572 , 
 n416573 , n416574 , n416575 , n94020 , n416577 , n416578 , n416579 , n94024 , n94025 , n94026 , 
 n416583 , n416584 , n416585 , n416586 , n416587 , n94032 , n416589 , n416590 , n416591 , n416592 , 
 n416593 , n94038 , n416595 , n416596 , n416597 , n416598 , n94043 , n416600 , n416601 , n416602 , 
 n416603 , n416604 , n416605 , n416606 , n94051 , n416608 , n94053 , n416610 , n416611 , n94056 , 
 n416613 , n416614 , n94059 , n94060 , n94061 , n416618 , n416619 , n94064 , n416621 , n416622 , 
 n94067 , n416624 , n416625 , n416626 , n416627 , n94072 , n416629 , n94074 , n416631 , n94076 , 
 n94077 , n94078 , n94079 , n416636 , n94081 , n94082 , n416639 , n416640 , n416641 , n94086 , 
 n94087 , n416644 , n416645 , n416646 , n416647 , n416648 , n416649 , n416650 , n416651 , n416652 , 
 n94097 , n416654 , n416655 , n94100 , n94101 , n416658 , n416659 , n416660 , n416661 , n94106 , 
 n416663 , n416664 , n416665 , n94110 , n416667 , n416668 , n94113 , n416670 , n416671 , n94116 , 
 n416673 , n416674 , n416675 , n416676 , n416677 , n416678 , n416679 , n416680 , n94125 , n416682 , 
 n416683 , n94128 , n416685 , n416686 , n416687 , n94132 , n94133 , n416690 , n416691 , n416692 , 
 n416693 , n416694 , n416695 , n94140 , n416697 , n416698 , n416699 , n416700 , n416701 , n94146 , 
 n416703 , n416704 , n416705 , n94150 , n416707 , n416708 , n416709 , n94154 , n94155 , n416712 , 
 n416713 , n94158 , n416715 , n416716 , n416717 , n94162 , n416719 , n416720 , n416721 , n416722 , 
 n416723 , n416724 , n416725 , n416726 , n416727 , n416728 , n416729 , n416730 , n416731 , n416732 , 
 n416733 , n416734 , n416735 , n416736 , n416737 , n416738 , n416739 , n416740 , n416741 , n416742 , 
 n416743 , n94188 , n416745 , n416746 , n94191 , n94192 , n416749 , n94194 , n416751 , n416752 , 
 n94197 , n416754 , n416755 , n94200 , n94201 , n416758 , n416759 , n94204 , n416761 , n94206 , 
 n416763 , n416764 , n94209 , n94210 , n416767 , n416768 , n416769 , n416770 , n94215 , n416772 , 
 n94217 , n416774 , n416775 , n416776 , n416777 , n416778 , n416779 , n416780 , n416781 , n94226 , 
 n416783 , n416784 , n416785 , n416786 , n416787 , n94232 , n94233 , n416790 , n416791 , n94236 , 
 n416793 , n416794 , n416795 , n416796 , n416797 , n416798 , n416799 , n416800 , n416801 , n94246 , 
 n416803 , n416804 , n416805 , n416806 , n94251 , n416808 , n416809 , n94254 , n416811 , n416812 , 
 n94257 , n94258 , n416815 , n416816 , n94261 , n416818 , n416819 , n416820 , n416821 , n416822 , 
 n416823 , n416824 , n416825 , n416826 , n94271 , n416828 , n416829 , n416830 , n416831 , n416832 , 
 n416833 , n416834 , n416835 , n416836 , n416837 , n416838 , n416839 , n416840 , n416841 , n94286 , 
 n416843 , n416844 , n416845 , n416846 , n416847 , n416848 , n416849 , n94294 , n416851 , n416852 , 
 n416853 , n416854 , n416855 , n416856 , n416857 , n416858 , n416859 , n416860 , n94305 , n416862 , 
 n416863 , n416864 , n416865 , n416866 , n94311 , n416868 , n416869 , n94314 , n416871 , n416872 , 
 n416873 , n416874 , n416875 , n416876 , n416877 , n416878 , n416879 , n416880 , n416881 , n416882 , 
 n416883 , n94328 , n416885 , n416886 , n94331 , n416888 , n416889 , n94334 , n416891 , n416892 , 
 n416893 , n416894 , n416895 , n416896 , n416897 , n94342 , n416899 , n416900 , n94345 , n416902 , 
 n416903 , n416904 , n94349 , n416906 , n416907 , n416908 , n416909 , n416910 , n416911 , n416912 , 
 n94357 , n94358 , n416915 , n416916 , n416917 , n416918 , n94363 , n416920 , n416921 , n94366 , 
 n416923 , n416924 , n94369 , n416926 , n416927 , n416928 , n416929 , n416930 , n416931 , n416932 , 
 n94377 , n94378 , n416935 , n416936 , n416937 , n416938 , n416939 , n416940 , n416941 , n94386 , 
 n416943 , n94388 , n416945 , n416946 , n416947 , n416948 , n416949 , n416950 , n94395 , n416952 , 
 n94397 , n94398 , n416955 , n94400 , n94401 , n94402 , n94403 , n416960 , n94405 , n416962 , 
 n416963 , n94408 , n416965 , n416966 , n416967 , n416968 , n416969 , n416970 , n94415 , n416972 , 
 n416973 , n416974 , n416975 , n94420 , n94421 , n416978 , n94423 , n416980 , n416981 , n94426 , 
 n94427 , n94428 , n416985 , n416986 , n416987 , n416988 , n416989 , n416990 , n416991 , n94436 , 
 n94437 , n416994 , n416995 , n416996 , n416997 , n416998 , n416999 , n417000 , n94445 , n417002 , 
 n417003 , n417004 , n417005 , n417006 , n417007 , n417008 , n94453 , n417010 , n417011 , n417012 , 
 n94457 , n417014 , n417015 , n94460 , n417017 , n94462 , n94463 , n417020 , n417021 , n417022 , 
 n94467 , n417024 , n417025 , n417026 , n417027 , n417028 , n417029 , n417030 , n417031 , n94476 , 
 n417033 , n417034 , n417035 , n417036 , n417037 , n417038 , n417039 , n417040 , n417041 , n417042 , 
 n417043 , n94488 , n94489 , n417046 , n94491 , n417048 , n417049 , n417050 , n94495 , n417052 , 
 n417053 , n94498 , n94499 , n417056 , n417057 , n417058 , n417059 , n417060 , n417061 , n94506 , 
 n94507 , n417064 , n94509 , n417066 , n94511 , n94512 , n94513 , n417070 , n417071 , n417072 , 
 n417073 , n94518 , n417075 , n417076 , n417077 , n417078 , n94523 , n94524 , n417081 , n417082 , 
 n417083 , n417084 , n417085 , n417086 , n417087 , n417088 , n94533 , n94534 , n94535 , n417092 , 
 n94537 , n94538 , n417095 , n417096 , n417097 , n417098 , n417099 , n417100 , n417101 , n417102 , 
 n417103 , n94548 , n417105 , n417106 , n94551 , n417108 , n417109 , n94554 , n94555 , n417112 , 
 n94557 , n417114 , n417115 , n417116 , n417117 , n417118 , n417119 , n417120 , n94565 , n417122 , 
 n417123 , n417124 , n94569 , n94570 , n94571 , n417128 , n417129 , n417130 , n417131 , n417132 , 
 n417133 , n417134 , n94579 , n417136 , n417137 , n417138 , n417139 , n417140 , n417141 , n417142 , 
 n94587 , n417144 , n94589 , n417146 , n417147 , n417148 , n417149 , n94594 , n417151 , n417152 , 
 n94597 , n94598 , n417155 , n417156 , n417157 , n417158 , n417159 , n417160 , n417161 , n417162 , 
 n94607 , n417164 , n417165 , n94610 , n94611 , n417168 , n94613 , n94614 , n417171 , n417172 , 
 n94616 , n417174 , n417175 , n417176 , n417177 , n417178 , n417179 , n417180 , n417181 , n94623 , 
 n417183 , n417184 , n417185 , n417186 , n417187 , n417188 , n417189 , n417190 , n417191 , n417192 , 
 n417193 , n417194 , n417195 , n417196 , n417197 , n94635 , n417199 , n417200 , n417201 , n417202 , 
 n94640 , n417204 , n417205 , n417206 , n417207 , n94645 , n94646 , n417210 , n417211 , n417212 , 
 n417213 , n417214 , n417215 , n417216 , n417217 , n417218 , n417219 , n94656 , n94657 , n94658 , 
 n417223 , n417224 , n417225 , n417226 , n417227 , n417228 , n417229 , n417230 , n417231 , n417232 , 
 n417233 , n417234 , n417235 , n417236 , n417237 , n417238 , n94668 , n417240 , n417241 , n417242 , 
 n417243 , n417244 , n417245 , n417246 , n417247 , n417248 , n417249 , n417250 , n417251 , n94678 , 
 n417253 , n417254 , n94681 , n417256 , n94683 , n417258 , n417259 , n417260 , n417261 , n417262 , 
 n417263 , n417264 , n417265 , n417266 , n417267 , n94690 , n417269 , n417270 , n417271 , n417272 , 
 n417273 , n417274 , n417275 , n417276 , n94695 , n417278 , n417279 , n417280 , n417281 , n417282 , 
 n417283 , n417284 , n417285 , n417286 , n417287 , n417288 , n417289 , n417290 , n417291 , n417292 , 
 n417293 , n417294 , n417295 , n417296 , n417297 , n417298 , n417299 , n417300 , n417301 , n417302 , 
 n417303 , n417304 , n417305 , n417306 , n417307 , n417308 , n417309 , n417310 , n417311 , n417312 , 
 n417313 , n417314 , n417315 , n417316 , n417317 , n417318 , n417319 , n417320 , n417321 , n417322 , 
 n417323 , n417324 , n417325 , n417326 , n417327 , n417328 , n417329 , n417330 , n417331 , n417332 , 
 n417333 , n417334 , n417335 , n417336 , n417337 , n417338 , n417339 , n417340 , n417341 , n417342 , 
 n417343 , n417344 , n417345 , n417346 , n417347 , n417348 , n417349 , n417350 , n417351 , n417352 , 
 n417353 , n417354 , n417355 , n417356 , n417357 , n417358 , n417359 , n417360 , n417361 , n417362 , 
 n417363 , n417364 , n417365 , n417366 , n417367 , n417368 , n417369 , n417370 , n417371 , n417372 , 
 n417373 , n417374 , n417375 , n417376 , n417377 , n417378 , n417379 , n417380 , n417381 , n417382 , 
 n417383 , n417384 , n417385 , n417386 , n417387 , n417388 , n417389 , n94698 , n94699 , n417392 , 
 n417393 , n417394 , n417395 , n417396 , n417397 , n417398 , n417399 , n94706 , n417401 , n94708 , 
 n94709 , n94710 , n417405 , n417406 , n94713 , n417408 , n417409 , n417410 , n417411 , n417412 , 
 n417413 , n94720 , n417415 , n417416 , n417417 , n417418 , n94725 , n94726 , n417421 , n417422 , 
 n417423 , n417424 , n417425 , n417426 , n417427 , n417428 , n417429 , n417430 , n417431 , n417432 , 
 n417433 , n417434 , n417435 , n417436 , n417437 , n417438 , n417439 , n417440 , n417441 , n417442 , 
 n417443 , n417444 , n417445 , n417446 , n417447 , n417448 , n417449 , n417450 , n417451 , n417452 , 
 n417453 , n417454 , n417455 , n417456 , n417457 , n417458 , n417459 , n417460 , n417461 , n417462 , 
 n417463 , n417464 , n417465 , n417466 , n417467 , n417468 , n417469 , n417470 , n417471 , n417472 , 
 n417473 , n417474 , n417475 , n417476 , n417477 , n417478 , n417479 , n417480 , n417481 , n417482 , 
 n417483 , n417484 , n417485 , n417486 , n417487 , n417488 , n417489 , n417490 , n417491 , n417492 , 
 n417493 , n417494 , n417495 , n417496 , n417497 , n417498 , n417499 , n417500 , n94732 , n417502 , 
 n417503 , n417504 , n417505 , n94737 , n94738 , n417508 , n417509 , n417510 , n417511 , n417512 , 
 n417513 , n417514 , n417515 , n417516 , n417517 , n417518 , n417519 , n417520 , n94740 , n94741 , 
 n417523 , n417524 , n417525 , n417526 , n417527 , n417528 , n417529 , n417530 , n94750 , n94751 , 
 n417533 , n417534 , n94754 , n417536 , n417537 , n417538 , n417539 , n417540 , n417541 , n417542 , 
 n94762 , n94763 , n417545 , n417546 , n417547 , n417548 , n94768 , n94769 , n417551 , n417552 , 
 n417553 , n417554 , n417555 , n417556 , n417557 , n417558 , n94774 , n417560 , n417561 , n94777 , 
 n417563 , n417564 , n94780 , n417566 , n417567 , n94783 , n417569 , n417570 , n94786 , n417572 , 
 n417573 , n94789 , n94790 , n94791 , n417577 , n417578 , n94794 , n94795 , n94796 , n417582 , 
 n417583 , n94799 , n94800 , n94801 , n417587 , n94803 , n417589 , n94805 , n417591 , n94807 , 
 n94808 , n417594 , n417595 , n94811 , n94812 , n417598 , n94814 , n94815 , n94816 , n94817 , 
 n417603 , n94819 , n417605 , n94821 , n94822 , n417608 , n417609 , n94825 , n417611 , n417612 , 
 n94828 , n417614 , n417615 , n417616 , n94831 , n417618 , n417619 , n417620 , n94833 , n417622 , 
 n417623 , n417624 , n417625 , n417626 , n94835 , n94836 , n94837 , n94838 , n94839 , n94840 , 
 n94841 , n94842 , n417635 , n94844 , n94845 , n94846 , n417639 , n417640 , n417641 , n417642 , 
 n417643 , n94850 , n417645 , n417646 , n94852 , n417648 , n417649 , n94855 , n417651 , n417652 , 
 n94858 , n417654 , n417655 , n94861 , n94862 , n417658 , n417659 , n94865 , n417661 , n417662 , 
 n94868 , n417664 , n417665 , n94871 , n417667 , n94873 , n417669 , n94875 , n94876 , n417672 , 
 n417673 , n94879 , n417675 , n417676 , n94882 , n417678 , n417679 , n94885 , n94886 , n94887 , 
 n94888 , n417684 , n417685 , n94891 , n94892 , n94893 , n417689 , n417690 , n94896 , n417692 , 
 n417693 , n94899 , n417695 , n417696 , n94900 , n94901 , n94902 , n417700 , n94903 , n94904 , 
 n94905 , n94906 , n94907 , n417706 , n417707 , n94910 , n417709 , n94912 , n94913 , n417712 , 
 n417713 , n94916 , n417715 , n417716 , n94918 , n417718 , n417719 , n94921 , n417721 , n94923 , 
 n94924 , n94925 , n94926 , n417726 , n94928 , n94929 , n417729 , n417730 , n94932 , n417732 , 
 n417733 , n94935 , n94936 , n417736 , n94938 , n94939 , n417739 , n417740 , n417741 , n417742 , 
 n417743 , n417744 , n417745 , n417746 , n417747 , n417748 , n417749 , n94948 , n94949 , n417752 , 
 n94951 , n417754 , n417755 , n417756 , n417757 , n94956 , n94957 , n417760 , n417761 , n417762 , 
 n417763 , n94962 , n417765 , n94964 , n417767 , n417768 , n417769 , n94968 , n417771 , n94970 , 
 n417773 , n94972 , n94973 , n417776 , n417777 , n94976 , n417779 , n417780 , n417781 , n94980 , 
 n417783 , n417784 , n417785 , n94984 , n94985 , n417788 , n417789 , n417790 , n94989 , n417792 , 
 n417793 , n94992 , n417795 , n94994 , n417797 , n417798 , n417799 , n417800 , n94999 , n417802 , 
 n417803 , n417804 , n417805 , n417806 , n95005 , n417808 , n417809 , n95008 , n417811 , n417812 , 
 n95011 , n417814 , n417815 , n95014 , n417817 , n95016 , n95017 , n95018 , n95019 , n417822 , 
 n417823 , n417824 , n417825 , n95023 , n95024 , n417828 , n95026 , n95027 , n417831 , n417832 , 
 n417833 , n95031 , n417835 , n95033 , n95034 , n417838 , n95036 , n417840 , n417841 , n417842 , 
 n95038 , n417844 , n95040 , n417846 , n417847 , n95043 , n417849 , n417850 , n95046 , n417852 , 
 n95048 , n95049 , n417855 , n417856 , n95051 , n417858 , n95053 , n95054 , n417861 , n417862 , 
 n417863 , n417864 , n417865 , n417866 , n417867 , n417868 , n417869 , n417870 , n417871 , n417872 , 
 n417873 , n417874 , n417875 , n417876 , n417877 , n417878 , n417879 , n417880 , n417881 , n417882 , 
 n417883 , n417884 , n417885 , n417886 , n417887 , n417888 , n417889 , n417890 , n417891 , n417892 , 
 n417893 , n417894 , n417895 , n417896 , n417897 , n417898 , n417899 , n417900 , n417901 , n417902 , 
 n417903 , n417904 , n417905 , n417906 , n417907 , n417908 , n417909 , n417910 , n417911 , n417912 , 
 n417913 , n417914 , n417915 , n417916 , n417917 , n417918 , n417919 , n417920 , n417921 , n417922 , 
 n417923 , n417924 , n417925 , n417926 , n417927 , n417928 , n417929 , n417930 , n417931 , n417932 , 
 n417933 , n417934 , n417935 , n417936 , n417937 , n417938 , n417939 , n417940 , n417941 , n417942 , 
 n417943 , n417944 , n417945 , n417946 , n417947 , n417948 , n417949 , n417950 , n417951 , n417952 , 
 n417953 , n417954 , n417955 , n417956 , n417957 , n417958 , n417959 , n417960 , n417961 , n417962 , 
 n417963 , n417964 , n417965 , n417966 , n417967 , n417968 , n417969 , n417970 , n417971 , n417972 , 
 n417973 , n417974 , n417975 , n417976 , n417977 , n417978 , n417979 , n417980 , n417981 , n417982 , 
 n417983 , n417984 , n417985 , n417986 , n417987 , n417988 , n417989 , n417990 , n417991 , n417992 , 
 n417993 , n417994 , n417995 , n417996 , n417997 , n417998 , n417999 , n418000 , n418001 , n418002 , 
 n418003 , n418004 , n418005 , n418006 , n418007 , n418008 , n418009 , n418010 , n418011 , n418012 , 
 n418013 , n418014 , n418015 , n418016 , n418017 , n418018 , n418019 , n418020 , n418021 , n418022 , 
 n418023 , n418024 , n418025 , n418026 , n418027 , n418028 , n418029 , n418030 , n418031 , n418032 , 
 n418033 , n418034 , n418035 , n418036 , n418037 , n418038 , n418039 , n418040 , n418041 , n418042 , 
 n418043 , n418044 , n418045 , n418046 , n418047 , n418048 , n418049 , n418050 , n418051 , n418052 , 
 n418053 , n418054 , n418055 , n418056 , n418057 , n418058 , n418059 , n418060 , n418061 , n418062 , 
 n418063 , n418064 , n418065 , n418066 , n418067 , n418068 , n418069 , n418070 , n418071 , n418072 , 
 n418073 , n418074 , n418075 , n418076 , n418077 , n418078 , n418079 , n418080 , n418081 , n418082 , 
 n418083 , n418084 , n418085 , n418086 , n418087 , n418088 , n418089 , n418090 , n418091 , n418092 , 
 n418093 , n418094 , n418095 , n418096 , n418097 , n418098 , n418099 , n418100 , n418101 , n418102 , 
 n418103 , n418104 , n418105 , n418106 , n418107 , n418108 , n418109 , n418110 , n418111 , n418112 , 
 n418113 , n418114 , n418115 , n418116 , n418117 , n418118 , n418119 , n418120 , n418121 , n418122 , 
 n418123 , n418124 , n418125 , n418126 , n418127 , n418128 , n418129 , n418130 , n418131 , n418132 , 
 n418133 , n418134 , n418135 , n418136 , n418137 , n418138 , n418139 , n418140 , n418141 , n418142 , 
 n418143 , n418144 , n418145 , n418146 , n418147 , n418148 , n418149 , n418150 , n418151 , n418152 , 
 n418153 , n418154 , n418155 , n418156 , n418157 , n418158 , n418159 , n418160 , n418161 , n418162 , 
 n418163 , n418164 , n418165 , n418166 , n418167 , n418168 , n418169 , n418170 , n418171 , n418172 , 
 n418173 , n418174 , n418175 , n418176 , n418177 , n418178 , n418179 , n418180 , n418181 , n418182 , 
 n418183 , n418184 , n418185 , n418186 , n418187 , n418188 , n418189 , n418190 , n418191 , n418192 , 
 n418193 , n418194 , n418195 , n418196 , n418197 , n418198 , n418199 , n418200 , n418201 , n418202 , 
 n418203 , n418204 , n418205 , n418206 , n418207 , n418208 , n418209 , n418210 , n418211 , n418212 , 
 n418213 , n418214 , n418215 , n418216 , n418217 , n418218 , n418219 , n418220 , n418221 , n418222 , 
 n418223 , n418224 , n418225 , n418226 , n418227 , n418228 , n418229 , n418230 , n418231 , n418232 , 
 n418233 , n418234 , n418235 , n418236 , n418237 , n418238 , n418239 , n418240 , n418241 , n418242 , 
 n418243 , n418244 , n418245 , n418246 , n418247 , n418248 , n418249 , n418250 , n418251 , n418252 , 
 n418253 , n418254 , n418255 , n418256 , n418257 , n418258 , n418259 , n418260 , n418261 , n418262 , 
 n418263 , n418264 , n418265 , n418266 , n418267 , n418268 , n418269 , n418270 , n418271 , n418272 , 
 n418273 , n418274 , n418275 , n418276 , n418277 , n418278 , n418279 , n418280 , n418281 , n418282 , 
 n418283 , n418284 , n418285 , n418286 , n418287 , n418288 , n418289 , n418290 , n418291 , n418292 , 
 n418293 , n418294 , n418295 , n418296 , n418297 , n418298 , n418299 , n418300 , n418301 , n418302 , 
 n418303 , n418304 , n418305 , n418306 , n418307 , n418308 , n418309 , n418310 , n418311 , n418312 , 
 n418313 , n418314 , n418315 , n418316 , n418317 , n418318 , n418319 , n418320 , n418321 , n418322 , 
 n418323 , n418324 , n418325 , n418326 , n418327 , n418328 , n418329 , n418330 , n418331 , n418332 , 
 n418333 , n418334 , n418335 , n418336 , n418337 , n418338 , n418339 , n418340 , n418341 , n418342 , 
 n418343 , n418344 , n418345 , n418346 , n418347 , n418348 , n418349 , n418350 , n418351 , n418352 , 
 n418353 , n418354 , n418355 , n418356 , n418357 , n418358 , n418359 , n418360 , n418361 , n418362 , 
 n418363 , n418364 , n418365 , n418366 , n418367 , n418368 , n418369 , n418370 , n418371 , n418372 , 
 n418373 , n418374 , n418375 , n418376 , n418377 , n418378 , n418379 , n418380 , n418381 , n418382 , 
 n418383 , n418384 , n418385 , n418386 , n418387 , n418388 , n418389 , n418390 , n418391 , n418392 , 
 n418393 , n418394 , n418395 , n418396 , n418397 , n418398 , n418399 , n418400 , n418401 , n418402 , 
 n418403 , n418404 , n418405 , n418406 , n418407 , n418408 , n418409 , n418410 , n418411 , n418412 , 
 n418413 , n418414 , n418415 , n418416 , n418417 , n418418 , n418419 , n418420 , n418421 , n418422 , 
 n418423 , n418424 , n418425 , n418426 , n418427 , n418428 , n418429 , n418430 , n418431 , n418432 , 
 n418433 , n418434 , n418435 , n418436 , n418437 , n418438 , n418439 , n418440 , n418441 , n418442 , 
 n418443 , n418444 , n418445 , n418446 , n418447 , n418448 , n418449 , n418450 , n418451 , n418452 , 
 n418453 , n418454 , n418455 , n418456 , n418457 , n418458 , n418459 , n418460 , n418461 , n418462 , 
 n418463 , n418464 , n418465 , n418466 , n418467 , n418468 , n418469 , n418470 , n418471 , n418472 , 
 n418473 , n418474 , n418475 , n418476 , n418477 , n418478 , n418479 , n418480 , n418481 , n418482 , 
 n418483 , n418484 , n418485 , n418486 , n418487 , n418488 , n418489 , n418490 , n418491 , n418492 , 
 n418493 , n418494 , n418495 , n418496 , n418497 , n418498 , n418499 , n418500 , n418501 , n418502 , 
 n418503 , n418504 , n418505 , n418506 , n418507 , n418508 , n418509 , n418510 , n418511 , n418512 , 
 n418513 , n418514 , n418515 , n418516 , n418517 , n418518 , n418519 , n418520 , n418521 , n418522 , 
 n418523 , n418524 , n418525 , n418526 , n418527 , n418528 , n418529 , n418530 , n418531 , n418532 , 
 n418533 , n418534 , n418535 , n418536 , n418537 , n418538 , n418539 , n418540 , n418541 , n418542 , 
 n418543 , n418544 , n418545 , n418546 , n418547 , n418548 , n418549 , n418550 , n418551 , n418552 , 
 n418553 , n418554 , n418555 , n418556 , n418557 , n418558 , n418559 , n418560 , n418561 , n418562 , 
 n418563 , n418564 , n418565 , n418566 , n418567 , n418568 , n418569 , n418570 , n418571 , n418572 , 
 n418573 , n418574 , n418575 , n418576 , n418577 , n418578 , n418579 , n418580 , n418581 , n418582 , 
 n418583 , n418584 , n418585 , n418586 , n418587 , n418588 , n418589 , n418590 , n418591 , n418592 , 
 n418593 , n418594 , n418595 , n418596 , n418597 , n418598 , n418599 , n418600 , n418601 , n418602 , 
 n418603 , n418604 , n418605 , n418606 , n418607 , n418608 , n418609 , n418610 , n418611 , n418612 , 
 n418613 , n418614 , n418615 , n418616 , n418617 , n418618 , n418619 , n418620 , n418621 , n418622 , 
 n418623 , n418624 , n418625 , n418626 , n418627 , n418628 , n418629 , n418630 , n418631 , n418632 , 
 n418633 , n418634 , n418635 , n418636 , n418637 , n418638 , n418639 , n418640 , n418641 , n418642 , 
 n418643 , n418644 , n418645 , n418646 , n418647 , n418648 , n418649 , n418650 , n418651 , n418652 , 
 n418653 , n418654 , n418655 , n418656 , n418657 , n418658 , n418659 , n418660 , n418661 , n418662 , 
 n418663 , n418664 , n418665 , n418666 , n418667 , n418668 , n418669 , n418670 , n418671 , n418672 , 
 n418673 , n418674 , n418675 , n418676 , n418677 , n418678 , n418679 , n418680 , n418681 , n418682 , 
 n418683 , n418684 , n418685 , n418686 , n418687 , n418688 , n418689 , n418690 , n418691 , n418692 , 
 n418693 , n418694 , n418695 , n418696 , n418697 , n418698 , n418699 , n418700 , n418701 , n418702 , 
 n418703 , n418704 , n418705 , n418706 , n418707 , n418708 , n418709 , n418710 , n418711 , n418712 , 
 n418713 , n418714 , n418715 , n418716 , n418717 , n418718 , n418719 , n418720 , n418721 , n418722 , 
 n418723 , n418724 , n418725 , n418726 , n418727 , n418728 , n418729 , n418730 , n418731 , n418732 , 
 n418733 , n418734 , n418735 , n418736 , n418737 , n418738 , n418739 , n418740 , n418741 , n418742 , 
 n418743 , n418744 , n418745 , n418746 , n418747 , n418748 , n418749 , n418750 , n418751 , n418752 , 
 n418753 , n418754 , n418755 , n418756 , n418757 , n418758 , n418759 , n418760 , n418761 , n418762 , 
 n418763 , n418764 , n418765 , n418766 , n418767 , n418768 , n418769 , n418770 , n418771 , n418772 , 
 n418773 , n418774 , n418775 , n418776 , n418777 , n418778 , n418779 , n418780 , n418781 , n418782 , 
 n418783 , n418784 , n418785 , n418786 , n418787 , n418788 , n418789 , n418790 , n418791 , n418792 , 
 n418793 , n418794 , n418795 , n418796 , n418797 , n418798 , n418799 , n418800 , n418801 , n418802 , 
 n418803 , n418804 , n418805 , n418806 , n418807 , n418808 , n418809 , n418810 , n418811 , n418812 , 
 n418813 , n418814 , n418815 , n418816 , n418817 , n418818 , n418819 , n418820 , n418821 , n418822 , 
 n418823 , n418824 , n418825 , n418826 , n418827 , n418828 , n418829 , n418830 , n418831 , n418832 , 
 n418833 , n418834 , n418835 , n418836 , n418837 , n418838 , n418839 , n418840 , n418841 , n418842 , 
 n418843 , n418844 , n418845 , n418846 , n418847 , n418848 , n418849 , n418850 , n418851 , n418852 , 
 n418853 , n418854 , n418855 , n418856 , n418857 , n418858 , n418859 , n418860 , n418861 , n418862 , 
 n418863 , n418864 , n418865 , n418866 , n418867 , n418868 , n418869 , n418870 , n418871 , n418872 , 
 n418873 , n418874 , n418875 , n418876 , n418877 , n418878 , n418879 , n418880 , n418881 , n418882 , 
 n418883 , n418884 , n418885 , n418886 , n418887 , n418888 , n418889 , n418890 , n418891 , n418892 , 
 n418893 , n418894 , n418895 , n418896 , n418897 , n418898 , n418899 , n418900 , n418901 , n418902 , 
 n418903 , n418904 , n418905 , n418906 , n418907 , n418908 , n418909 , n418910 , n418911 , n418912 , 
 n418913 , n418914 , n418915 , n418916 , n418917 , n418918 , n418919 , n418920 , n418921 , n418922 , 
 n418923 , n418924 , n418925 , n418926 , n418927 , n418928 , n418929 , n418930 , n418931 , n418932 , 
 n418933 , n418934 , n418935 , n418936 , n418937 , n418938 , n418939 , n418940 , n418941 , n418942 , 
 n418943 , n418944 , n418945 , n418946 , n418947 , n418948 , n418949 , n418950 , n418951 , n418952 , 
 n418953 , n418954 , n418955 , n418956 , n418957 , n418958 , n418959 , n418960 , n418961 , n418962 , 
 n418963 , n418964 , n418965 , n418966 , n418967 , n418968 , n418969 , n418970 , n418971 , n418972 , 
 n418973 , n418974 , n418975 , n418976 , n418977 , n418978 , n418979 , n418980 , n418981 , n418982 , 
 n418983 , n418984 , n418985 , n418986 , n418987 , n418988 , n418989 , n418990 , n418991 , n418992 , 
 n418993 , n418994 , n418995 , n418996 , n418997 , n418998 , n418999 , n419000 , n419001 , n419002 , 
 n419003 , n419004 , n419005 , n419006 , n419007 , n419008 , n419009 , n419010 , n419011 , n419012 , 
 n419013 , n419014 , n419015 , n419016 , n419017 , n419018 , n419019 , n419020 , n419021 , n419022 , 
 n419023 , n419024 , n419025 , n419026 , n419027 , n419028 , n419029 , n419030 , n419031 , n419032 , 
 n419033 , n419034 , n419035 , n419036 , n419037 , n419038 , n419039 , n419040 , n419041 , n419042 , 
 n419043 , n419044 , n419045 , n419046 , n419047 , n419048 , n419049 , n419050 , n419051 , n419052 , 
 n419053 , n419054 , n419055 , n419056 , n419057 , n419058 , n419059 , n419060 , n419061 , n419062 , 
 n419063 , n419064 , n419065 , n419066 , n419067 , n419068 , n419069 , n419070 , n419071 , n419072 , 
 n419073 , n419074 , n419075 , n419076 , n419077 , n419078 , n419079 , n419080 , n419081 , n419082 , 
 n419083 , n419084 , n419085 , n419086 , n419087 , n419088 , n419089 , n419090 , n419091 , n419092 , 
 n419093 , n419094 , n419095 , n419096 , n419097 , n419098 , n419099 , n419100 , n419101 , n419102 , 
 n419103 , n419104 , n419105 , n419106 , n419107 , n419108 , n419109 , n419110 , n419111 , n419112 , 
 n419113 , n419114 , n419115 , n419116 , n419117 , n419118 , n419119 , n419120 , n419121 , n419122 , 
 n419123 , n419124 , n419125 , n419126 , n419127 , n419128 , n419129 , n419130 , n419131 , n419132 , 
 n419133 , n419134 , n419135 , n419136 , n419137 , n419138 , n419139 , n419140 , n419141 , n419142 , 
 n419143 , n419144 , n419145 , n419146 , n419147 , n419148 , n419149 , n419150 , n419151 , n419152 , 
 n419153 , n419154 , n419155 , n419156 , n419157 , n419158 , n419159 , n419160 , n419161 , n419162 , 
 n419163 , n419164 , n419165 , n419166 , n419167 , n419168 , n419169 , n419170 , n419171 , n419172 , 
 n419173 , n419174 , n419175 , n419176 , n419177 , n419178 , n419179 , n419180 , n419181 , n419182 , 
 n419183 , n419184 , n419185 , n419186 , n419187 , n419188 , n419189 , n419190 , n419191 , n419192 , 
 n419193 , n419194 , n419195 , n419196 , n419197 , n419198 , n419199 , n419200 , n419201 , n419202 , 
 n419203 , n419204 , n419205 , n419206 , n419207 , n419208 , n419209 , n419210 , n419211 , n419212 , 
 n419213 , n419214 , n419215 , n419216 , n419217 , n419218 , n419219 , n419220 , n419221 , n419222 , 
 n419223 , n419224 , n419225 , n419226 , n419227 , n419228 , n419229 , n419230 , n419231 , n419232 , 
 n419233 , n419234 , n419235 , n419236 , n419237 , n419238 , n419239 , n419240 , n419241 , n419242 , 
 n419243 , n419244 , n419245 , n419246 , n419247 , n419248 , n419249 , n419250 , n419251 , n419252 , 
 n419253 , n419254 , n419255 , n419256 , n419257 , n419258 , n419259 , n419260 , n419261 , n419262 , 
 n419263 , n419264 , n419265 , n419266 , n419267 , n419268 , n419269 , n419270 , n419271 , n419272 , 
 n419273 , n419274 , n419275 , n419276 , n419277 , n419278 , n419279 , n419280 , n419281 , n419282 , 
 n419283 , n419284 , n419285 , n419286 , n419287 , n419288 , n419289 , n419290 , n419291 , n419292 , 
 n419293 , n419294 , n419295 , n419296 , n419297 , n419298 , n419299 , n419300 , n419301 , n419302 , 
 n419303 , n419304 , n419305 , n419306 , n419307 , n419308 , n419309 , n419310 , n419311 , n419312 , 
 n419313 , n419314 , n419315 , n419316 , n419317 , n419318 , n419319 , n419320 , n419321 , n419322 , 
 n419323 , n419324 , n419325 , n419326 , n419327 , n419328 , n419329 , n419330 , n419331 , n419332 , 
 n419333 , n419334 , n419335 , n419336 , n419337 , n419338 , n419339 , n419340 , n419341 , n419342 , 
 n419343 , n419344 , n419345 , n419346 , n419347 , n419348 , n419349 , n419350 , n419351 , n419352 , 
 n419353 , n419354 , n419355 , n419356 , n419357 , n419358 , n419359 , n419360 , n419361 , n419362 , 
 n419363 , n419364 , n419365 , n419366 , n419367 , n419368 , n419369 , n419370 , n419371 , n419372 , 
 n419373 , n419374 , n419375 , n419376 , n419377 , n419378 , n419379 , n419380 , n419381 , n419382 , 
 n419383 , n419384 , n419385 , n419386 , n419387 , n419388 , n419389 , n419390 , n419391 , n419392 , 
 n419393 , n419394 , n419395 , n419396 , n419397 , n419398 , n419399 , n419400 , n419401 , n419402 , 
 n419403 , n419404 , n419405 , n419406 , n419407 , n419408 , n419409 , n419410 , n419411 , n419412 , 
 n419413 , n419414 , n419415 , n419416 , n419417 , n419418 , n419419 , n419420 , n419421 , n419422 , 
 n419423 , n419424 , n419425 , n419426 , n419427 , n419428 , n419429 , n419430 , n419431 , n419432 , 
 n419433 , n419434 , n419435 , n419436 , n419437 , n419438 , n419439 , n419440 , n419441 , n419442 , 
 n419443 , n419444 , n419445 , n419446 , n419447 , n419448 , n419449 , n419450 , n419451 , n419452 , 
 n419453 , n419454 , n419455 , n419456 , n419457 , n419458 , n419459 , n419460 , n419461 , n419462 , 
 n419463 , n419464 , n419465 , n419466 , n419467 , n419468 , n419469 , n419470 , n419471 , n419472 , 
 n419473 , n419474 , n419475 , n419476 , n419477 , n419478 , n419479 , n419480 , n419481 , n419482 , 
 n419483 , n419484 , n419485 , n419486 , n419487 , n419488 , n419489 , n419490 , n419491 , n419492 , 
 n419493 , n419494 , n419495 , n419496 , n419497 , n419498 , n419499 , n419500 , n419501 , n419502 , 
 n419503 , n419504 , n419505 , n419506 , n419507 , n419508 , n419509 , n419510 , n419511 , n419512 , 
 n419513 , n419514 , n419515 , n419516 , n419517 , n419518 , n419519 , n419520 , n419521 , n419522 , 
 n419523 , n419524 , n419525 , n419526 , n419527 , n419528 , n419529 , n419530 , n419531 , n419532 , 
 n419533 , n419534 , n419535 , n419536 , n419537 , n419538 , n419539 , n419540 , n419541 , n419542 , 
 n419543 , n419544 , n419545 , n419546 , n419547 , n419548 , n419549 , n419550 , n419551 , n419552 , 
 n419553 , n419554 , n419555 , n419556 , n419557 , n419558 , n419559 , n419560 , n419561 , n419562 , 
 n419563 , n419564 , n419565 , n419566 , n419567 , n419568 , n419569 , n419570 , n419571 , n419572 , 
 n419573 , n419574 , n419575 , n419576 , n419577 , n419578 , n419579 , n419580 , n419581 , n419582 , 
 n419583 , n419584 , n419585 , n419586 , n419587 , n419588 , n419589 , n419590 , n419591 , n419592 , 
 n419593 , n419594 , n419595 , n419596 , n419597 , n419598 , n419599 , n419600 , n419601 , n419602 , 
 n419603 , n419604 , n419605 , n419606 , n419607 , n419608 , n419609 , n419610 , n419611 , n419612 , 
 n419613 , n419614 , n419615 , n419616 , n419617 , n419618 , n419619 , n419620 , n419621 , n419622 , 
 n419623 , n419624 , n419625 , n419626 , n419627 , n419628 , n419629 , n419630 , n419631 , n419632 , 
 n419633 , n419634 , n419635 , n419636 , n419637 , n419638 , n419639 , n419640 , n419641 , n419642 , 
 n419643 , n419644 , n419645 , n419646 , n419647 , n419648 , n419649 , n419650 , n419651 , n419652 , 
 n419653 , n419654 , n419655 , n419656 , n419657 , n419658 , n419659 , n419660 , n419661 , n419662 , 
 n419663 , n419664 , n419665 , n419666 , n419667 , n419668 , n419669 , n419670 , n419671 , n419672 , 
 n419673 , n419674 , n419675 , n419676 , n419677 , n419678 , n419679 , n419680 , n419681 , n419682 , 
 n419683 , n419684 , n419685 , n419686 , n419687 , n419688 , n419689 , n419690 , n419691 , n419692 , 
 n419693 , n419694 , n419695 , n419696 , n419697 , n419698 , n419699 , n419700 , n419701 , n419702 , 
 n419703 , n419704 , n419705 , n419706 , n419707 , n419708 , n419709 , n419710 , n419711 , n419712 , 
 n419713 , n419714 , n419715 , n419716 , n419717 , n419718 , n419719 , n419720 , n419721 , n419722 , 
 n419723 , n419724 , n419725 , n419726 , n419727 , n419728 , n419729 , n419730 , n419731 , n419732 , 
 n419733 , n419734 , n419735 , n419736 , n419737 , n419738 , n419739 , n419740 , n419741 , n419742 , 
 n419743 , n419744 , n419745 , n419746 , n419747 , n419748 , n419749 , n419750 , n419751 , n419752 , 
 n419753 , n419754 , n419755 , n419756 , n419757 , n419758 , n419759 , n419760 , n419761 , n419762 , 
 n419763 , n419764 , n419765 , n419766 , n419767 , n419768 , n419769 , n419770 , n419771 , n419772 , 
 n419773 , n419774 , n419775 , n419776 , n419777 , n419778 , n419779 , n419780 , n419781 , n419782 , 
 n419783 , n419784 , n419785 , n419786 , n419787 , n419788 , n419789 , n419790 , n419791 , n419792 , 
 n419793 , n419794 , n419795 , n419796 , n419797 , n419798 , n419799 , n419800 , n419801 , n419802 , 
 n419803 , n419804 , n419805 , n419806 , n419807 , n419808 , n419809 , n419810 , n419811 , n419812 , 
 n419813 , n419814 , n419815 , n419816 , n419817 , n419818 , n419819 , n419820 , n419821 , n419822 , 
 n419823 , n419824 , n419825 , n419826 , n419827 , n419828 , n419829 , n419830 , n419831 , n419832 , 
 n419833 , n419834 , n419835 , n419836 , n419837 , n419838 , n419839 , n419840 , n419841 , n419842 , 
 n419843 , n419844 , n419845 , n419846 , n419847 , n419848 , n419849 , n419850 , n419851 , n419852 , 
 n419853 , n419854 , n419855 , n419856 , n419857 , n419858 , n419859 , n419860 , n419861 , n419862 , 
 n419863 , n419864 , n419865 , n419866 , n419867 , n419868 , n419869 , n419870 , n419871 , n419872 , 
 n419873 , n419874 , n419875 , n419876 , n419877 , n419878 , n419879 , n419880 , n419881 , n419882 , 
 n419883 , n419884 , n419885 , n419886 , n419887 , n419888 , n419889 , n419890 , n419891 , n419892 , 
 n419893 , n419894 , n419895 , n419896 , n419897 , n419898 , n419899 , n419900 , n419901 , n419902 , 
 n419903 , n419904 , n419905 , n419906 , n419907 , n419908 , n419909 , n419910 , n419911 , n419912 , 
 n419913 , n419914 , n419915 , n419916 , n419917 , n419918 , n419919 , n419920 , n419921 , n419922 , 
 n419923 , n419924 , n419925 , n419926 , n419927 , n419928 , n419929 , n419930 , n419931 , n419932 , 
 n419933 , n419934 , n419935 , n419936 , n419937 , n419938 , n419939 , n419940 , n419941 , n419942 , 
 n419943 , n419944 , n419945 , n419946 , n419947 , n419948 , n419949 , n419950 , n419951 , n419952 , 
 n419953 , n419954 , n419955 , n419956 , n419957 , n419958 , n419959 , n419960 , n419961 , n419962 , 
 n419963 , n419964 , n419965 , n419966 , n419967 , n419968 , n419969 , n419970 , n419971 , n419972 , 
 n419973 , n419974 , n419975 , n419976 , n419977 , n419978 , n419979 , n419980 , n419981 , n419982 , 
 n419983 , n419984 , n419985 , n419986 , n419987 , n419988 , n419989 , n419990 , n419991 , n419992 , 
 n419993 , n419994 , n419995 , n419996 , n419997 , n419998 , n419999 , n420000 , n420001 , n420002 , 
 n420003 , n420004 , n420005 , n420006 , n420007 , n420008 , n420009 , n420010 , n420011 , n420012 , 
 n420013 , n420014 , n420015 , n420016 , n420017 , n420018 , n420019 , n420020 , n420021 , n420022 , 
 n420023 , n420024 , n420025 , n420026 , n420027 , n420028 , n420029 , n420030 , n420031 , n420032 , 
 n420033 , n420034 , n420035 , n420036 , n420037 , n420038 , n420039 , n420040 , n420041 , n420042 , 
 n420043 , n420044 , n420045 , n420046 , n420047 , n420048 , n420049 , n420050 , n420051 , n420052 , 
 n420053 , n420054 , n420055 , n420056 , n420057 , n420058 , n420059 , n420060 , n420061 , n420062 , 
 n420063 , n420064 , n420065 , n420066 , n420067 , n420068 , n420069 , n420070 , n420071 , n420072 , 
 n420073 , n420074 , n420075 , n420076 , n420077 , n420078 , n420079 , n420080 , n420081 , n420082 , 
 n420083 , n420084 , n420085 , n420086 , n420087 , n420088 , n420089 , n420090 , n420091 , n420092 , 
 n420093 , n420094 , n420095 , n420096 , n420097 , n420098 , n420099 , n420100 , n420101 , n420102 , 
 n420103 , n420104 , n420105 , n420106 , n420107 , n420108 , n420109 , n420110 , n420111 , n420112 , 
 n420113 , n420114 , n420115 , n420116 , n420117 , n420118 , n420119 , n420120 , n420121 , n420122 , 
 n420123 , n420124 , n420125 , n420126 , n420127 , n420128 , n420129 , n420130 , n420131 , n420132 , 
 n420133 , n420134 , n420135 , n420136 , n420137 , n420138 , n420139 , n420140 , n420141 , n420142 , 
 n420143 , n420144 , n420145 , n420146 , n420147 , n420148 , n420149 , n420150 , n420151 , n420152 , 
 n420153 , n420154 , n420155 , n420156 , n420157 , n420158 , n420159 , n420160 , n420161 , n420162 , 
 n420163 , n420164 , n420165 , n420166 , n420167 , n420168 , n420169 , n420170 , n420171 , n420172 , 
 n420173 , n420174 , n420175 , n420176 , n420177 , n420178 , n420179 , n420180 , n420181 , n420182 , 
 n420183 , n420184 , n420185 , n420186 , n420187 , n420188 , n420189 , n420190 , n420191 , n420192 , 
 n420193 , n420194 , n420195 , n420196 , n420197 , n420198 , n420199 , n420200 , n420201 , n420202 , 
 n420203 , n420204 , n420205 , n420206 , n420207 , n420208 , n420209 , n420210 , n420211 , n420212 , 
 n420213 , n420214 , n420215 , n420216 , n420217 , n420218 , n420219 , n420220 , n420221 , n420222 , 
 n420223 , n420224 , n420225 , n420226 , n420227 , n420228 , n420229 , n420230 , n420231 , n420232 , 
 n420233 , n420234 , n420235 , n420236 , n420237 , n420238 , n420239 , n420240 , n420241 , n420242 , 
 n420243 , n420244 , n420245 , n420246 , n420247 , n420248 , n420249 , n420250 , n420251 , n420252 , 
 n420253 , n420254 , n420255 , n420256 , n420257 , n420258 , n420259 , n420260 , n420261 , n420262 , 
 n420263 , n420264 , n420265 , n420266 , n420267 , n420268 , n420269 , n420270 , n420271 , n420272 , 
 n420273 , n420274 , n420275 , n420276 , n420277 , n420278 , n420279 , n420280 , n420281 , n420282 , 
 n420283 , n420284 , n420285 , n420286 , n420287 , n420288 , n420289 , n420290 , n420291 , n420292 , 
 n420293 , n420294 , n420295 , n420296 , n420297 , n420298 , n420299 , n420300 , n420301 , n420302 , 
 n420303 , n420304 , n420305 , n420306 , n420307 , n420308 , n420309 , n420310 , n420311 , n420312 , 
 n420313 , n420314 , n420315 , n420316 , n420317 , n420318 , n420319 , n420320 , n420321 , n420322 , 
 n420323 , n420324 , n420325 , n420326 , n420327 , n420328 , n420329 , n420330 , n420331 , n420332 , 
 n420333 , n420334 , n420335 , n420336 , n420337 , n420338 , n420339 , n420340 , n420341 , n420342 , 
 n420343 , n420344 , n420345 , n420346 , n420347 , n420348 , n420349 , n420350 , n420351 , n420352 , 
 n420353 , n420354 , n420355 , n420356 , n420357 , n420358 , n420359 , n420360 , n420361 , n420362 , 
 n420363 , n420364 , n420365 , n420366 , n420367 , n420368 , n420369 , n420370 , n420371 , n420372 , 
 n420373 , n420374 , n420375 , n420376 , n420377 , n420378 , n420379 , n420380 , n420381 , n420382 , 
 n420383 , n420384 , n420385 , n420386 , n420387 , n420388 , n420389 , n420390 , n420391 , n420392 , 
 n420393 , n420394 , n420395 , n420396 , n420397 , n420398 , n420399 , n420400 , n420401 , n420402 , 
 n420403 , n420404 , n420405 , n420406 , n420407 , n420408 , n420409 , n420410 , n420411 , n420412 , 
 n420413 , n420414 , n420415 , n420416 , n420417 , n420418 , n420419 , n420420 , n420421 , n420422 , 
 n420423 , n420424 , n420425 , n420426 , n420427 , n420428 , n420429 , n420430 , n420431 , n420432 , 
 n420433 , n420434 , n420435 , n420436 , n420437 , n420438 , n420439 , n420440 , n420441 , n420442 , 
 n420443 , n420444 , n420445 , n420446 , n420447 , n420448 , n420449 , n420450 , n420451 , n420452 , 
 n420453 , n420454 , n420455 , n420456 , n420457 , n420458 , n420459 , n420460 , n420461 , n420462 , 
 n420463 , n420464 , n420465 , n420466 , n420467 , n420468 , n420469 , n420470 , n420471 , n420472 , 
 n420473 , n420474 , n420475 , n420476 , n420477 , n420478 , n420479 , n420480 , n420481 , n420482 , 
 n420483 , n420484 , n420485 , n420486 , n420487 , n420488 , n420489 , n420490 , n420491 , n420492 , 
 n420493 , n420494 , n420495 , n420496 , n420497 , n420498 , n420499 , n420500 , n420501 , n420502 , 
 n420503 , n420504 , n420505 , n420506 , n420507 , n420508 , n420509 , n420510 , n420511 , n420512 , 
 n420513 , n420514 , n420515 , n420516 , n420517 , n420518 , n420519 , n420520 , n420521 , n420522 , 
 n420523 , n420524 , n420525 , n420526 , n420527 , n420528 , n420529 , n420530 , n420531 , n420532 , 
 n420533 , n420534 , n420535 , n420536 , n420537 , n420538 , n420539 , n420540 , n420541 , n420542 , 
 n420543 , n420544 , n420545 , n420546 , n420547 , n420548 , n420549 , n420550 , n420551 , n420552 , 
 n420553 , n420554 , n420555 , n420556 , n420557 , n420558 , n420559 , n420560 , n420561 , n420562 , 
 n420563 , n420564 , n420565 , n420566 , n420567 , n420568 , n420569 , n420570 , n420571 , n420572 , 
 n420573 , n420574 , n420575 , n420576 , n420577 , n420578 , n420579 , n420580 , n420581 , n420582 , 
 n420583 , n420584 , n420585 , n420586 , n420587 , n420588 , n420589 , n420590 , n420591 , n420592 , 
 n420593 , n420594 , n420595 , n420596 , n420597 , n420598 , n420599 , n420600 , n420601 , n420602 , 
 n420603 , n420604 , n420605 , n420606 , n420607 , n420608 , n420609 , n420610 , n420611 , n420612 , 
 n420613 , n420614 , n420615 , n420616 , n420617 , n420618 , n420619 , n420620 , n420621 , n420622 , 
 n420623 , n420624 , n420625 , n420626 , n420627 , n420628 , n420629 , n420630 , n420631 , n420632 , 
 n420633 , n420634 , n420635 , n420636 , n420637 , n420638 , n420639 , n420640 , n420641 , n420642 , 
 n420643 , n420644 , n420645 , n420646 , n420647 , n420648 , n420649 , n420650 , n420651 , n420652 , 
 n420653 , n420654 , n420655 , n420656 , n420657 , n420658 , n420659 , n420660 , n420661 , n420662 , 
 n420663 , n420664 , n420665 , n420666 , n420667 , n420668 , n420669 , n420670 , n420671 , n420672 , 
 n420673 , n420674 , n420675 , n420676 , n420677 , n420678 , n420679 , n420680 , n420681 , n420682 , 
 n420683 , n420684 , n420685 , n420686 , n420687 , n420688 , n420689 , n420690 , n420691 , n420692 , 
 n420693 , n420694 , n420695 , n420696 , n420697 , n420698 , n420699 , n420700 , n420701 , n420702 , 
 n420703 , n420704 , n420705 , n420706 , n420707 , n420708 , n420709 , n420710 , n420711 , n420712 , 
 n420713 , n420714 , n420715 , n420716 , n420717 , n420718 , n420719 , n420720 , n420721 , n420722 , 
 n420723 , n420724 , n420725 , n420726 , n420727 , n420728 , n420729 , n420730 , n420731 , n420732 , 
 n420733 , n420734 , n420735 , n420736 , n420737 , n420738 , n420739 , n420740 , n420741 , n420742 , 
 n420743 , n420744 , n420745 , n420746 , n420747 , n420748 , n420749 , n420750 , n420751 , n420752 , 
 n420753 , n420754 , n420755 , n420756 , n420757 , n420758 , n420759 , n420760 , n420761 , n420762 , 
 n420763 , n420764 , n420765 , n420766 , n420767 , n420768 , n420769 , n420770 , n420771 , n420772 , 
 n420773 , n420774 , n420775 , n420776 , n420777 , n420778 , n420779 , n420780 , n420781 , n420782 , 
 n420783 , n420784 , n420785 , n420786 , n420787 , n420788 , n420789 , n420790 , n420791 , n420792 , 
 n420793 , n420794 , n420795 , n420796 , n420797 , n420798 , n420799 , n420800 , n420801 , n420802 , 
 n420803 , n420804 , n420805 , n420806 , n420807 , n420808 , n420809 , n420810 , n420811 , n420812 , 
 n420813 , n420814 , n420815 , n420816 , n420817 , n420818 , n420819 , n420820 , n420821 , n420822 , 
 n420823 , n420824 , n420825 , n420826 , n420827 , n420828 , n420829 , n420830 , n420831 , n420832 , 
 n420833 , n420834 , n420835 , n420836 , n420837 , n420838 , n420839 , n420840 , n420841 , n420842 , 
 n420843 , n420844 , n420845 , n420846 , n420847 , n420848 , n420849 , n420850 , n420851 , n420852 , 
 n420853 , n420854 , n420855 , n420856 , n420857 , n420858 , n420859 , n420860 , n420861 , n420862 , 
 n420863 , n420864 , n420865 , n420866 , n420867 , n420868 , n420869 , n420870 , n420871 , n420872 , 
 n420873 , n420874 , n420875 , n420876 , n420877 , n420878 , n420879 , n420880 , n420881 , n420882 , 
 n420883 , n420884 , n420885 , n420886 , n420887 , n420888 , n420889 , n420890 , n420891 , n420892 , 
 n420893 , n420894 , n420895 , n420896 , n420897 , n420898 , n420899 , n420900 , n420901 , n420902 , 
 n420903 , n420904 , n420905 , n420906 , n420907 , n420908 , n420909 , n420910 , n420911 , n420912 , 
 n420913 , n420914 , n420915 , n420916 , n420917 , n420918 , n420919 , n420920 , n420921 , n420922 , 
 n420923 , n420924 , n420925 , n420926 , n420927 , n420928 , n420929 , n420930 , n420931 , n420932 , 
 n420933 , n420934 , n420935 , n420936 , n420937 , n420938 , n420939 , n420940 , n420941 , n420942 , 
 n420943 , n420944 , n420945 , n420946 , n420947 , n420948 , n420949 , n420950 , n420951 , n420952 , 
 n420953 , n420954 , n420955 , n420956 , n420957 , n420958 , n420959 , n420960 , n420961 , n420962 , 
 n420963 , n420964 , n420965 , n420966 , n420967 , n420968 , n420969 , n420970 , n420971 , n420972 , 
 n420973 , n420974 , n420975 , n420976 , n420977 , n420978 , n420979 , n420980 , n420981 , n420982 , 
 n420983 , n420984 , n420985 , n420986 , n420987 , n420988 , n420989 , n420990 , n420991 , n420992 , 
 n420993 , n420994 , n420995 , n420996 , n420997 , n420998 , n420999 , n421000 , n421001 , n421002 , 
 n421003 , n421004 , n421005 , n421006 , n421007 , n421008 , n421009 , n421010 , n421011 , n421012 , 
 n421013 , n421014 , n421015 , n421016 , n421017 , n421018 , n421019 , n421020 , n421021 , n421022 , 
 n421023 , n421024 , n421025 , n421026 , n421027 , n421028 , n421029 , n421030 , n421031 , n421032 , 
 n421033 , n421034 , n421035 , n421036 , n421037 , n421038 , n421039 , n421040 , n421041 , n421042 , 
 n421043 , n421044 , n421045 , n421046 , n421047 , n421048 , n421049 , n421050 , n421051 , n421052 , 
 n421053 , n421054 , n421055 , n421056 , n421057 , n421058 , n421059 , n421060 , n421061 , n421062 , 
 n421063 , n421064 , n421065 , n421066 , n421067 , n421068 , n421069 , n421070 , n421071 , n421072 , 
 n421073 , n421074 , n421075 , n421076 , n421077 , n421078 , n421079 , n421080 , n421081 , n421082 , 
 n421083 , n421084 , n421085 , n421086 , n421087 , n421088 , n421089 , n421090 , n421091 , n421092 , 
 n421093 , n421094 , n421095 , n421096 , n421097 , n421098 , n421099 , n421100 , n421101 , n421102 , 
 n421103 , n421104 , n421105 , n421106 , n421107 , n421108 , n421109 , n421110 , n421111 , n421112 , 
 n421113 , n421114 , n421115 , n421116 , n421117 , n421118 , n421119 , n421120 , n421121 , n421122 , 
 n421123 , n421124 , n421125 , n421126 , n421127 , n421128 , n421129 , n421130 , n421131 , n421132 , 
 n421133 , n421134 , n421135 , n421136 , n421137 , n421138 , n421139 , n421140 , n421141 , n421142 , 
 n421143 , n421144 , n421145 , n421146 , n421147 , n421148 , n421149 , n421150 , n421151 , n421152 , 
 n421153 , n421154 , n421155 , n421156 , n421157 , n421158 , n421159 , n421160 , n421161 , n421162 , 
 n421163 , n421164 , n421165 , n421166 , n421167 , n421168 , n421169 , n421170 , n421171 , n421172 , 
 n421173 , n421174 , n421175 , n421176 , n421177 , n421178 , n421179 , n421180 , n421181 , n421182 , 
 n421183 , n421184 , n421185 , n421186 , n421187 , n421188 , n421189 , n421190 , n421191 , n421192 , 
 n421193 , n421194 , n421195 , n421196 , n421197 , n421198 , n421199 , n421200 , n421201 , n421202 , 
 n421203 , n421204 , n421205 , n421206 , n421207 , n421208 , n421209 , n421210 , n421211 , n421212 , 
 n421213 , n421214 , n421215 , n421216 , n421217 , n421218 , n421219 , n421220 , n421221 , n421222 , 
 n421223 , n421224 , n421225 , n421226 , n421227 , n421228 , n421229 , n421230 , n421231 , n421232 , 
 n421233 , n421234 , n421235 , n421236 , n421237 , n421238 , n421239 , n421240 , n421241 , n421242 , 
 n421243 , n421244 , n421245 , n421246 , n421247 , n421248 , n421249 , n421250 , n421251 , n421252 , 
 n421253 , n421254 , n421255 , n421256 , n421257 , n421258 , n421259 , n421260 , n421261 , n421262 , 
 n421263 , n421264 , n421265 , n421266 , n421267 , n421268 , n421269 , n421270 , n421271 , n421272 , 
 n421273 , n421274 , n421275 , n421276 , n421277 , n421278 , n421279 , n421280 , n421281 , n421282 , 
 n421283 , n421284 , n421285 , n421286 , n421287 , n421288 , n421289 , n421290 , n421291 , n421292 , 
 n421293 , n421294 , n421295 , n421296 , n421297 , n421298 , n421299 , n421300 , n421301 , n421302 , 
 n421303 , n421304 , n421305 , n421306 , n421307 , n421308 , n421309 , n421310 , n421311 , n421312 , 
 n421313 , n421314 , n421315 , n421316 , n421317 , n421318 , n421319 , n421320 , n421321 , n421322 , 
 n421323 , n421324 , n421325 , n421326 , n421327 , n421328 , n421329 , n421330 , n421331 , n421332 , 
 n421333 , n421334 , n421335 , n421336 , n421337 , n421338 , n421339 , n421340 , n421341 , n421342 , 
 n421343 , n421344 , n421345 , n421346 , n421347 , n421348 , n421349 , n421350 , n421351 , n421352 , 
 n421353 , n421354 , n421355 , n421356 , n421357 , n421358 , n421359 , n421360 , n421361 , n421362 , 
 n421363 , n421364 , n421365 , n421366 , n421367 , n421368 , n421369 , n421370 , n421371 , n421372 , 
 n421373 , n421374 , n421375 , n421376 , n421377 , n421378 , n421379 , n421380 , n421381 , n421382 , 
 n421383 , n421384 , n421385 , n421386 , n421387 , n421388 , n421389 , n421390 , n421391 , n421392 , 
 n421393 , n421394 , n421395 , n421396 , n421397 , n421398 , n421399 , n421400 , n421401 , n421402 , 
 n421403 , n421404 , n421405 , n421406 , n421407 , n421408 , n421409 , n421410 , n421411 , n421412 , 
 n421413 , n421414 , n421415 , n421416 , n421417 , n421418 , n421419 , n421420 , n421421 , n421422 , 
 n421423 , n421424 , n421425 , n421426 , n421427 , n421428 , n421429 , n421430 , n421431 , n421432 , 
 n421433 , n421434 , n421435 , n421436 , n421437 , n421438 , n421439 , n421440 , n421441 , n421442 , 
 n421443 , n421444 , n421445 , n421446 , n421447 , n421448 , n421449 , n421450 , n421451 , n421452 , 
 n421453 , n421454 , n421455 , n421456 , n421457 , n421458 , n421459 , n421460 , n421461 , n421462 , 
 n421463 , n421464 , n421465 , n421466 , n421467 , n421468 , n421469 , n421470 , n421471 , n421472 , 
 n421473 , n421474 , n421475 , n421476 , n421477 , n421478 , n421479 , n421480 , n421481 , n421482 , 
 n421483 , n421484 , n421485 , n421486 , n421487 , n421488 , n421489 , n421490 , n421491 , n421492 , 
 n421493 , n421494 , n421495 , n421496 , n421497 , n421498 , n421499 , n421500 , n421501 , n421502 , 
 n421503 , n421504 , n421505 , n421506 , n421507 , n421508 , n421509 , n421510 , n421511 , n421512 , 
 n421513 , n421514 , n421515 , n421516 , n421517 , n421518 , n421519 , n421520 , n421521 , n421522 , 
 n421523 , n421524 , n421525 , n421526 , n421527 , n421528 , n421529 , n421530 , n421531 , n421532 , 
 n421533 , n421534 , n421535 , n421536 , n421537 , n421538 , n421539 , n421540 , n421541 , n421542 , 
 n421543 , n421544 , n421545 , n421546 , n421547 , n421548 , n421549 , n421550 , n421551 , n421552 , 
 n421553 , n421554 , n421555 , n421556 , n421557 , n421558 , n421559 , n421560 , n421561 , n421562 , 
 n421563 , n421564 , n421565 , n421566 , n421567 , n421568 , n421569 , n421570 , n421571 , n421572 , 
 n421573 , n421574 , n421575 , n421576 , n421577 , n421578 , n421579 , n421580 , n421581 , n421582 , 
 n421583 , n421584 , n421585 , n421586 , n421587 , n421588 , n421589 , n421590 , n421591 , n421592 , 
 n421593 , n421594 , n421595 , n421596 , n421597 , n421598 , n421599 , n421600 , n421601 , n421602 , 
 n421603 , n421604 , n421605 , n421606 , n421607 , n421608 , n421609 , n421610 , n421611 , n421612 , 
 n421613 , n421614 , n421615 , n421616 , n421617 , n421618 , n421619 , n421620 , n421621 , n421622 , 
 n421623 , n421624 , n421625 , n421626 , n421627 , n421628 , n421629 , n421630 , n421631 , n421632 , 
 n421633 , n421634 , n421635 , n421636 , n421637 , n421638 , n421639 , n421640 , n421641 , n421642 , 
 n421643 , n421644 , n421645 , n421646 , n421647 , n421648 , n421649 , n421650 , n421651 , n421652 , 
 n421653 , n421654 , n421655 , n421656 , n421657 , n421658 , n421659 , n421660 , n421661 , n421662 , 
 n421663 , n421664 , n421665 , n421666 , n421667 , n421668 , n421669 , n421670 , n421671 , n421672 , 
 n421673 , n421674 , n421675 , n421676 , n421677 , n421678 , n421679 , n421680 , n421681 , n421682 , 
 n421683 , n421684 , n421685 , n421686 , n421687 , n421688 , n421689 , n421690 , n421691 , n421692 , 
 n421693 , n421694 , n421695 , n421696 , n421697 , n421698 , n421699 , n421700 , n421701 , n421702 , 
 n421703 , n421704 , n421705 , n421706 , n421707 , n421708 , n421709 , n421710 , n421711 , n421712 , 
 n421713 , n421714 , n421715 , n421716 , n421717 , n421718 , n421719 , C0n , C0 , C1n , 
 C1 ;
buf ( n544 , n0 );
buf ( n545 , n1 );
buf ( n546 , n2 );
buf ( n547 , n3 );
buf ( n548 , n4 );
buf ( n549 , n5 );
buf ( n550 , n6 );
buf ( n551 , n7 );
buf ( n552 , n8 );
buf ( n553 , n9 );
buf ( n554 , n10 );
buf ( n555 , n11 );
buf ( n556 , n12 );
buf ( n557 , n13 );
buf ( n558 , n14 );
buf ( n559 , n15 );
buf ( n560 , n16 );
buf ( n561 , n17 );
buf ( n562 , n18 );
buf ( n563 , n19 );
buf ( n564 , n20 );
buf ( n565 , n21 );
buf ( n566 , n22 );
buf ( n567 , n23 );
buf ( n568 , n24 );
buf ( n569 , n25 );
buf ( n570 , n26 );
buf ( n571 , n27 );
buf ( n572 , n28 );
buf ( n573 , n29 );
buf ( n574 , n30 );
buf ( n575 , n31 );
buf ( n576 , n32 );
buf ( n577 , n33 );
buf ( n578 , n34 );
buf ( n579 , n35 );
buf ( n580 , n36 );
buf ( n581 , n37 );
buf ( n582 , n38 );
buf ( n583 , n39 );
buf ( n584 , n40 );
buf ( n585 , n41 );
buf ( n586 , n42 );
buf ( n587 , n43 );
buf ( n588 , n44 );
buf ( n589 , n45 );
buf ( n590 , n46 );
buf ( n591 , n47 );
buf ( n592 , n48 );
buf ( n593 , n49 );
buf ( n594 , n50 );
buf ( n595 , n51 );
buf ( n596 , n52 );
buf ( n597 , n53 );
buf ( n598 , n54 );
buf ( n599 , n55 );
buf ( n600 , n56 );
buf ( n601 , n57 );
buf ( n602 , n58 );
buf ( n603 , n59 );
buf ( n604 , n60 );
buf ( n605 , n61 );
buf ( n606 , n62 );
buf ( n607 , n63 );
buf ( n608 , n64 );
buf ( n609 , n65 );
buf ( n610 , n66 );
buf ( n611 , n67 );
buf ( n612 , n68 );
buf ( n613 , n69 );
buf ( n614 , n70 );
buf ( n615 , n71 );
buf ( n616 , n72 );
buf ( n617 , n73 );
buf ( n618 , n74 );
buf ( n619 , n75 );
buf ( n620 , n76 );
buf ( n621 , n77 );
buf ( n622 , n78 );
buf ( n623 , n79 );
buf ( n80 , n624 );
buf ( n81 , n625 );
buf ( n82 , n626 );
buf ( n83 , n627 );
buf ( n84 , n628 );
buf ( n85 , n629 );
buf ( n86 , n630 );
buf ( n87 , n631 );
buf ( n88 , n632 );
buf ( n89 , n633 );
buf ( n90 , n634 );
buf ( n91 , n635 );
buf ( n92 , n636 );
buf ( n93 , n637 );
buf ( n94 , n638 );
buf ( n95 , n639 );
buf ( n96 , n640 );
buf ( n97 , n641 );
buf ( n98 , n642 );
buf ( n99 , n643 );
buf ( n100 , n644 );
buf ( n101 , n645 );
buf ( n102 , n646 );
buf ( n103 , n647 );
buf ( n104 , n648 );
buf ( n105 , n649 );
buf ( n106 , n650 );
buf ( n107 , n651 );
buf ( n108 , n652 );
buf ( n109 , n653 );
buf ( n110 , n654 );
buf ( n111 , n655 );
buf ( n112 , n656 );
buf ( n113 , n657 );
buf ( n114 , n658 );
buf ( n115 , n659 );
buf ( n116 , n660 );
buf ( n117 , n661 );
buf ( n118 , n662 );
buf ( n119 , n663 );
buf ( n120 , n664 );
buf ( n121 , n665 );
buf ( n122 , n666 );
buf ( n123 , n667 );
buf ( n124 , n668 );
buf ( n125 , n669 );
buf ( n126 , n670 );
buf ( n127 , n671 );
buf ( n128 , n672 );
buf ( n129 , n673 );
buf ( n130 , n674 );
buf ( n131 , n675 );
buf ( n132 , n676 );
buf ( n133 , n677 );
buf ( n134 , n678 );
buf ( n135 , n679 );
buf ( n136 , n680 );
buf ( n137 , n681 );
buf ( n138 , n682 );
buf ( n139 , n683 );
buf ( n140 , n684 );
buf ( n141 , n685 );
buf ( n142 , n686 );
buf ( n143 , n687 );
buf ( n144 , n688 );
buf ( n145 , n689 );
buf ( n146 , n690 );
buf ( n147 , n691 );
buf ( n148 , n692 );
buf ( n149 , n693 );
buf ( n150 , n694 );
buf ( n151 , n695 );
buf ( n152 , n696 );
buf ( n153 , n697 );
buf ( n154 , n698 );
buf ( n155 , n699 );
buf ( n156 , n700 );
buf ( n157 , n701 );
buf ( n158 , n702 );
buf ( n159 , n703 );
buf ( n160 , n704 );
buf ( n161 , n705 );
buf ( n162 , n706 );
buf ( n163 , n707 );
buf ( n164 , n708 );
buf ( n165 , n709 );
buf ( n166 , n710 );
buf ( n167 , n711 );
buf ( n168 , n712 );
buf ( n169 , n713 );
buf ( n170 , n714 );
buf ( n171 , n715 );
buf ( n172 , n716 );
buf ( n173 , n717 );
buf ( n174 , n718 );
buf ( n175 , n719 );
buf ( n176 , n720 );
buf ( n177 , n721 );
buf ( n178 , n722 );
buf ( n179 , n723 );
buf ( n180 , n724 );
buf ( n181 , n725 );
buf ( n182 , n726 );
buf ( n183 , n727 );
buf ( n184 , n728 );
buf ( n185 , n729 );
buf ( n186 , n730 );
buf ( n187 , n731 );
buf ( n188 , n732 );
buf ( n189 , n733 );
buf ( n190 , n734 );
buf ( n191 , n735 );
buf ( n192 , n736 );
buf ( n193 , n737 );
buf ( n194 , n738 );
buf ( n195 , n739 );
buf ( n196 , n740 );
buf ( n197 , n741 );
buf ( n198 , n742 );
buf ( n199 , n743 );
buf ( n200 , n744 );
buf ( n201 , n745 );
buf ( n202 , n746 );
buf ( n203 , n747 );
buf ( n204 , n748 );
buf ( n205 , n749 );
buf ( n206 , n750 );
buf ( n207 , n751 );
buf ( n208 , n752 );
buf ( n209 , n753 );
buf ( n210 , n754 );
buf ( n211 , n755 );
buf ( n212 , n756 );
buf ( n213 , n757 );
buf ( n214 , n758 );
buf ( n215 , n759 );
buf ( n216 , n760 );
buf ( n217 , n761 );
buf ( n218 , n762 );
buf ( n219 , n763 );
buf ( n220 , n764 );
buf ( n221 , n765 );
buf ( n222 , n766 );
buf ( n223 , n767 );
buf ( n224 , n768 );
buf ( n225 , n769 );
buf ( n226 , n770 );
buf ( n227 , n771 );
buf ( n228 , n772 );
buf ( n229 , n773 );
buf ( n230 , n774 );
buf ( n231 , n775 );
buf ( n232 , n776 );
buf ( n233 , n777 );
buf ( n234 , n778 );
buf ( n235 , n779 );
buf ( n236 , n780 );
buf ( n237 , n781 );
buf ( n238 , n782 );
buf ( n239 , n783 );
buf ( n240 , n784 );
buf ( n241 , n785 );
buf ( n242 , n786 );
buf ( n243 , n787 );
buf ( n244 , n788 );
buf ( n245 , n789 );
buf ( n246 , n790 );
buf ( n247 , n791 );
buf ( n248 , n792 );
buf ( n249 , n793 );
buf ( n250 , n794 );
buf ( n251 , n795 );
buf ( n252 , n796 );
buf ( n253 , n797 );
buf ( n254 , n798 );
buf ( n255 , n799 );
buf ( n256 , n800 );
buf ( n257 , n801 );
buf ( n258 , n802 );
buf ( n259 , n803 );
buf ( n260 , n804 );
buf ( n261 , n805 );
buf ( n262 , n806 );
buf ( n263 , n807 );
buf ( n264 , n808 );
buf ( n265 , n809 );
buf ( n266 , n810 );
buf ( n267 , n811 );
buf ( n268 , n812 );
buf ( n269 , n813 );
buf ( n270 , n814 );
buf ( n271 , n815 );
buf ( n624 , n421595 );
buf ( n625 , n343349 );
buf ( n626 , n343357 );
buf ( n627 , n343360 );
buf ( n628 , n343363 );
buf ( n629 , n343366 );
buf ( n630 , n23519 );
buf ( n631 , n343512 );
buf ( n632 , n343508 );
buf ( n633 , n343500 );
buf ( n634 , n343399 );
buf ( n635 , n343402 );
buf ( n636 , n421607 );
buf ( n637 , n421604 );
buf ( n638 , n421601 );
buf ( n639 , n421598 );
buf ( n640 , n343405 );
buf ( n641 , n343408 );
buf ( n642 , n343411 );
buf ( n643 , n421587 );
buf ( n644 , n343423 );
buf ( n645 , n343435 );
buf ( n646 , n343438 );
buf ( n647 , n343446 );
buf ( n648 , n23463 );
buf ( n649 , n23475 );
buf ( n650 , n343473 );
buf ( n651 , n421645 );
buf ( n652 , n343476 );
buf ( n653 , n421615 );
buf ( n654 , n421612 );
buf ( n655 , n321494 );
buf ( n656 , n421591 );
buf ( n657 , n352666 );
buf ( n658 , n352674 );
buf ( n659 , n352818 );
buf ( n660 , n421579 );
buf ( n661 , n352822 );
buf ( n662 , n352692 );
buf ( n663 , n352695 );
buf ( n664 , n352698 );
buf ( n665 , n352701 );
buf ( n666 , n352704 );
buf ( n667 , n32674 );
buf ( n668 , n352710 );
buf ( n669 , n352713 );
buf ( n670 , n352716 );
buf ( n671 , n352728 );
buf ( n672 , n421719 );
buf ( n673 , n421544 );
buf ( n674 , n352731 );
buf ( n675 , n352739 );
buf ( n676 , n352751 );
buf ( n677 , n352759 );
buf ( n678 , n352767 );
buf ( n679 , n352775 );
buf ( n680 , n421550 );
buf ( n681 , n352783 );
buf ( n682 , n352786 );
buf ( n683 , n352789 );
buf ( n684 , n352792 );
buf ( n685 , n352795 );
buf ( n686 , n352798 );
buf ( n687 , n352427 );
buf ( n688 , n421450 );
buf ( n689 , n421450 );
buf ( n690 , n421450 );
buf ( n691 , n421450 );
buf ( n692 , n421450 );
buf ( n693 , n421450 );
buf ( n694 , n421450 );
buf ( n695 , n421450 );
buf ( n696 , n421450 );
buf ( n697 , n421450 );
buf ( n698 , n421450 );
buf ( n699 , n421450 );
buf ( n700 , n421450 );
buf ( n701 , n421450 );
buf ( n702 , n421450 );
buf ( n703 , n421450 );
buf ( n704 , n421450 );
buf ( n705 , n421450 );
buf ( n706 , n421450 );
buf ( n707 , n421450 );
buf ( n708 , n421450 );
buf ( n709 , n421450 );
buf ( n710 , n421450 );
buf ( n711 , n421450 );
buf ( n712 , n421450 );
buf ( n713 , n421450 );
buf ( n714 , n421450 );
buf ( n715 , n421450 );
buf ( n716 , n421454 );
buf ( n717 , n421359 );
buf ( n718 , n421325 );
buf ( n719 , n421243 );
buf ( n720 , n420118 );
buf ( n721 , n419623 );
buf ( n722 , n419717 );
buf ( n723 , n421462 );
buf ( n724 , n419732 );
buf ( n725 , n419673 );
buf ( n726 , n421500 );
buf ( n727 , n419651 );
buf ( n728 , n421437 );
buf ( n729 , n421640 );
buf ( n730 , n419754 );
buf ( n731 , n419774 );
buf ( n732 , n421202 );
buf ( n733 , n421432 );
buf ( n734 , n421410 );
buf ( n735 , n421395 );
buf ( n736 , n421399 );
buf ( n737 , n421512 );
buf ( n738 , n421663 );
buf ( n739 , n421527 );
buf ( n740 , n421650 );
buf ( n741 , n421628 );
buf ( n742 , n421266 );
buf ( n743 , n421676 );
buf ( n744 , n421533 );
buf ( n745 , n420244 );
buf ( n746 , n421276 );
buf ( n747 , n420203 );
buf ( n748 , n421196 );
buf ( n749 , n421381 );
buf ( n750 , n421489 );
buf ( n751 , n421475 );
buf ( n752 , n419996 );
buf ( n753 , n420175 );
buf ( n754 , n420145 );
buf ( n755 , n421296 );
buf ( n756 , n421300 );
buf ( n757 , n421342 );
buf ( n758 , n419860 );
buf ( n759 , n419888 );
buf ( n760 , n421385 );
buf ( n761 , n419937 );
buf ( n762 , n421184 );
buf ( n763 , n420305 );
buf ( n764 , n420316 );
buf ( n765 , n421703 );
buf ( n766 , n421711 );
buf ( n767 , n420284 );
buf ( n768 , n420331 );
buf ( n769 , n420343 );
buf ( n770 , n420362 );
buf ( n771 , n421541 );
buf ( n772 , n420398 );
buf ( n773 , n420413 );
buf ( n774 , n420439 );
buf ( n775 , n420465 );
buf ( n776 , n420480 );
buf ( n777 , n420497 );
buf ( n778 , n421718 );
buf ( n779 , n420539 );
buf ( n780 , n420562 );
buf ( n781 , n420576 );
buf ( n782 , n421147 );
buf ( n783 , n421151 );
buf ( n784 , n421573 );
buf ( n785 , n421688 );
buf ( n786 , n421155 );
buf ( n787 , n421163 );
buf ( n788 , n421167 );
buf ( n789 , n421171 );
buf ( n790 , n420596 );
buf ( n791 , n420599 );
buf ( n792 , n420602 );
buf ( n793 , n420623 );
buf ( n794 , n421565 );
buf ( n795 , n421175 );
buf ( n796 , n421180 );
buf ( n797 , n420660 );
buf ( n798 , n421188 );
buf ( n799 , n421192 );
buf ( n800 , n421559 );
buf ( n801 , n420701 );
buf ( n802 , n420715 );
buf ( n803 , n420729 );
buf ( n804 , n420742 );
buf ( n805 , n420787 );
buf ( n806 , n420799 );
buf ( n807 , n420832 );
buf ( n808 , n421610 );
buf ( n809 , n420859 );
buf ( n810 , n421032 );
buf ( n811 , n421053 );
buf ( n812 , n421060 );
buf ( n813 , n421071 );
buf ( n814 , n421074 );
buf ( n815 , n421139 );
buf ( n320434 , n555 );
buf ( n320435 , n574 );
xor ( n320436 , n320434 , n320435 );
buf ( n320437 , n320436 );
not ( n320438 , n320437 );
not ( n320439 , n575 );
nand ( n320440 , n320439 , n574 );
not ( n320441 , n320440 );
not ( n320442 , n320441 );
or ( n320443 , n320438 , n320442 );
not ( n320444 , n554 );
and ( n320445 , n574 , n320444 );
not ( n320446 , n574 );
and ( n320447 , n320446 , n554 );
or ( n320448 , n320445 , n320447 );
buf ( n320449 , n320448 );
buf ( n320450 , n575 );
nand ( n320451 , n320449 , n320450 );
buf ( n320452 , n320451 );
nand ( n320453 , n320443 , n320452 );
buf ( n320454 , n559 );
buf ( n320455 , n571 );
or ( n320456 , n320454 , n320455 );
buf ( n320457 , n572 );
nand ( n320458 , n320456 , n320457 );
buf ( n320459 , n320458 );
buf ( n320460 , n559 );
buf ( n320461 , n571 );
nand ( n320462 , n320460 , n320461 );
buf ( n320463 , n320462 );
and ( n320464 , n320459 , n320463 , n570 );
nand ( n320465 , n320453 , n320464 );
buf ( n320466 , n558 );
buf ( n320467 , n570 );
xor ( n320468 , n320466 , n320467 );
buf ( n320469 , n320468 );
buf ( n320470 , n320469 );
not ( n320471 , n320470 );
xor ( n320472 , n571 , n570 );
not ( n320473 , n320472 );
xor ( n320474 , n571 , n572 );
nor ( n320475 , n320473 , n320474 );
buf ( n320476 , n320475 );
buf ( n320477 , n320476 );
not ( n320478 , n320477 );
or ( n320479 , n320471 , n320478 );
xor ( n320480 , n571 , n572 );
buf ( n320481 , n320480 );
buf ( n320482 , n320481 );
buf ( n320483 , n320482 );
buf ( n320484 , n320483 );
buf ( n320485 , n557 );
buf ( n320486 , n570 );
xor ( n320487 , n320485 , n320486 );
buf ( n320488 , n320487 );
buf ( n320489 , n320488 );
nand ( n320490 , n320484 , n320489 );
buf ( n320491 , n320490 );
buf ( n320492 , n320491 );
nand ( n320493 , n320479 , n320492 );
buf ( n320494 , n320493 );
xor ( n320495 , n320465 , n320494 );
xor ( n320496 , n569 , n570 );
buf ( n320497 , n320496 );
buf ( n320498 , n320497 );
buf ( n320499 , n320498 );
buf ( n320500 , n320499 );
buf ( n320501 , n559 );
and ( n320502 , n320500 , n320501 );
buf ( n320503 , n320502 );
buf ( n320504 , n320503 );
not ( n320505 , n320441 );
not ( n320506 , n320448 );
or ( n320507 , n320505 , n320506 );
not ( n320508 , n553 );
not ( n320509 , n574 );
not ( n320510 , n320509 );
or ( n320511 , n320508 , n320510 );
not ( n320512 , n553 );
nand ( n320513 , n320512 , n574 );
nand ( n320514 , n320511 , n320513 );
nand ( n320515 , n320514 , n575 );
nand ( n320516 , n320507 , n320515 );
buf ( n320517 , n320516 );
xor ( n320518 , n320504 , n320517 );
buf ( n320519 , n556 );
buf ( n320520 , n572 );
xor ( n320521 , n320519 , n320520 );
buf ( n320522 , n320521 );
buf ( n320523 , n320522 );
not ( n320524 , n320523 );
xor ( n320525 , n573 , n574 );
not ( n320526 , n320525 );
xor ( n320527 , n573 , n572 );
nand ( n320528 , n320526 , n320527 );
buf ( n320529 , n320528 );
not ( n320530 , n320529 );
buf ( n320531 , n320530 );
buf ( n320532 , n320531 );
not ( n320533 , n320532 );
or ( n320534 , n320524 , n320533 );
xor ( n320535 , n573 , n574 );
buf ( n320536 , n320535 );
buf ( n320537 , n555 );
buf ( n320538 , n572 );
xor ( n320539 , n320537 , n320538 );
buf ( n320540 , n320539 );
buf ( n320541 , n320540 );
nand ( n320542 , n320536 , n320541 );
buf ( n320543 , n320542 );
buf ( n320544 , n320543 );
nand ( n320545 , n320534 , n320544 );
buf ( n320546 , n320545 );
buf ( n320547 , n320546 );
xor ( n320548 , n320518 , n320547 );
buf ( n320549 , n320548 );
xnor ( n320550 , n320495 , n320549 );
buf ( n320551 , n320550 );
buf ( n320552 , n320474 );
buf ( n320553 , n559 );
and ( n320554 , n320552 , n320553 );
buf ( n320555 , n320554 );
buf ( n320556 , n320555 );
buf ( n320557 , n556 );
buf ( n320558 , n574 );
xor ( n320559 , n320557 , n320558 );
buf ( n320560 , n320559 );
buf ( n320561 , n320560 );
not ( n823 , n320561 );
buf ( n320563 , n320441 );
not ( n825 , n320563 );
or ( n320565 , n823 , n825 );
buf ( n320566 , n320437 );
buf ( n320567 , n575 );
nand ( n829 , n320566 , n320567 );
buf ( n320569 , n829 );
buf ( n320570 , n320569 );
nand ( n832 , n320565 , n320570 );
buf ( n833 , n832 );
buf ( n320573 , n833 );
xor ( n835 , n320556 , n320573 );
xor ( n320575 , n572 , n558 );
buf ( n320576 , n320575 );
not ( n838 , n320576 );
buf ( n320578 , n320531 );
not ( n320579 , n320578 );
or ( n841 , n838 , n320579 );
buf ( n320581 , n320535 );
buf ( n843 , n557 );
buf ( n320583 , n572 );
xor ( n320584 , n843 , n320583 );
buf ( n320585 , n320584 );
buf ( n320586 , n320585 );
nand ( n320587 , n320581 , n320586 );
buf ( n320588 , n320587 );
buf ( n320589 , n320588 );
nand ( n320590 , n841 , n320589 );
buf ( n320591 , n320590 );
buf ( n320592 , n320591 );
and ( n320593 , n835 , n320592 );
and ( n855 , n320556 , n320573 );
or ( n320595 , n320593 , n855 );
buf ( n320596 , n320595 );
buf ( n858 , n320596 );
and ( n320598 , n587 , n588 );
not ( n860 , n587 );
not ( n320600 , n588 );
and ( n320601 , n860 , n320600 );
nor ( n863 , n320598 , n320601 );
and ( n320603 , n863 , n559 );
buf ( n320604 , n320603 );
buf ( n320605 , n556 );
buf ( n320606 , n590 );
xor ( n320607 , n320605 , n320606 );
buf ( n320608 , n320607 );
buf ( n320609 , n320608 );
not ( n320610 , n320609 );
not ( n320611 , n591 );
and ( n873 , n320611 , n590 );
buf ( n320613 , n873 );
not ( n875 , n320613 );
or ( n876 , n320610 , n875 );
buf ( n320616 , n555 );
buf ( n320617 , n590 );
xor ( n879 , n320616 , n320617 );
buf ( n320619 , n879 );
buf ( n320620 , n320619 );
buf ( n320621 , n591 );
nand ( n883 , n320620 , n320621 );
buf ( n320623 , n883 );
buf ( n320624 , n320623 );
nand ( n886 , n876 , n320624 );
buf ( n320626 , n886 );
buf ( n320627 , n320626 );
xor ( n320628 , n320604 , n320627 );
buf ( n890 , n558 );
buf ( n891 , n588 );
xor ( n892 , n890 , n891 );
buf ( n893 , n892 );
buf ( n320633 , n893 );
not ( n895 , n320633 );
xnor ( n320635 , n589 , n590 );
xor ( n320636 , n589 , n588 );
and ( n898 , n320635 , n320636 );
buf ( n320638 , n898 );
not ( n900 , n320638 );
or ( n320640 , n895 , n900 );
xor ( n902 , n589 , n590 );
buf ( n320642 , n902 );
buf ( n320643 , n320642 );
buf ( n320644 , n557 );
buf ( n320645 , n588 );
xor ( n320646 , n320644 , n320645 );
buf ( n320647 , n320646 );
buf ( n320648 , n320647 );
nand ( n320649 , n320643 , n320648 );
buf ( n320650 , n320649 );
buf ( n320651 , n320650 );
nand ( n320652 , n320640 , n320651 );
buf ( n320653 , n320652 );
buf ( n320654 , n320653 );
and ( n320655 , n320628 , n320654 );
and ( n320656 , n320604 , n320627 );
or ( n320657 , n320655 , n320656 );
buf ( n320658 , n320657 );
buf ( n320659 , n320658 );
xor ( n921 , n858 , n320659 );
buf ( n320661 , n320647 );
not ( n923 , n320661 );
not ( n320663 , n902 );
nand ( n320664 , n320663 , n320636 );
not ( n926 , n320664 );
buf ( n320666 , n926 );
not ( n928 , n320666 );
or ( n929 , n923 , n928 );
buf ( n320669 , n320642 );
buf ( n320670 , n556 );
buf ( n320671 , n588 );
xor ( n933 , n320670 , n320671 );
buf ( n320673 , n933 );
buf ( n320674 , n320673 );
nand ( n320675 , n320669 , n320674 );
buf ( n320676 , n320675 );
buf ( n320677 , n320676 );
nand ( n320678 , n929 , n320677 );
buf ( n320679 , n320678 );
buf ( n320680 , n320679 );
buf ( n320681 , n559 );
buf ( n320682 , n586 );
xor ( n944 , n320681 , n320682 );
buf ( n320684 , n944 );
buf ( n320685 , n320684 );
not ( n947 , n320685 );
xnor ( n320687 , n587 , n586 );
xor ( n320688 , n587 , n588 );
nor ( n320689 , n320687 , n320688 );
buf ( n320690 , n320689 );
buf ( n320691 , n320690 );
buf ( n320692 , n320691 );
buf ( n320693 , n320692 );
not ( n320694 , n320693 );
or ( n320695 , n947 , n320694 );
not ( n320696 , n320688 );
buf ( n320697 , n320696 );
not ( n959 , n320697 );
buf ( n320699 , n959 );
buf ( n320700 , n320699 );
buf ( n320701 , n558 );
buf ( n320702 , n586 );
xor ( n320703 , n320701 , n320702 );
buf ( n320704 , n320703 );
buf ( n320705 , n320704 );
nand ( n320706 , n320700 , n320705 );
buf ( n320707 , n320706 );
buf ( n320708 , n320707 );
nand ( n970 , n320695 , n320708 );
buf ( n971 , n970 );
buf ( n320711 , n971 );
xor ( n973 , n320680 , n320711 );
buf ( n320713 , n559 );
buf ( n320714 , n587 );
or ( n976 , n320713 , n320714 );
buf ( n320716 , n588 );
nand ( n320717 , n976 , n320716 );
buf ( n320718 , n320717 );
buf ( n320719 , n320718 );
buf ( n320720 , n559 );
buf ( n320721 , n587 );
nand ( n983 , n320720 , n320721 );
buf ( n320723 , n983 );
buf ( n320724 , n320723 );
buf ( n320725 , n586 );
and ( n987 , n320719 , n320724 , n320725 );
buf ( n320727 , n987 );
buf ( n320728 , n320727 );
buf ( n320729 , n320619 );
not ( n991 , n320729 );
nand ( n992 , n320611 , n590 );
not ( n320732 , n992 );
buf ( n320733 , n320732 );
not ( n995 , n320733 );
or ( n320735 , n991 , n995 );
and ( n320736 , n554 , n590 );
not ( n998 , n554 );
buf ( n320738 , n590 );
not ( n320739 , n320738 );
buf ( n320740 , n320739 );
and ( n320741 , n998 , n320740 );
nor ( n1003 , n320736 , n320741 );
nand ( n320743 , n1003 , n591 );
buf ( n320744 , n320743 );
nand ( n320745 , n320735 , n320744 );
buf ( n320746 , n320745 );
buf ( n320747 , n320746 );
xor ( n320748 , n320728 , n320747 );
buf ( n320749 , n320748 );
buf ( n320750 , n320749 );
xor ( n320751 , n973 , n320750 );
buf ( n320752 , n320751 );
buf ( n320753 , n320752 );
and ( n320754 , n921 , n320753 );
and ( n320755 , n858 , n320659 );
or ( n1017 , n320754 , n320755 );
buf ( n320757 , n1017 );
buf ( n1019 , n320757 );
xor ( n1020 , n320551 , n1019 );
not ( n320760 , n320585 );
not ( n320761 , n320527 );
nor ( n1023 , n320761 , n320525 );
not ( n1024 , n1023 );
or ( n1025 , n320760 , n1024 );
buf ( n1026 , n320525 );
buf ( n320766 , n1026 );
buf ( n320767 , n320522 );
nand ( n1029 , n320766 , n320767 );
buf ( n320769 , n1029 );
nand ( n1031 , n1025 , n320769 );
buf ( n320771 , n1031 );
not ( n1033 , n320771 );
xor ( n1034 , n320464 , n320453 );
buf ( n320774 , n1034 );
not ( n1036 , n320774 );
or ( n320776 , n1033 , n1036 );
or ( n320777 , n1034 , n1031 );
buf ( n320778 , n559 );
buf ( n320779 , n570 );
xor ( n1041 , n320778 , n320779 );
buf ( n320781 , n1041 );
buf ( n320782 , n320781 );
not ( n320783 , n320782 );
buf ( n320784 , n320476 );
not ( n1046 , n320784 );
or ( n320786 , n320783 , n1046 );
buf ( n320787 , n320483 );
buf ( n320788 , n320469 );
nand ( n320789 , n320787 , n320788 );
buf ( n320790 , n320789 );
buf ( n320791 , n320790 );
nand ( n1053 , n320786 , n320791 );
buf ( n320793 , n1053 );
nand ( n320794 , n320777 , n320793 );
buf ( n320795 , n320794 );
nand ( n320796 , n320776 , n320795 );
buf ( n320797 , n320796 );
buf ( n320798 , n320797 );
xor ( n320799 , n320680 , n320711 );
and ( n320800 , n320799 , n320750 );
and ( n1062 , n320680 , n320711 );
or ( n320802 , n320800 , n1062 );
buf ( n320803 , n320802 );
buf ( n320804 , n320803 );
xor ( n320805 , n320798 , n320804 );
buf ( n320806 , n320704 );
not ( n320807 , n320806 );
buf ( n320808 , n320692 );
not ( n1070 , n320808 );
or ( n1071 , n320807 , n1070 );
buf ( n1072 , n320699 );
buf ( n320812 , n557 );
buf ( n320813 , n586 );
xor ( n320814 , n320812 , n320813 );
buf ( n320815 , n320814 );
buf ( n1077 , n320815 );
nand ( n1078 , n1072 , n1077 );
buf ( n1079 , n1078 );
buf ( n320819 , n1079 );
nand ( n1081 , n1071 , n320819 );
buf ( n1082 , n1081 );
buf ( n320822 , n1082 );
and ( n1084 , n320728 , n320747 );
buf ( n320824 , n1084 );
buf ( n1086 , n320824 );
buf ( n320826 , n1086 );
xor ( n1088 , n320822 , n320826 );
xor ( n1089 , n585 , n586 );
and ( n1090 , n559 , n1089 );
buf ( n320830 , n1090 );
not ( n320831 , n1003 );
not ( n1093 , n320732 );
or ( n1094 , n320831 , n1093 );
and ( n1095 , n553 , n590 );
not ( n1096 , n553 );
not ( n1097 , n590 );
and ( n320837 , n1096 , n1097 );
nor ( n320838 , n1095 , n320837 );
nand ( n320839 , n320838 , n591 );
nand ( n1101 , n1094 , n320839 );
buf ( n320841 , n1101 );
xor ( n320842 , n320830 , n320841 );
buf ( n1104 , n320673 );
not ( n1105 , n1104 );
buf ( n320845 , n926 );
not ( n1107 , n320845 );
or ( n320847 , n1105 , n1107 );
buf ( n320848 , n320642 );
buf ( n320849 , n555 );
buf ( n320850 , n588 );
xor ( n1112 , n320849 , n320850 );
buf ( n320852 , n1112 );
buf ( n320853 , n320852 );
nand ( n320854 , n320848 , n320853 );
buf ( n320855 , n320854 );
buf ( n320856 , n320855 );
nand ( n320857 , n320847 , n320856 );
buf ( n320858 , n320857 );
buf ( n320859 , n320858 );
xor ( n320860 , n320842 , n320859 );
buf ( n320861 , n320860 );
buf ( n320862 , n320861 );
xor ( n320863 , n1088 , n320862 );
buf ( n320864 , n320863 );
buf ( n320865 , n320864 );
xor ( n320866 , n320805 , n320865 );
buf ( n320867 , n320866 );
buf ( n320868 , n320867 );
xor ( n1130 , n1020 , n320868 );
buf ( n320870 , n1130 );
buf ( n320871 , n320870 );
not ( n320872 , n320871 );
not ( n1134 , n320793 );
not ( n320874 , n1034 );
or ( n320875 , n1134 , n320874 );
or ( n1137 , n320793 , n1034 );
nand ( n320877 , n320875 , n1137 );
buf ( n320878 , n320877 );
buf ( n320879 , n1031 );
not ( n1141 , n320879 );
buf ( n320881 , n1141 );
buf ( n320882 , n320881 );
and ( n320883 , n320878 , n320882 );
not ( n1145 , n320878 );
buf ( n320885 , n1031 );
buf ( n320886 , n320885 );
and ( n320887 , n1145 , n320886 );
nor ( n1149 , n320883 , n320887 );
buf ( n320889 , n1149 );
buf ( n1151 , n320889 );
xor ( n320891 , n574 , n557 );
buf ( n320892 , n320891 );
not ( n1154 , n320892 );
buf ( n320894 , n320441 );
not ( n320895 , n320894 );
or ( n1157 , n1154 , n320895 );
buf ( n320897 , n320560 );
buf ( n320898 , n575 );
nand ( n1160 , n320897 , n320898 );
buf ( n1161 , n1160 );
buf ( n320901 , n1161 );
nand ( n320902 , n1157 , n320901 );
buf ( n320903 , n320902 );
buf ( n320904 , n320903 );
buf ( n320905 , n559 );
buf ( n320906 , n573 );
or ( n1168 , n320905 , n320906 );
buf ( n320908 , n574 );
nand ( n1170 , n1168 , n320908 );
buf ( n320910 , n1170 );
buf ( n320911 , n320910 );
buf ( n320912 , n559 );
buf ( n320913 , n573 );
nand ( n1175 , n320912 , n320913 );
buf ( n320915 , n1175 );
buf ( n320916 , n320915 );
buf ( n320917 , n572 );
nand ( n1179 , n320911 , n320916 , n320917 );
buf ( n320919 , n1179 );
buf ( n1181 , n320919 );
not ( n320921 , n1181 );
buf ( n320922 , n320921 );
buf ( n320923 , n320922 );
and ( n320924 , n320904 , n320923 );
buf ( n320925 , n320924 );
buf ( n320926 , n320925 );
or ( n320927 , n559 , n589 );
nand ( n320928 , n320927 , n590 );
buf ( n320929 , n559 );
buf ( n320930 , n589 );
nand ( n320931 , n320929 , n320930 );
buf ( n320932 , n320931 );
and ( n320933 , n320928 , n320932 , n588 );
and ( n1195 , n557 , n320740 );
not ( n320935 , n557 );
and ( n1197 , n320935 , n590 );
or ( n1198 , n1195 , n1197 );
not ( n1199 , n1198 );
not ( n1200 , n873 );
or ( n320940 , n1199 , n1200 );
buf ( n320941 , n591 );
buf ( n320942 , n320608 );
nand ( n1204 , n320941 , n320942 );
buf ( n320944 , n1204 );
nand ( n320945 , n320940 , n320944 );
and ( n320946 , n320933 , n320945 );
buf ( n320947 , n320946 );
xor ( n320948 , n320926 , n320947 );
xor ( n320949 , n320604 , n320627 );
xor ( n1211 , n320949 , n320654 );
buf ( n320951 , n1211 );
buf ( n320952 , n320951 );
and ( n1214 , n320948 , n320952 );
and ( n1215 , n320926 , n320947 );
or ( n1216 , n1214 , n1215 );
buf ( n320956 , n1216 );
buf ( n320957 , n320956 );
xor ( n1219 , n1151 , n320957 );
xor ( n1220 , n858 , n320659 );
xor ( n1221 , n1220 , n320753 );
buf ( n320961 , n1221 );
buf ( n320962 , n320961 );
and ( n320963 , n1219 , n320962 );
and ( n320964 , n1151 , n320957 );
or ( n1226 , n320963 , n320964 );
buf ( n320966 , n1226 );
buf ( n320967 , n320966 );
not ( n1229 , n320967 );
buf ( n320969 , n1229 );
buf ( n320970 , n320969 );
nand ( n1232 , n320872 , n320970 );
buf ( n320972 , n1232 );
not ( n1234 , n320972 );
xor ( n320974 , n320551 , n1019 );
and ( n320975 , n320974 , n320868 );
and ( n320976 , n320551 , n1019 );
or ( n320977 , n320975 , n320976 );
buf ( n320978 , n320977 );
buf ( n320979 , n320978 );
xor ( n320980 , n320798 , n320804 );
and ( n1242 , n320980 , n320865 );
and ( n1243 , n320798 , n320804 );
or ( n320983 , n1242 , n1243 );
buf ( n320984 , n320983 );
not ( n1246 , n320984 );
nand ( n320986 , n320441 , n320514 );
not ( n320987 , n552 );
not ( n1249 , n320509 );
or ( n320989 , n320987 , n1249 );
not ( n320990 , n552 );
nand ( n1252 , n320990 , n574 );
nand ( n320992 , n320989 , n1252 );
nand ( n320993 , n320992 , n575 );
nand ( n320994 , n320986 , n320993 );
buf ( n320995 , n320994 );
not ( n1257 , n320995 );
buf ( n320997 , n559 );
buf ( n320998 , n569 );
or ( n1260 , n320997 , n320998 );
buf ( n321000 , n570 );
nand ( n1262 , n1260 , n321000 );
buf ( n1263 , n1262 );
buf ( n321003 , n1263 );
buf ( n321004 , n559 );
buf ( n321005 , n569 );
nand ( n321006 , n321004 , n321005 );
buf ( n321007 , n321006 );
buf ( n1269 , n321007 );
buf ( n321009 , n568 );
nand ( n321010 , n321003 , n1269 , n321009 );
buf ( n321011 , n321010 );
buf ( n321012 , n321011 );
not ( n321013 , n321012 );
and ( n321014 , n1257 , n321013 );
buf ( n321015 , n320994 );
buf ( n321016 , n321011 );
and ( n321017 , n321015 , n321016 );
nor ( n1279 , n321014 , n321017 );
buf ( n321019 , n1279 );
xor ( n1281 , n320504 , n320517 );
and ( n321021 , n1281 , n320547 );
and ( n321022 , n320504 , n320517 );
or ( n1284 , n321021 , n321022 );
buf ( n321024 , n1284 );
xor ( n1286 , n321019 , n321024 );
buf ( n321026 , n1286 );
not ( n321027 , n321026 );
buf ( n321028 , n321027 );
not ( n1290 , n321028 );
not ( n1291 , n320488 );
not ( n321031 , n320472 );
nor ( n321032 , n320474 , n321031 );
not ( n1294 , n321032 );
or ( n321034 , n1291 , n1294 );
buf ( n321035 , n320480 );
buf ( n321036 , n556 );
buf ( n321037 , n570 );
xor ( n321038 , n321036 , n321037 );
buf ( n321039 , n321038 );
buf ( n1301 , n321039 );
nand ( n1302 , n321035 , n1301 );
buf ( n1303 , n1302 );
nand ( n321043 , n321034 , n1303 );
not ( n1305 , n321043 );
not ( n321045 , n1023 );
not ( n1307 , n320540 );
or ( n321047 , n321045 , n1307 );
buf ( n321048 , n1026 );
buf ( n321049 , n554 );
buf ( n321050 , n572 );
xor ( n1312 , n321049 , n321050 );
buf ( n321052 , n1312 );
buf ( n1314 , n321052 );
nand ( n1315 , n321048 , n1314 );
buf ( n1316 , n1315 );
nand ( n321056 , n321047 , n1316 );
xor ( n1318 , n1305 , n321056 );
buf ( n321058 , n559 );
buf ( n321059 , n568 );
xor ( n321060 , n321058 , n321059 );
buf ( n321061 , n321060 );
buf ( n321062 , n321061 );
not ( n321063 , n321062 );
not ( n321064 , n320496 );
xor ( n1326 , n568 , n569 );
nand ( n321066 , n321064 , n1326 );
buf ( n1328 , n321066 );
not ( n321068 , n1328 );
buf ( n321069 , n321068 );
buf ( n321070 , n321069 );
buf ( n1332 , n321070 );
buf ( n321072 , n1332 );
buf ( n321073 , n321072 );
not ( n1335 , n321073 );
or ( n321075 , n321063 , n1335 );
buf ( n1337 , n320496 );
buf ( n1338 , n1337 );
buf ( n1339 , n1338 );
buf ( n321079 , n1339 );
buf ( n321080 , n558 );
buf ( n321081 , n568 );
xor ( n321082 , n321080 , n321081 );
buf ( n321083 , n321082 );
buf ( n321084 , n321083 );
nand ( n1346 , n321079 , n321084 );
buf ( n321086 , n1346 );
buf ( n321087 , n321086 );
nand ( n1349 , n321075 , n321087 );
buf ( n321089 , n1349 );
buf ( n321090 , n321089 );
buf ( n1352 , n321090 );
buf ( n321092 , n1352 );
xnor ( n1354 , n1318 , n321092 );
buf ( n321094 , n1354 );
not ( n321095 , n321094 );
buf ( n321096 , n321095 );
not ( n321097 , n321096 );
or ( n321098 , n1290 , n321097 );
nand ( n1360 , n1286 , n1354 );
nand ( n321100 , n321098 , n1360 );
not ( n321101 , n321100 );
not ( n1363 , n321101 );
or ( n1364 , n1246 , n1363 );
not ( n321104 , n320984 );
nand ( n321105 , n321100 , n321104 );
nand ( n1367 , n1364 , n321105 );
xor ( n321107 , n320822 , n320826 );
and ( n321108 , n321107 , n320862 );
and ( n1370 , n320822 , n320826 );
or ( n321110 , n321108 , n1370 );
buf ( n321111 , n321110 );
not ( n1373 , n320549 );
not ( n1374 , n320494 );
nand ( n321114 , n1374 , n320465 );
not ( n1376 , n321114 );
or ( n321116 , n1373 , n1376 );
not ( n1378 , n320465 );
nand ( n1379 , n1378 , n320494 );
nand ( n321119 , n321116 , n1379 );
xor ( n321120 , n321111 , n321119 );
buf ( n321121 , n559 );
buf ( n321122 , n585 );
or ( n321123 , n321121 , n321122 );
buf ( n321124 , n586 );
nand ( n1386 , n321123 , n321124 );
buf ( n321126 , n1386 );
buf ( n321127 , n559 );
buf ( n321128 , n585 );
nand ( n1390 , n321127 , n321128 );
buf ( n321130 , n1390 );
and ( n321131 , n321126 , n321130 , n584 );
buf ( n321132 , n320838 );
not ( n321133 , n321132 );
buf ( n321134 , n320732 );
not ( n1396 , n321134 );
or ( n321136 , n321133 , n1396 );
and ( n1398 , n590 , n552 );
not ( n1399 , n590 );
and ( n321139 , n1399 , n320990 );
nor ( n321140 , n1398 , n321139 );
buf ( n321141 , n321140 );
buf ( n321142 , n591 );
nand ( n321143 , n321141 , n321142 );
buf ( n321144 , n321143 );
buf ( n321145 , n321144 );
nand ( n1407 , n321136 , n321145 );
buf ( n321147 , n1407 );
xor ( n321148 , n321131 , n321147 );
xor ( n321149 , n320830 , n320841 );
and ( n1411 , n321149 , n320859 );
and ( n321151 , n320830 , n320841 );
or ( n321152 , n1411 , n321151 );
buf ( n321153 , n321152 );
xor ( n321154 , n321148 , n321153 );
buf ( n321155 , n320852 );
not ( n1417 , n321155 );
buf ( n321157 , n898 );
not ( n321158 , n321157 );
or ( n1420 , n1417 , n321158 );
buf ( n1421 , n320642 );
buf ( n321161 , n554 );
buf ( n321162 , n588 );
xor ( n321163 , n321161 , n321162 );
buf ( n321164 , n321163 );
buf ( n321165 , n321164 );
nand ( n321166 , n1421 , n321165 );
buf ( n321167 , n321166 );
buf ( n321168 , n321167 );
nand ( n1430 , n1420 , n321168 );
buf ( n321170 , n1430 );
buf ( n321171 , n320815 );
not ( n1433 , n321171 );
buf ( n321173 , n320692 );
not ( n321174 , n321173 );
or ( n1436 , n1433 , n321174 );
buf ( n321176 , n320699 );
buf ( n321177 , n556 );
buf ( n321178 , n586 );
xor ( n1440 , n321177 , n321178 );
buf ( n1441 , n1440 );
buf ( n321181 , n1441 );
nand ( n1443 , n321176 , n321181 );
buf ( n321183 , n1443 );
buf ( n321184 , n321183 );
nand ( n321185 , n1436 , n321184 );
buf ( n321186 , n321185 );
xor ( n1448 , n321170 , n321186 );
buf ( n321188 , n559 );
buf ( n321189 , n584 );
xor ( n1451 , n321188 , n321189 );
buf ( n321191 , n1451 );
buf ( n321192 , n321191 );
not ( n1454 , n321192 );
not ( n321194 , n1089 );
not ( n321195 , n584 );
not ( n1457 , n585 );
not ( n321197 , n1457 );
or ( n321198 , n321195 , n321197 );
not ( n321199 , n584 );
nand ( n321200 , n321199 , n585 );
nand ( n1462 , n321198 , n321200 );
nand ( n321202 , n321194 , n1462 );
not ( n321203 , n321202 );
buf ( n321204 , n321203 );
not ( n1466 , n321204 );
or ( n321206 , n1454 , n1466 );
not ( n321207 , n1089 );
not ( n1469 , n321207 );
buf ( n321209 , n1469 );
buf ( n1471 , n321209 );
buf ( n1472 , n558 );
buf ( n1473 , n584 );
xor ( n1474 , n1472 , n1473 );
buf ( n1475 , n1474 );
buf ( n321215 , n1475 );
nand ( n321216 , n1471 , n321215 );
buf ( n321217 , n321216 );
buf ( n321218 , n321217 );
nand ( n321219 , n321206 , n321218 );
buf ( n321220 , n321219 );
xor ( n321221 , n1448 , n321220 );
xor ( n321222 , n321154 , n321221 );
xor ( n1484 , n321120 , n321222 );
and ( n321224 , n1367 , n1484 );
not ( n321225 , n1367 );
not ( n1487 , n1484 );
and ( n321227 , n321225 , n1487 );
nor ( n1489 , n321224 , n321227 );
buf ( n321229 , n1489 );
nor ( n321230 , n320979 , n321229 );
buf ( n321231 , n321230 );
nor ( n321232 , n1234 , n321231 );
not ( n1494 , n321232 );
xor ( n1495 , n320556 , n320573 );
xor ( n321235 , n1495 , n320592 );
buf ( n321236 , n321235 );
buf ( n321237 , n321236 );
buf ( n321238 , n559 );
buf ( n321239 , n588 );
xor ( n1501 , n321238 , n321239 );
buf ( n1502 , n1501 );
buf ( n321242 , n1502 );
not ( n1504 , n321242 );
buf ( n321244 , n898 );
not ( n321245 , n321244 );
or ( n321246 , n1504 , n321245 );
buf ( n321247 , n320642 );
buf ( n321248 , n893 );
nand ( n321249 , n321247 , n321248 );
buf ( n321250 , n321249 );
buf ( n321251 , n321250 );
nand ( n321252 , n321246 , n321251 );
buf ( n321253 , n321252 );
buf ( n321254 , n321253 );
xor ( n1516 , n572 , n559 );
buf ( n321256 , n1516 );
not ( n1518 , n321256 );
buf ( n321258 , n1023 );
not ( n321259 , n321258 );
or ( n321260 , n1518 , n321259 );
buf ( n321261 , n320535 );
buf ( n321262 , n320575 );
nand ( n321263 , n321261 , n321262 );
buf ( n321264 , n321263 );
buf ( n321265 , n321264 );
nand ( n321266 , n321260 , n321265 );
buf ( n321267 , n321266 );
buf ( n321268 , n321267 );
buf ( n1530 , n321268 );
buf ( n1531 , n1530 );
buf ( n321271 , n1531 );
or ( n1533 , n321254 , n321271 );
xor ( n321273 , n320933 , n320945 );
buf ( n321274 , n321273 );
nand ( n321275 , n1533 , n321274 );
buf ( n321276 , n321275 );
buf ( n321277 , n321276 );
buf ( n321278 , n1531 );
buf ( n321279 , n321253 );
nand ( n1541 , n321278 , n321279 );
buf ( n1542 , n1541 );
buf ( n1543 , n1542 );
nand ( n1544 , n321277 , n1543 );
buf ( n1545 , n1544 );
buf ( n321285 , n1545 );
xor ( n321286 , n321237 , n321285 );
xor ( n1548 , n320926 , n320947 );
xor ( n321288 , n1548 , n320952 );
buf ( n321289 , n321288 );
buf ( n321290 , n321289 );
and ( n321291 , n321286 , n321290 );
and ( n321292 , n321237 , n321285 );
or ( n1554 , n321291 , n321292 );
buf ( n321294 , n1554 );
buf ( n321295 , n321294 );
not ( n1557 , n321295 );
buf ( n1558 , n1557 );
not ( n321298 , n1558 );
xor ( n1560 , n1151 , n320957 );
xor ( n321300 , n1560 , n320962 );
buf ( n321301 , n321300 );
buf ( n321302 , n321301 );
not ( n321303 , n321302 );
buf ( n321304 , n321303 );
not ( n321305 , n321304 );
or ( n1567 , n321298 , n321305 );
xor ( n1568 , n321237 , n321285 );
xor ( n1569 , n1568 , n321290 );
buf ( n321309 , n1569 );
buf ( n321310 , n320903 );
buf ( n321311 , n320922 );
and ( n321312 , n321310 , n321311 );
not ( n1574 , n321310 );
buf ( n321314 , n320919 );
and ( n1576 , n1574 , n321314 );
nor ( n1577 , n321312 , n1576 );
buf ( n321317 , n1577 );
buf ( n321318 , n321317 );
not ( n1580 , n321318 );
buf ( n321320 , n558 );
buf ( n321321 , n590 );
xor ( n321322 , n321320 , n321321 );
buf ( n321323 , n321322 );
buf ( n321324 , n321323 );
not ( n321325 , n321324 );
buf ( n321326 , n873 );
not ( n1588 , n321326 );
or ( n321328 , n321325 , n1588 );
buf ( n321329 , n1198 );
buf ( n321330 , n591 );
nand ( n321331 , n321329 , n321330 );
buf ( n321332 , n321331 );
buf ( n321333 , n321332 );
nand ( n1595 , n321328 , n321333 );
buf ( n321335 , n1595 );
buf ( n321336 , n321335 );
buf ( n321337 , n1026 );
buf ( n321338 , n559 );
and ( n1600 , n321337 , n321338 );
buf ( n321340 , n1600 );
buf ( n321341 , n321340 );
nand ( n1603 , n321336 , n321341 );
buf ( n321343 , n1603 );
buf ( n321344 , n321343 );
nand ( n1606 , n1580 , n321344 );
buf ( n321346 , n1606 );
buf ( n321347 , n321346 );
not ( n1609 , n321347 );
buf ( n321349 , n321267 );
not ( n1611 , n321349 );
buf ( n321351 , n1611 );
buf ( n321352 , n321351 );
buf ( n321353 , n321273 );
and ( n1615 , n321352 , n321353 );
not ( n1616 , n321352 );
buf ( n321356 , n321273 );
not ( n1618 , n321356 );
buf ( n321358 , n1618 );
buf ( n321359 , n321358 );
and ( n1621 , n1616 , n321359 );
nor ( n1622 , n1615 , n1621 );
buf ( n321362 , n1622 );
buf ( n321363 , n321362 );
buf ( n321364 , n321253 );
and ( n1626 , n321363 , n321364 );
not ( n1627 , n321363 );
buf ( n321367 , n321253 );
not ( n1629 , n321367 );
buf ( n321369 , n1629 );
buf ( n321370 , n321369 );
and ( n1632 , n1627 , n321370 );
nor ( n1633 , n1626 , n1632 );
buf ( n321373 , n1633 );
buf ( n321374 , n321373 );
not ( n1636 , n321374 );
buf ( n321376 , n1636 );
buf ( n321377 , n321376 );
not ( n1639 , n321377 );
or ( n1640 , n1609 , n1639 );
buf ( n321380 , n321343 );
not ( n1642 , n321380 );
buf ( n321382 , n321317 );
nand ( n1644 , n1642 , n321382 );
buf ( n321384 , n1644 );
buf ( n321385 , n321384 );
nand ( n1647 , n1640 , n321385 );
buf ( n321387 , n1647 );
nand ( n1649 , n321309 , n321387 );
not ( n1650 , n1649 );
nand ( n1651 , n1567 , n1650 );
buf ( n321391 , n321301 );
buf ( n321392 , n321294 );
nand ( n1654 , n321391 , n321392 );
buf ( n321394 , n1654 );
nand ( n1656 , n1651 , n321394 );
not ( n1657 , n1656 );
xnor ( n1658 , n321343 , n321317 );
buf ( n321398 , n1658 );
not ( n1660 , n321398 );
buf ( n321400 , n1660 );
buf ( n321401 , n321400 );
not ( n1663 , n321401 );
buf ( n321403 , n321373 );
not ( n1665 , n321403 );
buf ( n321405 , n1665 );
buf ( n321406 , n321405 );
not ( n1668 , n321406 );
or ( n1669 , n1663 , n1668 );
buf ( n321409 , n321373 );
buf ( n321410 , n1658 );
nand ( n1672 , n321409 , n321410 );
buf ( n321412 , n1672 );
buf ( n321413 , n321412 );
nand ( n1675 , n1669 , n321413 );
buf ( n321415 , n1675 );
buf ( n321416 , n320441 );
not ( n1678 , n321416 );
and ( n1679 , n574 , n558 );
not ( n1680 , n574 );
not ( n1681 , n558 );
and ( n1682 , n1680 , n1681 );
nor ( n1683 , n1679 , n1682 );
buf ( n321423 , n1683 );
not ( n1685 , n321423 );
or ( n1686 , n1678 , n1685 );
buf ( n321426 , n575 );
buf ( n321427 , n320891 );
nand ( n1689 , n321426 , n321427 );
buf ( n321429 , n1689 );
buf ( n321430 , n321429 );
nand ( n1692 , n1686 , n321430 );
buf ( n321432 , n1692 );
not ( n1694 , n321432 );
buf ( n321434 , n320642 );
buf ( n321435 , n559 );
and ( n1697 , n321434 , n321435 );
buf ( n321437 , n1697 );
not ( n1699 , n321437 );
nand ( n1700 , n1694 , n1699 );
not ( n1701 , n1700 );
xor ( n1702 , n321340 , n321335 );
not ( n1703 , n1702 );
or ( n1704 , n1701 , n1703 );
nand ( n1705 , n321437 , n321432 );
nand ( n1706 , n1704 , n1705 );
nand ( n1707 , n321415 , n1706 );
buf ( n321447 , n1707 );
not ( n1709 , n321447 );
buf ( n321449 , n1709 );
not ( n1711 , n321449 );
buf ( n321451 , n559 );
buf ( n321452 , n591 );
nand ( n1714 , n321451 , n321452 );
buf ( n321454 , n1714 );
buf ( n321455 , n321454 );
buf ( n321456 , n590 );
and ( n1718 , n321455 , n321456 );
buf ( n321458 , n1718 );
buf ( n321459 , n321458 );
buf ( n321460 , n559 );
buf ( n321461 , n575 );
nand ( n1723 , n321460 , n321461 );
buf ( n321463 , n1723 );
buf ( n321464 , n321463 );
buf ( n321465 , n574 );
and ( n1727 , n321464 , n321465 );
buf ( n321467 , n1727 );
buf ( n321468 , n321467 );
or ( n1730 , n321459 , n321468 );
buf ( n321470 , n1730 );
not ( n1732 , n321470 );
not ( n1733 , n591 );
not ( n1734 , n321323 );
or ( n1735 , n1733 , n1734 );
not ( n1736 , n559 );
nand ( n1737 , n1736 , n873 );
nand ( n1738 , n1735 , n1737 );
not ( n1739 , n1738 );
or ( n1740 , n1732 , n1739 );
buf ( n321480 , n321467 );
buf ( n321481 , n321458 );
nand ( n1743 , n321480 , n321481 );
buf ( n321483 , n1743 );
nand ( n1745 , n1740 , n321483 );
xor ( n1746 , n321432 , n1699 );
xnor ( n1747 , n1746 , n1702 );
nand ( n1748 , n1745 , n1747 );
buf ( n321488 , n1748 );
not ( n1750 , n321488 );
buf ( n321490 , n1750 );
buf ( n321491 , n559 );
buf ( n321492 , n575 );
and ( n1754 , n321491 , n321492 );
buf ( n321494 , n1754 );
buf ( n321495 , n321494 );
buf ( n321496 , n559 );
buf ( n321497 , n591 );
and ( n1759 , n321496 , n321497 );
buf ( n321499 , n1759 );
buf ( n321500 , n321499 );
and ( n1762 , n321495 , n321500 );
buf ( n321502 , n1762 );
not ( n1764 , n321502 );
not ( n1765 , n575 );
not ( n1766 , n1683 );
or ( n1767 , n1765 , n1766 );
not ( n1768 , n559 );
not ( n1769 , n575 );
nand ( n1770 , n1768 , n1769 , n574 );
nand ( n1771 , n1767 , n1770 );
not ( n1772 , n1771 );
nand ( n1773 , n1764 , n1772 );
not ( n1774 , n1773 );
xor ( n1775 , n321467 , n321458 );
xor ( n1776 , n1775 , n1738 );
not ( n1777 , n1776 );
or ( n1778 , n1774 , n1777 );
nand ( n1779 , n321502 , n1771 );
nand ( n1780 , n1778 , n1779 );
buf ( n321520 , n1780 );
not ( n1782 , n321520 );
buf ( n321522 , n1747 );
buf ( n321523 , n1745 );
nor ( n1785 , n321522 , n321523 );
buf ( n321525 , n1785 );
buf ( n321526 , n321525 );
nor ( n1788 , n1782 , n321526 );
buf ( n321528 , n1788 );
or ( n1790 , n321490 , n321528 );
buf ( n321530 , n321415 );
not ( n1792 , n321530 );
buf ( n321532 , n1792 );
buf ( n321533 , n1706 );
not ( n1795 , n321533 );
buf ( n321535 , n1795 );
nand ( n1797 , n321532 , n321535 );
nand ( n1798 , n1790 , n1797 );
nand ( n1799 , n1711 , n1798 );
buf ( n321539 , n1799 );
buf ( n1801 , n321539 );
buf ( n321541 , n1801 );
buf ( n321542 , n321301 );
buf ( n321543 , n321294 );
nor ( n1805 , n321542 , n321543 );
buf ( n321545 , n1805 );
not ( n1807 , n321545 );
buf ( n321547 , n321309 );
not ( n1809 , n321547 );
buf ( n321549 , n1809 );
buf ( n321550 , n321549 );
buf ( n321551 , n321387 );
not ( n1813 , n321551 );
buf ( n321553 , n1813 );
buf ( n321554 , n321553 );
nand ( n1816 , n321550 , n321554 );
buf ( n321556 , n1816 );
nand ( n1818 , n321541 , n1807 , n321556 );
nand ( n1819 , n1657 , n1818 );
not ( n1820 , n1819 );
or ( n1821 , n1494 , n1820 );
buf ( n321561 , n320870 );
buf ( n1823 , n321561 );
buf ( n321563 , n1823 );
buf ( n1825 , n320966 );
nand ( n1826 , n321563 , n1825 );
not ( n1827 , n1826 );
not ( n1828 , n321231 );
and ( n1829 , n1827 , n1828 );
and ( n1830 , n1489 , n320978 );
nor ( n1831 , n1829 , n1830 );
nand ( n1832 , n1821 , n1831 );
not ( n1833 , n1832 );
not ( n1834 , n1833 );
not ( n1835 , n1834 );
buf ( n321575 , n559 );
buf ( n321576 , n564 );
xor ( n1838 , n321575 , n321576 );
buf ( n321578 , n1838 );
buf ( n321579 , n321578 );
not ( n1841 , n321579 );
not ( n1842 , n566 );
not ( n1843 , n1842 );
not ( n1844 , n564 );
nor ( n1845 , n1844 , n565 );
not ( n1846 , n1845 );
or ( n1847 , n1843 , n1846 );
not ( n1848 , n564 );
nand ( n1849 , n1848 , n566 , n565 );
nand ( n1850 , n1847 , n1849 );
buf ( n321590 , n1850 );
buf ( n1852 , n321590 );
buf ( n321592 , n1852 );
buf ( n321593 , n321592 );
not ( n1855 , n321593 );
or ( n1856 , n1841 , n1855 );
xor ( n1857 , n565 , n566 );
buf ( n321597 , n1857 );
buf ( n321598 , n558 );
buf ( n321599 , n564 );
xor ( n1861 , n321598 , n321599 );
buf ( n321601 , n1861 );
buf ( n321602 , n321601 );
nand ( n1864 , n321597 , n321602 );
buf ( n321604 , n1864 );
buf ( n321605 , n321604 );
nand ( n1867 , n1856 , n321605 );
buf ( n321607 , n1867 );
buf ( n321608 , n321607 );
buf ( n321609 , n553 );
buf ( n321610 , n570 );
xor ( n1872 , n321609 , n321610 );
buf ( n321612 , n1872 );
buf ( n321613 , n321612 );
not ( n1875 , n321613 );
buf ( n321615 , n320476 );
not ( n1877 , n321615 );
or ( n1878 , n1875 , n1877 );
buf ( n321618 , n320483 );
buf ( n321619 , n552 );
buf ( n321620 , n570 );
xor ( n1882 , n321619 , n321620 );
buf ( n321622 , n1882 );
buf ( n321623 , n321622 );
nand ( n1885 , n321618 , n321623 );
buf ( n321625 , n1885 );
buf ( n321626 , n321625 );
nand ( n1888 , n1878 , n321626 );
buf ( n321628 , n1888 );
buf ( n321629 , n321628 );
xor ( n1891 , n321608 , n321629 );
buf ( n321631 , n551 );
buf ( n321632 , n572 );
xor ( n1894 , n321631 , n321632 );
buf ( n321634 , n1894 );
buf ( n321635 , n321634 );
not ( n321636 , n321635 );
buf ( n321637 , n320531 );
not ( n321638 , n321637 );
or ( n321639 , n321636 , n321638 );
buf ( n321640 , n320535 );
buf ( n321641 , n550 );
buf ( n321642 , n572 );
xor ( n321643 , n321641 , n321642 );
buf ( n321644 , n321643 );
buf ( n321645 , n321644 );
nand ( n321646 , n321640 , n321645 );
buf ( n321647 , n321646 );
buf ( n321648 , n321647 );
nand ( n321649 , n321639 , n321648 );
buf ( n321650 , n321649 );
buf ( n321651 , n559 );
buf ( n321652 , n565 );
or ( n321653 , n321651 , n321652 );
buf ( n321654 , n566 );
nand ( n321655 , n321653 , n321654 );
buf ( n321656 , n321655 );
buf ( n321657 , n321656 );
buf ( n321658 , n559 );
buf ( n321659 , n565 );
nand ( n321660 , n321658 , n321659 );
buf ( n321661 , n321660 );
buf ( n321662 , n321661 );
buf ( n321663 , n564 );
nand ( n321664 , n321657 , n321662 , n321663 );
buf ( n321665 , n321664 );
xnor ( n321666 , n321650 , n321665 );
buf ( n321667 , n321666 );
xor ( n321668 , n1891 , n321667 );
buf ( n321669 , n321668 );
buf ( n321670 , n321669 );
buf ( n321671 , n559 );
buf ( n321672 , n567 );
or ( n321673 , n321671 , n321672 );
buf ( n321674 , n568 );
nand ( n321675 , n321673 , n321674 );
buf ( n321676 , n321675 );
buf ( n1900 , n321676 );
buf ( n321678 , n559 );
buf ( n321679 , n567 );
nand ( n321680 , n321678 , n321679 );
buf ( n321681 , n321680 );
buf ( n321682 , n321681 );
buf ( n321683 , n566 );
and ( n321684 , n1900 , n321682 , n321683 );
buf ( n321685 , n321684 );
buf ( n321686 , n321685 );
buf ( n1910 , n553 );
buf ( n321688 , n572 );
xor ( n1912 , n1910 , n321688 );
buf ( n1913 , n1912 );
buf ( n321691 , n1913 );
not ( n1914 , n321691 );
buf ( n321693 , n320531 );
not ( n321694 , n321693 );
or ( n321695 , n1914 , n321694 );
buf ( n321696 , n1026 );
buf ( n321697 , n552 );
buf ( n321698 , n572 );
xor ( n321699 , n321697 , n321698 );
buf ( n321700 , n321699 );
buf ( n321701 , n321700 );
nand ( n321702 , n321696 , n321701 );
buf ( n321703 , n321702 );
buf ( n321704 , n321703 );
nand ( n321705 , n321695 , n321704 );
buf ( n321706 , n321705 );
buf ( n321707 , n321706 );
and ( n321708 , n321686 , n321707 );
buf ( n321709 , n321708 );
buf ( n321710 , n321709 );
buf ( n1929 , n550 );
buf ( n1930 , n574 );
xor ( n1931 , n1929 , n1930 );
buf ( n1932 , n1931 );
not ( n321715 , n1932 );
not ( n1934 , n575 );
or ( n1935 , n321715 , n1934 );
and ( n321718 , n551 , n574 );
not ( n1937 , n551 );
and ( n321720 , n1937 , n320509 );
nor ( n321721 , n321718 , n321720 );
nand ( n1940 , n321721 , n320441 );
nand ( n1941 , n1935 , n1940 );
not ( n321724 , n1941 );
xor ( n1943 , n568 , n557 );
buf ( n321726 , n1943 );
not ( n1945 , n321726 );
buf ( n321728 , n321069 );
not ( n1947 , n321728 );
or ( n1948 , n1945 , n1947 );
buf ( n321731 , n1339 );
buf ( n321732 , n556 );
buf ( n321733 , n568 );
xor ( n1952 , n321732 , n321733 );
buf ( n321735 , n1952 );
buf ( n321736 , n321735 );
nand ( n1955 , n321731 , n321736 );
buf ( n321738 , n1955 );
buf ( n321739 , n321738 );
nand ( n1958 , n1948 , n321739 );
buf ( n321741 , n1958 );
not ( n1960 , n321741 );
or ( n1961 , n321724 , n1960 );
or ( n1962 , n321741 , n1941 );
buf ( n321745 , n559 );
buf ( n321746 , n566 );
xor ( n1965 , n321745 , n321746 );
buf ( n321748 , n1965 );
not ( n1967 , n321748 );
not ( n321750 , n566 );
nor ( n321751 , n567 , n568 );
not ( n1970 , n321751 );
or ( n321753 , n321750 , n1970 );
not ( n1972 , n566 );
nand ( n321755 , n1972 , n567 , n568 );
nand ( n321756 , n321753 , n321755 );
buf ( n1975 , n321756 );
not ( n1976 , n1975 );
or ( n321759 , n1967 , n1976 );
buf ( n321760 , n558 );
buf ( n321761 , n566 );
xor ( n321762 , n321760 , n321761 );
buf ( n321763 , n321762 );
buf ( n321764 , n321763 );
buf ( n1983 , n567 );
buf ( n321766 , n568 );
xor ( n321767 , n1983 , n321766 );
buf ( n321768 , n321767 );
buf ( n321769 , n321768 );
buf ( n321770 , n321769 );
buf ( n321771 , n321770 );
buf ( n321772 , n321771 );
nand ( n321773 , n321764 , n321772 );
buf ( n321774 , n321773 );
nand ( n321775 , n321759 , n321774 );
nand ( n321776 , n1962 , n321775 );
nand ( n321777 , n1961 , n321776 );
buf ( n1996 , n321777 );
xor ( n1997 , n321710 , n1996 );
buf ( n321780 , n1857 );
buf ( n1999 , n559 );
and ( n2000 , n321780 , n1999 );
buf ( n321783 , n2000 );
buf ( n2002 , n321783 );
buf ( n321785 , n321735 );
not ( n2004 , n321785 );
buf ( n321787 , n321069 );
not ( n2006 , n321787 );
or ( n2007 , n2004 , n2006 );
buf ( n321790 , n320499 );
buf ( n2009 , n555 );
buf ( n2010 , n568 );
xor ( n2011 , n2009 , n2010 );
buf ( n2012 , n2011 );
buf ( n321795 , n2012 );
nand ( n321796 , n321790 , n321795 );
buf ( n321797 , n321796 );
buf ( n321798 , n321797 );
nand ( n2017 , n2007 , n321798 );
buf ( n321800 , n2017 );
buf ( n321801 , n321800 );
xor ( n2020 , n2002 , n321801 );
buf ( n321803 , n321700 );
not ( n2022 , n321803 );
buf ( n321805 , n320531 );
not ( n321806 , n321805 );
or ( n321807 , n2022 , n321806 );
buf ( n321808 , n1026 );
buf ( n321809 , n321634 );
nand ( n321810 , n321808 , n321809 );
buf ( n321811 , n321810 );
buf ( n321812 , n321811 );
nand ( n321813 , n321807 , n321812 );
buf ( n321814 , n321813 );
buf ( n321815 , n321814 );
xor ( n321816 , n2020 , n321815 );
buf ( n321817 , n321816 );
buf ( n2036 , n321817 );
and ( n2037 , n1997 , n2036 );
and ( n321820 , n321710 , n1996 );
or ( n2039 , n2037 , n321820 );
buf ( n321822 , n2039 );
buf ( n321823 , n321822 );
xor ( n2042 , n321670 , n321823 );
xor ( n2043 , n2002 , n321801 );
and ( n321826 , n2043 , n321815 );
and ( n2045 , n2002 , n321801 );
or ( n321828 , n321826 , n2045 );
buf ( n321829 , n321828 );
buf ( n321830 , n320441 );
not ( n321831 , n321830 );
buf ( n321832 , n549 );
buf ( n321833 , n574 );
xor ( n321834 , n321832 , n321833 );
buf ( n321835 , n321834 );
buf ( n321836 , n321835 );
not ( n321837 , n321836 );
or ( n2056 , n321831 , n321837 );
buf ( n321839 , n548 );
buf ( n321840 , n574 );
xor ( n2059 , n321839 , n321840 );
buf ( n321842 , n2059 );
buf ( n321843 , n321842 );
buf ( n321844 , n575 );
nand ( n2063 , n321843 , n321844 );
buf ( n321846 , n2063 );
buf ( n321847 , n321846 );
nand ( n2066 , n2056 , n321847 );
buf ( n321849 , n2066 );
buf ( n321850 , n321849 );
buf ( n321851 , n2012 );
not ( n321852 , n321851 );
buf ( n321853 , n321069 );
not ( n321854 , n321853 );
or ( n2073 , n321852 , n321854 );
buf ( n321856 , n1339 );
buf ( n321857 , n554 );
buf ( n321858 , n568 );
xor ( n321859 , n321857 , n321858 );
buf ( n321860 , n321859 );
buf ( n321861 , n321860 );
nand ( n321862 , n321856 , n321861 );
buf ( n321863 , n321862 );
buf ( n321864 , n321863 );
nand ( n321865 , n2073 , n321864 );
buf ( n321866 , n321865 );
buf ( n2085 , n321866 );
xor ( n2086 , n321850 , n2085 );
buf ( n321869 , n556 );
buf ( n321870 , n566 );
not ( n2089 , n321870 );
xor ( n321872 , n321869 , n2089 );
buf ( n321873 , n321872 );
buf ( n321874 , n321873 );
not ( n2093 , n321874 );
buf ( n321876 , n321771 );
nand ( n2095 , n2093 , n321876 );
buf ( n321878 , n2095 );
buf ( n321879 , n557 );
buf ( n321880 , n566 );
xor ( n2099 , n321879 , n321880 );
buf ( n321882 , n2099 );
and ( n321883 , n566 , n321751 );
not ( n2102 , n566 );
and ( n321885 , n567 , n568 );
and ( n2104 , n2102 , n321885 );
or ( n2105 , n321883 , n2104 );
nand ( n2106 , n321882 , n2105 );
nand ( n321889 , n321878 , n2106 );
buf ( n321890 , n321889 );
xor ( n321891 , n2086 , n321890 );
buf ( n321892 , n321891 );
xor ( n2111 , n321829 , n321892 );
buf ( n321894 , n320441 );
not ( n2113 , n321894 );
buf ( n321896 , n1932 );
not ( n321897 , n321896 );
or ( n2116 , n2113 , n321897 );
buf ( n321899 , n321835 );
buf ( n321900 , n575 );
nand ( n2119 , n321899 , n321900 );
buf ( n2120 , n2119 );
buf ( n321903 , n2120 );
nand ( n2122 , n2116 , n321903 );
buf ( n2123 , n2122 );
buf ( n321906 , n2123 );
buf ( n321907 , n554 );
buf ( n321908 , n570 );
xor ( n321909 , n321907 , n321908 );
buf ( n321910 , n321909 );
buf ( n321911 , n321910 );
not ( n321912 , n321911 );
buf ( n321913 , n320476 );
not ( n321914 , n321913 );
or ( n321915 , n321912 , n321914 );
buf ( n321916 , n320483 );
buf ( n321917 , n321612 );
nand ( n321918 , n321916 , n321917 );
buf ( n321919 , n321918 );
buf ( n321920 , n321919 );
nand ( n321921 , n321915 , n321920 );
buf ( n321922 , n321921 );
buf ( n321923 , n321922 );
xor ( n2142 , n321906 , n321923 );
buf ( n321925 , n321763 );
not ( n321926 , n321925 );
buf ( n321927 , n1975 );
not ( n321928 , n321927 );
or ( n2147 , n321926 , n321928 );
buf ( n321930 , n321771 );
buf ( n321931 , n321882 );
nand ( n2150 , n321930 , n321931 );
buf ( n321933 , n2150 );
buf ( n321934 , n321933 );
nand ( n321935 , n2147 , n321934 );
buf ( n321936 , n321935 );
buf ( n321937 , n321936 );
and ( n321938 , n2142 , n321937 );
and ( n2157 , n321906 , n321923 );
or ( n321940 , n321938 , n2157 );
buf ( n321941 , n321940 );
xor ( n2160 , n2111 , n321941 );
buf ( n321943 , n2160 );
xor ( n321944 , n2042 , n321943 );
buf ( n321945 , n321944 );
and ( n321946 , n320986 , n320993 );
nor ( n321947 , n321946 , n321011 );
buf ( n321948 , n321052 );
not ( n321949 , n321948 );
buf ( n321950 , n320531 );
not ( n2169 , n321950 );
or ( n321952 , n321949 , n2169 );
buf ( n321953 , n1026 );
buf ( n321954 , n1913 );
nand ( n321955 , n321953 , n321954 );
buf ( n321956 , n321955 );
buf ( n321957 , n321956 );
nand ( n2176 , n321952 , n321957 );
buf ( n321959 , n2176 );
or ( n2178 , n321947 , n321959 );
buf ( n321961 , n321039 );
not ( n2180 , n321961 );
buf ( n321963 , n320476 );
not ( n2182 , n321963 );
or ( n2183 , n2180 , n2182 );
buf ( n321966 , n320483 );
buf ( n321967 , n555 );
buf ( n321968 , n570 );
xor ( n321969 , n321967 , n321968 );
buf ( n321970 , n321969 );
buf ( n321971 , n321970 );
nand ( n321972 , n321966 , n321971 );
buf ( n321973 , n321972 );
buf ( n321974 , n321973 );
nand ( n2193 , n2183 , n321974 );
buf ( n321976 , n2193 );
nand ( n2195 , n2178 , n321976 );
buf ( n321978 , n2195 );
buf ( n321979 , n321011 );
not ( n2198 , n321979 );
buf ( n321981 , n320994 );
nand ( n321982 , n2198 , n321981 );
buf ( n321983 , n321982 );
buf ( n321984 , n321983 );
not ( n321985 , n321984 );
buf ( n321986 , n321985 );
buf ( n321987 , n321986 );
buf ( n321988 , n321959 );
nand ( n321989 , n321987 , n321988 );
buf ( n321990 , n321989 );
buf ( n2209 , n321990 );
nand ( n321992 , n321978 , n2209 );
buf ( n321993 , n321992 );
buf ( n321994 , n321993 );
buf ( n321995 , n321741 );
not ( n2214 , n321995 );
buf ( n321997 , n1941 );
not ( n2216 , n321997 );
buf ( n321999 , n2216 );
buf ( n322000 , n321999 );
not ( n2219 , n322000 );
and ( n2220 , n2214 , n2219 );
buf ( n322003 , n321741 );
buf ( n322004 , n321999 );
and ( n2223 , n322003 , n322004 );
nor ( n2224 , n2220 , n2223 );
buf ( n322007 , n2224 );
xnor ( n2226 , n321775 , n322007 );
buf ( n322009 , n2226 );
xor ( n2228 , n321994 , n322009 );
buf ( n322011 , n321970 );
not ( n2230 , n322011 );
buf ( n322013 , n320476 );
not ( n2232 , n322013 );
or ( n2233 , n2230 , n2232 );
buf ( n322016 , n320483 );
buf ( n322017 , n321910 );
nand ( n2236 , n322016 , n322017 );
buf ( n322019 , n2236 );
buf ( n322020 , n322019 );
nand ( n2239 , n2233 , n322020 );
buf ( n322022 , n2239 );
buf ( n322023 , n322022 );
xor ( n2242 , n321686 , n321707 );
buf ( n322025 , n2242 );
buf ( n322026 , n322025 );
xor ( n2245 , n322023 , n322026 );
nand ( n2246 , n321771 , n559 );
buf ( n322029 , n2246 );
not ( n2248 , n322029 );
not ( n2249 , n575 );
not ( n2250 , n321721 );
or ( n2251 , n2249 , n2250 );
nand ( n2252 , n320992 , n1769 , n574 );
nand ( n2253 , n2251 , n2252 );
not ( n2254 , n2253 );
buf ( n322037 , n2254 );
not ( n2256 , n322037 );
or ( n2257 , n2248 , n2256 );
buf ( n322040 , n321083 );
not ( n2259 , n322040 );
buf ( n322042 , n321069 );
not ( n2261 , n322042 );
or ( n2262 , n2259 , n2261 );
buf ( n322045 , n1339 );
buf ( n322046 , n1943 );
nand ( n2265 , n322045 , n322046 );
buf ( n322048 , n2265 );
buf ( n322049 , n322048 );
nand ( n2268 , n2262 , n322049 );
buf ( n322051 , n2268 );
buf ( n322052 , n322051 );
nand ( n2271 , n2257 , n322052 );
buf ( n322054 , n2271 );
buf ( n322055 , n322054 );
buf ( n322056 , n2253 );
not ( n2275 , n2246 );
buf ( n322058 , n2275 );
nand ( n2277 , n322056 , n322058 );
buf ( n322060 , n2277 );
buf ( n322061 , n322060 );
nand ( n2280 , n322055 , n322061 );
buf ( n322063 , n2280 );
buf ( n322064 , n322063 );
xor ( n2283 , n2245 , n322064 );
buf ( n322066 , n2283 );
buf ( n322067 , n322066 );
and ( n2286 , n2228 , n322067 );
and ( n2287 , n321994 , n322009 );
or ( n2288 , n2286 , n2287 );
buf ( n322071 , n2288 );
buf ( n322072 , n322071 );
buf ( n322073 , n321164 );
not ( n2292 , n322073 );
buf ( n322075 , n898 );
not ( n2294 , n322075 );
or ( n2295 , n2292 , n2294 );
buf ( n322078 , n320642 );
buf ( n322079 , n553 );
buf ( n322080 , n588 );
xor ( n2299 , n322079 , n322080 );
buf ( n322082 , n2299 );
buf ( n322083 , n322082 );
nand ( n2302 , n322078 , n322083 );
buf ( n322085 , n2302 );
buf ( n322086 , n322085 );
nand ( n2305 , n2295 , n322086 );
buf ( n322088 , n2305 );
buf ( n322089 , n322088 );
buf ( n322090 , n1441 );
not ( n2309 , n322090 );
buf ( n322092 , n320692 );
not ( n2311 , n322092 );
or ( n2312 , n2309 , n2311 );
buf ( n322095 , n320699 );
buf ( n322096 , n555 );
buf ( n322097 , n586 );
xor ( n2316 , n322096 , n322097 );
buf ( n322099 , n2316 );
buf ( n322100 , n322099 );
nand ( n2319 , n322095 , n322100 );
buf ( n322102 , n2319 );
buf ( n322103 , n322102 );
nand ( n322104 , n2312 , n322103 );
buf ( n322105 , n322104 );
buf ( n322106 , n322105 );
xor ( n322107 , n322089 , n322106 );
and ( n322108 , n321131 , n321147 );
buf ( n322109 , n322108 );
and ( n322110 , n322107 , n322109 );
and ( n322111 , n322089 , n322106 );
or ( n322112 , n322110 , n322111 );
buf ( n322113 , n322112 );
buf ( n322114 , n322113 );
and ( n322115 , n551 , n590 );
not ( n322116 , n551 );
and ( n322117 , n322116 , n1097 );
nor ( n322118 , n322115 , n322117 );
buf ( n322119 , n322118 );
not ( n322120 , n322119 );
buf ( n322121 , n873 );
not ( n2320 , n322121 );
or ( n322123 , n322120 , n2320 );
buf ( n322124 , n550 );
buf ( n322125 , n590 );
xor ( n322126 , n322124 , n322125 );
buf ( n322127 , n322126 );
buf ( n322128 , n322127 );
buf ( n322129 , n591 );
nand ( n2324 , n322128 , n322129 );
buf ( n322131 , n2324 );
buf ( n322132 , n322131 );
nand ( n322133 , n322123 , n322132 );
buf ( n322134 , n322133 );
buf ( n322135 , n322134 );
buf ( n322136 , n559 );
buf ( n322137 , n582 );
xor ( n322138 , n322136 , n322137 );
buf ( n322139 , n322138 );
buf ( n322140 , n322139 );
not ( n322141 , n322140 );
xnor ( n322142 , n583 , n582 );
xor ( n322143 , n583 , n584 );
nor ( n322144 , n322142 , n322143 );
not ( n322145 , n322144 );
not ( n2327 , n322145 );
buf ( n322147 , n2327 );
not ( n2329 , n322147 );
or ( n322149 , n322141 , n2329 );
not ( n2330 , n322143 );
not ( n2331 , n2330 );
buf ( n322152 , n2331 );
buf ( n322153 , n558 );
buf ( n322154 , n582 );
xor ( n2335 , n322153 , n322154 );
buf ( n322156 , n2335 );
buf ( n322157 , n322156 );
nand ( n2338 , n322152 , n322157 );
buf ( n322159 , n2338 );
buf ( n322160 , n322159 );
nand ( n322161 , n322149 , n322160 );
buf ( n322162 , n322161 );
buf ( n322163 , n322162 );
xor ( n2342 , n322135 , n322163 );
buf ( n322165 , n557 );
buf ( n322166 , n584 );
xor ( n2345 , n322165 , n322166 );
buf ( n322168 , n2345 );
buf ( n322169 , n322168 );
not ( n2347 , n322169 );
buf ( n322171 , n321202 );
buf ( n2349 , n322171 );
buf ( n322173 , n2349 );
buf ( n322174 , n322173 );
not ( n2352 , n322174 );
buf ( n322176 , n2352 );
buf ( n322177 , n322176 );
not ( n2355 , n322177 );
or ( n2356 , n2347 , n2355 );
buf ( n322180 , n321209 );
buf ( n322181 , n556 );
buf ( n322182 , n584 );
xor ( n2360 , n322181 , n322182 );
buf ( n2361 , n2360 );
buf ( n322185 , n2361 );
nand ( n2363 , n322180 , n322185 );
buf ( n2364 , n2363 );
buf ( n322188 , n2364 );
nand ( n2366 , n2356 , n322188 );
buf ( n322190 , n2366 );
buf ( n322191 , n322190 );
xor ( n322192 , n2342 , n322191 );
buf ( n322193 , n322192 );
buf ( n322194 , n322193 );
xor ( n322195 , n322114 , n322194 );
buf ( n322196 , n322099 );
not ( n322197 , n322196 );
buf ( n322198 , n320692 );
not ( n2376 , n322198 );
or ( n322200 , n322197 , n2376 );
buf ( n322201 , n320699 );
buf ( n322202 , n554 );
buf ( n322203 , n586 );
xor ( n322204 , n322202 , n322203 );
buf ( n322205 , n322204 );
buf ( n322206 , n322205 );
nand ( n2381 , n322201 , n322206 );
buf ( n322208 , n2381 );
buf ( n322209 , n322208 );
nand ( n2384 , n322200 , n322209 );
buf ( n322211 , n2384 );
buf ( n322212 , n322211 );
buf ( n322213 , n559 );
buf ( n322214 , n583 );
or ( n2389 , n322213 , n322214 );
buf ( n322216 , n584 );
nand ( n2391 , n2389 , n322216 );
buf ( n322218 , n2391 );
buf ( n322219 , n559 );
buf ( n322220 , n583 );
nand ( n322221 , n322219 , n322220 );
buf ( n322222 , n322221 );
nand ( n322223 , n322218 , n322222 , n582 );
not ( n2398 , n322223 );
not ( n322225 , n322082 );
not ( n322226 , n926 );
or ( n2401 , n322225 , n322226 );
buf ( n322228 , n320642 );
buf ( n322229 , n552 );
buf ( n322230 , n588 );
xor ( n322231 , n322229 , n322230 );
buf ( n322232 , n322231 );
buf ( n322233 , n322232 );
nand ( n322234 , n322228 , n322233 );
buf ( n322235 , n322234 );
nand ( n322236 , n2401 , n322235 );
not ( n322237 , n322236 );
or ( n2412 , n2398 , n322237 );
or ( n322239 , n322223 , n322236 );
nand ( n322240 , n2412 , n322239 );
buf ( n322241 , n322240 );
xor ( n322242 , n322212 , n322241 );
not ( n322243 , n320732 );
not ( n2418 , n321140 );
or ( n322245 , n322243 , n2418 );
nand ( n322246 , n322118 , n591 );
nand ( n322247 , n322245 , n322246 );
buf ( n322248 , n322247 );
buf ( n322249 , n2331 );
buf ( n322250 , n559 );
and ( n2425 , n322249 , n322250 );
buf ( n322252 , n2425 );
buf ( n322253 , n322252 );
xor ( n322254 , n322248 , n322253 );
buf ( n322255 , n1475 );
not ( n2430 , n322255 );
buf ( n322257 , n321203 );
not ( n322258 , n322257 );
or ( n2433 , n2430 , n322258 );
buf ( n322260 , n321209 );
buf ( n322261 , n322168 );
nand ( n2436 , n322260 , n322261 );
buf ( n2437 , n2436 );
buf ( n322264 , n2437 );
nand ( n2439 , n2433 , n322264 );
buf ( n2440 , n2439 );
buf ( n322267 , n2440 );
and ( n322268 , n322254 , n322267 );
and ( n2443 , n322248 , n322253 );
or ( n322270 , n322268 , n2443 );
buf ( n322271 , n322270 );
buf ( n322272 , n322271 );
xor ( n322273 , n322242 , n322272 );
buf ( n322274 , n322273 );
buf ( n322275 , n322274 );
and ( n322276 , n322195 , n322275 );
and ( n2451 , n322114 , n322194 );
or ( n322278 , n322276 , n2451 );
buf ( n322279 , n322278 );
buf ( n322280 , n322279 );
xor ( n322281 , n322072 , n322280 );
buf ( n322282 , n322205 );
not ( n322283 , n322282 );
buf ( n322284 , n320692 );
not ( n2459 , n322284 );
or ( n2460 , n322283 , n2459 );
buf ( n322287 , n320699 );
buf ( n322288 , n553 );
buf ( n322289 , n586 );
xor ( n322290 , n322288 , n322289 );
buf ( n322291 , n322290 );
buf ( n322292 , n322291 );
nand ( n322293 , n322287 , n322292 );
buf ( n322294 , n322293 );
buf ( n322295 , n322294 );
nand ( n2470 , n2460 , n322295 );
buf ( n2471 , n2470 );
buf ( n322298 , n2471 );
buf ( n322299 , n322156 );
not ( n322300 , n322299 );
buf ( n322301 , n2327 );
not ( n2476 , n322301 );
or ( n322303 , n322300 , n2476 );
buf ( n2478 , n2331 );
buf ( n2479 , n557 );
buf ( n322306 , n582 );
xor ( n322307 , n2479 , n322306 );
buf ( n322308 , n322307 );
buf ( n322309 , n322308 );
nand ( n2484 , n2478 , n322309 );
buf ( n322311 , n2484 );
buf ( n322312 , n322311 );
nand ( n2487 , n322303 , n322312 );
buf ( n322314 , n2487 );
buf ( n322315 , n322127 );
not ( n322316 , n322315 );
buf ( n322317 , n873 );
not ( n322318 , n322317 );
or ( n2493 , n322316 , n322318 );
buf ( n322320 , n549 );
buf ( n2495 , n590 );
xor ( n2496 , n322320 , n2495 );
buf ( n2497 , n2496 );
buf ( n322324 , n2497 );
buf ( n322325 , n591 );
nand ( n322326 , n322324 , n322325 );
buf ( n322327 , n322326 );
buf ( n322328 , n322327 );
nand ( n322329 , n2493 , n322328 );
buf ( n322330 , n322329 );
xor ( n322331 , n322314 , n322330 );
buf ( n322332 , n322331 );
xor ( n2504 , n322298 , n322332 );
buf ( n322334 , n2504 );
buf ( n322335 , n322334 );
xor ( n2505 , n322212 , n322241 );
and ( n2506 , n2505 , n322272 );
and ( n322338 , n322212 , n322241 );
or ( n2508 , n2506 , n322338 );
buf ( n322340 , n2508 );
buf ( n322341 , n322340 );
xor ( n322342 , n322335 , n322341 );
and ( n322343 , n322218 , n322222 , n582 );
and ( n2513 , n322343 , n322236 );
buf ( n322345 , n2513 );
xor ( n322346 , n581 , n582 );
buf ( n322347 , n322346 );
buf ( n322348 , n559 );
and ( n2518 , n322347 , n322348 );
buf ( n2519 , n2518 );
buf ( n322351 , n2519 );
buf ( n322352 , n2361 );
not ( n322353 , n322352 );
buf ( n322354 , n321207 );
buf ( n322355 , n1462 );
nand ( n322356 , n322354 , n322355 );
buf ( n322357 , n322356 );
buf ( n322358 , n322357 );
not ( n322359 , n322358 );
buf ( n322360 , n322359 );
buf ( n322361 , n322360 );
not ( n322362 , n322361 );
or ( n322363 , n322353 , n322362 );
buf ( n322364 , n1469 );
buf ( n2534 , n555 );
buf ( n322366 , n584 );
xor ( n322367 , n2534 , n322366 );
buf ( n322368 , n322367 );
buf ( n322369 , n322368 );
nand ( n2539 , n322364 , n322369 );
buf ( n322371 , n2539 );
buf ( n322372 , n322371 );
nand ( n322373 , n322363 , n322372 );
buf ( n322374 , n322373 );
buf ( n322375 , n322374 );
xor ( n2544 , n322351 , n322375 );
buf ( n322377 , n322232 );
not ( n2546 , n322377 );
buf ( n322379 , n926 );
not ( n2548 , n322379 );
or ( n322381 , n2546 , n2548 );
buf ( n322382 , n320642 );
buf ( n322383 , n551 );
buf ( n322384 , n588 );
xor ( n2549 , n322383 , n322384 );
buf ( n322386 , n2549 );
buf ( n322387 , n322386 );
nand ( n322388 , n322382 , n322387 );
buf ( n322389 , n322388 );
buf ( n322390 , n322389 );
nand ( n322391 , n322381 , n322390 );
buf ( n322392 , n322391 );
buf ( n322393 , n322392 );
xor ( n322394 , n2544 , n322393 );
buf ( n322395 , n322394 );
buf ( n322396 , n322395 );
xor ( n2561 , n322345 , n322396 );
xor ( n2562 , n322135 , n322163 );
and ( n322399 , n2562 , n322191 );
and ( n2564 , n322135 , n322163 );
or ( n2565 , n322399 , n2564 );
buf ( n322402 , n2565 );
buf ( n322403 , n322402 );
xor ( n2568 , n2561 , n322403 );
buf ( n322405 , n2568 );
buf ( n322406 , n322405 );
xor ( n322407 , n322342 , n322406 );
buf ( n322408 , n322407 );
buf ( n322409 , n322408 );
and ( n322410 , n322281 , n322409 );
and ( n2570 , n322072 , n322280 );
or ( n322412 , n322410 , n2570 );
buf ( n322413 , n322412 );
xor ( n322414 , n321945 , n322413 );
xor ( n322415 , n321906 , n321923 );
xor ( n2575 , n322415 , n321937 );
buf ( n322417 , n2575 );
buf ( n322418 , n322417 );
xor ( n2578 , n322023 , n322026 );
and ( n2579 , n2578 , n322064 );
and ( n322421 , n322023 , n322026 );
or ( n322422 , n2579 , n322421 );
buf ( n322423 , n322422 );
buf ( n322424 , n322423 );
xor ( n322425 , n322418 , n322424 );
xor ( n2585 , n321710 , n1996 );
xor ( n322427 , n2585 , n2036 );
buf ( n322428 , n322427 );
buf ( n322429 , n322428 );
and ( n2589 , n322425 , n322429 );
and ( n2590 , n322418 , n322424 );
or ( n2591 , n2589 , n2590 );
buf ( n322433 , n2591 );
xor ( n322434 , n322335 , n322341 );
and ( n2594 , n322434 , n322406 );
and ( n322436 , n322335 , n322341 );
or ( n322437 , n2594 , n322436 );
buf ( n322438 , n322437 );
xor ( n322439 , n322433 , n322438 );
buf ( n322440 , n322291 );
not ( n2600 , n322440 );
buf ( n322442 , n320692 );
not ( n322443 , n322442 );
or ( n322444 , n2600 , n322443 );
buf ( n322445 , n320699 );
buf ( n322446 , n552 );
buf ( n322447 , n586 );
xor ( n2607 , n322446 , n322447 );
buf ( n322449 , n2607 );
buf ( n322450 , n322449 );
nand ( n322451 , n322445 , n322450 );
buf ( n322452 , n322451 );
buf ( n322453 , n322452 );
nand ( n322454 , n322444 , n322453 );
buf ( n322455 , n322454 );
buf ( n322456 , n559 );
buf ( n322457 , n580 );
xor ( n322458 , n322456 , n322457 );
buf ( n322459 , n322458 );
buf ( n322460 , n322459 );
not ( n322461 , n322460 );
not ( n2621 , n580 );
nor ( n322463 , n581 , n582 );
not ( n322464 , n322463 );
or ( n322465 , n2621 , n322464 );
not ( n2625 , n580 );
nand ( n322467 , n2625 , n581 , n582 );
nand ( n322468 , n322465 , n322467 );
buf ( n322469 , n322468 );
not ( n322470 , n322469 );
or ( n322471 , n322461 , n322470 );
buf ( n322472 , n322346 );
buf ( n322473 , n322472 );
buf ( n322474 , n322473 );
buf ( n322475 , n322474 );
xor ( n322476 , n580 , n558 );
buf ( n322477 , n322476 );
nand ( n322478 , n322475 , n322477 );
buf ( n322479 , n322478 );
buf ( n322480 , n322479 );
nand ( n2640 , n322471 , n322480 );
buf ( n322482 , n2640 );
not ( n2642 , n322482 );
xor ( n2643 , n322455 , n2642 );
not ( n322485 , n322386 );
not ( n322486 , n926 );
or ( n2646 , n322485 , n322486 );
buf ( n322488 , n320642 );
buf ( n322489 , n550 );
buf ( n322490 , n588 );
xor ( n322491 , n322489 , n322490 );
buf ( n322492 , n322491 );
buf ( n322493 , n322492 );
nand ( n2653 , n322488 , n322493 );
buf ( n322495 , n2653 );
nand ( n322496 , n2646 , n322495 );
buf ( n322497 , n559 );
buf ( n322498 , n581 );
or ( n2658 , n322497 , n322498 );
buf ( n322500 , n582 );
nand ( n322501 , n2658 , n322500 );
buf ( n322502 , n322501 );
buf ( n322503 , n559 );
buf ( n322504 , n581 );
nand ( n322505 , n322503 , n322504 );
buf ( n322506 , n322505 );
nand ( n322507 , n322502 , n322506 , n580 );
and ( n322508 , n322496 , n322507 );
not ( n2668 , n322496 );
not ( n322510 , n322507 );
and ( n322511 , n2668 , n322510 );
nor ( n2671 , n322508 , n322511 );
xor ( n2672 , n2643 , n2671 );
buf ( n322514 , n2672 );
xor ( n322515 , n322345 , n322396 );
and ( n2675 , n322515 , n322403 );
and ( n322517 , n322345 , n322396 );
or ( n322518 , n2675 , n322517 );
buf ( n322519 , n322518 );
buf ( n322520 , n322519 );
xor ( n322521 , n322514 , n322520 );
buf ( n322522 , n322314 );
buf ( n322523 , n322330 );
or ( n322524 , n322522 , n322523 );
buf ( n322525 , n2471 );
nand ( n322526 , n322524 , n322525 );
buf ( n322527 , n322526 );
buf ( n322528 , n322527 );
buf ( n322529 , n322314 );
buf ( n322530 , n322330 );
nand ( n2690 , n322529 , n322530 );
buf ( n2691 , n2690 );
buf ( n2692 , n2691 );
nand ( n2693 , n322528 , n2692 );
buf ( n2694 , n2693 );
buf ( n322536 , n2694 );
xor ( n2696 , n322351 , n322375 );
and ( n322538 , n2696 , n322393 );
and ( n2698 , n322351 , n322375 );
or ( n322540 , n322538 , n2698 );
buf ( n322541 , n322540 );
buf ( n322542 , n322541 );
xor ( n322543 , n322536 , n322542 );
not ( n322544 , n320732 );
not ( n2704 , n2497 );
or ( n322546 , n322544 , n2704 );
xor ( n322547 , n590 , n548 );
buf ( n322548 , n322547 );
buf ( n322549 , n591 );
nand ( n322550 , n322548 , n322549 );
buf ( n322551 , n322550 );
nand ( n322552 , n322546 , n322551 );
not ( n2711 , n322308 );
not ( n322554 , n322145 );
not ( n322555 , n322554 );
or ( n2714 , n2711 , n322555 );
buf ( n2715 , n322143 );
buf ( n322558 , n2715 );
xor ( n322559 , n582 , n556 );
buf ( n322560 , n322559 );
nand ( n2719 , n322558 , n322560 );
buf ( n322562 , n2719 );
nand ( n322563 , n2714 , n322562 );
xor ( n2722 , n322552 , n322563 );
buf ( n322565 , n321209 );
buf ( n322566 , n554 );
buf ( n322567 , n584 );
xor ( n2726 , n322566 , n322567 );
buf ( n322569 , n2726 );
buf ( n322570 , n322569 );
nand ( n2729 , n322565 , n322570 );
buf ( n322572 , n2729 );
nand ( n2731 , n321203 , n322368 );
nand ( n2732 , n322572 , n2731 );
xor ( n322575 , n2722 , n2732 );
buf ( n322576 , n322575 );
xor ( n322577 , n322543 , n322576 );
buf ( n322578 , n322577 );
buf ( n322579 , n322578 );
xor ( n322580 , n322521 , n322579 );
buf ( n322581 , n322580 );
xor ( n2740 , n322439 , n322581 );
xor ( n322583 , n322414 , n2740 );
buf ( n322584 , n322583 );
xor ( n322585 , n322418 , n322424 );
xor ( n322586 , n322585 , n322429 );
buf ( n322587 , n322586 );
buf ( n322588 , n322587 );
and ( n322589 , n2246 , n2253 );
not ( n322590 , n2246 );
and ( n2749 , n322590 , n2254 );
nor ( n322592 , n322589 , n2749 );
xor ( n322593 , n322051 , n322592 );
not ( n2752 , n322593 );
buf ( n322595 , n2752 );
not ( n322596 , n322595 );
buf ( n322597 , n321043 );
buf ( n322598 , n321089 );
nor ( n322599 , n322597 , n322598 );
buf ( n322600 , n322599 );
buf ( n322601 , n322600 );
not ( n2760 , n321056 );
buf ( n322603 , n2760 );
or ( n322604 , n322601 , n322603 );
buf ( n2763 , n321043 );
buf ( n322606 , n321089 );
nand ( n2765 , n2763 , n322606 );
buf ( n322608 , n2765 );
buf ( n322609 , n322608 );
nand ( n2768 , n322604 , n322609 );
buf ( n322611 , n2768 );
buf ( n322612 , n322611 );
not ( n322613 , n322612 );
or ( n2772 , n322596 , n322613 );
not ( n2773 , n322611 );
nand ( n322616 , n2773 , n322593 );
xnor ( n322617 , n321976 , n321959 );
buf ( n322618 , n322617 );
buf ( n322619 , n321983 );
and ( n322620 , n322618 , n322619 );
not ( n2779 , n322618 );
buf ( n322622 , n321986 );
and ( n322623 , n2779 , n322622 );
nor ( n322624 , n322620 , n322623 );
buf ( n322625 , n322624 );
nand ( n322626 , n322616 , n322625 );
buf ( n2785 , n322626 );
nand ( n2786 , n2772 , n2785 );
buf ( n2787 , n2786 );
buf ( n322630 , n2787 );
xor ( n2789 , n322248 , n322253 );
xor ( n322632 , n2789 , n322267 );
buf ( n322633 , n322632 );
buf ( n322634 , n322633 );
xor ( n2793 , n321170 , n321186 );
and ( n2794 , n2793 , n321220 );
and ( n322637 , n321170 , n321186 );
or ( n322638 , n2794 , n322637 );
buf ( n322639 , n322638 );
xor ( n2798 , n322634 , n322639 );
xor ( n322641 , n322089 , n322106 );
xor ( n322642 , n322641 , n322109 );
buf ( n322643 , n322642 );
buf ( n322644 , n322643 );
and ( n322645 , n2798 , n322644 );
and ( n2804 , n322634 , n322639 );
or ( n2805 , n322645 , n2804 );
buf ( n322648 , n2805 );
buf ( n322649 , n322648 );
xor ( n322650 , n322630 , n322649 );
xor ( n2809 , n322114 , n322194 );
xor ( n2810 , n2809 , n322275 );
buf ( n322653 , n2810 );
buf ( n322654 , n322653 );
and ( n2813 , n322650 , n322654 );
and ( n322656 , n322630 , n322649 );
or ( n322657 , n2813 , n322656 );
buf ( n322658 , n322657 );
buf ( n322659 , n322658 );
xor ( n322660 , n322588 , n322659 );
xor ( n322661 , n322072 , n322280 );
xor ( n2820 , n322661 , n322409 );
buf ( n322663 , n2820 );
buf ( n322664 , n322663 );
and ( n2823 , n322660 , n322664 );
and ( n322666 , n322588 , n322659 );
or ( n322667 , n2823 , n322666 );
buf ( n322668 , n322667 );
buf ( n322669 , n322668 );
nor ( n322670 , n322584 , n322669 );
buf ( n322671 , n322670 );
buf ( n322672 , n322671 );
xor ( n322673 , n322588 , n322659 );
xor ( n2832 , n322673 , n322664 );
buf ( n322675 , n2832 );
buf ( n322676 , n322675 );
xor ( n2835 , n321994 , n322009 );
xor ( n322678 , n2835 , n322067 );
buf ( n322679 , n322678 );
buf ( n322680 , n322679 );
not ( n322681 , n321024 );
nand ( n2840 , n322681 , n321019 );
not ( n2841 , n2840 );
not ( n2842 , n1354 );
or ( n2843 , n2841 , n2842 );
buf ( n322686 , n321019 );
not ( n2845 , n322686 );
buf ( n322688 , n321024 );
nand ( n2847 , n2845 , n322688 );
buf ( n322690 , n2847 );
nand ( n322691 , n2843 , n322690 );
buf ( n322692 , n322691 );
not ( n322693 , n321221 );
not ( n322694 , n321153 );
buf ( n2853 , n321148 );
not ( n322696 , n2853 );
nand ( n2855 , n322694 , n322696 );
not ( n322698 , n2855 );
or ( n322699 , n322693 , n322698 );
nand ( n322700 , n321153 , n2853 );
nand ( n322701 , n322699 , n322700 );
buf ( n322702 , n322701 );
xor ( n322703 , n322692 , n322702 );
xor ( n322704 , n322634 , n322639 );
xor ( n322705 , n322704 , n322644 );
buf ( n322706 , n322705 );
buf ( n322707 , n322706 );
and ( n322708 , n322703 , n322707 );
and ( n2867 , n322692 , n322702 );
or ( n322710 , n322708 , n2867 );
buf ( n322711 , n322710 );
buf ( n322712 , n322711 );
xor ( n322713 , n322680 , n322712 );
xor ( n2872 , n322630 , n322649 );
xor ( n322715 , n2872 , n322654 );
buf ( n322716 , n322715 );
buf ( n322717 , n322716 );
and ( n322718 , n322713 , n322717 );
and ( n322719 , n322680 , n322712 );
or ( n2878 , n322718 , n322719 );
buf ( n322721 , n2878 );
buf ( n322722 , n322721 );
nor ( n2881 , n322676 , n322722 );
buf ( n2882 , n2881 );
buf ( n322725 , n2882 );
nor ( n2884 , n322672 , n322725 );
buf ( n322727 , n2884 );
buf ( n322728 , n322727 );
xor ( n322729 , n322680 , n322712 );
xor ( n322730 , n322729 , n322717 );
buf ( n322731 , n322730 );
buf ( n322732 , n322731 );
buf ( n322733 , n322611 );
buf ( n322734 , n2752 );
and ( n322735 , n322733 , n322734 );
not ( n2893 , n322733 );
buf ( n322737 , n322593 );
and ( n2895 , n2893 , n322737 );
nor ( n322739 , n322735 , n2895 );
buf ( n322740 , n322739 );
buf ( n322741 , n322740 );
buf ( n322742 , n322625 );
xor ( n2900 , n322741 , n322742 );
buf ( n322744 , n2900 );
buf ( n322745 , n322744 );
xor ( n2903 , n321111 , n321119 );
and ( n2904 , n2903 , n321222 );
and ( n2905 , n321111 , n321119 );
or ( n322749 , n2904 , n2905 );
buf ( n322750 , n322749 );
xor ( n2908 , n322745 , n322750 );
xor ( n2909 , n322692 , n322702 );
xor ( n322753 , n2909 , n322707 );
buf ( n322754 , n322753 );
buf ( n322755 , n322754 );
and ( n2913 , n2908 , n322755 );
and ( n2914 , n322745 , n322750 );
or ( n2915 , n2913 , n2914 );
buf ( n322759 , n2915 );
buf ( n322760 , n322759 );
nor ( n322761 , n322732 , n322760 );
buf ( n322762 , n322761 );
buf ( n322763 , n322762 );
xor ( n2921 , n322745 , n322750 );
xor ( n2922 , n2921 , n322755 );
buf ( n322766 , n2922 );
buf ( n322767 , n322766 );
nand ( n2925 , n321101 , n321104 );
not ( n2926 , n2925 );
not ( n2927 , n1484 );
or ( n2928 , n2926 , n2927 );
nand ( n2929 , n321100 , n320984 );
nand ( n2930 , n2928 , n2929 );
buf ( n322774 , n2930 );
nor ( n2932 , n322767 , n322774 );
buf ( n322776 , n2932 );
buf ( n322777 , n322776 );
nor ( n2935 , n322763 , n322777 );
buf ( n322779 , n2935 );
buf ( n322780 , n322779 );
and ( n2938 , n322728 , n322780 );
buf ( n322782 , n2938 );
not ( n2940 , n322782 );
or ( n2941 , n1835 , n2940 );
not ( n2942 , n322727 );
buf ( n322786 , n322766 );
buf ( n322787 , n2930 );
nand ( n2945 , n322786 , n322787 );
buf ( n322789 , n2945 );
or ( n2947 , n322762 , n322789 );
buf ( n322791 , n322731 );
buf ( n322792 , n322759 );
nand ( n2950 , n322791 , n322792 );
buf ( n322794 , n2950 );
nand ( n2952 , n2947 , n322794 );
not ( n2953 , n2952 );
or ( n2954 , n2942 , n2953 );
not ( n2955 , n322583 );
buf ( n322799 , n322668 );
not ( n2957 , n322799 );
buf ( n322801 , n2957 );
nand ( n2959 , n2955 , n322801 );
buf ( n322803 , n322675 );
buf ( n322804 , n322721 );
and ( n2962 , n322803 , n322804 );
buf ( n322806 , n2962 );
and ( n2964 , n2959 , n322806 );
and ( n2965 , n322583 , n322668 );
nor ( n2966 , n2964 , n2965 );
nand ( n2967 , n2954 , n2966 );
buf ( n322811 , n2967 );
not ( n2969 , n322811 );
buf ( n322813 , n2969 );
nand ( n2971 , n2941 , n322813 );
not ( n2972 , n2971 );
buf ( n322816 , n547 );
buf ( n322817 , n572 );
xor ( n2975 , n322816 , n322817 );
buf ( n322819 , n2975 );
buf ( n322820 , n322819 );
not ( n2978 , n322820 );
buf ( n322822 , n1023 );
not ( n2980 , n322822 );
or ( n2981 , n2978 , n2980 );
buf ( n322825 , n1026 );
xor ( n2983 , n572 , n546 );
buf ( n322827 , n2983 );
nand ( n2985 , n322825 , n322827 );
buf ( n322829 , n2985 );
buf ( n322830 , n322829 );
nand ( n2988 , n2981 , n322830 );
buf ( n322832 , n2988 );
buf ( n322833 , n559 );
buf ( n322834 , n560 );
xor ( n2992 , n322833 , n322834 );
buf ( n322836 , n2992 );
buf ( n322837 , n322836 );
not ( n2995 , n322837 );
and ( n2996 , n560 , n561 );
not ( n2997 , n560 );
not ( n2998 , n561 );
and ( n2999 , n2997 , n2998 );
nor ( n3000 , n2996 , n2999 );
not ( n3001 , n3000 );
buf ( n322845 , n561 );
buf ( n322846 , n562 );
xor ( n3004 , n322845 , n322846 );
buf ( n322848 , n3004 );
nor ( n3006 , n3001 , n322848 );
buf ( n322850 , n3006 );
not ( n3008 , n322850 );
or ( n3009 , n2995 , n3008 );
xor ( n3010 , n562 , n561 );
buf ( n322854 , n3010 );
buf ( n322855 , n558 );
buf ( n322856 , n560 );
xor ( n3014 , n322855 , n322856 );
buf ( n322858 , n3014 );
buf ( n322859 , n322858 );
nand ( n3017 , n322854 , n322859 );
buf ( n322861 , n3017 );
buf ( n322862 , n322861 );
nand ( n3020 , n3009 , n322862 );
buf ( n322864 , n3020 );
buf ( n322865 , n322864 );
not ( n3023 , n322865 );
buf ( n322867 , n3023 );
xor ( n3025 , n322832 , n322867 );
xor ( n3026 , n568 , n551 );
buf ( n322870 , n3026 );
not ( n3028 , n322870 );
buf ( n322872 , n321069 );
not ( n3030 , n322872 );
or ( n3031 , n3028 , n3030 );
buf ( n322875 , n1339 );
buf ( n322876 , n550 );
buf ( n322877 , n568 );
xor ( n3035 , n322876 , n322877 );
buf ( n322879 , n3035 );
buf ( n322880 , n322879 );
nand ( n3038 , n322875 , n322880 );
buf ( n322882 , n3038 );
buf ( n322883 , n322882 );
nand ( n3041 , n3031 , n322883 );
buf ( n322885 , n3041 );
xor ( n3043 , n3025 , n322885 );
buf ( n322887 , n3043 );
xor ( n3045 , n566 , n554 );
not ( n3046 , n3045 );
not ( n3047 , n1975 );
or ( n3048 , n3046 , n3047 );
buf ( n322892 , n321771 );
buf ( n322893 , n553 );
buf ( n322894 , n566 );
xor ( n3052 , n322893 , n322894 );
buf ( n322896 , n3052 );
buf ( n322897 , n322896 );
nand ( n3055 , n322892 , n322897 );
buf ( n322899 , n3055 );
nand ( n3057 , n3048 , n322899 );
not ( n3058 , n3057 );
xor ( n3059 , n568 , n552 );
and ( n3060 , n321072 , n3059 );
and ( n3061 , n1339 , n3026 );
nor ( n3062 , n3060 , n3061 );
not ( n3063 , n3062 );
not ( n3064 , n3063 );
or ( n3065 , n3058 , n3064 );
not ( n3066 , n3062 );
buf ( n322910 , n3057 );
not ( n3068 , n322910 );
buf ( n322912 , n3068 );
not ( n3070 , n322912 );
or ( n3071 , n3066 , n3070 );
buf ( n322915 , n550 );
buf ( n322916 , n570 );
xor ( n3074 , n322915 , n322916 );
buf ( n322918 , n3074 );
not ( n3076 , n322918 );
not ( n3077 , n321032 );
or ( n3078 , n3076 , n3077 );
buf ( n322922 , n320483 );
xor ( n3080 , n570 , n549 );
buf ( n322924 , n3080 );
nand ( n3082 , n322922 , n322924 );
buf ( n322926 , n3082 );
nand ( n3084 , n3078 , n322926 );
nand ( n3085 , n3071 , n3084 );
nand ( n3086 , n3065 , n3085 );
buf ( n322930 , n3086 );
xor ( n3088 , n322887 , n322930 );
not ( n3089 , n565 );
nand ( n3090 , n1842 , n3089 , n564 );
nand ( n3091 , n1849 , n3090 );
not ( n3092 , n3091 );
buf ( n322936 , n555 );
buf ( n322937 , n564 );
xor ( n3095 , n322936 , n322937 );
buf ( n322939 , n3095 );
not ( n3097 , n322939 );
or ( n3098 , n3092 , n3097 );
buf ( n322942 , n1857 );
buf ( n322943 , n554 );
buf ( n322944 , n564 );
xor ( n3102 , n322943 , n322944 );
buf ( n322946 , n3102 );
buf ( n322947 , n322946 );
nand ( n3105 , n322942 , n322947 );
buf ( n322949 , n3105 );
nand ( n3107 , n3098 , n322949 );
buf ( n322951 , n3107 );
not ( n3109 , n3080 );
nor ( n3110 , n321031 , n320480 );
not ( n3111 , n3110 );
or ( n3112 , n3109 , n3111 );
buf ( n322956 , n320480 );
xor ( n3114 , n570 , n548 );
buf ( n322958 , n3114 );
nand ( n3116 , n322956 , n322958 );
buf ( n322960 , n3116 );
nand ( n3118 , n3112 , n322960 );
buf ( n322962 , n3118 );
xor ( n3120 , n322951 , n322962 );
not ( n3121 , n321771 );
and ( n3122 , n566 , n552 );
not ( n3123 , n566 );
and ( n3124 , n3123 , n320990 );
nor ( n3125 , n3122 , n3124 );
not ( n3126 , n3125 );
or ( n3127 , n3121 , n3126 );
buf ( n322971 , n1975 );
not ( n3129 , n322971 );
buf ( n322973 , n3129 );
buf ( n322974 , n322896 );
not ( n3132 , n322974 );
buf ( n322976 , n3132 );
or ( n3134 , n322973 , n322976 );
nand ( n3135 , n3127 , n3134 );
buf ( n322979 , n3135 );
xor ( n3137 , n3120 , n322979 );
buf ( n322981 , n3137 );
buf ( n322982 , n322981 );
xor ( n3140 , n3088 , n322982 );
buf ( n322984 , n3140 );
buf ( n322985 , n322984 );
buf ( n322986 , n558 );
buf ( n322987 , n562 );
xor ( n3145 , n322986 , n322987 );
buf ( n322989 , n3145 );
not ( n3147 , n322989 );
buf ( n322991 , n562 );
buf ( n322992 , n563 );
xnor ( n3150 , n322991 , n322992 );
buf ( n322994 , n3150 );
buf ( n322995 , n563 );
buf ( n322996 , n564 );
xor ( n3154 , n322995 , n322996 );
buf ( n322998 , n3154 );
nor ( n3156 , n322994 , n322998 );
buf ( n3157 , n3156 );
not ( n3158 , n3157 );
or ( n3159 , n3147 , n3158 );
buf ( n323003 , n563 );
buf ( n323004 , n564 );
xor ( n3162 , n323003 , n323004 );
buf ( n323006 , n3162 );
buf ( n323007 , n323006 );
buf ( n3165 , n323007 );
buf ( n323009 , n3165 );
buf ( n323010 , n323009 );
buf ( n323011 , n557 );
buf ( n323012 , n562 );
xor ( n3170 , n323011 , n323012 );
buf ( n323014 , n3170 );
buf ( n323015 , n323014 );
nand ( n3173 , n323010 , n323015 );
buf ( n323017 , n3173 );
nand ( n3175 , n3159 , n323017 );
buf ( n323019 , n3175 );
buf ( n323020 , n556 );
buf ( n323021 , n564 );
xor ( n3179 , n323020 , n323021 );
buf ( n323023 , n3179 );
buf ( n323024 , n323023 );
not ( n3182 , n323024 );
buf ( n323026 , n321592 );
not ( n3184 , n323026 );
or ( n3185 , n3182 , n3184 );
buf ( n3186 , n1857 );
buf ( n323030 , n3186 );
buf ( n323031 , n322939 );
nand ( n3189 , n323030 , n323031 );
buf ( n323033 , n3189 );
buf ( n323034 , n323033 );
nand ( n3192 , n3185 , n323034 );
buf ( n323036 , n3192 );
buf ( n323037 , n323036 );
xor ( n3195 , n323019 , n323037 );
buf ( n323039 , n559 );
buf ( n323040 , n563 );
or ( n3198 , n323039 , n323040 );
buf ( n323042 , n564 );
nand ( n3200 , n3198 , n323042 );
buf ( n323044 , n3200 );
buf ( n323045 , n323044 );
buf ( n323046 , n559 );
buf ( n323047 , n563 );
nand ( n3205 , n323046 , n323047 );
buf ( n323049 , n3205 );
buf ( n323050 , n323049 );
buf ( n323051 , n562 );
and ( n3209 , n323045 , n323050 , n323051 );
buf ( n323053 , n3209 );
buf ( n323054 , n323053 );
buf ( n323055 , n547 );
buf ( n323056 , n574 );
xor ( n3214 , n323055 , n323056 );
buf ( n323058 , n3214 );
buf ( n323059 , n323058 );
not ( n3217 , n323059 );
buf ( n323061 , n320441 );
not ( n3219 , n323061 );
or ( n3220 , n3217 , n3219 );
buf ( n323064 , n546 );
buf ( n323065 , n574 );
xor ( n3223 , n323064 , n323065 );
buf ( n323067 , n3223 );
buf ( n323068 , n323067 );
buf ( n323069 , n575 );
nand ( n3227 , n323068 , n323069 );
buf ( n323071 , n3227 );
buf ( n323072 , n323071 );
nand ( n3230 , n3220 , n323072 );
buf ( n323074 , n3230 );
buf ( n323075 , n323074 );
and ( n3233 , n323054 , n323075 );
buf ( n323077 , n3233 );
buf ( n323078 , n323077 );
xor ( n3236 , n3195 , n323078 );
buf ( n323080 , n3236 );
buf ( n323081 , n323080 );
xor ( n3239 , n3084 , n3063 );
xor ( n3240 , n3239 , n3057 );
buf ( n323084 , n3240 );
xor ( n3242 , n323081 , n323084 );
xor ( n3243 , n323054 , n323075 );
buf ( n323087 , n3243 );
buf ( n323088 , n323087 );
buf ( n323089 , n321842 );
not ( n3247 , n323089 );
buf ( n323091 , n320441 );
not ( n3249 , n323091 );
or ( n3250 , n3247 , n3249 );
buf ( n323094 , n323058 );
buf ( n323095 , n575 );
nand ( n3253 , n323094 , n323095 );
buf ( n323097 , n3253 );
buf ( n323098 , n323097 );
nand ( n3256 , n3250 , n323098 );
buf ( n323100 , n3256 );
buf ( n323101 , n323100 );
buf ( n323102 , n321601 );
not ( n3260 , n323102 );
buf ( n323104 , n1850 );
not ( n3262 , n323104 );
or ( n3263 , n3260 , n3262 );
buf ( n323107 , n1857 );
buf ( n323108 , n557 );
buf ( n323109 , n564 );
xor ( n3267 , n323108 , n323109 );
buf ( n323111 , n3267 );
buf ( n323112 , n323111 );
nand ( n3270 , n323107 , n323112 );
buf ( n323114 , n3270 );
buf ( n323115 , n323114 );
nand ( n3273 , n3263 , n323115 );
buf ( n323117 , n3273 );
buf ( n323118 , n323117 );
xor ( n3276 , n323101 , n323118 );
buf ( n323120 , n322973 );
buf ( n323121 , n321873 );
or ( n3279 , n323120 , n323121 );
buf ( n323123 , n321771 );
buf ( n323124 , n555 );
buf ( n323125 , n566 );
xor ( n3283 , n323124 , n323125 );
buf ( n323127 , n3283 );
buf ( n323128 , n323127 );
nand ( n3286 , n323123 , n323128 );
buf ( n323130 , n3286 );
buf ( n323131 , n323130 );
nand ( n3289 , n3279 , n323131 );
buf ( n323133 , n3289 );
buf ( n323134 , n323133 );
and ( n3292 , n3276 , n323134 );
and ( n3293 , n323101 , n323118 );
or ( n3294 , n3292 , n3293 );
buf ( n323138 , n3294 );
buf ( n323139 , n323138 );
xor ( n3297 , n323088 , n323139 );
nand ( n3298 , n323006 , n559 );
not ( n3299 , n3298 );
not ( n3300 , n321644 );
nor ( n3301 , n320761 , n320525 );
not ( n3302 , n3301 );
or ( n3303 , n3300 , n3302 );
not ( n3304 , n320535 );
not ( n3305 , n3304 );
buf ( n323149 , n549 );
buf ( n323150 , n572 );
xor ( n3308 , n323149 , n323150 );
buf ( n323152 , n3308 );
nand ( n3310 , n3305 , n323152 );
nand ( n3311 , n3303 , n3310 );
not ( n3312 , n3311 );
not ( n3313 , n3312 );
or ( n3314 , n3299 , n3313 );
not ( n3315 , n321860 );
not ( n3316 , n321069 );
or ( n3317 , n3315 , n3316 );
buf ( n323161 , n1339 );
buf ( n323162 , n553 );
buf ( n323163 , n568 );
xor ( n3321 , n323162 , n323163 );
buf ( n323165 , n3321 );
buf ( n323166 , n323165 );
nand ( n3324 , n323161 , n323166 );
buf ( n323168 , n3324 );
nand ( n3326 , n3317 , n323168 );
nand ( n3327 , n3314 , n3326 );
not ( n3328 , n3298 );
nand ( n3329 , n3328 , n3311 );
nand ( n3330 , n3327 , n3329 );
buf ( n323174 , n3330 );
and ( n3332 , n3297 , n323174 );
and ( n3333 , n323088 , n323139 );
or ( n3334 , n3332 , n3333 );
buf ( n323178 , n3334 );
buf ( n323179 , n323178 );
and ( n3337 , n3242 , n323179 );
and ( n3338 , n323081 , n323084 );
or ( n3339 , n3337 , n3338 );
buf ( n323183 , n3339 );
buf ( n323184 , n323183 );
xor ( n3342 , n322985 , n323184 );
xor ( n3343 , n323019 , n323037 );
and ( n3344 , n3343 , n323078 );
and ( n3345 , n323019 , n323037 );
or ( n3346 , n3344 , n3345 );
buf ( n323190 , n3346 );
buf ( n323191 , n323190 );
not ( n3349 , n323014 );
not ( n3350 , n3156 );
or ( n3351 , n3349 , n3350 );
buf ( n323195 , n323009 );
xor ( n3353 , n562 , n556 );
buf ( n323197 , n3353 );
nand ( n3355 , n323195 , n323197 );
buf ( n323199 , n3355 );
nand ( n3357 , n3351 , n323199 );
buf ( n323201 , n559 );
buf ( n323202 , n561 );
or ( n3360 , n323201 , n323202 );
buf ( n323204 , n562 );
nand ( n3362 , n3360 , n323204 );
buf ( n323206 , n3362 );
buf ( n323207 , n323206 );
buf ( n323208 , n559 );
buf ( n323209 , n561 );
nand ( n3367 , n323208 , n323209 );
buf ( n323211 , n3367 );
buf ( n323212 , n323211 );
buf ( n323213 , n560 );
nand ( n3371 , n323207 , n323212 , n323213 );
buf ( n323215 , n3371 );
buf ( n323216 , n545 );
buf ( n323217 , n574 );
xor ( n3375 , n323216 , n323217 );
buf ( n323219 , n3375 );
not ( n3377 , n323219 );
not ( n3378 , n320441 );
or ( n323222 , n3377 , n3378 );
xor ( n323223 , n574 , n544 );
buf ( n323224 , n323223 );
buf ( n323225 , n575 );
nand ( n323226 , n323224 , n323225 );
buf ( n323227 , n323226 );
nand ( n3385 , n323222 , n323227 );
xnor ( n323229 , n323215 , n3385 );
xor ( n323230 , n3357 , n323229 );
buf ( n323231 , n548 );
buf ( n323232 , n572 );
xor ( n323233 , n323231 , n323232 );
buf ( n323234 , n323233 );
buf ( n323235 , n323234 );
not ( n3393 , n323235 );
buf ( n323237 , n320531 );
not ( n3395 , n323237 );
or ( n323239 , n3393 , n3395 );
buf ( n3397 , n320535 );
buf ( n323241 , n322819 );
nand ( n323242 , n3397 , n323241 );
buf ( n323243 , n323242 );
buf ( n323244 , n323243 );
nand ( n323245 , n323239 , n323244 );
buf ( n323246 , n323245 );
not ( n3404 , n323246 );
buf ( n323248 , n323067 );
not ( n323249 , n323248 );
buf ( n323250 , n320441 );
not ( n3408 , n323250 );
or ( n323252 , n323249 , n3408 );
buf ( n323253 , n323219 );
buf ( n323254 , n575 );
nand ( n323255 , n323253 , n323254 );
buf ( n323256 , n323255 );
buf ( n323257 , n323256 );
nand ( n323258 , n323252 , n323257 );
buf ( n323259 , n323258 );
not ( n323260 , n323259 );
buf ( n323261 , n322848 );
buf ( n323262 , n559 );
and ( n323263 , n323261 , n323262 );
buf ( n323264 , n323263 );
not ( n3422 , n323264 );
nand ( n3423 , n323260 , n3422 );
not ( n3424 , n3423 );
or ( n3425 , n3404 , n3424 );
nand ( n3426 , n323264 , n323259 );
nand ( n3427 , n3425 , n3426 );
xor ( n3428 , n323230 , n3427 );
buf ( n323272 , n3428 );
xor ( n323273 , n323191 , n323272 );
buf ( n323274 , n559 );
buf ( n323275 , n562 );
xor ( n3433 , n323274 , n323275 );
buf ( n323277 , n3433 );
buf ( n323278 , n323277 );
not ( n3436 , n323278 );
buf ( n3437 , n322994 );
buf ( n323281 , n322998 );
nor ( n323282 , n3437 , n323281 );
buf ( n323283 , n323282 );
buf ( n323284 , n323283 );
not ( n323285 , n323284 );
or ( n3443 , n3436 , n323285 );
buf ( n323287 , n323006 );
buf ( n3445 , n322989 );
nand ( n3446 , n323287 , n3445 );
buf ( n3447 , n3446 );
buf ( n3448 , n3447 );
nand ( n3449 , n3443 , n3448 );
buf ( n3450 , n3449 );
not ( n323294 , n3450 );
buf ( n323295 , n323111 );
not ( n323296 , n323295 );
buf ( n323297 , n1850 );
not ( n323298 , n323297 );
or ( n3456 , n323296 , n323298 );
buf ( n323300 , n1857 );
buf ( n323301 , n323023 );
nand ( n323302 , n323300 , n323301 );
buf ( n323303 , n323302 );
buf ( n323304 , n323303 );
nand ( n323305 , n3456 , n323304 );
buf ( n323306 , n323305 );
not ( n3464 , n323306 );
nand ( n323308 , n323294 , n3464 );
not ( n323309 , n323308 );
buf ( n323310 , n551 );
buf ( n323311 , n570 );
xor ( n323312 , n323310 , n323311 );
buf ( n323313 , n323312 );
buf ( n323314 , n323313 );
not ( n323315 , n323314 );
buf ( n323316 , n320476 );
not ( n3474 , n323316 );
or ( n323318 , n323315 , n3474 );
buf ( n3476 , n320483 );
buf ( n323320 , n322918 );
nand ( n323321 , n3476 , n323320 );
buf ( n323322 , n323321 );
buf ( n323323 , n323322 );
nand ( n323324 , n323318 , n323323 );
buf ( n323325 , n323324 );
not ( n3483 , n323325 );
or ( n323327 , n323309 , n3483 );
nand ( n323328 , n323306 , n3450 );
nand ( n323329 , n323327 , n323328 );
not ( n3487 , n323329 );
not ( n323331 , n323264 );
not ( n3489 , n323260 );
or ( n3490 , n323331 , n3489 );
nand ( n323334 , n323259 , n3422 );
nand ( n323335 , n3490 , n323334 );
xor ( n323336 , n323335 , n323246 );
not ( n3494 , n323336 );
or ( n323338 , n3487 , n3494 );
nor ( n323339 , n323336 , n323329 );
buf ( n323340 , n323165 );
not ( n323341 , n323340 );
buf ( n323342 , n321069 );
not ( n3500 , n323342 );
or ( n323344 , n323341 , n3500 );
buf ( n323345 , n1339 );
buf ( n323346 , n3059 );
nand ( n3504 , n323345 , n323346 );
buf ( n323348 , n3504 );
buf ( n323349 , n323348 );
nand ( n323350 , n323344 , n323349 );
buf ( n323351 , n323350 );
buf ( n323352 , n323351 );
buf ( n323353 , n322973 );
buf ( n323354 , n323127 );
not ( n3512 , n323354 );
buf ( n323356 , n3512 );
buf ( n323357 , n323356 );
or ( n3515 , n323353 , n323357 );
buf ( n323359 , n321771 );
buf ( n323360 , n3045 );
nand ( n3518 , n323359 , n323360 );
buf ( n323362 , n3518 );
buf ( n323363 , n323362 );
nand ( n3521 , n3515 , n323363 );
buf ( n323365 , n3521 );
buf ( n323366 , n323365 );
xor ( n3524 , n323352 , n323366 );
buf ( n323368 , n323152 );
not ( n3526 , n323368 );
buf ( n323370 , n1023 );
not ( n323371 , n323370 );
or ( n3529 , n3526 , n323371 );
buf ( n323373 , n1026 );
buf ( n323374 , n323234 );
nand ( n3532 , n323373 , n323374 );
buf ( n323376 , n3532 );
buf ( n323377 , n323376 );
nand ( n323378 , n3529 , n323377 );
buf ( n323379 , n323378 );
buf ( n323380 , n323379 );
and ( n3538 , n3524 , n323380 );
and ( n323382 , n323352 , n323366 );
or ( n3540 , n3538 , n323382 );
buf ( n323384 , n3540 );
buf ( n323385 , n323384 );
not ( n3543 , n323385 );
buf ( n323387 , n3543 );
or ( n323388 , n323339 , n323387 );
nand ( n3546 , n323338 , n323388 );
buf ( n323390 , n3546 );
xor ( n323391 , n323273 , n323390 );
buf ( n323392 , n323391 );
buf ( n323393 , n323392 );
xnor ( n323394 , n3342 , n323393 );
buf ( n323395 , n323394 );
buf ( n323396 , n323395 );
xor ( n323397 , n323088 , n323139 );
xor ( n3555 , n323397 , n323174 );
buf ( n323399 , n3555 );
buf ( n323400 , n323399 );
xor ( n323401 , n323101 , n323118 );
xor ( n323402 , n323401 , n323134 );
buf ( n323403 , n323402 );
xor ( n323404 , n3298 , n3311 );
xnor ( n3562 , n323404 , n3326 );
or ( n323406 , n323403 , n3562 );
not ( n323407 , n323406 );
xor ( n323408 , n321608 , n321629 );
and ( n3566 , n323408 , n321667 );
and ( n323410 , n321608 , n321629 );
or ( n323411 , n3566 , n323410 );
buf ( n323412 , n323411 );
not ( n323413 , n323412 );
or ( n3571 , n323407 , n323413 );
nand ( n323415 , n323403 , n3562 );
nand ( n3573 , n3571 , n323415 );
buf ( n323417 , n3573 );
xor ( n323418 , n323400 , n323417 );
not ( n323419 , n3464 );
not ( n3577 , n3450 );
or ( n323421 , n323419 , n3577 );
nand ( n323422 , n323294 , n323306 );
nand ( n323423 , n323421 , n323422 );
and ( n3581 , n323423 , n323325 );
not ( n323425 , n323423 );
not ( n323426 , n323325 );
and ( n3584 , n323425 , n323426 );
nor ( n323428 , n3581 , n3584 );
buf ( n323429 , n323428 );
xor ( n3587 , n323352 , n323366 );
xor ( n3588 , n3587 , n323380 );
buf ( n323432 , n3588 );
buf ( n323433 , n323432 );
xor ( n3591 , n323429 , n323433 );
buf ( n323435 , n321622 );
not ( n323436 , n323435 );
buf ( n323437 , n320476 );
not ( n323438 , n323437 );
or ( n3596 , n323436 , n323438 );
buf ( n323440 , n320480 );
buf ( n323441 , n323313 );
nand ( n3599 , n323440 , n323441 );
buf ( n323443 , n3599 );
buf ( n323444 , n323443 );
nand ( n3602 , n3596 , n323444 );
buf ( n323446 , n3602 );
buf ( n323447 , n323446 );
not ( n323448 , n323447 );
buf ( n323449 , n323448 );
buf ( n3607 , n323449 );
not ( n3608 , n3607 );
buf ( n323452 , n321665 );
not ( n323453 , n323452 );
buf ( n323454 , n321650 );
nand ( n323455 , n323453 , n323454 );
buf ( n323456 , n323455 );
buf ( n323457 , n323456 );
not ( n3615 , n323457 );
or ( n323459 , n3608 , n3615 );
xor ( n323460 , n321850 , n2085 );
and ( n3618 , n323460 , n321890 );
and ( n3619 , n321850 , n2085 );
or ( n323463 , n3618 , n3619 );
buf ( n323464 , n323463 );
buf ( n323465 , n323464 );
nand ( n3623 , n323459 , n323465 );
buf ( n3624 , n3623 );
buf ( n323468 , n3624 );
buf ( n323469 , n323456 );
not ( n323470 , n323469 );
buf ( n323471 , n323446 );
nand ( n3629 , n323470 , n323471 );
buf ( n3630 , n3629 );
buf ( n323474 , n3630 );
nand ( n323475 , n323468 , n323474 );
buf ( n323476 , n323475 );
buf ( n323477 , n323476 );
xor ( n3635 , n3591 , n323477 );
buf ( n323479 , n3635 );
buf ( n323480 , n323479 );
and ( n3638 , n323418 , n323480 );
and ( n323482 , n323400 , n323417 );
or ( n323483 , n3638 , n323482 );
buf ( n323484 , n323483 );
buf ( n323485 , n323484 );
buf ( n323486 , n559 );
buf ( n323487 , n579 );
or ( n323488 , n323486 , n323487 );
buf ( n323489 , n580 );
nand ( n323490 , n323488 , n323489 );
buf ( n323491 , n323490 );
buf ( n323492 , n323491 );
buf ( n323493 , n559 );
buf ( n323494 , n579 );
nand ( n3652 , n323493 , n323494 );
buf ( n3653 , n3652 );
buf ( n3654 , n3653 );
buf ( n323498 , n578 );
and ( n323499 , n323492 , n3654 , n323498 );
buf ( n323500 , n323499 );
buf ( n323501 , n323500 );
not ( n323502 , n591 );
buf ( n323503 , n546 );
buf ( n323504 , n590 );
xor ( n3662 , n323503 , n323504 );
buf ( n323506 , n3662 );
not ( n3664 , n323506 );
or ( n323508 , n323502 , n3664 );
xor ( n3666 , n590 , n547 );
nand ( n3667 , n873 , n3666 );
nand ( n323511 , n323508 , n3667 );
buf ( n323512 , n323511 );
xor ( n323513 , n323501 , n323512 );
buf ( n323514 , n323513 );
buf ( n323515 , n323514 );
buf ( n323516 , n322547 );
not ( n3674 , n323516 );
buf ( n323518 , n320732 );
not ( n323519 , n323518 );
or ( n3677 , n3674 , n323519 );
buf ( n323521 , n3666 );
buf ( n323522 , n591 );
nand ( n3680 , n323521 , n323522 );
buf ( n323524 , n3680 );
buf ( n323525 , n323524 );
nand ( n3683 , n3677 , n323525 );
buf ( n323527 , n3683 );
buf ( n323528 , n323527 );
buf ( n323529 , n322476 );
not ( n323530 , n323529 );
not ( n323531 , n322463 );
not ( n3689 , n580 );
or ( n323533 , n323531 , n3689 );
nand ( n323534 , n323533 , n322467 );
buf ( n323535 , n323534 );
not ( n3693 , n323535 );
or ( n3694 , n323530 , n3693 );
buf ( n323538 , n322346 );
xor ( n3696 , n580 , n557 );
buf ( n323540 , n3696 );
nand ( n3698 , n323538 , n323540 );
buf ( n323542 , n3698 );
buf ( n323543 , n323542 );
nand ( n3701 , n3694 , n323543 );
buf ( n3702 , n3701 );
buf ( n3703 , n3702 );
xor ( n3704 , n323528 , n3703 );
buf ( n323548 , n322559 );
not ( n323549 , n323548 );
not ( n323550 , n322145 );
buf ( n323551 , n323550 );
not ( n323552 , n323551 );
or ( n3710 , n323549 , n323552 );
and ( n323554 , n584 , n583 );
not ( n323555 , n584 );
not ( n323556 , n583 );
and ( n3714 , n323555 , n323556 );
nor ( n323558 , n323554 , n3714 );
not ( n323559 , n323558 );
buf ( n323560 , n323559 );
not ( n323561 , n323560 );
buf ( n323562 , n323561 );
buf ( n323563 , n323562 );
xor ( n3721 , n582 , n555 );
buf ( n323565 , n3721 );
nand ( n3723 , n323563 , n323565 );
buf ( n323567 , n3723 );
buf ( n323568 , n323567 );
nand ( n3726 , n3710 , n323568 );
buf ( n3727 , n3726 );
buf ( n323571 , n3727 );
and ( n3729 , n3704 , n323571 );
and ( n323573 , n323528 , n3703 );
or ( n323574 , n3729 , n323573 );
buf ( n323575 , n323574 );
buf ( n323576 , n323575 );
xor ( n323577 , n323515 , n323576 );
and ( n3735 , n579 , n580 );
not ( n323579 , n579 );
and ( n323580 , n323579 , n2625 );
nor ( n3738 , n3735 , n323580 );
buf ( n323582 , n3738 );
buf ( n323583 , n559 );
and ( n3741 , n323582 , n323583 );
buf ( n323585 , n3741 );
buf ( n323586 , n323585 );
buf ( n323587 , n322569 );
not ( n323588 , n323587 );
buf ( n323589 , n322357 );
not ( n323590 , n323589 );
buf ( n323591 , n323590 );
buf ( n323592 , n323591 );
not ( n3750 , n323592 );
or ( n323594 , n323588 , n3750 );
not ( n3752 , n321207 );
buf ( n323596 , n3752 );
buf ( n3754 , n553 );
buf ( n3755 , n584 );
xor ( n3756 , n3754 , n3755 );
buf ( n3757 , n3756 );
buf ( n323601 , n3757 );
nand ( n323602 , n323596 , n323601 );
buf ( n323603 , n323602 );
buf ( n323604 , n323603 );
nand ( n323605 , n323594 , n323604 );
buf ( n323606 , n323605 );
buf ( n323607 , n323606 );
xor ( n323608 , n323586 , n323607 );
buf ( n323609 , n322492 );
not ( n323610 , n323609 );
buf ( n323611 , n898 );
not ( n323612 , n323611 );
or ( n3770 , n323610 , n323612 );
buf ( n323614 , n320642 );
buf ( n323615 , n549 );
buf ( n323616 , n588 );
xor ( n323617 , n323615 , n323616 );
buf ( n323618 , n323617 );
buf ( n323619 , n323618 );
nand ( n323620 , n323614 , n323619 );
buf ( n323621 , n323620 );
buf ( n323622 , n323621 );
nand ( n323623 , n3770 , n323622 );
buf ( n323624 , n323623 );
buf ( n323625 , n323624 );
and ( n323626 , n323608 , n323625 );
and ( n323627 , n323586 , n323607 );
or ( n3785 , n323626 , n323627 );
buf ( n323629 , n3785 );
buf ( n323630 , n323629 );
xor ( n3788 , n323577 , n323630 );
buf ( n323632 , n3788 );
buf ( n323633 , n323632 );
xor ( n3791 , n323586 , n323607 );
xor ( n3792 , n3791 , n323625 );
buf ( n323636 , n3792 );
buf ( n323637 , n323636 );
xor ( n3795 , n323528 , n3703 );
xor ( n323639 , n3795 , n323571 );
buf ( n323640 , n323639 );
buf ( n323641 , n323640 );
xor ( n3799 , n323637 , n323641 );
not ( n323643 , n322455 );
not ( n3801 , n323643 );
not ( n3802 , n2642 );
or ( n323646 , n3801 , n3802 );
not ( n323647 , n2671 );
nand ( n323648 , n323646 , n323647 );
not ( n3806 , n323643 );
nand ( n323650 , n322482 , n3806 );
nand ( n323651 , n323648 , n323650 );
buf ( n323652 , n323651 );
and ( n323653 , n3799 , n323652 );
and ( n323654 , n323637 , n323641 );
or ( n3812 , n323653 , n323654 );
buf ( n323656 , n3812 );
buf ( n323657 , n323656 );
xor ( n323658 , n323633 , n323657 );
buf ( n323659 , n3696 );
not ( n323660 , n323659 );
buf ( n323661 , n323534 );
not ( n3819 , n323661 );
or ( n323663 , n323660 , n3819 );
buf ( n3821 , n322346 );
buf ( n323665 , n556 );
buf ( n323666 , n580 );
xor ( n323667 , n323665 , n323666 );
buf ( n323668 , n323667 );
buf ( n323669 , n323668 );
nand ( n323670 , n3821 , n323669 );
buf ( n323671 , n323670 );
buf ( n323672 , n323671 );
nand ( n323673 , n323663 , n323672 );
buf ( n323674 , n323673 );
buf ( n323675 , n323674 );
buf ( n3833 , n551 );
buf ( n3834 , n586 );
xor ( n3835 , n3833 , n3834 );
buf ( n3836 , n3835 );
buf ( n323680 , n3836 );
not ( n3838 , n323680 );
buf ( n323682 , n320692 );
not ( n323683 , n323682 );
or ( n3841 , n3838 , n323683 );
buf ( n323685 , n320699 );
xor ( n3843 , n586 , n550 );
buf ( n323687 , n3843 );
nand ( n3845 , n323685 , n323687 );
buf ( n323689 , n3845 );
buf ( n323690 , n323689 );
nand ( n323691 , n3841 , n323690 );
buf ( n323692 , n323691 );
buf ( n323693 , n323692 );
xor ( n3851 , n323675 , n323693 );
buf ( n323695 , n559 );
buf ( n323696 , n578 );
xor ( n3854 , n323695 , n323696 );
buf ( n323698 , n3854 );
buf ( n323699 , n323698 );
not ( n3857 , n323699 );
xor ( n3858 , n579 , n580 );
not ( n3859 , n3858 );
buf ( n323703 , n578 );
buf ( n323704 , n579 );
xor ( n323705 , n323703 , n323704 );
buf ( n323706 , n323705 );
nand ( n323707 , n3859 , n323706 );
not ( n3865 , n323707 );
buf ( n323709 , n3865 );
not ( n3867 , n323709 );
or ( n3868 , n3857 , n3867 );
not ( n3869 , n3858 );
buf ( n323713 , n3869 );
not ( n323714 , n323713 );
buf ( n323715 , n323714 );
buf ( n323716 , n323715 );
buf ( n3874 , n558 );
buf ( n3875 , n578 );
xor ( n3876 , n3874 , n3875 );
buf ( n323720 , n3876 );
buf ( n323721 , n323720 );
nand ( n3879 , n323716 , n323721 );
buf ( n3880 , n3879 );
buf ( n323724 , n3880 );
nand ( n3882 , n3868 , n323724 );
buf ( n3883 , n3882 );
buf ( n323727 , n3883 );
xor ( n323728 , n3851 , n323727 );
buf ( n323729 , n323728 );
buf ( n323730 , n323729 );
buf ( n323731 , n323618 );
not ( n323732 , n323731 );
buf ( n323733 , n898 );
not ( n323734 , n323733 );
or ( n3892 , n323732 , n323734 );
buf ( n323736 , n320642 );
buf ( n3894 , n548 );
buf ( n3895 , n588 );
xor ( n3896 , n3894 , n3895 );
buf ( n3897 , n3896 );
buf ( n323741 , n3897 );
nand ( n323742 , n323736 , n323741 );
buf ( n323743 , n323742 );
buf ( n323744 , n323743 );
nand ( n323745 , n3892 , n323744 );
buf ( n323746 , n323745 );
buf ( n323747 , n323746 );
buf ( n323748 , n3721 );
not ( n3906 , n323748 );
buf ( n323750 , n323550 );
not ( n3908 , n323750 );
or ( n323752 , n3906 , n3908 );
buf ( n323753 , n323559 );
not ( n3911 , n323753 );
buf ( n323755 , n3911 );
buf ( n3913 , n323755 );
buf ( n323757 , n554 );
buf ( n323758 , n582 );
xor ( n323759 , n323757 , n323758 );
buf ( n323760 , n323759 );
buf ( n323761 , n323760 );
nand ( n323762 , n3913 , n323761 );
buf ( n323763 , n323762 );
buf ( n323764 , n323763 );
nand ( n323765 , n323752 , n323764 );
buf ( n323766 , n323765 );
buf ( n323767 , n323766 );
xor ( n323768 , n323747 , n323767 );
buf ( n323769 , n3757 );
not ( n3927 , n323769 );
buf ( n323771 , n322176 );
not ( n3929 , n323771 );
or ( n3930 , n3927 , n3929 );
buf ( n323774 , n321209 );
buf ( n323775 , n552 );
buf ( n323776 , n584 );
xor ( n323777 , n323775 , n323776 );
buf ( n323778 , n323777 );
buf ( n323779 , n323778 );
nand ( n3937 , n323774 , n323779 );
buf ( n323781 , n3937 );
buf ( n323782 , n323781 );
nand ( n323783 , n3930 , n323782 );
buf ( n323784 , n323783 );
buf ( n323785 , n323784 );
xor ( n323786 , n323768 , n323785 );
buf ( n323787 , n323786 );
buf ( n323788 , n323787 );
xor ( n323789 , n323730 , n323788 );
buf ( n323790 , n322449 );
not ( n3948 , n323790 );
buf ( n323792 , n320692 );
not ( n323793 , n323792 );
or ( n3951 , n3948 , n323793 );
buf ( n323795 , n320699 );
buf ( n323796 , n3836 );
nand ( n3954 , n323795 , n323796 );
buf ( n323798 , n3954 );
buf ( n323799 , n323798 );
nand ( n323800 , n3951 , n323799 );
buf ( n323801 , n323800 );
buf ( n323802 , n323801 );
and ( n323803 , n322496 , n322510 );
buf ( n323804 , n323803 );
xor ( n323805 , n323802 , n323804 );
xor ( n3963 , n322552 , n322563 );
and ( n323807 , n3963 , n2732 );
and ( n323808 , n322552 , n322563 );
or ( n3966 , n323807 , n323808 );
buf ( n323810 , n3966 );
and ( n323811 , n323805 , n323810 );
and ( n3969 , n323802 , n323804 );
or ( n323813 , n323811 , n3969 );
buf ( n323814 , n323813 );
buf ( n323815 , n323814 );
xor ( n3973 , n323789 , n323815 );
buf ( n323817 , n3973 );
buf ( n323818 , n323817 );
and ( n323819 , n323658 , n323818 );
and ( n3977 , n323633 , n323657 );
or ( n3978 , n323819 , n3977 );
buf ( n323822 , n3978 );
buf ( n323823 , n323822 );
xor ( n323824 , n323485 , n323823 );
buf ( n323825 , n577 );
buf ( n323826 , n578 );
xor ( n3984 , n323825 , n323826 );
buf ( n323828 , n3984 );
buf ( n323829 , n323828 );
buf ( n323830 , n559 );
and ( n323831 , n323829 , n323830 );
buf ( n323832 , n323831 );
buf ( n323833 , n323832 );
buf ( n323834 , n323506 );
not ( n323835 , n323834 );
buf ( n323836 , n320732 );
not ( n3994 , n323836 );
or ( n323838 , n323835 , n3994 );
buf ( n323839 , n545 );
buf ( n323840 , n590 );
xor ( n323841 , n323839 , n323840 );
buf ( n323842 , n323841 );
buf ( n323843 , n323842 );
buf ( n323844 , n591 );
nand ( n323845 , n323843 , n323844 );
buf ( n323846 , n323845 );
buf ( n323847 , n323846 );
nand ( n4005 , n323838 , n323847 );
buf ( n323849 , n4005 );
buf ( n323850 , n323849 );
xor ( n4008 , n323833 , n323850 );
buf ( n323852 , n3897 );
not ( n4010 , n323852 );
buf ( n323854 , n926 );
not ( n4012 , n323854 );
or ( n4013 , n4010 , n4012 );
buf ( n323857 , n320642 );
buf ( n323858 , n547 );
buf ( n323859 , n588 );
xor ( n4017 , n323858 , n323859 );
buf ( n323861 , n4017 );
buf ( n323862 , n323861 );
nand ( n4020 , n323857 , n323862 );
buf ( n323864 , n4020 );
buf ( n323865 , n323864 );
nand ( n4023 , n4013 , n323865 );
buf ( n323867 , n4023 );
buf ( n323868 , n323867 );
xor ( n4026 , n4008 , n323868 );
buf ( n323870 , n4026 );
buf ( n323871 , n323870 );
xor ( n4029 , n323675 , n323693 );
and ( n323873 , n4029 , n323727 );
and ( n4031 , n323675 , n323693 );
or ( n323875 , n323873 , n4031 );
buf ( n323876 , n323875 );
buf ( n323877 , n323876 );
xor ( n323878 , n323871 , n323877 );
xor ( n323879 , n323747 , n323767 );
and ( n323880 , n323879 , n323785 );
and ( n4038 , n323747 , n323767 );
or ( n323882 , n323880 , n4038 );
buf ( n323883 , n323882 );
buf ( n323884 , n323883 );
xor ( n4042 , n323878 , n323884 );
buf ( n323886 , n4042 );
buf ( n323887 , n323886 );
buf ( n323888 , n323668 );
not ( n4046 , n323888 );
buf ( n323890 , n322468 );
not ( n323891 , n323890 );
or ( n323892 , n4046 , n323891 );
buf ( n323893 , n322474 );
buf ( n323894 , n555 );
buf ( n323895 , n580 );
xor ( n323896 , n323894 , n323895 );
buf ( n323897 , n323896 );
buf ( n323898 , n323897 );
nand ( n323899 , n323893 , n323898 );
buf ( n323900 , n323899 );
buf ( n323901 , n323900 );
nand ( n4059 , n323892 , n323901 );
buf ( n323903 , n4059 );
buf ( n323904 , n323903 );
buf ( n323905 , n323720 );
not ( n4063 , n323905 );
buf ( n323907 , n3865 );
not ( n323908 , n323907 );
or ( n323909 , n4063 , n323908 );
buf ( n323910 , n323715 );
buf ( n323911 , n557 );
buf ( n323912 , n578 );
xor ( n323913 , n323911 , n323912 );
buf ( n323914 , n323913 );
buf ( n323915 , n323914 );
nand ( n323916 , n323910 , n323915 );
buf ( n323917 , n323916 );
buf ( n323918 , n323917 );
nand ( n4076 , n323909 , n323918 );
buf ( n323920 , n4076 );
buf ( n323921 , n323920 );
xor ( n4079 , n323904 , n323921 );
and ( n4080 , n323501 , n323512 );
buf ( n323924 , n4080 );
buf ( n323925 , n323924 );
xor ( n323926 , n4079 , n323925 );
buf ( n323927 , n323926 );
buf ( n323928 , n323927 );
buf ( n323929 , n323778 );
not ( n323930 , n323929 );
buf ( n323931 , n321203 );
not ( n4089 , n323931 );
or ( n323933 , n323930 , n4089 );
buf ( n4091 , n1469 );
buf ( n323935 , n551 );
buf ( n323936 , n584 );
xor ( n323937 , n323935 , n323936 );
buf ( n323938 , n323937 );
buf ( n323939 , n323938 );
nand ( n323940 , n4091 , n323939 );
buf ( n323941 , n323940 );
buf ( n323942 , n323941 );
nand ( n323943 , n323933 , n323942 );
buf ( n323944 , n323943 );
buf ( n323945 , n323760 );
not ( n4103 , n323945 );
and ( n4104 , n583 , n582 );
not ( n323948 , n583 );
not ( n323949 , n582 );
and ( n323950 , n323948 , n323949 );
nor ( n4108 , n4104 , n323950 );
not ( n323952 , n4108 );
nor ( n323953 , n323952 , n322143 );
buf ( n323954 , n323953 );
not ( n323955 , n323954 );
or ( n4113 , n4103 , n323955 );
buf ( n4114 , n322143 );
buf ( n323958 , n4114 );
buf ( n323959 , n323958 );
buf ( n323960 , n323959 );
buf ( n323961 , n553 );
buf ( n323962 , n582 );
xor ( n4120 , n323961 , n323962 );
buf ( n323964 , n4120 );
buf ( n323965 , n323964 );
nand ( n4123 , n323960 , n323965 );
buf ( n323967 , n4123 );
buf ( n323968 , n323967 );
nand ( n323969 , n4113 , n323968 );
buf ( n323970 , n323969 );
xor ( n4128 , n323944 , n323970 );
buf ( n323972 , n3843 );
not ( n4130 , n323972 );
buf ( n323974 , n320692 );
not ( n323975 , n323974 );
or ( n323976 , n4130 , n323975 );
buf ( n323977 , n320699 );
xor ( n323978 , n586 , n549 );
buf ( n323979 , n323978 );
nand ( n4137 , n323977 , n323979 );
buf ( n323981 , n4137 );
buf ( n323982 , n323981 );
nand ( n4140 , n323976 , n323982 );
buf ( n323984 , n4140 );
xor ( n4142 , n4128 , n323984 );
buf ( n323986 , n4142 );
xor ( n323987 , n323928 , n323986 );
xor ( n323988 , n323515 , n323576 );
and ( n4146 , n323988 , n323630 );
and ( n4147 , n323515 , n323576 );
or ( n4148 , n4146 , n4147 );
buf ( n323992 , n4148 );
buf ( n323993 , n323992 );
xor ( n323994 , n323987 , n323993 );
buf ( n323995 , n323994 );
buf ( n323996 , n323995 );
xor ( n4154 , n323887 , n323996 );
xor ( n4155 , n323730 , n323788 );
and ( n4156 , n4155 , n323815 );
and ( n324000 , n323730 , n323788 );
or ( n324001 , n4156 , n324000 );
buf ( n324002 , n324001 );
buf ( n324003 , n324002 );
xor ( n4161 , n4154 , n324003 );
buf ( n324005 , n4161 );
buf ( n324006 , n324005 );
and ( n4164 , n323824 , n324006 );
and ( n324008 , n323485 , n323823 );
or ( n4166 , n4164 , n324008 );
buf ( n324010 , n4166 );
buf ( n324011 , n324010 );
xor ( n324012 , n323396 , n324011 );
xor ( n324013 , n323429 , n323433 );
and ( n4171 , n324013 , n323477 );
and ( n324015 , n323429 , n323433 );
or ( n324016 , n4171 , n324015 );
buf ( n324017 , n324016 );
buf ( n324018 , n324017 );
not ( n324019 , n324018 );
not ( n324020 , n323329 );
not ( n4178 , n324020 );
not ( n324022 , n323387 );
or ( n4180 , n4178 , n324022 );
nand ( n4181 , n323384 , n323329 );
nand ( n324025 , n4180 , n4181 );
and ( n324026 , n324025 , n323336 );
not ( n4184 , n324025 );
buf ( n324028 , n323336 );
not ( n324029 , n324028 );
buf ( n324030 , n324029 );
and ( n4188 , n4184 , n324030 );
nor ( n324032 , n324026 , n4188 );
buf ( n324033 , n324032 );
not ( n4191 , n324033 );
buf ( n4192 , n4191 );
buf ( n324036 , n4192 );
not ( n324037 , n324036 );
or ( n324038 , n324019 , n324037 );
buf ( n324039 , n4192 );
buf ( n324040 , n324017 );
or ( n324041 , n324039 , n324040 );
xor ( n4199 , n323081 , n323084 );
xor ( n4200 , n4199 , n323179 );
buf ( n324044 , n4200 );
buf ( n324045 , n324044 );
nand ( n324046 , n324041 , n324045 );
buf ( n324047 , n324046 );
buf ( n324048 , n324047 );
nand ( n324049 , n324038 , n324048 );
buf ( n324050 , n324049 );
buf ( n324051 , n324050 );
xor ( n324052 , n323887 , n323996 );
and ( n4210 , n324052 , n324003 );
and ( n324054 , n323887 , n323996 );
or ( n324055 , n4210 , n324054 );
buf ( n324056 , n324055 );
buf ( n4214 , n324056 );
xor ( n4215 , n324051 , n4214 );
not ( n324059 , n323897 );
not ( n324060 , n322468 );
or ( n4218 , n324059 , n324060 );
buf ( n324062 , n554 );
buf ( n324063 , n580 );
xor ( n4221 , n324062 , n324063 );
buf ( n4222 , n4221 );
nand ( n324066 , n322474 , n4222 );
nand ( n4224 , n4218 , n324066 );
buf ( n4225 , n323978 );
not ( n4226 , n4225 );
buf ( n4227 , n320692 );
not ( n4228 , n4227 );
or ( n4229 , n4226 , n4228 );
buf ( n4230 , n320699 );
xor ( n4231 , n586 , n548 );
buf ( n324075 , n4231 );
nand ( n324076 , n4230 , n324075 );
buf ( n324077 , n324076 );
buf ( n324078 , n324077 );
nand ( n4236 , n4229 , n324078 );
buf ( n4237 , n4236 );
xor ( n324081 , n4224 , n4237 );
buf ( n324082 , n323964 );
not ( n324083 , n324082 );
buf ( n324084 , n2327 );
not ( n4242 , n324084 );
or ( n324086 , n324083 , n4242 );
buf ( n324087 , n323562 );
buf ( n324088 , n552 );
buf ( n324089 , n582 );
xor ( n324090 , n324088 , n324089 );
buf ( n324091 , n324090 );
buf ( n324092 , n324091 );
nand ( n4250 , n324087 , n324092 );
buf ( n324094 , n4250 );
buf ( n324095 , n324094 );
nand ( n4253 , n324086 , n324095 );
buf ( n324097 , n4253 );
xor ( n4255 , n324081 , n324097 );
not ( n4256 , n4255 );
not ( n4257 , n4256 );
buf ( n324101 , n323861 );
not ( n4259 , n324101 );
buf ( n324103 , n926 );
not ( n4261 , n324103 );
or ( n324105 , n4259 , n4261 );
buf ( n324106 , n320642 );
buf ( n324107 , n546 );
buf ( n324108 , n588 );
xor ( n324109 , n324107 , n324108 );
buf ( n324110 , n324109 );
buf ( n324111 , n324110 );
nand ( n4269 , n324106 , n324111 );
buf ( n324113 , n4269 );
buf ( n324114 , n324113 );
nand ( n324115 , n324105 , n324114 );
buf ( n324116 , n324115 );
buf ( n4274 , n559 );
buf ( n4275 , n576 );
xor ( n4276 , n4274 , n4275 );
buf ( n4277 , n4276 );
buf ( n324121 , n4277 );
not ( n324122 , n324121 );
buf ( n324123 , n576 );
buf ( n324124 , n577 );
xnor ( n324125 , n324123 , n324124 );
buf ( n324126 , n324125 );
buf ( n324127 , n324126 );
buf ( n324128 , n323828 );
nor ( n4286 , n324127 , n324128 );
buf ( n324130 , n4286 );
buf ( n324131 , n324130 );
not ( n4289 , n324131 );
or ( n324133 , n324122 , n4289 );
buf ( n4291 , n323828 );
buf ( n324135 , n558 );
buf ( n324136 , n576 );
xor ( n324137 , n324135 , n324136 );
buf ( n324138 , n324137 );
buf ( n324139 , n324138 );
nand ( n324140 , n4291 , n324139 );
buf ( n324141 , n324140 );
buf ( n324142 , n324141 );
nand ( n324143 , n324133 , n324142 );
buf ( n324144 , n324143 );
xor ( n324145 , n324116 , n324144 );
buf ( n324146 , n323938 );
not ( n4304 , n324146 );
buf ( n324148 , n323591 );
not ( n4306 , n324148 );
or ( n4307 , n4304 , n4306 );
buf ( n324151 , n3752 );
buf ( n324152 , n550 );
buf ( n324153 , n584 );
xor ( n324154 , n324152 , n324153 );
buf ( n324155 , n324154 );
buf ( n324156 , n324155 );
nand ( n324157 , n324151 , n324156 );
buf ( n324158 , n324157 );
buf ( n324159 , n324158 );
nand ( n324160 , n4307 , n324159 );
buf ( n324161 , n324160 );
xor ( n4319 , n324145 , n324161 );
not ( n324163 , n323970 );
not ( n324164 , n323984 );
or ( n4322 , n324163 , n324164 );
nand ( n4323 , n321203 , n323778 );
not ( n4324 , n4323 );
not ( n4325 , n323941 );
or ( n4326 , n4324 , n4325 );
or ( n4327 , n323984 , n323970 );
nand ( n324171 , n4326 , n4327 );
nand ( n4329 , n4322 , n324171 );
and ( n324173 , n4319 , n4329 );
not ( n4331 , n4319 );
not ( n4332 , n4329 );
and ( n4333 , n4331 , n4332 );
nor ( n324177 , n324173 , n4333 );
not ( n324178 , n324177 );
or ( n4336 , n4257 , n324178 );
or ( n324180 , n324177 , n4256 );
nand ( n324181 , n4336 , n324180 );
buf ( n324182 , n324181 );
xor ( n4340 , n323928 , n323986 );
and ( n324184 , n4340 , n323993 );
and ( n324185 , n323928 , n323986 );
or ( n4343 , n324184 , n324185 );
buf ( n324187 , n4343 );
buf ( n324188 , n324187 );
xor ( n4346 , n324182 , n324188 );
xor ( n324190 , n323904 , n323921 );
and ( n324191 , n324190 , n323925 );
and ( n4349 , n323904 , n323921 );
or ( n324193 , n324191 , n4349 );
buf ( n324194 , n324193 );
buf ( n324195 , n324194 );
buf ( n324196 , n323914 );
not ( n4354 , n324196 );
buf ( n324198 , n3865 );
not ( n324199 , n324198 );
or ( n4357 , n4354 , n324199 );
buf ( n324201 , n323715 );
buf ( n324202 , n556 );
buf ( n324203 , n578 );
xor ( n4361 , n324202 , n324203 );
buf ( n324205 , n4361 );
buf ( n324206 , n324205 );
nand ( n4364 , n324201 , n324206 );
buf ( n324208 , n4364 );
buf ( n324209 , n324208 );
nand ( n4367 , n4357 , n324209 );
buf ( n324211 , n4367 );
buf ( n324212 , n324211 );
buf ( n324213 , n559 );
buf ( n324214 , n577 );
or ( n324215 , n324213 , n324214 );
buf ( n324216 , n578 );
nand ( n324217 , n324215 , n324216 );
buf ( n324218 , n324217 );
buf ( n324219 , n324218 );
buf ( n324220 , n559 );
buf ( n324221 , n577 );
nand ( n4379 , n324220 , n324221 );
buf ( n4380 , n4379 );
buf ( n324224 , n4380 );
buf ( n324225 , n576 );
and ( n4383 , n324219 , n324224 , n324225 );
buf ( n324227 , n4383 );
buf ( n324228 , n324227 );
buf ( n324229 , n323842 );
not ( n324230 , n324229 );
buf ( n324231 , n873 );
not ( n324232 , n324231 );
or ( n4390 , n324230 , n324232 );
buf ( n324234 , n544 );
buf ( n324235 , n590 );
xor ( n324236 , n324234 , n324235 );
buf ( n324237 , n324236 );
buf ( n324238 , n324237 );
buf ( n324239 , n591 );
nand ( n324240 , n324238 , n324239 );
buf ( n324241 , n324240 );
buf ( n324242 , n324241 );
nand ( n324243 , n4390 , n324242 );
buf ( n324244 , n324243 );
buf ( n324245 , n324244 );
xor ( n324246 , n324228 , n324245 );
buf ( n324247 , n324246 );
buf ( n324248 , n324247 );
xor ( n324249 , n324212 , n324248 );
xor ( n4407 , n323833 , n323850 );
and ( n324251 , n4407 , n323868 );
and ( n4409 , n323833 , n323850 );
or ( n4410 , n324251 , n4409 );
buf ( n324254 , n4410 );
buf ( n324255 , n324254 );
xor ( n324256 , n324249 , n324255 );
buf ( n324257 , n324256 );
buf ( n324258 , n324257 );
xor ( n4416 , n324195 , n324258 );
xor ( n4417 , n323871 , n323877 );
and ( n4418 , n4417 , n323884 );
and ( n4419 , n323871 , n323877 );
or ( n324263 , n4418 , n4419 );
buf ( n324264 , n324263 );
buf ( n324265 , n324264 );
xor ( n324266 , n4416 , n324265 );
buf ( n324267 , n324266 );
buf ( n324268 , n324267 );
xor ( n4426 , n4346 , n324268 );
buf ( n324270 , n4426 );
buf ( n324271 , n324270 );
xor ( n324272 , n4215 , n324271 );
buf ( n324273 , n324272 );
buf ( n324274 , n324273 );
xor ( n324275 , n324012 , n324274 );
buf ( n324276 , n324275 );
buf ( n324277 , n324276 );
xor ( n4435 , n324032 , n324017 );
xnor ( n4436 , n4435 , n324044 );
buf ( n324280 , n4436 );
not ( n324281 , n323456 );
not ( n324282 , n324281 );
not ( n4440 , n323446 );
or ( n324284 , n324282 , n4440 );
nand ( n4442 , n323449 , n323456 );
nand ( n4443 , n324284 , n4442 );
buf ( n4444 , n323464 );
and ( n4445 , n4443 , n4444 );
not ( n4446 , n4443 );
not ( n4447 , n4444 );
and ( n324291 , n4446 , n4447 );
nor ( n324292 , n4445 , n324291 );
not ( n324293 , n324292 );
buf ( n324294 , n324293 );
not ( n324295 , n324294 );
not ( n324296 , n321829 );
not ( n4454 , n321892 );
or ( n324298 , n324296 , n4454 );
not ( n4456 , n321829 );
not ( n4457 , n4456 );
not ( n324301 , n321892 );
not ( n4459 , n324301 );
or ( n324303 , n4457 , n4459 );
nand ( n4461 , n324303 , n321941 );
nand ( n324305 , n324298 , n4461 );
buf ( n324306 , n324305 );
not ( n324307 , n324306 );
or ( n324308 , n324295 , n324307 );
buf ( n324309 , n324292 );
not ( n4467 , n324309 );
buf ( n324311 , n324305 );
not ( n4469 , n324311 );
buf ( n324313 , n4469 );
buf ( n324314 , n324313 );
not ( n4472 , n324314 );
or ( n4473 , n4467 , n4472 );
not ( n4474 , n323403 );
xor ( n4475 , n3562 , n4474 );
xnor ( n4476 , n4475 , n323412 );
buf ( n324320 , n4476 );
nand ( n324321 , n4473 , n324320 );
buf ( n324322 , n324321 );
buf ( n324323 , n324322 );
nand ( n4481 , n324308 , n324323 );
buf ( n324325 , n4481 );
xor ( n324326 , n323802 , n323804 );
xor ( n324327 , n324326 , n323810 );
buf ( n324328 , n324327 );
buf ( n324329 , n324328 );
xor ( n4487 , n322536 , n322542 );
and ( n4488 , n4487 , n322576 );
and ( n4489 , n322536 , n322542 );
or ( n4490 , n4488 , n4489 );
buf ( n324334 , n4490 );
buf ( n324335 , n324334 );
xor ( n4493 , n324329 , n324335 );
xor ( n4494 , n323637 , n323641 );
xor ( n4495 , n4494 , n323652 );
buf ( n324339 , n4495 );
buf ( n324340 , n324339 );
and ( n4498 , n4493 , n324340 );
and ( n324342 , n324329 , n324335 );
or ( n324343 , n4498 , n324342 );
buf ( n324344 , n324343 );
xor ( n324345 , n324325 , n324344 );
xor ( n4503 , n323633 , n323657 );
xor ( n4504 , n4503 , n323818 );
buf ( n324348 , n4504 );
and ( n4506 , n324345 , n324348 );
and ( n4507 , n324325 , n324344 );
or ( n324351 , n4506 , n4507 );
buf ( n324352 , n324351 );
xor ( n324353 , n324280 , n324352 );
xor ( n4511 , n323485 , n323823 );
xor ( n324355 , n4511 , n324006 );
buf ( n324356 , n324355 );
buf ( n324357 , n324356 );
and ( n324358 , n324353 , n324357 );
and ( n4516 , n324280 , n324352 );
or ( n4517 , n324358 , n4516 );
buf ( n324361 , n4517 );
buf ( n324362 , n324361 );
nor ( n4520 , n324277 , n324362 );
buf ( n324364 , n4520 );
buf ( n324365 , n324364 );
xor ( n4523 , n324280 , n324352 );
xor ( n4524 , n4523 , n324357 );
buf ( n324368 , n4524 );
buf ( n324369 , n324368 );
xor ( n4527 , n323400 , n323417 );
xor ( n4528 , n4527 , n323480 );
buf ( n324372 , n4528 );
xor ( n324373 , n322514 , n322520 );
and ( n324374 , n324373 , n322579 );
and ( n4532 , n322514 , n322520 );
or ( n324376 , n324374 , n4532 );
buf ( n324377 , n324376 );
buf ( n324378 , n324377 );
xor ( n324379 , n321670 , n321823 );
and ( n324380 , n324379 , n321943 );
and ( n4538 , n321670 , n321823 );
or ( n324382 , n324380 , n4538 );
buf ( n324383 , n324382 );
buf ( n324384 , n324383 );
xor ( n324385 , n324378 , n324384 );
xor ( n4543 , n324329 , n324335 );
xor ( n324387 , n4543 , n324340 );
buf ( n324388 , n324387 );
buf ( n324389 , n324388 );
and ( n4547 , n324385 , n324389 );
and ( n324391 , n324378 , n324384 );
or ( n324392 , n4547 , n324391 );
buf ( n324393 , n324392 );
xor ( n324394 , n324372 , n324393 );
xor ( n4552 , n324325 , n324344 );
xor ( n4553 , n4552 , n324348 );
and ( n4554 , n324394 , n4553 );
and ( n4555 , n324372 , n324393 );
or ( n4556 , n4554 , n4555 );
buf ( n324400 , n4556 );
nor ( n324401 , n324369 , n324400 );
buf ( n324402 , n324401 );
buf ( n324403 , n324402 );
nor ( n4561 , n324365 , n324403 );
buf ( n324405 , n4561 );
xor ( n4563 , n324372 , n324393 );
xor ( n324407 , n4563 , n4553 );
buf ( n324408 , n324407 );
not ( n324409 , n324408 );
buf ( n324410 , n324409 );
buf ( n324411 , n324410 );
not ( n4569 , n321829 );
not ( n4570 , n321892 );
or ( n324414 , n4569 , n4570 );
nand ( n324415 , n324414 , n4461 );
xor ( n324416 , n324292 , n324415 );
xnor ( n4574 , n324416 , n4476 );
buf ( n324418 , n4574 );
xor ( n324419 , n322433 , n322438 );
and ( n4577 , n324419 , n322581 );
and ( n324421 , n322433 , n322438 );
or ( n324422 , n4577 , n324421 );
buf ( n324423 , n324422 );
xor ( n324424 , n324418 , n324423 );
xor ( n4582 , n324378 , n324384 );
xor ( n324426 , n4582 , n324389 );
buf ( n324427 , n324426 );
buf ( n324428 , n324427 );
and ( n4586 , n324424 , n324428 );
and ( n4587 , n324418 , n324423 );
or ( n4588 , n4586 , n4587 );
buf ( n4589 , n4588 );
buf ( n324433 , n4589 );
not ( n4591 , n324433 );
buf ( n324435 , n4591 );
buf ( n324436 , n324435 );
nand ( n4594 , n324411 , n324436 );
buf ( n324438 , n4594 );
buf ( n324439 , n324438 );
xor ( n4597 , n324418 , n324423 );
xor ( n324441 , n4597 , n324428 );
buf ( n324442 , n324441 );
buf ( n324443 , n324442 );
not ( n324444 , n324443 );
buf ( n324445 , n324444 );
buf ( n324446 , n324445 );
xor ( n324447 , n321945 , n322413 );
and ( n4605 , n324447 , n2740 );
and ( n324449 , n321945 , n322413 );
or ( n324450 , n4605 , n324449 );
buf ( n324451 , n324450 );
not ( n324452 , n324451 );
buf ( n324453 , n324452 );
buf ( n324454 , n324453 );
nand ( n4612 , n324446 , n324454 );
buf ( n324456 , n4612 );
buf ( n324457 , n324456 );
and ( n4615 , n324439 , n324457 );
buf ( n324459 , n4615 );
and ( n4617 , n324405 , n324459 );
not ( n4618 , n4617 );
or ( n4619 , n2972 , n4618 );
buf ( n324463 , n324402 );
not ( n4621 , n324463 );
buf ( n324465 , n324407 );
buf ( n324466 , n4589 );
or ( n324467 , n324465 , n324466 );
buf ( n324468 , n324467 );
buf ( n324469 , n324468 );
nand ( n4627 , n324407 , n4589 );
buf ( n324471 , n324442 );
buf ( n324472 , n324450 );
nand ( n324473 , n324471 , n324472 );
buf ( n324474 , n324473 );
nand ( n324475 , n4627 , n324474 );
buf ( n324476 , n324475 );
nand ( n324477 , n4621 , n324469 , n324476 );
buf ( n324478 , n324477 );
not ( n324479 , n324478 );
not ( n4637 , n324361 );
not ( n4638 , n324276 );
or ( n4639 , n4637 , n4638 );
buf ( n324483 , n324368 );
buf ( n324484 , n4556 );
nand ( n4642 , n324483 , n324484 );
buf ( n324486 , n4642 );
nand ( n4644 , n4639 , n324486 );
not ( n4645 , n4644 );
not ( n4646 , n4645 );
or ( n4647 , n324479 , n4646 );
buf ( n324491 , n324364 );
not ( n4649 , n324491 );
buf ( n324493 , n4649 );
nand ( n4651 , n4647 , n324493 );
nand ( n4652 , n4619 , n4651 );
not ( n4653 , n4652 );
not ( n4654 , n4653 );
buf ( n324498 , n4654 );
not ( n4656 , n324498 );
xor ( n4657 , n570 , n544 );
not ( n4658 , n4657 );
not ( n4659 , n320476 );
or ( n4660 , n4658 , n4659 );
buf ( n324504 , n320483 );
buf ( n324505 , n570 );
nand ( n4663 , n324504 , n324505 );
buf ( n324507 , n4663 );
nand ( n4665 , n4660 , n324507 );
buf ( n324509 , n4665 );
not ( n4667 , n324509 );
buf ( n324511 , n4667 );
buf ( n324512 , n324511 );
buf ( n324513 , n556 );
buf ( n324514 , n560 );
and ( n4672 , n324513 , n324514 );
buf ( n324516 , n4672 );
buf ( n324517 , n324516 );
buf ( n324518 , n547 );
buf ( n324519 , n568 );
xor ( n4677 , n324518 , n324519 );
buf ( n324521 , n4677 );
buf ( n324522 , n324521 );
not ( n4680 , n324522 );
xnor ( n4681 , n568 , n569 );
nor ( n4682 , n4681 , n320496 );
buf ( n324526 , n4682 );
not ( n4684 , n324526 );
or ( n324528 , n4680 , n4684 );
buf ( n324529 , n320499 );
buf ( n4687 , n546 );
buf ( n324531 , n568 );
xor ( n324532 , n4687 , n324531 );
buf ( n324533 , n324532 );
buf ( n324534 , n324533 );
nand ( n324535 , n324529 , n324534 );
buf ( n324536 , n324535 );
buf ( n324537 , n324536 );
nand ( n4695 , n324528 , n324537 );
buf ( n324539 , n4695 );
buf ( n324540 , n324539 );
xor ( n4698 , n324517 , n324540 );
xor ( n4699 , n564 , n551 );
buf ( n324543 , n4699 );
not ( n4701 , n324543 );
buf ( n324545 , n1850 );
not ( n4703 , n324545 );
or ( n4704 , n4701 , n4703 );
buf ( n324548 , n1857 );
buf ( n324549 , n550 );
buf ( n324550 , n564 );
xor ( n324551 , n324549 , n324550 );
buf ( n324552 , n324551 );
buf ( n324553 , n324552 );
nand ( n324554 , n324548 , n324553 );
buf ( n324555 , n324554 );
buf ( n324556 , n324555 );
nand ( n324557 , n4704 , n324556 );
buf ( n324558 , n324557 );
buf ( n324559 , n324558 );
and ( n4717 , n4698 , n324559 );
and ( n4718 , n324517 , n324540 );
or ( n4719 , n4717 , n4718 );
buf ( n324563 , n4719 );
buf ( n324564 , n324563 );
xor ( n4722 , n324512 , n324564 );
xor ( n4723 , n570 , n545 );
not ( n4724 , n4723 );
not ( n4725 , n3110 );
or ( n4726 , n4724 , n4725 );
nand ( n4727 , n320480 , n4657 );
nand ( n4728 , n4726 , n4727 );
not ( n4729 , n3304 );
not ( n4730 , n320528 );
or ( n4731 , n4729 , n4730 );
nand ( n4732 , n4731 , n572 );
xor ( n4733 , n4728 , n4732 );
buf ( n324577 , n549 );
buf ( n324578 , n566 );
xor ( n4736 , n324577 , n324578 );
buf ( n324580 , n4736 );
buf ( n324581 , n324580 );
not ( n4739 , n324581 );
buf ( n324583 , n1975 );
not ( n324584 , n324583 );
or ( n324585 , n4739 , n324584 );
buf ( n324586 , n548 );
buf ( n324587 , n566 );
xor ( n4742 , n324586 , n324587 );
buf ( n324589 , n4742 );
buf ( n324590 , n324589 );
buf ( n324591 , n321771 );
nand ( n4746 , n324590 , n324591 );
buf ( n324593 , n4746 );
buf ( n324594 , n324593 );
nand ( n4749 , n324585 , n324594 );
buf ( n324596 , n4749 );
and ( n4751 , n4733 , n324596 );
and ( n4752 , n4728 , n4732 );
or ( n4753 , n4751 , n4752 );
buf ( n324600 , n4753 );
xor ( n4755 , n4722 , n324600 );
buf ( n324602 , n4755 );
buf ( n324603 , n557 );
buf ( n324604 , n560 );
and ( n4759 , n324603 , n324604 );
buf ( n324606 , n4759 );
buf ( n324607 , n324606 );
not ( n4762 , n321756 );
buf ( n324609 , n550 );
buf ( n324610 , n566 );
xor ( n4765 , n324609 , n324610 );
buf ( n324612 , n4765 );
not ( n4767 , n324612 );
or ( n4768 , n4762 , n4767 );
buf ( n324615 , n324580 );
buf ( n324616 , n321768 );
nand ( n4771 , n324615 , n324616 );
buf ( n324618 , n4771 );
nand ( n4773 , n4768 , n324618 );
buf ( n324620 , n4773 );
xor ( n4775 , n324607 , n324620 );
buf ( n324622 , n546 );
buf ( n324623 , n570 );
xor ( n4778 , n324622 , n324623 );
buf ( n324625 , n4778 );
not ( n4780 , n324625 );
not ( n324627 , n321032 );
or ( n4782 , n4780 , n324627 );
nand ( n324629 , n320480 , n4723 );
nand ( n4784 , n4782 , n324629 );
buf ( n324631 , n4784 );
and ( n4786 , n4775 , n324631 );
and ( n4787 , n324607 , n324620 );
or ( n4788 , n4786 , n4787 );
buf ( n324635 , n4788 );
buf ( n324636 , n324635 );
xor ( n4791 , n562 , n554 );
buf ( n324638 , n4791 );
not ( n4793 , n324638 );
buf ( n324640 , n323283 );
not ( n4795 , n324640 );
or ( n4796 , n4793 , n4795 );
buf ( n324643 , n323006 );
buf ( n324644 , n553 );
buf ( n324645 , n562 );
xor ( n4800 , n324644 , n324645 );
buf ( n324647 , n4800 );
buf ( n4802 , n324647 );
nand ( n4803 , n324643 , n4802 );
buf ( n4804 , n4803 );
buf ( n324651 , n4804 );
nand ( n324652 , n4796 , n324651 );
buf ( n324653 , n324652 );
buf ( n324654 , n324653 );
not ( n324655 , n324654 );
xor ( n324656 , n568 , n548 );
buf ( n324657 , n324656 );
not ( n324658 , n324657 );
buf ( n324659 , n4682 );
not ( n4814 , n324659 );
or ( n4815 , n324658 , n4814 );
buf ( n324662 , n320499 );
buf ( n324663 , n324521 );
nand ( n4818 , n324662 , n324663 );
buf ( n324665 , n4818 );
buf ( n324666 , n324665 );
nand ( n324667 , n4815 , n324666 );
buf ( n324668 , n324667 );
buf ( n324669 , n324668 );
not ( n324670 , n324669 );
or ( n4825 , n324655 , n324670 );
buf ( n324672 , n324668 );
buf ( n324673 , n324653 );
or ( n324674 , n324672 , n324673 );
xor ( n324675 , n564 , n552 );
not ( n4830 , n324675 );
not ( n324677 , n3091 );
or ( n4832 , n4830 , n324677 );
buf ( n324679 , n1857 );
buf ( n324680 , n4699 );
nand ( n4835 , n324679 , n324680 );
buf ( n4836 , n4835 );
nand ( n324683 , n4832 , n4836 );
buf ( n324684 , n324683 );
nand ( n4839 , n324674 , n324684 );
buf ( n324686 , n4839 );
buf ( n324687 , n324686 );
nand ( n324688 , n4825 , n324687 );
buf ( n324689 , n324688 );
buf ( n324690 , n324689 );
xor ( n324691 , n324636 , n324690 );
xor ( n324692 , n4728 , n4732 );
xor ( n4847 , n324692 , n324596 );
buf ( n324694 , n4847 );
and ( n324695 , n324691 , n324694 );
and ( n4850 , n324636 , n324690 );
or ( n324697 , n324695 , n4850 );
buf ( n324698 , n324697 );
xor ( n324699 , n324602 , n324698 );
buf ( n324700 , n324647 );
not ( n324701 , n324700 );
buf ( n324702 , n323283 );
not ( n4857 , n324702 );
or ( n324704 , n324701 , n4857 );
buf ( n4859 , n323006 );
buf ( n324706 , n552 );
buf ( n324707 , n562 );
xor ( n324708 , n324706 , n324707 );
buf ( n324709 , n324708 );
buf ( n324710 , n324709 );
nand ( n324711 , n4859 , n324710 );
buf ( n324712 , n324711 );
buf ( n324713 , n324712 );
nand ( n324714 , n324704 , n324713 );
buf ( n324715 , n324714 );
buf ( n324716 , n324715 );
not ( n324717 , n324716 );
buf ( n324718 , n324717 );
buf ( n324719 , n324718 );
not ( n324720 , n324719 );
buf ( n324721 , n555 );
buf ( n324722 , n560 );
xor ( n324723 , n324721 , n324722 );
buf ( n324724 , n324723 );
buf ( n324725 , n324724 );
not ( n4880 , n324725 );
not ( n324727 , n322848 );
and ( n324728 , n324727 , n3000 );
buf ( n324729 , n324728 );
not ( n4884 , n324729 );
or ( n324731 , n4880 , n4884 );
buf ( n4886 , n3010 );
buf ( n324733 , n554 );
buf ( n324734 , n560 );
xor ( n324735 , n324733 , n324734 );
buf ( n324736 , n324735 );
buf ( n324737 , n324736 );
nand ( n324738 , n4886 , n324737 );
buf ( n324739 , n324738 );
buf ( n324740 , n324739 );
nand ( n4895 , n324731 , n324740 );
buf ( n4896 , n4895 );
buf ( n324743 , n4896 );
not ( n4898 , n324743 );
buf ( n4899 , n4898 );
buf ( n324746 , n4899 );
not ( n4901 , n324746 );
or ( n324748 , n324720 , n4901 );
buf ( n324749 , n544 );
buf ( n324750 , n572 );
xor ( n324751 , n324749 , n324750 );
buf ( n324752 , n324751 );
buf ( n324753 , n324752 );
not ( n4908 , n324753 );
buf ( n324755 , n320531 );
not ( n4910 , n324755 );
or ( n4911 , n4908 , n4910 );
buf ( n324758 , n320535 );
buf ( n324759 , n572 );
nand ( n4914 , n324758 , n324759 );
buf ( n324761 , n4914 );
buf ( n324762 , n324761 );
nand ( n4917 , n4911 , n324762 );
buf ( n324764 , n4917 );
buf ( n324765 , n324764 );
nand ( n324766 , n324748 , n324765 );
buf ( n324767 , n324766 );
buf ( n324768 , n324767 );
buf ( n324769 , n4896 );
buf ( n324770 , n324715 );
nand ( n4925 , n324769 , n324770 );
buf ( n324772 , n4925 );
buf ( n324773 , n324772 );
nand ( n324774 , n324768 , n324773 );
buf ( n324775 , n324774 );
buf ( n324776 , n324775 );
buf ( n324777 , n324709 );
not ( n324778 , n324777 );
buf ( n324779 , n322994 );
buf ( n324780 , n322998 );
nor ( n324781 , n324779 , n324780 );
buf ( n324782 , n324781 );
buf ( n324783 , n324782 );
not ( n4938 , n324783 );
or ( n4939 , n324778 , n4938 );
buf ( n324786 , n323006 );
buf ( n324787 , n551 );
buf ( n324788 , n562 );
xor ( n324789 , n324787 , n324788 );
buf ( n324790 , n324789 );
buf ( n324791 , n324790 );
nand ( n324792 , n324786 , n324791 );
buf ( n324793 , n324792 );
buf ( n324794 , n324793 );
nand ( n324795 , n4939 , n324794 );
buf ( n324796 , n324795 );
not ( n4951 , n4682 );
not ( n4952 , n324533 );
or ( n4953 , n4951 , n4952 );
buf ( n324800 , n320499 );
buf ( n324801 , n545 );
buf ( n324802 , n568 );
xor ( n4957 , n324801 , n324802 );
buf ( n324804 , n4957 );
buf ( n324805 , n324804 );
nand ( n4960 , n324800 , n324805 );
buf ( n324807 , n4960 );
nand ( n324808 , n4953 , n324807 );
not ( n324809 , n3091 );
not ( n4964 , n324552 );
or ( n324811 , n324809 , n4964 );
buf ( n324812 , n1857 );
buf ( n324813 , n549 );
buf ( n324814 , n564 );
xor ( n4969 , n324813 , n324814 );
buf ( n324816 , n4969 );
buf ( n324817 , n324816 );
nand ( n324818 , n324812 , n324817 );
buf ( n324819 , n324818 );
nand ( n324820 , n324811 , n324819 );
xor ( n4975 , n324808 , n324820 );
xor ( n4976 , n324796 , n4975 );
buf ( n324823 , n4976 );
xor ( n4978 , n324776 , n324823 );
buf ( n324825 , n555 );
buf ( n324826 , n560 );
and ( n324827 , n324825 , n324826 );
buf ( n324828 , n324827 );
buf ( n324829 , n324828 );
buf ( n324830 , n324589 );
not ( n324831 , n324830 );
buf ( n324832 , n1975 );
not ( n324833 , n324832 );
or ( n324834 , n324831 , n324833 );
buf ( n324835 , n547 );
buf ( n324836 , n566 );
xor ( n324837 , n324835 , n324836 );
buf ( n324838 , n324837 );
buf ( n324839 , n324838 );
buf ( n324840 , n321771 );
nand ( n4995 , n324839 , n324840 );
buf ( n324842 , n4995 );
buf ( n324843 , n324842 );
nand ( n4998 , n324834 , n324843 );
buf ( n324845 , n4998 );
buf ( n5000 , n324845 );
xor ( n5001 , n324829 , n5000 );
buf ( n324848 , n324736 );
not ( n5003 , n324848 );
buf ( n324850 , n324728 );
not ( n5005 , n324850 );
or ( n324852 , n5003 , n5005 );
buf ( n5007 , n3010 );
buf ( n5008 , n5007 );
buf ( n324855 , n5008 );
buf ( n324856 , n324855 );
buf ( n324857 , n553 );
buf ( n324858 , n560 );
xor ( n324859 , n324857 , n324858 );
buf ( n324860 , n324859 );
buf ( n324861 , n324860 );
nand ( n324862 , n324856 , n324861 );
buf ( n324863 , n324862 );
buf ( n5018 , n324863 );
nand ( n5019 , n324852 , n5018 );
buf ( n5020 , n5019 );
buf ( n324867 , n5020 );
xor ( n324868 , n5001 , n324867 );
buf ( n324869 , n324868 );
buf ( n324870 , n324869 );
xor ( n324871 , n4978 , n324870 );
buf ( n324872 , n324871 );
and ( n324873 , n324699 , n324872 );
and ( n5028 , n324602 , n324698 );
or ( n324875 , n324873 , n5028 );
not ( n324876 , n324875 );
xor ( n5031 , n324829 , n5000 );
and ( n324878 , n5031 , n324867 );
and ( n5033 , n324829 , n5000 );
or ( n5034 , n324878 , n5033 );
buf ( n324881 , n5034 );
buf ( n5036 , n324881 );
buf ( n324883 , n324790 );
not ( n5038 , n324883 );
buf ( n324885 , n3157 );
not ( n324886 , n324885 );
or ( n5041 , n5038 , n324886 );
buf ( n324888 , n323009 );
buf ( n324889 , n550 );
buf ( n324890 , n562 );
xor ( n324891 , n324889 , n324890 );
buf ( n324892 , n324891 );
buf ( n324893 , n324892 );
nand ( n324894 , n324888 , n324893 );
buf ( n324895 , n324894 );
buf ( n324896 , n324895 );
nand ( n324897 , n5041 , n324896 );
buf ( n324898 , n324897 );
buf ( n324899 , n324838 );
not ( n5054 , n324899 );
buf ( n324901 , n1975 );
not ( n5056 , n324901 );
or ( n5057 , n5054 , n5056 );
buf ( n324904 , n546 );
buf ( n324905 , n566 );
xor ( n5060 , n324904 , n324905 );
buf ( n324907 , n5060 );
buf ( n324908 , n324907 );
buf ( n324909 , n321771 );
nand ( n5064 , n324908 , n324909 );
buf ( n5065 , n5064 );
buf ( n324912 , n5065 );
nand ( n324913 , n5057 , n324912 );
buf ( n324914 , n324913 );
not ( n5069 , n324914 );
xor ( n324916 , n324898 , n5069 );
xor ( n324917 , n561 , n560 );
and ( n5072 , n324727 , n324860 , n324917 );
buf ( n324919 , n552 );
buf ( n324920 , n560 );
xor ( n5075 , n324919 , n324920 );
buf ( n324922 , n5075 );
and ( n5077 , n324855 , n324922 );
nor ( n324924 , n5072 , n5077 );
xor ( n324925 , n324916 , n324924 );
buf ( n5080 , n324925 );
xor ( n5081 , n5036 , n5080 );
buf ( n324928 , n320483 );
buf ( n324929 , n320475 );
or ( n5084 , n324928 , n324929 );
buf ( n324931 , n570 );
nand ( n5086 , n5084 , n324931 );
buf ( n324933 , n5086 );
buf ( n5088 , n324933 );
buf ( n324935 , n324816 );
not ( n5090 , n324935 );
buf ( n324937 , n321592 );
not ( n5092 , n324937 );
or ( n5093 , n5090 , n5092 );
buf ( n324940 , n3186 );
buf ( n324941 , n548 );
buf ( n324942 , n564 );
xor ( n5097 , n324941 , n324942 );
buf ( n324944 , n5097 );
buf ( n324945 , n324944 );
nand ( n5100 , n324940 , n324945 );
buf ( n324947 , n5100 );
buf ( n324948 , n324947 );
nand ( n5103 , n5093 , n324948 );
buf ( n324950 , n5103 );
not ( n5105 , n324950 );
xor ( n5106 , n5088 , n5105 );
buf ( n324953 , n324804 );
not ( n5108 , n324953 );
buf ( n324955 , n321072 );
not ( n5110 , n324955 );
or ( n5111 , n5108 , n5110 );
buf ( n324958 , n1339 );
buf ( n324959 , n544 );
buf ( n324960 , n568 );
xor ( n5115 , n324959 , n324960 );
buf ( n324962 , n5115 );
buf ( n324963 , n324962 );
nand ( n5118 , n324958 , n324963 );
buf ( n324965 , n5118 );
buf ( n324966 , n324965 );
nand ( n5121 , n5111 , n324966 );
buf ( n324968 , n5121 );
not ( n5123 , n324968 );
not ( n324970 , n5123 );
xnor ( n324971 , n5106 , n324970 );
buf ( n324972 , n324971 );
xor ( n5127 , n5081 , n324972 );
buf ( n324974 , n5127 );
not ( n324975 , n324974 );
buf ( n324976 , n554 );
buf ( n324977 , n560 );
and ( n5132 , n324976 , n324977 );
buf ( n324979 , n5132 );
buf ( n5134 , n324979 );
buf ( n5135 , n4665 );
xor ( n5136 , n5134 , n5135 );
or ( n324983 , n324796 , n324808 );
nand ( n5138 , n324983 , n324820 );
nand ( n5139 , n324796 , n324808 );
nand ( n5140 , n5138 , n5139 );
buf ( n324987 , n5140 );
xor ( n5142 , n5136 , n324987 );
buf ( n324989 , n5142 );
buf ( n324990 , n324989 );
xor ( n5145 , n324512 , n324564 );
and ( n324992 , n5145 , n324600 );
and ( n324993 , n324512 , n324564 );
or ( n5148 , n324992 , n324993 );
buf ( n324995 , n5148 );
buf ( n324996 , n324995 );
xor ( n5151 , n324990 , n324996 );
xor ( n324998 , n324776 , n324823 );
and ( n324999 , n324998 , n324870 );
and ( n5154 , n324776 , n324823 );
or ( n325001 , n324999 , n5154 );
buf ( n325002 , n325001 );
buf ( n325003 , n325002 );
xor ( n5158 , n5151 , n325003 );
buf ( n325005 , n5158 );
nand ( n325006 , n324876 , n324975 , n325005 );
not ( n325007 , n324875 );
not ( n5162 , n325005 );
nand ( n325009 , n325007 , n5162 , n324974 );
nand ( n5164 , n5162 , n324875 , n324975 );
nand ( n5165 , n324974 , n325005 , n324875 );
nand ( n5166 , n325006 , n325009 , n5164 , n5165 );
xor ( n5167 , n560 , n556 );
buf ( n325014 , n5167 );
not ( n5169 , n325014 );
buf ( n325016 , n324728 );
not ( n5171 , n325016 );
or ( n325018 , n5169 , n5171 );
buf ( n325019 , n3010 );
buf ( n325020 , n324724 );
nand ( n5175 , n325019 , n325020 );
buf ( n325022 , n5175 );
buf ( n325023 , n325022 );
nand ( n5178 , n325018 , n325023 );
buf ( n325025 , n5178 );
buf ( n325026 , n325025 );
not ( n5181 , n325026 );
buf ( n325028 , n5181 );
buf ( n325029 , n325028 );
not ( n5184 , n325029 );
buf ( n325031 , n549 );
buf ( n325032 , n568 );
xor ( n5187 , n325031 , n325032 );
buf ( n325034 , n5187 );
buf ( n325035 , n325034 );
not ( n5190 , n325035 );
buf ( n325037 , n321069 );
not ( n5192 , n325037 );
or ( n5193 , n5190 , n5192 );
buf ( n325040 , n1339 );
buf ( n325041 , n324656 );
nand ( n5196 , n325040 , n325041 );
buf ( n325043 , n5196 );
buf ( n325044 , n325043 );
nand ( n5199 , n5193 , n325044 );
buf ( n325046 , n5199 );
buf ( n325047 , n325046 );
not ( n5202 , n325047 );
buf ( n325049 , n5202 );
buf ( n325050 , n325049 );
not ( n5205 , n325050 );
or ( n5206 , n5184 , n5205 );
not ( n5207 , n324764 );
buf ( n325054 , n5207 );
nand ( n5209 , n5206 , n325054 );
buf ( n325056 , n5209 );
buf ( n325057 , n325056 );
buf ( n325058 , n325046 );
buf ( n325059 , n325025 );
nand ( n5214 , n325058 , n325059 );
buf ( n325061 , n5214 );
buf ( n325062 , n325061 );
nand ( n5217 , n325057 , n325062 );
buf ( n325064 , n5217 );
buf ( n325065 , n325064 );
xor ( n5220 , n324517 , n324540 );
xor ( n5221 , n5220 , n324559 );
buf ( n325068 , n5221 );
buf ( n325069 , n325068 );
xor ( n5224 , n325065 , n325069 );
buf ( n325071 , n324715 );
not ( n5226 , n325071 );
buf ( n325073 , n4899 );
not ( n5228 , n325073 );
or ( n5229 , n5226 , n5228 );
buf ( n325076 , n324718 );
buf ( n325077 , n4896 );
nand ( n5232 , n325076 , n325077 );
buf ( n325079 , n5232 );
buf ( n325080 , n325079 );
nand ( n5235 , n5229 , n325080 );
buf ( n325082 , n5235 );
buf ( n325083 , n325082 );
buf ( n325084 , n324764 );
and ( n5239 , n325083 , n325084 );
not ( n5240 , n325083 );
buf ( n325087 , n5207 );
and ( n5242 , n5240 , n325087 );
nor ( n5243 , n5239 , n5242 );
buf ( n325090 , n5243 );
buf ( n325091 , n325090 );
and ( n5246 , n5224 , n325091 );
and ( n5247 , n325065 , n325069 );
or ( n5248 , n5246 , n5247 );
buf ( n325095 , n5248 );
not ( n5250 , n325095 );
xor ( n5251 , n324668 , n324683 );
not ( n5252 , n5251 );
not ( n5253 , n324653 );
or ( n5254 , n5252 , n5253 );
not ( n5255 , n5251 );
not ( n5256 , n324653 );
nand ( n5257 , n5255 , n5256 );
nand ( n5258 , n5254 , n5257 );
not ( n5259 , n5258 );
not ( n5260 , n5259 );
buf ( n325107 , n558 );
buf ( n325108 , n560 );
and ( n5263 , n325107 , n325108 );
buf ( n325110 , n5263 );
buf ( n325111 , n325110 );
buf ( n325112 , n574 );
not ( n5267 , n325112 );
buf ( n325114 , n5267 );
buf ( n325115 , n325114 );
xor ( n5270 , n325111 , n325115 );
xor ( n5271 , n560 , n557 );
buf ( n325118 , n5271 );
not ( n5273 , n325118 );
buf ( n325120 , n3006 );
not ( n5275 , n325120 );
or ( n5276 , n5273 , n5275 );
buf ( n325123 , n3010 );
buf ( n325124 , n5167 );
nand ( n5279 , n325123 , n325124 );
buf ( n325126 , n5279 );
buf ( n325127 , n325126 );
nand ( n5282 , n5276 , n325127 );
buf ( n325129 , n5282 );
buf ( n325130 , n325129 );
and ( n5285 , n5270 , n325130 );
and ( n5286 , n325111 , n325115 );
or ( n5287 , n5285 , n5286 );
buf ( n325134 , n5287 );
not ( n5289 , n325134 );
or ( n5290 , n5260 , n5289 );
buf ( n325137 , n325134 );
not ( n5292 , n325137 );
buf ( n325139 , n5292 );
not ( n5294 , n325139 );
not ( n5295 , n5258 );
or ( n5296 , n5294 , n5295 );
buf ( n325143 , n547 );
buf ( n325144 , n570 );
xor ( n5299 , n325143 , n325144 );
buf ( n325146 , n5299 );
not ( n5301 , n325146 );
not ( n5302 , n3110 );
or ( n5303 , n5301 , n5302 );
buf ( n325150 , n320474 );
buf ( n325151 , n324625 );
nand ( n5306 , n325150 , n325151 );
buf ( n325153 , n5306 );
nand ( n5308 , n5303 , n325153 );
buf ( n325155 , n5308 );
not ( n5310 , n325155 );
xor ( n5311 , n566 , n551 );
buf ( n325158 , n5311 );
not ( n5313 , n325158 );
buf ( n325160 , n321756 );
not ( n5315 , n325160 );
or ( n5316 , n5313 , n5315 );
buf ( n325163 , n321768 );
buf ( n325164 , n324612 );
nand ( n5319 , n325163 , n325164 );
buf ( n325166 , n5319 );
buf ( n325167 , n325166 );
nand ( n5322 , n5316 , n325167 );
buf ( n325169 , n5322 );
buf ( n325170 , n325169 );
not ( n5325 , n325170 );
or ( n5326 , n5310 , n5325 );
buf ( n325173 , n325169 );
buf ( n325174 , n5308 );
or ( n5329 , n325173 , n325174 );
xor ( n5330 , n572 , n545 );
buf ( n325177 , n5330 );
not ( n5332 , n325177 );
buf ( n325179 , n3301 );
not ( n5334 , n325179 );
or ( n5335 , n5332 , n5334 );
buf ( n325182 , n320525 );
buf ( n325183 , n324752 );
nand ( n5338 , n325182 , n325183 );
buf ( n325185 , n5338 );
buf ( n325186 , n325185 );
nand ( n5341 , n5335 , n325186 );
buf ( n325188 , n5341 );
buf ( n325189 , n325188 );
nand ( n5344 , n5329 , n325189 );
buf ( n325191 , n5344 );
buf ( n325192 , n325191 );
nand ( n5347 , n5326 , n325192 );
buf ( n325194 , n5347 );
nand ( n5349 , n5296 , n325194 );
nand ( n5350 , n5290 , n5349 );
buf ( n325197 , n5350 );
xor ( n5352 , n324636 , n324690 );
xor ( n5353 , n5352 , n324694 );
buf ( n325200 , n5353 );
buf ( n325201 , n325200 );
xor ( n5356 , n325197 , n325201 );
buf ( n325203 , n559 );
buf ( n325204 , n560 );
and ( n5359 , n325203 , n325204 );
buf ( n325206 , n5359 );
buf ( n325207 , n325206 );
buf ( n325208 , n323223 );
not ( n5363 , n325208 );
buf ( n325210 , n320441 );
not ( n5365 , n325210 );
or ( n5366 , n5363 , n5365 );
buf ( n325213 , n574 );
buf ( n325214 , n575 );
nand ( n5369 , n325213 , n325214 );
buf ( n325216 , n5369 );
buf ( n325217 , n325216 );
nand ( n5372 , n5366 , n325217 );
buf ( n325219 , n5372 );
buf ( n325220 , n325219 );
xor ( n5375 , n325207 , n325220 );
buf ( n325222 , n2983 );
not ( n325223 , n325222 );
buf ( n325224 , n3301 );
not ( n325225 , n325224 );
or ( n325226 , n325223 , n325225 );
buf ( n325227 , n320525 );
buf ( n325228 , n5330 );
nand ( n5383 , n325227 , n325228 );
buf ( n325230 , n5383 );
buf ( n325231 , n325230 );
nand ( n325232 , n325226 , n325231 );
buf ( n325233 , n325232 );
buf ( n325234 , n325233 );
and ( n325235 , n5375 , n325234 );
and ( n325236 , n325207 , n325220 );
or ( n5391 , n325235 , n325236 );
buf ( n325238 , n5391 );
buf ( n325239 , n325238 );
not ( n5394 , n322879 );
not ( n5395 , n4682 );
or ( n5396 , n5394 , n5395 );
buf ( n325243 , n320499 );
buf ( n325244 , n325034 );
nand ( n5399 , n325243 , n325244 );
buf ( n325246 , n5399 );
nand ( n5401 , n5396 , n325246 );
not ( n5402 , n5401 );
not ( n5403 , n3125 );
not ( n5404 , n2105 );
or ( n5405 , n5403 , n5404 );
nand ( n5406 , n5311 , n321768 );
nand ( n5407 , n5405 , n5406 );
not ( n325254 , n5407 );
or ( n5409 , n5402 , n325254 );
nor ( n5410 , n5401 , n5407 );
and ( n5411 , n3006 , n322858 );
buf ( n5412 , n3010 );
buf ( n5413 , n5271 );
and ( n5414 , n5412 , n5413 );
buf ( n5415 , n5414 );
nor ( n325262 , n5411 , n5415 );
or ( n5417 , n5410 , n325262 );
nand ( n325264 , n5409 , n5417 );
buf ( n325265 , n325264 );
xor ( n325266 , n325239 , n325265 );
buf ( n325267 , n322946 );
not ( n5422 , n325267 );
buf ( n325269 , n1850 );
not ( n325270 , n325269 );
or ( n325271 , n5422 , n325270 );
buf ( n325272 , n1857 );
xor ( n325273 , n564 , n553 );
buf ( n325274 , n325273 );
nand ( n5429 , n325272 , n325274 );
buf ( n5430 , n5429 );
buf ( n325277 , n5430 );
nand ( n5432 , n325271 , n325277 );
buf ( n5433 , n5432 );
not ( n325280 , n5433 );
buf ( n325281 , n3353 );
not ( n325282 , n325281 );
buf ( n325283 , n3156 );
not ( n5438 , n325283 );
or ( n325285 , n325282 , n5438 );
buf ( n325286 , n323006 );
xor ( n325287 , n562 , n555 );
buf ( n325288 , n325287 );
nand ( n5443 , n325286 , n325288 );
buf ( n325290 , n5443 );
buf ( n325291 , n325290 );
nand ( n5445 , n325285 , n325291 );
buf ( n325293 , n5445 );
not ( n5447 , n325293 );
or ( n5448 , n325280 , n5447 );
not ( n5449 , n3114 );
not ( n5450 , n321032 );
or ( n5451 , n5449 , n5450 );
buf ( n325299 , n320480 );
buf ( n325300 , n325146 );
nand ( n5454 , n325299 , n325300 );
buf ( n325302 , n5454 );
nand ( n325303 , n5451 , n325302 );
buf ( n325304 , n325303 );
not ( n325305 , n325304 );
buf ( n325306 , n325305 );
buf ( n325307 , n5433 );
buf ( n325308 , n325293 );
nor ( n325309 , n325307 , n325308 );
buf ( n325310 , n325309 );
or ( n325311 , n325306 , n325310 );
nand ( n325312 , n5448 , n325311 );
buf ( n325313 , n325312 );
and ( n5467 , n325266 , n325313 );
and ( n325315 , n325239 , n325265 );
or ( n325316 , n5467 , n325315 );
buf ( n325317 , n325316 );
buf ( n325318 , n325317 );
xor ( n325319 , n324607 , n324620 );
xor ( n5473 , n325319 , n324631 );
buf ( n325321 , n5473 );
buf ( n325322 , n325321 );
nor ( n325323 , n325318 , n325322 );
buf ( n325324 , n325323 );
buf ( n325325 , n325324 );
xnor ( n325326 , n325025 , n325049 );
buf ( n325327 , n325326 );
buf ( n325328 , n324764 );
and ( n325329 , n325327 , n325328 );
not ( n325330 , n325327 );
buf ( n325331 , n5207 );
and ( n325332 , n325330 , n325331 );
nor ( n5486 , n325329 , n325332 );
buf ( n325334 , n5486 );
buf ( n325335 , n325334 );
or ( n5489 , n325325 , n325335 );
buf ( n325337 , n325317 );
buf ( n325338 , n325321 );
nand ( n325339 , n325337 , n325338 );
buf ( n325340 , n325339 );
buf ( n325341 , n325340 );
nand ( n325342 , n5489 , n325341 );
buf ( n325343 , n325342 );
buf ( n325344 , n325343 );
and ( n325345 , n5356 , n325344 );
and ( n5499 , n325197 , n325201 );
or ( n5500 , n325345 , n5499 );
buf ( n325348 , n5500 );
not ( n325349 , n325348 );
or ( n5503 , n5250 , n325349 );
or ( n325351 , n325348 , n325095 );
xor ( n325352 , n324602 , n324698 );
xor ( n5506 , n325352 , n324872 );
nand ( n325354 , n325351 , n5506 );
nand ( n325355 , n5503 , n325354 );
buf ( n5509 , n325355 );
buf ( n325357 , n555 );
buf ( n325358 , n576 );
and ( n325359 , n325357 , n325358 );
buf ( n325360 , n325359 );
buf ( n325361 , n325360 );
xor ( n5515 , n582 , n548 );
buf ( n325363 , n5515 );
not ( n5516 , n325363 );
buf ( n325365 , n322554 );
not ( n325366 , n325365 );
or ( n5519 , n5516 , n325366 );
buf ( n325368 , n323755 );
buf ( n325369 , n547 );
buf ( n325370 , n582 );
xor ( n5523 , n325369 , n325370 );
buf ( n325372 , n5523 );
buf ( n325373 , n325372 );
nand ( n5526 , n325368 , n325373 );
buf ( n325375 , n5526 );
buf ( n325376 , n325375 );
nand ( n325377 , n5519 , n325376 );
buf ( n325378 , n325377 );
buf ( n325379 , n325378 );
xor ( n5532 , n325361 , n325379 );
buf ( n325381 , n554 );
buf ( n5534 , n576 );
xor ( n5535 , n325381 , n5534 );
buf ( n325384 , n5535 );
buf ( n325385 , n325384 );
not ( n5538 , n325385 );
buf ( n325387 , n324126 );
buf ( n325388 , n323828 );
nor ( n325389 , n325387 , n325388 );
buf ( n325390 , n325389 );
buf ( n325391 , n325390 );
not ( n325392 , n325391 );
or ( n5545 , n5538 , n325392 );
buf ( n325394 , n323828 );
not ( n5547 , n325394 );
buf ( n325396 , n5547 );
buf ( n325397 , n325396 );
not ( n5550 , n325397 );
buf ( n325399 , n5550 );
buf ( n325400 , n325399 );
buf ( n325401 , n553 );
buf ( n325402 , n576 );
xor ( n5555 , n325401 , n325402 );
buf ( n325404 , n5555 );
buf ( n325405 , n325404 );
nand ( n5558 , n325400 , n325405 );
buf ( n325407 , n5558 );
buf ( n325408 , n325407 );
nand ( n5561 , n5545 , n325408 );
buf ( n325410 , n5561 );
buf ( n325411 , n325410 );
and ( n5564 , n5532 , n325411 );
and ( n5565 , n325361 , n325379 );
or ( n5566 , n5564 , n5565 );
buf ( n325415 , n5566 );
buf ( n325416 , n325415 );
buf ( n325417 , n325404 );
not ( n5570 , n325417 );
buf ( n325419 , n324126 );
buf ( n325420 , n323828 );
nor ( n325421 , n325419 , n325420 );
buf ( n325422 , n325421 );
buf ( n325423 , n325422 );
not ( n5576 , n325423 );
or ( n325425 , n5570 , n5576 );
buf ( n325426 , n323828 );
buf ( n5579 , n325426 );
buf ( n5580 , n5579 );
buf ( n325429 , n5580 );
buf ( n325430 , n552 );
buf ( n325431 , n576 );
xor ( n325432 , n325430 , n325431 );
buf ( n325433 , n325432 );
buf ( n325434 , n325433 );
nand ( n325435 , n325429 , n325434 );
buf ( n325436 , n325435 );
buf ( n325437 , n325436 );
nand ( n5590 , n325425 , n325437 );
buf ( n325439 , n5590 );
buf ( n325440 , n325439 );
buf ( n325441 , n551 );
buf ( n325442 , n578 );
xor ( n5595 , n325441 , n325442 );
buf ( n325444 , n5595 );
buf ( n325445 , n325444 );
not ( n5598 , n325445 );
buf ( n325447 , n3865 );
not ( n5600 , n325447 );
or ( n325449 , n5598 , n5600 );
buf ( n325450 , n323715 );
buf ( n325451 , n550 );
buf ( n325452 , n578 );
xor ( n325453 , n325451 , n325452 );
buf ( n325454 , n325453 );
buf ( n325455 , n325454 );
nand ( n325456 , n325450 , n325455 );
buf ( n325457 , n325456 );
buf ( n325458 , n325457 );
nand ( n325459 , n325449 , n325458 );
buf ( n325460 , n325459 );
buf ( n325461 , n325460 );
xor ( n325462 , n325440 , n325461 );
buf ( n325463 , n325372 );
not ( n325464 , n325463 );
buf ( n325465 , n322554 );
not ( n325466 , n325465 );
or ( n325467 , n325464 , n325466 );
buf ( n325468 , n323562 );
buf ( n325469 , n546 );
buf ( n325470 , n582 );
xor ( n5623 , n325469 , n325470 );
buf ( n325472 , n5623 );
buf ( n325473 , n325472 );
nand ( n5626 , n325468 , n325473 );
buf ( n5627 , n5626 );
buf ( n325476 , n5627 );
nand ( n5629 , n325467 , n325476 );
buf ( n5630 , n5629 );
buf ( n325479 , n5630 );
xor ( n325480 , n325462 , n325479 );
buf ( n325481 , n325480 );
buf ( n325482 , n325481 );
xor ( n325483 , n325416 , n325482 );
buf ( n325484 , n320692 );
buf ( n325485 , n320699 );
or ( n325486 , n325484 , n325485 );
buf ( n325487 , n586 );
nand ( n325488 , n325486 , n325487 );
buf ( n325489 , n325488 );
buf ( n325490 , n325489 );
buf ( n325491 , n549 );
buf ( n325492 , n580 );
xor ( n325493 , n325491 , n325492 );
buf ( n325494 , n325493 );
buf ( n325495 , n325494 );
not ( n325496 , n325495 );
not ( n325497 , n322468 );
not ( n5650 , n325497 );
buf ( n325499 , n5650 );
not ( n5652 , n325499 );
or ( n325501 , n325496 , n5652 );
buf ( n325502 , n322474 );
buf ( n325503 , n548 );
buf ( n325504 , n580 );
xor ( n5657 , n325503 , n325504 );
buf ( n325506 , n5657 );
buf ( n325507 , n325506 );
nand ( n5660 , n325502 , n325507 );
buf ( n325509 , n5660 );
buf ( n325510 , n325509 );
nand ( n5663 , n325501 , n325510 );
buf ( n325512 , n5663 );
buf ( n325513 , n325512 );
xor ( n325514 , n325490 , n325513 );
buf ( n325515 , n545 );
buf ( n325516 , n584 );
xor ( n325517 , n325515 , n325516 );
buf ( n325518 , n325517 );
buf ( n325519 , n325518 );
not ( n5672 , n325519 );
buf ( n325521 , n322176 );
not ( n5674 , n325521 );
or ( n5675 , n5672 , n5674 );
buf ( n325524 , n321209 );
buf ( n325525 , n544 );
buf ( n325526 , n584 );
xor ( n5679 , n325525 , n325526 );
buf ( n325528 , n5679 );
buf ( n325529 , n325528 );
nand ( n325530 , n325524 , n325529 );
buf ( n325531 , n325530 );
buf ( n325532 , n325531 );
nand ( n325533 , n5675 , n325532 );
buf ( n325534 , n325533 );
buf ( n325535 , n325534 );
xor ( n325536 , n325514 , n325535 );
buf ( n325537 , n325536 );
buf ( n325538 , n325537 );
xor ( n5691 , n325483 , n325538 );
buf ( n325540 , n5691 );
buf ( n325541 , n325540 );
not ( n325542 , n863 );
buf ( n5695 , n544 );
buf ( n5696 , n586 );
xor ( n5697 , n5695 , n5696 );
buf ( n5698 , n5697 );
not ( n325547 , n5698 );
or ( n5700 , n325542 , n325547 );
and ( n325549 , n587 , n586 );
not ( n5702 , n587 );
not ( n5703 , n586 );
and ( n5704 , n5702 , n5703 );
nor ( n325553 , n325549 , n5704 );
not ( n325554 , n863 );
and ( n5707 , n545 , n586 );
not ( n325556 , n545 );
not ( n325557 , n586 );
and ( n5710 , n325556 , n325557 );
nor ( n325559 , n5707 , n5710 );
nand ( n5712 , n325553 , n325554 , n325559 );
nand ( n325561 , n5700 , n5712 );
not ( n325562 , n325561 );
nand ( n325563 , n589 , n590 );
and ( n5716 , n325563 , n588 );
and ( n325565 , n325562 , n5716 );
not ( n5718 , n325562 );
not ( n5719 , n5716 );
and ( n325568 , n5718 , n5719 );
nor ( n5721 , n325565 , n325568 );
buf ( n325570 , n5721 );
xor ( n5723 , n582 , n549 );
buf ( n325572 , n5723 );
not ( n325573 , n325572 );
buf ( n325574 , n323953 );
not ( n325575 , n325574 );
or ( n325576 , n325573 , n325575 );
buf ( n325577 , n323959 );
buf ( n325578 , n5515 );
nand ( n5731 , n325577 , n325578 );
buf ( n325580 , n5731 );
buf ( n325581 , n325580 );
nand ( n5734 , n325576 , n325581 );
buf ( n325583 , n5734 );
buf ( n325584 , n325583 );
not ( n325585 , n325584 );
buf ( n325586 , n325585 );
buf ( n325587 , n325586 );
and ( n325588 , n325570 , n325587 );
not ( n5741 , n325570 );
buf ( n325590 , n325583 );
and ( n325591 , n5741 , n325590 );
nor ( n5744 , n325588 , n325591 );
buf ( n325593 , n5744 );
not ( n5746 , n325593 );
not ( n5747 , n5746 );
buf ( n325596 , n546 );
buf ( n325597 , n586 );
xor ( n5750 , n325596 , n325597 );
buf ( n325599 , n5750 );
not ( n5752 , n325599 );
not ( n5753 , n320692 );
or ( n5754 , n5752 , n5753 );
buf ( n325603 , n320699 );
buf ( n325604 , n325559 );
nand ( n325605 , n325603 , n325604 );
buf ( n325606 , n325605 );
nand ( n5759 , n5754 , n325606 );
not ( n325608 , n5759 );
and ( n5761 , n582 , n550 );
not ( n5762 , n582 );
not ( n5763 , n550 );
and ( n5764 , n5762 , n5763 );
nor ( n325613 , n5761 , n5764 );
buf ( n325614 , n325613 );
not ( n325615 , n325614 );
buf ( n325616 , n323953 );
not ( n325617 , n325616 );
or ( n325618 , n325615 , n325617 );
buf ( n325619 , n322143 );
buf ( n325620 , n5723 );
nand ( n5773 , n325619 , n325620 );
buf ( n325622 , n5773 );
buf ( n325623 , n325622 );
nand ( n5776 , n325618 , n325623 );
buf ( n325625 , n5776 );
buf ( n325626 , n557 );
buf ( n325627 , n576 );
nand ( n325628 , n325626 , n325627 );
buf ( n325629 , n325628 );
buf ( n325630 , n325629 );
not ( n325631 , n325630 );
buf ( n325632 , n325631 );
or ( n5785 , n325625 , n325632 );
not ( n5786 , n5785 );
or ( n5787 , n325608 , n5786 );
buf ( n325636 , n325625 );
buf ( n325637 , n325632 );
nand ( n5790 , n325636 , n325637 );
buf ( n325639 , n5790 );
nand ( n5792 , n5787 , n325639 );
not ( n5793 , n5792 );
or ( n5794 , n5747 , n5793 );
not ( n5795 , n5792 );
not ( n5796 , n5795 );
not ( n5797 , n325593 );
or ( n5798 , n5796 , n5797 );
xor ( n325647 , n584 , n548 );
buf ( n325648 , n325647 );
not ( n325649 , n325648 );
buf ( n325650 , n321203 );
not ( n325651 , n325650 );
or ( n325652 , n325649 , n325651 );
buf ( n325653 , n3752 );
xor ( n325654 , n584 , n547 );
buf ( n325655 , n325654 );
nand ( n5808 , n325653 , n325655 );
buf ( n325657 , n5808 );
buf ( n325658 , n325657 );
nand ( n5811 , n325652 , n325658 );
buf ( n325660 , n5811 );
buf ( n325661 , n325660 );
not ( n5814 , n325661 );
xor ( n325663 , n580 , n551 );
and ( n325664 , n322346 , n325663 );
not ( n5817 , n322346 );
xor ( n325666 , n580 , n552 );
and ( n5819 , n581 , n580 );
not ( n5820 , n581 );
not ( n5821 , n580 );
and ( n5822 , n5820 , n5821 );
nor ( n325671 , n5819 , n5822 );
and ( n325672 , n325666 , n325671 );
and ( n325673 , n5817 , n325672 );
or ( n5826 , n325664 , n325673 );
buf ( n325675 , n5826 );
not ( n325676 , n325675 );
or ( n5829 , n5814 , n325676 );
buf ( n325678 , n325660 );
buf ( n325679 , n5826 );
or ( n5832 , n325678 , n325679 );
xor ( n325681 , n578 , n554 );
buf ( n325682 , n325681 );
not ( n325683 , n325682 );
not ( n5836 , n323706 );
nor ( n325685 , n5836 , n3738 );
buf ( n325686 , n325685 );
not ( n5839 , n325686 );
or ( n325688 , n325683 , n5839 );
buf ( n325689 , n3738 );
and ( n5842 , n578 , n553 );
not ( n325691 , n578 );
and ( n325692 , n325691 , n320512 );
nor ( n5845 , n5842 , n325692 );
buf ( n325694 , n5845 );
nand ( n5847 , n325689 , n325694 );
buf ( n325696 , n5847 );
buf ( n325697 , n325696 );
nand ( n5850 , n325688 , n325697 );
buf ( n325699 , n5850 );
buf ( n325700 , n325699 );
nand ( n325701 , n5832 , n325700 );
buf ( n325702 , n325701 );
buf ( n325703 , n325702 );
nand ( n325704 , n5829 , n325703 );
buf ( n325705 , n325704 );
nand ( n325706 , n5798 , n325705 );
nand ( n325707 , n5794 , n325706 );
buf ( n325708 , n325707 );
buf ( n325709 , n5698 );
not ( n325710 , n325709 );
buf ( n325711 , n320692 );
not ( n325712 , n325711 );
or ( n325713 , n325710 , n325712 );
buf ( n325714 , n320699 );
buf ( n325715 , n586 );
nand ( n5868 , n325714 , n325715 );
buf ( n325717 , n5868 );
buf ( n325718 , n325717 );
nand ( n5871 , n325713 , n325718 );
buf ( n325720 , n5871 );
buf ( n325721 , n325720 );
not ( n5874 , n325721 );
buf ( n325723 , n5874 );
buf ( n5876 , n325723 );
nor ( n325725 , n325561 , n325583 );
or ( n5878 , n325725 , n5716 );
nand ( n325727 , n325583 , n325561 );
nand ( n5880 , n5878 , n325727 );
buf ( n325729 , n5880 );
not ( n325730 , n325729 );
buf ( n325731 , n325730 );
buf ( n325732 , n325731 );
xor ( n5885 , n5876 , n325732 );
buf ( n325734 , n556 );
buf ( n325735 , n576 );
nand ( n5888 , n325734 , n325735 );
buf ( n325737 , n5888 );
not ( n325738 , n325737 );
buf ( n325739 , n325654 );
not ( n5892 , n325739 );
buf ( n325741 , n323591 );
not ( n325742 , n325741 );
or ( n5895 , n5892 , n325742 );
buf ( n325744 , n3752 );
buf ( n325745 , n546 );
buf ( n325746 , n584 );
xor ( n325747 , n325745 , n325746 );
buf ( n325748 , n325747 );
buf ( n325749 , n325748 );
nand ( n325750 , n325744 , n325749 );
buf ( n325751 , n325750 );
buf ( n325752 , n325751 );
nand ( n325753 , n5895 , n325752 );
buf ( n325754 , n325753 );
not ( n325755 , n325754 );
not ( n5908 , n325755 );
or ( n5909 , n325738 , n5908 );
not ( n325758 , n325663 );
not ( n325759 , n322468 );
or ( n5912 , n325758 , n325759 );
buf ( n325761 , n322474 );
buf ( n325762 , n550 );
buf ( n325763 , n580 );
xor ( n325764 , n325762 , n325763 );
buf ( n325765 , n325764 );
buf ( n325766 , n325765 );
nand ( n5919 , n325761 , n325766 );
buf ( n325768 , n5919 );
nand ( n5921 , n5912 , n325768 );
nand ( n325770 , n5909 , n5921 );
not ( n325771 , n325737 );
nand ( n5924 , n325771 , n325754 );
nand ( n5925 , n325770 , n5924 );
buf ( n325774 , n5925 );
xnor ( n325775 , n5885 , n325774 );
buf ( n325776 , n325775 );
buf ( n325777 , n325776 );
xor ( n5930 , n325708 , n325777 );
buf ( n325779 , n555 );
buf ( n325780 , n576 );
xor ( n5933 , n325779 , n325780 );
buf ( n325782 , n5933 );
buf ( n325783 , n325782 );
not ( n5936 , n325783 );
buf ( n325785 , n325422 );
not ( n5938 , n325785 );
or ( n5939 , n5936 , n5938 );
buf ( n5940 , n323828 );
buf ( n325789 , n325384 );
nand ( n5942 , n5940 , n325789 );
buf ( n325791 , n5942 );
buf ( n325792 , n325791 );
nand ( n325793 , n5939 , n325792 );
buf ( n325794 , n325793 );
xor ( n5947 , n588 , n544 );
not ( n5948 , n5947 );
not ( n5949 , n926 );
or ( n5950 , n5948 , n5949 );
nand ( n325799 , n588 , n320642 );
nand ( n325800 , n5950 , n325799 );
or ( n5953 , n325794 , n325800 );
not ( n325802 , n5845 );
not ( n5955 , n325685 );
or ( n325804 , n325802 , n5955 );
buf ( n325805 , n552 );
buf ( n325806 , n578 );
xor ( n325807 , n325805 , n325806 );
buf ( n325808 , n325807 );
nand ( n325809 , n323715 , n325808 );
nand ( n5962 , n325804 , n325809 );
nand ( n325811 , n5953 , n5962 );
buf ( n325812 , n325811 );
nand ( n5965 , n325794 , n325800 );
buf ( n325814 , n5965 );
nand ( n325815 , n325812 , n325814 );
buf ( n325816 , n325815 );
buf ( n325817 , n325816 );
buf ( n325818 , n325765 );
not ( n325819 , n325818 );
buf ( n325820 , n323534 );
not ( n5973 , n325820 );
or ( n325822 , n325819 , n5973 );
buf ( n325823 , n322346 );
buf ( n325824 , n325494 );
nand ( n5977 , n325823 , n325824 );
buf ( n325826 , n5977 );
buf ( n325827 , n325826 );
nand ( n5980 , n325822 , n325827 );
buf ( n325829 , n5980 );
buf ( n325830 , n325829 );
buf ( n325831 , n325808 );
not ( n325832 , n325831 );
buf ( n325833 , n325685 );
not ( n325834 , n325833 );
or ( n325835 , n325832 , n325834 );
buf ( n325836 , n3738 );
buf ( n325837 , n325444 );
nand ( n5990 , n325836 , n325837 );
buf ( n325839 , n5990 );
buf ( n325840 , n325839 );
nand ( n5993 , n325835 , n325840 );
buf ( n325842 , n5993 );
buf ( n5995 , n325842 );
xor ( n5996 , n325830 , n5995 );
buf ( n325845 , n325748 );
not ( n325846 , n325845 );
buf ( n325847 , n321203 );
not ( n6000 , n325847 );
or ( n325849 , n325846 , n6000 );
buf ( n325850 , n321209 );
buf ( n325851 , n325518 );
nand ( n325852 , n325850 , n325851 );
buf ( n325853 , n325852 );
buf ( n325854 , n325853 );
nand ( n6007 , n325849 , n325854 );
buf ( n325856 , n6007 );
buf ( n325857 , n325856 );
xor ( n325858 , n5996 , n325857 );
buf ( n325859 , n325858 );
buf ( n325860 , n325859 );
xor ( n6013 , n325817 , n325860 );
xor ( n325862 , n325361 , n325379 );
xor ( n6015 , n325862 , n325411 );
buf ( n325864 , n6015 );
buf ( n325865 , n325864 );
xor ( n6018 , n6013 , n325865 );
buf ( n325867 , n6018 );
buf ( n325868 , n325867 );
and ( n6021 , n5930 , n325868 );
and ( n6022 , n325708 , n325777 );
or ( n325871 , n6021 , n6022 );
buf ( n325872 , n325871 );
buf ( n6025 , n325872 );
xor ( n6026 , n325541 , n6025 );
buf ( n325875 , n325720 );
not ( n325876 , n325875 );
buf ( n325877 , n325731 );
not ( n325878 , n325877 );
or ( n325879 , n325876 , n325878 );
buf ( n325880 , n5925 );
nand ( n325881 , n325879 , n325880 );
buf ( n325882 , n325881 );
buf ( n325883 , n325882 );
buf ( n325884 , n5880 );
buf ( n325885 , n325723 );
nand ( n6038 , n325884 , n325885 );
buf ( n325887 , n6038 );
buf ( n325888 , n325887 );
nand ( n6041 , n325883 , n325888 );
buf ( n325890 , n6041 );
buf ( n325891 , n325890 );
buf ( n325892 , n554 );
buf ( n6045 , n576 );
and ( n6046 , n325892 , n6045 );
buf ( n6047 , n6046 );
buf ( n325896 , n6047 );
buf ( n325897 , n325720 );
xor ( n325898 , n325896 , n325897 );
xor ( n325899 , n325830 , n5995 );
and ( n6052 , n325899 , n325857 );
and ( n325901 , n325830 , n5995 );
or ( n325902 , n6052 , n325901 );
buf ( n325903 , n325902 );
buf ( n325904 , n325903 );
xor ( n325905 , n325898 , n325904 );
buf ( n325906 , n325905 );
buf ( n325907 , n325906 );
xor ( n325908 , n325891 , n325907 );
xor ( n6061 , n325817 , n325860 );
and ( n6062 , n6061 , n325865 );
and ( n325911 , n325817 , n325860 );
or ( n6064 , n6062 , n325911 );
buf ( n325913 , n6064 );
buf ( n325914 , n325913 );
xor ( n6067 , n325908 , n325914 );
buf ( n325916 , n6067 );
buf ( n325917 , n325916 );
xor ( n6070 , n6026 , n325917 );
buf ( n325919 , n6070 );
buf ( n325920 , n325919 );
xor ( n325921 , n5509 , n325920 );
xor ( n6074 , n325737 , n5921 );
xor ( n325923 , n6074 , n325754 );
buf ( n325924 , n325923 );
not ( n6077 , n325924 );
not ( n325926 , n325800 );
buf ( n6079 , n549 );
buf ( n325928 , n584 );
xor ( n6081 , n6079 , n325928 );
buf ( n325930 , n6081 );
buf ( n325931 , n325930 );
not ( n6084 , n325931 );
buf ( n325933 , n321203 );
not ( n325934 , n325933 );
or ( n325935 , n6084 , n325934 );
buf ( n325936 , n1469 );
buf ( n325937 , n325647 );
nand ( n325938 , n325936 , n325937 );
buf ( n325939 , n325938 );
buf ( n325940 , n325939 );
nand ( n325941 , n325935 , n325940 );
buf ( n325942 , n325941 );
xor ( n325943 , n325926 , n325942 );
buf ( n325944 , n556 );
buf ( n325945 , n576 );
xor ( n325946 , n325944 , n325945 );
buf ( n325947 , n325946 );
buf ( n325948 , n325947 );
not ( n6101 , n325948 );
buf ( n325950 , n325422 );
buf ( n325951 , n325950 );
buf ( n325952 , n325951 );
buf ( n325953 , n325952 );
not ( n6106 , n325953 );
or ( n325955 , n6101 , n6106 );
buf ( n325956 , n5580 );
buf ( n325957 , n325782 );
nand ( n325958 , n325956 , n325957 );
buf ( n325959 , n325958 );
buf ( n325960 , n325959 );
nand ( n325961 , n325955 , n325960 );
buf ( n325962 , n325961 );
and ( n6115 , n325943 , n325962 );
and ( n325964 , n325926 , n325942 );
or ( n6117 , n6115 , n325964 );
not ( n6118 , n6117 );
buf ( n325967 , n6118 );
not ( n6120 , n325967 );
or ( n6121 , n6077 , n6120 );
xnor ( n325970 , n5962 , n325794 );
xnor ( n6123 , n325970 , n325800 );
buf ( n325972 , n6123 );
nand ( n6125 , n6121 , n325972 );
buf ( n6126 , n6125 );
buf ( n325975 , n6126 );
buf ( n325976 , n325923 );
not ( n325977 , n325976 );
buf ( n325978 , n6117 );
nand ( n6131 , n325977 , n325978 );
buf ( n325980 , n6131 );
buf ( n6133 , n325980 );
nand ( n6134 , n325975 , n6133 );
buf ( n6135 , n6134 );
buf ( n325984 , n6135 );
xor ( n6137 , n325708 , n325777 );
xor ( n325986 , n6137 , n325868 );
buf ( n325987 , n325986 );
buf ( n325988 , n325987 );
xor ( n6141 , n325984 , n325988 );
buf ( n325990 , n558 );
buf ( n325991 , n576 );
and ( n325992 , n325990 , n325991 );
buf ( n325993 , n325992 );
buf ( n325994 , n325993 );
buf ( n325995 , n320740 );
xor ( n6148 , n325994 , n325995 );
buf ( n325997 , n557 );
buf ( n325998 , n576 );
xor ( n325999 , n325997 , n325998 );
buf ( n326000 , n325999 );
buf ( n326001 , n326000 );
not ( n6154 , n326001 );
buf ( n326003 , n325390 );
not ( n6156 , n326003 );
or ( n6157 , n6154 , n6156 );
buf ( n326006 , n325399 );
buf ( n326007 , n325947 );
nand ( n6160 , n326006 , n326007 );
buf ( n326009 , n6160 );
buf ( n326010 , n326009 );
nand ( n6163 , n6157 , n326010 );
buf ( n326012 , n6163 );
buf ( n326013 , n326012 );
and ( n6166 , n6148 , n326013 );
and ( n6167 , n325994 , n325995 );
or ( n6168 , n6166 , n6167 );
buf ( n326017 , n6168 );
buf ( n326018 , n326017 );
xor ( n6171 , n586 , n547 );
buf ( n326020 , n6171 );
not ( n6173 , n326020 );
buf ( n326022 , n320692 );
not ( n6175 , n326022 );
or ( n6176 , n6173 , n6175 );
buf ( n326025 , n320699 );
buf ( n326026 , n325599 );
nand ( n6179 , n326025 , n326026 );
buf ( n326028 , n6179 );
buf ( n326029 , n326028 );
nand ( n6182 , n6176 , n326029 );
buf ( n326031 , n6182 );
not ( n6184 , n326031 );
buf ( n326033 , n551 );
buf ( n326034 , n582 );
xor ( n326035 , n326033 , n326034 );
buf ( n326036 , n326035 );
not ( n326037 , n326036 );
not ( n6190 , n322144 );
or ( n326039 , n326037 , n6190 );
nand ( n6192 , n323558 , n325613 );
nand ( n6193 , n326039 , n6192 );
not ( n326042 , n6193 );
buf ( n326043 , n545 );
buf ( n326044 , n588 );
xor ( n326045 , n326043 , n326044 );
buf ( n326046 , n326045 );
not ( n6199 , n326046 );
not ( n326048 , n926 );
or ( n6201 , n6199 , n326048 );
buf ( n326050 , n320642 );
buf ( n6203 , n5947 );
nand ( n6204 , n326050 , n6203 );
buf ( n6205 , n6204 );
nand ( n326054 , n6201 , n6205 );
not ( n326055 , n326054 );
nand ( n6208 , n326042 , n326055 );
not ( n326057 , n6208 );
or ( n6210 , n6184 , n326057 );
buf ( n326059 , n6193 );
buf ( n326060 , n326054 );
nand ( n6213 , n326059 , n326060 );
buf ( n6214 , n6213 );
nand ( n326063 , n6210 , n6214 );
buf ( n326064 , n326063 );
xor ( n6217 , n326018 , n326064 );
xor ( n326066 , n5826 , n325699 );
xor ( n6219 , n326066 , n325660 );
buf ( n326068 , n6219 );
and ( n326069 , n6217 , n326068 );
and ( n6222 , n326018 , n326064 );
or ( n326071 , n326069 , n6222 );
buf ( n326072 , n326071 );
buf ( n326073 , n326072 );
xor ( n6226 , n5792 , n325705 );
xor ( n326075 , n6226 , n5746 );
buf ( n326076 , n326075 );
xor ( n326077 , n326073 , n326076 );
xor ( n326078 , n325625 , n5759 );
xnor ( n326079 , n326078 , n325629 );
buf ( n326080 , n326079 );
xor ( n326081 , n325926 , n325942 );
xor ( n6234 , n326081 , n325962 );
buf ( n326083 , n6234 );
xor ( n6236 , n326080 , n326083 );
not ( n326085 , n4231 );
not ( n6238 , n320692 );
or ( n6239 , n326085 , n6238 );
nand ( n326088 , n6171 , n863 );
nand ( n326089 , n6239 , n326088 );
not ( n6242 , n326089 );
not ( n326091 , n4222 );
not ( n326092 , n323534 );
or ( n326093 , n326091 , n326092 );
buf ( n326094 , n322346 );
buf ( n326095 , n553 );
buf ( n326096 , n580 );
xor ( n6249 , n326095 , n326096 );
buf ( n6250 , n6249 );
buf ( n326099 , n6250 );
nand ( n6252 , n326094 , n326099 );
buf ( n326101 , n6252 );
nand ( n6254 , n326093 , n326101 );
not ( n6255 , n6254 );
or ( n6256 , n6242 , n6255 );
buf ( n326105 , n4222 );
not ( n6258 , n326105 );
buf ( n326107 , n323534 );
not ( n326108 , n326107 );
or ( n6261 , n6258 , n326108 );
buf ( n326110 , n326101 );
nand ( n6263 , n6261 , n326110 );
buf ( n326112 , n6263 );
or ( n6265 , n326089 , n326112 );
buf ( n326114 , n324205 );
not ( n6267 , n326114 );
buf ( n326116 , n325685 );
not ( n6269 , n326116 );
or ( n6270 , n6267 , n6269 );
buf ( n326119 , n3738 );
buf ( n326120 , n555 );
buf ( n326121 , n578 );
xor ( n6274 , n326120 , n326121 );
buf ( n326123 , n6274 );
buf ( n326124 , n326123 );
nand ( n326125 , n326119 , n326124 );
buf ( n326126 , n326125 );
buf ( n326127 , n326126 );
nand ( n6280 , n6270 , n326127 );
buf ( n326129 , n6280 );
nand ( n6282 , n6265 , n326129 );
nand ( n326131 , n6256 , n6282 );
buf ( n326132 , n326131 );
buf ( n326133 , n559 );
buf ( n326134 , n576 );
nand ( n6287 , n326133 , n326134 );
buf ( n326136 , n6287 );
buf ( n326137 , n326136 );
not ( n6290 , n326137 );
buf ( n326139 , n324237 );
not ( n6292 , n326139 );
buf ( n326141 , n320732 );
not ( n6294 , n326141 );
or ( n6295 , n6292 , n6294 );
buf ( n6296 , n590 );
buf ( n326145 , n591 );
nand ( n326146 , n6296 , n326145 );
buf ( n326147 , n326146 );
buf ( n326148 , n326147 );
nand ( n326149 , n6295 , n326148 );
buf ( n326150 , n326149 );
buf ( n326151 , n326150 );
not ( n6304 , n326151 );
buf ( n326153 , n6304 );
buf ( n326154 , n326153 );
not ( n6307 , n326154 );
or ( n6308 , n6290 , n6307 );
buf ( n326157 , n324110 );
not ( n6310 , n326157 );
buf ( n326159 , n898 );
not ( n6312 , n326159 );
or ( n6313 , n6310 , n6312 );
buf ( n326162 , n320642 );
buf ( n326163 , n326046 );
nand ( n326164 , n326162 , n326163 );
buf ( n326165 , n326164 );
buf ( n326166 , n326165 );
nand ( n326167 , n6313 , n326166 );
buf ( n326168 , n326167 );
buf ( n326169 , n326168 );
nand ( n326170 , n6308 , n326169 );
buf ( n326171 , n326170 );
buf ( n326172 , n326171 );
buf ( n326173 , n326136 );
not ( n326174 , n326173 );
buf ( n6327 , n326150 );
nand ( n6328 , n326174 , n6327 );
buf ( n6329 , n6328 );
buf ( n326178 , n6329 );
nand ( n6331 , n326172 , n326178 );
buf ( n6332 , n6331 );
buf ( n6333 , n6332 );
xor ( n6334 , n326132 , n6333 );
buf ( n326183 , n324091 );
not ( n326184 , n326183 );
buf ( n326185 , n2327 );
not ( n326186 , n326185 );
or ( n326187 , n326184 , n326186 );
buf ( n326188 , n2331 );
buf ( n326189 , n326036 );
nand ( n6342 , n326188 , n326189 );
buf ( n326191 , n6342 );
buf ( n326192 , n326191 );
nand ( n6345 , n326187 , n326192 );
buf ( n326194 , n6345 );
not ( n6347 , n326194 );
buf ( n326196 , n324155 );
not ( n6349 , n326196 );
buf ( n326198 , n321203 );
not ( n326199 , n326198 );
or ( n6352 , n6349 , n326199 );
buf ( n326201 , n1469 );
buf ( n326202 , n325930 );
nand ( n326203 , n326201 , n326202 );
buf ( n326204 , n326203 );
buf ( n326205 , n326204 );
nand ( n326206 , n6352 , n326205 );
buf ( n326207 , n326206 );
not ( n6360 , n326207 );
or ( n326209 , n6347 , n6360 );
buf ( n326210 , n326194 );
buf ( n326211 , n326207 );
nor ( n326212 , n326210 , n326211 );
buf ( n326213 , n326212 );
buf ( n326214 , n324138 );
not ( n326215 , n326214 );
buf ( n326216 , n324130 );
not ( n326217 , n326216 );
or ( n6370 , n326215 , n326217 );
buf ( n6371 , n323828 );
buf ( n326220 , n326000 );
nand ( n326221 , n6371 , n326220 );
buf ( n326222 , n326221 );
buf ( n326223 , n326222 );
nand ( n6376 , n6370 , n326223 );
buf ( n326225 , n6376 );
buf ( n326226 , n326225 );
not ( n326227 , n326226 );
buf ( n326228 , n326227 );
or ( n6381 , n326213 , n326228 );
nand ( n326230 , n326209 , n6381 );
buf ( n326231 , n326230 );
and ( n6384 , n6334 , n326231 );
and ( n326233 , n326132 , n6333 );
or ( n6386 , n6384 , n326233 );
buf ( n326235 , n6386 );
buf ( n326236 , n326235 );
and ( n6389 , n6236 , n326236 );
and ( n326238 , n326080 , n326083 );
or ( n6391 , n6389 , n326238 );
buf ( n326240 , n6391 );
buf ( n326241 , n326240 );
and ( n326242 , n326077 , n326241 );
and ( n326243 , n326073 , n326076 );
or ( n6396 , n326242 , n326243 );
buf ( n326245 , n6396 );
buf ( n6398 , n326245 );
and ( n6399 , n6141 , n6398 );
and ( n326248 , n325984 , n325988 );
or ( n6401 , n6399 , n326248 );
buf ( n326250 , n6401 );
buf ( n326251 , n326250 );
xor ( n6404 , n325921 , n326251 );
buf ( n326253 , n6404 );
xor ( n6406 , n5166 , n326253 );
xor ( n6407 , n325065 , n325069 );
xor ( n6408 , n6407 , n325091 );
buf ( n326257 , n6408 );
buf ( n326258 , n326257 );
buf ( n326259 , n325287 );
not ( n6412 , n326259 );
buf ( n326261 , n3157 );
not ( n326262 , n326261 );
or ( n326263 , n6412 , n326262 );
buf ( n326264 , n323009 );
buf ( n326265 , n4791 );
nand ( n6418 , n326264 , n326265 );
buf ( n326267 , n6418 );
buf ( n326268 , n326267 );
nand ( n6421 , n326263 , n326268 );
buf ( n326270 , n6421 );
buf ( n326271 , n326270 );
buf ( n326272 , n325273 );
not ( n6425 , n326272 );
buf ( n326274 , n321592 );
not ( n6427 , n326274 );
or ( n326276 , n6425 , n6427 );
buf ( n326277 , n3186 );
buf ( n326278 , n324675 );
nand ( n6431 , n326277 , n326278 );
buf ( n326280 , n6431 );
buf ( n326281 , n326280 );
nand ( n6434 , n326276 , n326281 );
buf ( n326283 , n6434 );
buf ( n326284 , n326283 );
xor ( n6437 , n326271 , n326284 );
buf ( n326286 , n325049 );
and ( n6439 , n6437 , n326286 );
and ( n6440 , n326271 , n326284 );
or ( n6441 , n6439 , n6440 );
buf ( n326290 , n6441 );
buf ( n326291 , n326290 );
not ( n6444 , n326291 );
and ( n6445 , n325194 , n325139 );
not ( n6446 , n325194 );
and ( n6447 , n6446 , n325134 );
nor ( n6448 , n6445 , n6447 );
not ( n6449 , n324653 );
not ( n326298 , n5251 );
or ( n6451 , n6449 , n326298 );
nand ( n326300 , n6451 , n5257 );
and ( n326301 , n6448 , n326300 );
not ( n6454 , n6448 );
not ( n326303 , n326300 );
and ( n6456 , n6454 , n326303 );
nor ( n326305 , n326301 , n6456 );
buf ( n326306 , n326305 );
not ( n6459 , n326306 );
or ( n6460 , n6444 , n6459 );
xor ( n6461 , n325111 , n325115 );
xor ( n6462 , n6461 , n325130 );
buf ( n326311 , n6462 );
not ( n6464 , n326311 );
buf ( n326313 , n325188 );
not ( n6466 , n326313 );
buf ( n326315 , n6466 );
xor ( n6468 , n5308 , n326315 );
not ( n6469 , n325169 );
xor ( n6470 , n6468 , n6469 );
not ( n6471 , n6470 );
or ( n6472 , n6464 , n6471 );
not ( n326321 , n326311 );
not ( n6474 , n326321 );
not ( n326323 , n6470 );
not ( n326324 , n326323 );
or ( n326325 , n6474 , n326324 );
not ( n6478 , n322885 );
not ( n6479 , n322864 );
or ( n326328 , n6478 , n6479 );
or ( n6481 , n322885 , n322864 );
nand ( n6482 , n6481 , n322832 );
nand ( n326331 , n326328 , n6482 );
not ( n326332 , n326331 );
not ( n326333 , n323215 );
nand ( n6486 , n326333 , n3385 );
nand ( n326335 , n326332 , n6486 );
not ( n326336 , n326335 );
xor ( n6489 , n322951 , n322962 );
and ( n326338 , n6489 , n322979 );
and ( n326339 , n322951 , n322962 );
or ( n6492 , n326338 , n326339 );
buf ( n326341 , n6492 );
not ( n326342 , n326341 );
or ( n326343 , n326336 , n326342 );
or ( n6496 , n326332 , n6486 );
nand ( n326345 , n326343 , n6496 );
nand ( n6498 , n326325 , n326345 );
nand ( n6499 , n6472 , n6498 );
buf ( n6500 , n326290 );
not ( n326349 , n6500 );
buf ( n326350 , n326349 );
not ( n6503 , n326305 );
nand ( n326352 , n326350 , n6503 );
nand ( n326353 , n6499 , n326352 );
buf ( n326354 , n326353 );
nand ( n326355 , n6460 , n326354 );
buf ( n326356 , n326355 );
buf ( n326357 , n326356 );
xor ( n326358 , n326258 , n326357 );
xor ( n326359 , n325197 , n325201 );
xor ( n6512 , n326359 , n325344 );
buf ( n326361 , n6512 );
buf ( n326362 , n326361 );
and ( n6515 , n326358 , n326362 );
and ( n326364 , n326258 , n326357 );
or ( n326365 , n6515 , n326364 );
buf ( n326366 , n326365 );
buf ( n326367 , n326366 );
xor ( n6520 , n325984 , n325988 );
xor ( n6521 , n6520 , n6398 );
buf ( n326370 , n6521 );
buf ( n326371 , n326370 );
xor ( n6524 , n326367 , n326371 );
and ( n6525 , n325923 , n6117 );
not ( n6526 , n325923 );
and ( n6527 , n6526 , n6118 );
or ( n6528 , n6525 , n6527 );
and ( n6529 , n6528 , n6123 );
not ( n6530 , n6528 );
not ( n326379 , n6123 );
and ( n326380 , n6530 , n326379 );
nor ( n326381 , n6529 , n326380 );
buf ( n326382 , n326381 );
buf ( n326383 , n326123 );
not ( n326384 , n326383 );
buf ( n326385 , n3865 );
not ( n326386 , n326385 );
or ( n6539 , n326384 , n326386 );
buf ( n326388 , n323715 );
buf ( n326389 , n325681 );
nand ( n6542 , n326388 , n326389 );
buf ( n326391 , n6542 );
buf ( n326392 , n326391 );
nand ( n326393 , n6539 , n326392 );
buf ( n326394 , n326393 );
buf ( n326395 , n326394 );
buf ( n326396 , n6250 );
not ( n326397 , n326396 );
buf ( n326398 , n322468 );
not ( n326399 , n326398 );
or ( n6552 , n326397 , n326399 );
buf ( n326401 , n322474 );
buf ( n326402 , n325666 );
nand ( n6555 , n326401 , n326402 );
buf ( n326404 , n6555 );
buf ( n326405 , n326404 );
nand ( n6558 , n6552 , n326405 );
buf ( n326407 , n6558 );
buf ( n326408 , n326407 );
xor ( n6561 , n326395 , n326408 );
buf ( n326410 , n325942 );
not ( n326411 , n326410 );
buf ( n326412 , n326411 );
buf ( n326413 , n326412 );
and ( n326414 , n6561 , n326413 );
and ( n6567 , n326395 , n326408 );
or ( n326416 , n326414 , n6567 );
buf ( n326417 , n326416 );
buf ( n326418 , n326417 );
xor ( n6571 , n326018 , n326064 );
xor ( n6572 , n6571 , n326068 );
buf ( n326421 , n6572 );
buf ( n326422 , n326421 );
xor ( n326423 , n326418 , n326422 );
xor ( n6576 , n325994 , n325995 );
xor ( n6577 , n6576 , n326013 );
buf ( n326426 , n6577 );
buf ( n326427 , n326426 );
not ( n326428 , n326031 );
not ( n326429 , n326428 );
not ( n6582 , n326055 );
not ( n326431 , n6193 );
or ( n326432 , n6582 , n326431 );
or ( n6585 , n6193 , n326055 );
nand ( n6586 , n326432 , n6585 );
not ( n6587 , n6586 );
or ( n6588 , n326429 , n6587 );
or ( n6589 , n6586 , n326428 );
nand ( n6590 , n6588 , n6589 );
buf ( n326439 , n6590 );
xor ( n6592 , n326427 , n326439 );
and ( n6593 , n324228 , n324245 );
buf ( n326442 , n6593 );
buf ( n326443 , n326442 );
xor ( n326444 , n324116 , n324144 );
and ( n326445 , n326444 , n324161 );
and ( n6598 , n324116 , n324144 );
or ( n326447 , n326445 , n6598 );
buf ( n326448 , n326447 );
xor ( n326449 , n326443 , n326448 );
xor ( n6602 , n4224 , n4237 );
and ( n326451 , n6602 , n324097 );
and ( n6604 , n4224 , n4237 );
or ( n6605 , n326451 , n6604 );
buf ( n326454 , n6605 );
and ( n326455 , n326449 , n326454 );
and ( n326456 , n326443 , n326448 );
or ( n6609 , n326455 , n326456 );
buf ( n326458 , n6609 );
buf ( n326459 , n326458 );
and ( n6612 , n6592 , n326459 );
and ( n326461 , n326427 , n326439 );
or ( n326462 , n6612 , n326461 );
buf ( n326463 , n326462 );
buf ( n326464 , n326463 );
and ( n6617 , n326423 , n326464 );
and ( n326466 , n326418 , n326422 );
or ( n6619 , n6617 , n326466 );
buf ( n326468 , n6619 );
buf ( n326469 , n326468 );
xor ( n6622 , n326382 , n326469 );
xor ( n326471 , n326073 , n326076 );
xor ( n326472 , n326471 , n326241 );
buf ( n326473 , n326472 );
buf ( n326474 , n326473 );
and ( n326475 , n6622 , n326474 );
and ( n326476 , n326382 , n326469 );
or ( n6629 , n326475 , n326476 );
buf ( n326478 , n6629 );
buf ( n326479 , n326478 );
and ( n6632 , n6524 , n326479 );
and ( n326481 , n326367 , n326371 );
or ( n326482 , n6632 , n326481 );
buf ( n326483 , n326482 );
xor ( n6636 , n6406 , n326483 );
not ( n326485 , n6636 );
xor ( n6638 , n5506 , n325095 );
xor ( n326487 , n6638 , n325348 );
buf ( n6640 , n326487 );
not ( n6641 , n6503 );
not ( n6642 , n326290 );
or ( n326491 , n6641 , n6642 );
nand ( n326492 , n326350 , n326305 );
nand ( n6645 , n326491 , n326492 );
xor ( n6646 , n6645 , n6499 );
not ( n326495 , n6646 );
xor ( n6648 , n326271 , n326284 );
xor ( n326497 , n6648 , n326286 );
buf ( n326498 , n326497 );
buf ( n326499 , n326498 );
xor ( n6652 , n325239 , n325265 );
xor ( n326501 , n6652 , n325313 );
buf ( n326502 , n326501 );
buf ( n326503 , n326502 );
xor ( n6656 , n326499 , n326503 );
xor ( n6657 , n5433 , n325306 );
xor ( n326506 , n6657 , n325293 );
buf ( n326507 , n326506 );
not ( n326508 , n326507 );
buf ( n326509 , n326508 );
not ( n6662 , n326509 );
xor ( n6663 , n325207 , n325220 );
xor ( n6664 , n6663 , n325234 );
buf ( n326513 , n6664 );
not ( n326514 , n326513 );
or ( n6667 , n6662 , n326514 );
buf ( n326516 , n326513 );
not ( n6669 , n326516 );
buf ( n326518 , n6669 );
not ( n6671 , n326518 );
not ( n6672 , n326506 );
or ( n6673 , n6671 , n6672 );
buf ( n326522 , n325262 );
not ( n6675 , n326522 );
not ( n6676 , n5407 );
not ( n6677 , n5401 );
not ( n6678 , n6677 );
or ( n326527 , n6676 , n6678 );
or ( n6680 , n6677 , n5407 );
nand ( n326529 , n326527 , n6680 );
buf ( n326530 , n326529 );
not ( n326531 , n326530 );
or ( n6684 , n6675 , n326531 );
buf ( n326533 , n326529 );
buf ( n326534 , n325262 );
or ( n326535 , n326533 , n326534 );
buf ( n326536 , n326535 );
buf ( n326537 , n326536 );
nand ( n6690 , n6684 , n326537 );
buf ( n6691 , n6690 );
nand ( n326540 , n6673 , n6691 );
nand ( n6693 , n6667 , n326540 );
buf ( n326542 , n6693 );
and ( n326543 , n6656 , n326542 );
and ( n326544 , n326499 , n326503 );
or ( n326545 , n326543 , n326544 );
buf ( n326546 , n326545 );
buf ( n326547 , n326546 );
not ( n326548 , n326547 );
buf ( n326549 , n325321 );
buf ( n326550 , n325334 );
xor ( n326551 , n326549 , n326550 );
buf ( n326552 , n325317 );
xor ( n6705 , n326551 , n326552 );
buf ( n326554 , n6705 );
buf ( n6707 , n326554 );
nand ( n6708 , n326548 , n6707 );
buf ( n6709 , n6708 );
not ( n6710 , n6709 );
or ( n6711 , n326495 , n6710 );
buf ( n326560 , n326546 );
buf ( n326561 , n326554 );
not ( n326562 , n326561 );
buf ( n326563 , n326562 );
buf ( n326564 , n326563 );
nand ( n6717 , n326560 , n326564 );
buf ( n326566 , n6717 );
nand ( n6719 , n6711 , n326566 );
buf ( n326568 , n6719 );
xor ( n326569 , n326080 , n326083 );
xor ( n326570 , n326569 , n326236 );
buf ( n326571 , n326570 );
xor ( n326572 , n326395 , n326408 );
xor ( n6725 , n326572 , n326413 );
buf ( n326574 , n6725 );
buf ( n326575 , n326225 );
buf ( n326576 , n326194 );
xor ( n326577 , n326575 , n326576 );
buf ( n326578 , n326207 );
xnor ( n326579 , n326577 , n326578 );
buf ( n326580 , n326579 );
buf ( n326581 , n326580 );
not ( n6734 , n326581 );
buf ( n326583 , n6734 );
not ( n6736 , n326583 );
xor ( n326585 , n326136 , n326150 );
xor ( n6738 , n326585 , n326168 );
buf ( n326587 , n6738 );
not ( n6740 , n326587 );
buf ( n326589 , n6740 );
not ( n6742 , n326589 );
or ( n326591 , n6736 , n6742 );
buf ( n326592 , n6738 );
not ( n6745 , n326592 );
buf ( n326594 , n326580 );
not ( n326595 , n326594 );
or ( n6748 , n6745 , n326595 );
buf ( n6749 , n326089 );
not ( n6750 , n6749 );
buf ( n326599 , n326129 );
not ( n6752 , n326599 );
buf ( n326601 , n326112 );
not ( n6754 , n326601 );
buf ( n326603 , n6754 );
buf ( n326604 , n326603 );
not ( n6757 , n326604 );
and ( n6758 , n6752 , n6757 );
buf ( n326607 , n326129 );
buf ( n326608 , n326603 );
and ( n6761 , n326607 , n326608 );
nor ( n326610 , n6758 , n6761 );
buf ( n326611 , n326610 );
not ( n326612 , n326611 );
or ( n6765 , n6750 , n326612 );
or ( n326614 , n326611 , n6749 );
nand ( n326615 , n6765 , n326614 );
buf ( n326616 , n326615 );
nand ( n326617 , n6748 , n326616 );
buf ( n326618 , n326617 );
nand ( n6771 , n326591 , n326618 );
xor ( n326620 , n326574 , n6771 );
xor ( n326621 , n326132 , n6333 );
xor ( n6774 , n326621 , n326231 );
buf ( n326623 , n6774 );
and ( n6776 , n326620 , n326623 );
and ( n6777 , n326574 , n6771 );
or ( n326626 , n6776 , n6777 );
xor ( n326627 , n326571 , n326626 );
xor ( n326628 , n326418 , n326422 );
xor ( n6781 , n326628 , n326464 );
buf ( n326630 , n6781 );
and ( n326631 , n326627 , n326630 );
and ( n6784 , n326571 , n326626 );
or ( n326633 , n326631 , n6784 );
buf ( n326634 , n326633 );
xor ( n6787 , n326568 , n326634 );
xor ( n326636 , n326382 , n326469 );
xor ( n326637 , n326636 , n326474 );
buf ( n326638 , n326637 );
buf ( n326639 , n326638 );
and ( n6792 , n6787 , n326639 );
and ( n6793 , n326568 , n326634 );
or ( n6794 , n6792 , n6793 );
buf ( n326643 , n6794 );
buf ( n326644 , n326643 );
xor ( n326645 , n6640 , n326644 );
xor ( n326646 , n326367 , n326371 );
xor ( n6799 , n326646 , n326479 );
buf ( n326648 , n6799 );
buf ( n326649 , n326648 );
and ( n6802 , n326645 , n326649 );
and ( n6803 , n6640 , n326644 );
or ( n6804 , n6802 , n6803 );
buf ( n326653 , n6804 );
buf ( n326654 , n326653 );
not ( n6807 , n326654 );
buf ( n326656 , n6807 );
nand ( n6809 , n326485 , n326656 );
buf ( n6810 , n324962 );
not ( n6811 , n6810 );
buf ( n6812 , n321072 );
not ( n6813 , n6812 );
or ( n6814 , n6811 , n6813 );
buf ( n6815 , n1339 );
buf ( n326664 , n568 );
nand ( n326665 , n6815 , n326664 );
buf ( n326666 , n326665 );
buf ( n326667 , n326666 );
nand ( n326668 , n6814 , n326667 );
buf ( n326669 , n326668 );
not ( n326670 , n326669 );
not ( n326671 , n326670 );
buf ( n326672 , n324892 );
not ( n326673 , n326672 );
buf ( n326674 , n3157 );
not ( n326675 , n326674 );
or ( n6828 , n326673 , n326675 );
buf ( n326677 , n323009 );
buf ( n326678 , n549 );
buf ( n326679 , n562 );
xor ( n6832 , n326678 , n326679 );
buf ( n326681 , n6832 );
buf ( n326682 , n326681 );
nand ( n326683 , n326677 , n326682 );
buf ( n326684 , n326683 );
buf ( n326685 , n326684 );
nand ( n6838 , n6828 , n326685 );
buf ( n326687 , n6838 );
buf ( n326688 , n324922 );
not ( n6841 , n326688 );
buf ( n326690 , n324728 );
not ( n6843 , n326690 );
or ( n6844 , n6841 , n6843 );
buf ( n326693 , n324855 );
buf ( n326694 , n551 );
buf ( n326695 , n560 );
xor ( n6848 , n326694 , n326695 );
buf ( n6849 , n6848 );
buf ( n326698 , n6849 );
nand ( n6851 , n326693 , n326698 );
buf ( n326700 , n6851 );
buf ( n326701 , n326700 );
nand ( n6854 , n6844 , n326701 );
buf ( n326703 , n6854 );
xor ( n6856 , n326687 , n326703 );
not ( n6857 , n6856 );
or ( n6858 , n326671 , n6857 );
or ( n6859 , n6856 , n326670 );
nand ( n6860 , n6858 , n6859 );
not ( n6861 , n324898 );
not ( n6862 , n324914 );
or ( n6863 , n6861 , n6862 );
not ( n326712 , n324898 );
not ( n6865 , n326712 );
not ( n326714 , n5069 );
or ( n6867 , n6865 , n326714 );
not ( n326716 , n324924 );
nand ( n6869 , n6867 , n326716 );
nand ( n326718 , n6863 , n6869 );
or ( n326719 , n6860 , n326718 );
not ( n6872 , n5088 );
not ( n6873 , n6872 );
not ( n6874 , n5123 );
or ( n6875 , n6873 , n6874 );
not ( n326724 , n5105 );
nand ( n326725 , n6875 , n326724 );
nand ( n6878 , n324970 , n5088 );
nand ( n326727 , n326725 , n6878 );
nand ( n326728 , n326719 , n326727 );
nand ( n6881 , n6860 , n326718 );
nand ( n326730 , n326728 , n6881 );
buf ( n6883 , n326730 );
buf ( n6884 , n553 );
buf ( n6885 , n560 );
nand ( n6886 , n6884 , n6885 );
buf ( n6887 , n6886 );
buf ( n6888 , n6887 );
not ( n6889 , n6888 );
buf ( n6890 , n6889 );
buf ( n326739 , n6890 );
not ( n6892 , n326739 );
buf ( n326741 , n324907 );
not ( n326742 , n326741 );
buf ( n326743 , n1975 );
not ( n326744 , n326743 );
or ( n326745 , n326742 , n326744 );
buf ( n326746 , n321771 );
buf ( n326747 , n545 );
buf ( n326748 , n566 );
xor ( n6901 , n326747 , n326748 );
buf ( n326750 , n6901 );
buf ( n326751 , n326750 );
nand ( n6904 , n326746 , n326751 );
buf ( n326753 , n6904 );
buf ( n326754 , n326753 );
nand ( n6907 , n326745 , n326754 );
buf ( n326756 , n6907 );
buf ( n326757 , n326756 );
not ( n6910 , n326757 );
buf ( n326759 , n6910 );
buf ( n326760 , n326759 );
not ( n6913 , n326760 );
or ( n6914 , n6892 , n6913 );
buf ( n326763 , n6887 );
not ( n6916 , n326763 );
buf ( n326765 , n326756 );
not ( n6918 , n326765 );
or ( n6919 , n6916 , n6918 );
buf ( n326768 , n324944 );
not ( n6921 , n326768 );
buf ( n326770 , n321592 );
not ( n6923 , n326770 );
or ( n6924 , n6921 , n6923 );
buf ( n326773 , n3186 );
buf ( n326774 , n547 );
buf ( n326775 , n564 );
xor ( n6928 , n326774 , n326775 );
buf ( n326777 , n6928 );
buf ( n326778 , n326777 );
nand ( n6931 , n326773 , n326778 );
buf ( n326780 , n6931 );
buf ( n326781 , n326780 );
nand ( n6934 , n6924 , n326781 );
buf ( n326783 , n6934 );
buf ( n326784 , n326783 );
nand ( n6937 , n6919 , n326784 );
buf ( n326786 , n6937 );
buf ( n326787 , n326786 );
nand ( n6940 , n6914 , n326787 );
buf ( n326789 , n6940 );
buf ( n326790 , n326789 );
buf ( n326791 , n326681 );
not ( n6944 , n326791 );
buf ( n326793 , n3157 );
not ( n6946 , n326793 );
or ( n6947 , n6944 , n6946 );
buf ( n326796 , n323009 );
buf ( n326797 , n548 );
buf ( n326798 , n562 );
xor ( n6951 , n326797 , n326798 );
buf ( n326800 , n6951 );
buf ( n326801 , n326800 );
nand ( n6954 , n326796 , n326801 );
buf ( n326803 , n6954 );
buf ( n326804 , n326803 );
nand ( n6957 , n6947 , n326804 );
buf ( n326806 , n6957 );
buf ( n326807 , n326806 );
buf ( n326808 , n1339 );
buf ( n326809 , n321072 );
or ( n6962 , n326808 , n326809 );
buf ( n326811 , n568 );
nand ( n6964 , n6962 , n326811 );
buf ( n326813 , n6964 );
buf ( n326814 , n326813 );
xor ( n6967 , n326807 , n326814 );
buf ( n326816 , n326750 );
not ( n6969 , n326816 );
buf ( n326818 , n1975 );
not ( n6971 , n326818 );
or ( n6972 , n6969 , n6971 );
buf ( n326821 , n321771 );
buf ( n326822 , n544 );
buf ( n326823 , n566 );
xor ( n6976 , n326822 , n326823 );
buf ( n326825 , n6976 );
buf ( n326826 , n326825 );
nand ( n6979 , n326821 , n326826 );
buf ( n326828 , n6979 );
buf ( n326829 , n326828 );
nand ( n6982 , n6972 , n326829 );
buf ( n326831 , n6982 );
buf ( n326832 , n326831 );
xor ( n6985 , n6967 , n326832 );
buf ( n326834 , n6985 );
buf ( n326835 , n326834 );
xor ( n6988 , n326790 , n326835 );
buf ( n326837 , n326756 );
buf ( n326838 , n326687 );
not ( n6991 , n326838 );
buf ( n326840 , n326669 );
not ( n6993 , n326840 );
or ( n6994 , n6991 , n6993 );
buf ( n326843 , n326669 );
buf ( n326844 , n326687 );
or ( n6997 , n326843 , n326844 );
buf ( n326846 , n326703 );
nand ( n6999 , n6997 , n326846 );
buf ( n326848 , n6999 );
buf ( n326849 , n326848 );
nand ( n7002 , n6994 , n326849 );
buf ( n326851 , n7002 );
buf ( n326852 , n326851 );
xor ( n7005 , n326837 , n326852 );
buf ( n326854 , n552 );
buf ( n326855 , n560 );
and ( n7008 , n326854 , n326855 );
buf ( n326857 , n7008 );
buf ( n326858 , n326857 );
buf ( n326859 , n326777 );
not ( n7012 , n326859 );
buf ( n326861 , n321592 );
not ( n7014 , n326861 );
or ( n7015 , n7012 , n7014 );
buf ( n326864 , n1857 );
buf ( n326865 , n546 );
buf ( n326866 , n564 );
xor ( n7019 , n326865 , n326866 );
buf ( n326868 , n7019 );
buf ( n326869 , n326868 );
nand ( n7022 , n326864 , n326869 );
buf ( n326871 , n7022 );
buf ( n326872 , n326871 );
nand ( n7025 , n7015 , n326872 );
buf ( n326874 , n7025 );
buf ( n326875 , n326874 );
xor ( n7028 , n326858 , n326875 );
buf ( n326877 , n6849 );
not ( n7030 , n326877 );
and ( n7031 , n324727 , n324917 );
buf ( n326880 , n7031 );
not ( n7033 , n326880 );
or ( n7034 , n7030 , n7033 );
buf ( n326883 , n324855 );
buf ( n326884 , n550 );
buf ( n326885 , n560 );
xor ( n7038 , n326884 , n326885 );
buf ( n326887 , n7038 );
buf ( n326888 , n326887 );
nand ( n7041 , n326883 , n326888 );
buf ( n326890 , n7041 );
buf ( n326891 , n326890 );
nand ( n7044 , n7034 , n326891 );
buf ( n326893 , n7044 );
buf ( n326894 , n326893 );
xor ( n7047 , n7028 , n326894 );
buf ( n326896 , n7047 );
buf ( n326897 , n326896 );
xor ( n7050 , n7005 , n326897 );
buf ( n326899 , n7050 );
buf ( n326900 , n326899 );
xor ( n7053 , n6988 , n326900 );
buf ( n326902 , n7053 );
buf ( n326903 , n326902 );
xor ( n7056 , n6883 , n326903 );
xor ( n7057 , n5134 , n5135 );
and ( n7058 , n7057 , n324987 );
and ( n7059 , n5134 , n5135 );
or ( n7060 , n7058 , n7059 );
buf ( n326909 , n7060 );
buf ( n326910 , n326909 );
not ( n7063 , n326910 );
buf ( n326912 , n7063 );
buf ( n326913 , n326912 );
xor ( n7066 , n6890 , n326783 );
buf ( n326915 , n7066 );
buf ( n326916 , n326756 );
and ( n7069 , n326915 , n326916 );
not ( n7070 , n326915 );
buf ( n326919 , n326759 );
and ( n7072 , n7070 , n326919 );
nor ( n7073 , n7069 , n7072 );
buf ( n326922 , n7073 );
buf ( n326923 , n326922 );
nand ( n7076 , n326913 , n326923 );
buf ( n326925 , n7076 );
buf ( n326926 , n326925 );
not ( n7079 , n326926 );
xor ( n7080 , n5036 , n5080 );
and ( n7081 , n7080 , n324972 );
and ( n7082 , n5036 , n5080 );
or ( n7083 , n7081 , n7082 );
buf ( n326932 , n7083 );
buf ( n326933 , n326932 );
not ( n7086 , n326933 );
or ( n7087 , n7079 , n7086 );
buf ( n326936 , n326909 );
buf ( n326937 , n326922 );
not ( n7090 , n326937 );
buf ( n326939 , n7090 );
buf ( n326940 , n326939 );
nand ( n7093 , n326936 , n326940 );
buf ( n326942 , n7093 );
buf ( n326943 , n326942 );
nand ( n7096 , n7087 , n326943 );
buf ( n326945 , n7096 );
buf ( n326946 , n326945 );
xor ( n7099 , n7056 , n326946 );
buf ( n326948 , n7099 );
not ( n7101 , n325005 );
not ( n7102 , n324974 );
or ( n7103 , n7101 , n7102 );
or ( n7104 , n325005 , n324974 );
nand ( n7105 , n7104 , n324875 );
nand ( n7106 , n7103 , n7105 );
xor ( n7107 , n325541 , n6025 );
and ( n7108 , n7107 , n325917 );
and ( n7109 , n325541 , n6025 );
or ( n7110 , n7108 , n7109 );
buf ( n326959 , n7110 );
xor ( n7112 , n7106 , n326959 );
xor ( n7113 , n325440 , n325461 );
and ( n7114 , n7113 , n325479 );
and ( n7115 , n325440 , n325461 );
or ( n7116 , n7114 , n7115 );
buf ( n326965 , n7116 );
buf ( n326966 , n326965 );
buf ( n326967 , n325433 );
not ( n7120 , n326967 );
buf ( n326969 , n325390 );
not ( n7122 , n326969 );
or ( n7123 , n7120 , n7122 );
buf ( n326972 , n325399 );
buf ( n326973 , n551 );
buf ( n326974 , n576 );
xor ( n7127 , n326973 , n326974 );
buf ( n326976 , n7127 );
buf ( n326977 , n326976 );
nand ( n7130 , n326972 , n326977 );
buf ( n326979 , n7130 );
buf ( n326980 , n326979 );
nand ( n7133 , n7123 , n326980 );
buf ( n326982 , n7133 );
not ( n7135 , n325528 );
not ( n7136 , n321203 );
or ( n7137 , n7135 , n7136 );
buf ( n326986 , n3752 );
buf ( n326987 , n584 );
nand ( n7140 , n326986 , n326987 );
buf ( n326989 , n7140 );
nand ( n7142 , n7137 , n326989 );
xor ( n7143 , n326982 , n7142 );
buf ( n326992 , n325454 );
not ( n7145 , n326992 );
buf ( n326994 , n3865 );
not ( n7147 , n326994 );
or ( n7148 , n7145 , n7147 );
buf ( n326997 , n323715 );
buf ( n326998 , n549 );
buf ( n326999 , n578 );
xor ( n7152 , n326998 , n326999 );
buf ( n327001 , n7152 );
buf ( n327002 , n327001 );
nand ( n7155 , n326997 , n327002 );
buf ( n327004 , n7155 );
buf ( n327005 , n327004 );
nand ( n7158 , n7148 , n327005 );
buf ( n327007 , n7158 );
and ( n7160 , n7143 , n327007 );
not ( n7161 , n7143 );
not ( n7162 , n327007 );
and ( n7163 , n7161 , n7162 );
nor ( n7164 , n7160 , n7163 );
buf ( n327013 , n7164 );
xor ( n7166 , n326966 , n327013 );
xor ( n7167 , n325490 , n325513 );
and ( n7168 , n7167 , n325535 );
and ( n7169 , n325490 , n325513 );
or ( n7170 , n7168 , n7169 );
buf ( n327019 , n7170 );
buf ( n327020 , n327019 );
xor ( n7173 , n7166 , n327020 );
buf ( n327022 , n7173 );
buf ( n327023 , n327022 );
xor ( n7176 , n325891 , n325907 );
and ( n7177 , n7176 , n325914 );
and ( n7178 , n325891 , n325907 );
or ( n7179 , n7177 , n7178 );
buf ( n327028 , n7179 );
buf ( n327029 , n327028 );
xor ( n7182 , n327023 , n327029 );
buf ( n327031 , n553 );
buf ( n327032 , n576 );
and ( n7185 , n327031 , n327032 );
buf ( n327034 , n7185 );
buf ( n327035 , n327034 );
buf ( n327036 , n325506 );
not ( n7189 , n327036 );
buf ( n327038 , n5650 );
not ( n7191 , n327038 );
or ( n7192 , n7189 , n7191 );
buf ( n327041 , n322474 );
buf ( n327042 , n547 );
buf ( n327043 , n580 );
xor ( n7196 , n327042 , n327043 );
buf ( n327045 , n7196 );
buf ( n327046 , n327045 );
nand ( n7199 , n327041 , n327046 );
buf ( n327048 , n7199 );
buf ( n327049 , n327048 );
nand ( n7202 , n7192 , n327049 );
buf ( n327051 , n7202 );
buf ( n327052 , n327051 );
xor ( n7205 , n327035 , n327052 );
buf ( n327054 , n325472 );
not ( n7207 , n327054 );
buf ( n327056 , n323550 );
not ( n7209 , n327056 );
or ( n7210 , n7207 , n7209 );
buf ( n327059 , n323562 );
buf ( n327060 , n545 );
buf ( n327061 , n582 );
xor ( n7214 , n327060 , n327061 );
buf ( n327063 , n7214 );
buf ( n327064 , n327063 );
nand ( n7217 , n327059 , n327064 );
buf ( n327066 , n7217 );
buf ( n327067 , n327066 );
nand ( n7220 , n7210 , n327067 );
buf ( n327069 , n7220 );
buf ( n327070 , n327069 );
not ( n7223 , n327070 );
buf ( n327072 , n7223 );
buf ( n327073 , n327072 );
xor ( n7226 , n7205 , n327073 );
buf ( n327075 , n7226 );
buf ( n327076 , n327075 );
xor ( n7229 , n325896 , n325897 );
and ( n7230 , n7229 , n325904 );
and ( n7231 , n325896 , n325897 );
or ( n7232 , n7230 , n7231 );
buf ( n327081 , n7232 );
buf ( n327082 , n327081 );
xor ( n7235 , n327076 , n327082 );
xor ( n7236 , n325416 , n325482 );
and ( n7237 , n7236 , n325538 );
and ( n7238 , n325416 , n325482 );
or ( n7239 , n7237 , n7238 );
buf ( n327088 , n7239 );
buf ( n327089 , n327088 );
xor ( n7242 , n7235 , n327089 );
buf ( n327091 , n7242 );
buf ( n327092 , n327091 );
xor ( n7245 , n7182 , n327092 );
buf ( n327094 , n7245 );
and ( n7247 , n7112 , n327094 );
and ( n7248 , n7106 , n326959 );
or ( n7249 , n7247 , n7248 );
xor ( n7250 , n326948 , n7249 );
xor ( n7251 , n326966 , n327013 );
and ( n7252 , n7251 , n327020 );
and ( n7253 , n326966 , n327013 );
or ( n7254 , n7252 , n7253 );
buf ( n327103 , n7254 );
buf ( n327104 , n327103 );
xor ( n7257 , n327035 , n327052 );
and ( n7258 , n7257 , n327073 );
and ( n7259 , n327035 , n327052 );
or ( n7260 , n7258 , n7259 );
buf ( n327109 , n7260 );
buf ( n327110 , n327109 );
buf ( n327111 , n327063 );
not ( n7264 , n327111 );
buf ( n327113 , n323550 );
not ( n7266 , n327113 );
or ( n7267 , n7264 , n7266 );
buf ( n327116 , n323562 );
buf ( n327117 , n544 );
buf ( n327118 , n582 );
xor ( n7271 , n327117 , n327118 );
buf ( n327120 , n7271 );
buf ( n327121 , n327120 );
nand ( n7274 , n327116 , n327121 );
buf ( n327123 , n7274 );
buf ( n327124 , n327123 );
nand ( n7277 , n7267 , n327124 );
buf ( n327126 , n7277 );
buf ( n327127 , n327126 );
buf ( n327128 , n327001 );
not ( n7281 , n327128 );
buf ( n327130 , n3865 );
not ( n7283 , n327130 );
or ( n7284 , n7281 , n7283 );
buf ( n327133 , n323715 );
buf ( n327134 , n548 );
buf ( n327135 , n578 );
xor ( n7288 , n327134 , n327135 );
buf ( n327137 , n7288 );
buf ( n327138 , n327137 );
nand ( n7291 , n327133 , n327138 );
buf ( n327140 , n7291 );
buf ( n327141 , n327140 );
nand ( n7294 , n7284 , n327141 );
buf ( n327143 , n7294 );
buf ( n327144 , n327143 );
xor ( n7297 , n327127 , n327144 );
buf ( n327146 , n322176 );
buf ( n327147 , n321209 );
or ( n7300 , n327146 , n327147 );
buf ( n327149 , n584 );
nand ( n7302 , n7300 , n327149 );
buf ( n327151 , n7302 );
buf ( n327152 , n327151 );
xor ( n7305 , n7297 , n327152 );
buf ( n327154 , n7305 );
buf ( n327155 , n327154 );
xor ( n7308 , n327110 , n327155 );
buf ( n327157 , n327069 );
not ( n7310 , n7142 );
not ( n7311 , n326982 );
or ( n7312 , n7310 , n7311 );
or ( n7313 , n326982 , n7142 );
nand ( n7314 , n7313 , n327007 );
nand ( n7315 , n7312 , n7314 );
buf ( n327164 , n7315 );
xor ( n7317 , n327157 , n327164 );
buf ( n327166 , n552 );
buf ( n327167 , n576 );
and ( n7320 , n327166 , n327167 );
buf ( n327169 , n7320 );
buf ( n327170 , n327169 );
buf ( n327171 , n326976 );
not ( n7324 , n327171 );
buf ( n327173 , n324130 );
not ( n7326 , n327173 );
or ( n7327 , n7324 , n7326 );
buf ( n327176 , n5580 );
buf ( n327177 , n550 );
buf ( n327178 , n576 );
xor ( n7331 , n327177 , n327178 );
buf ( n327180 , n7331 );
buf ( n327181 , n327180 );
nand ( n7334 , n327176 , n327181 );
buf ( n327183 , n7334 );
buf ( n327184 , n327183 );
nand ( n7337 , n7327 , n327184 );
buf ( n327186 , n7337 );
buf ( n327187 , n327186 );
xor ( n7340 , n327170 , n327187 );
buf ( n327189 , n327045 );
not ( n7342 , n327189 );
buf ( n327191 , n322468 );
not ( n7344 , n327191 );
or ( n7345 , n7342 , n7344 );
buf ( n327194 , n322474 );
buf ( n327195 , n546 );
buf ( n327196 , n580 );
xor ( n7349 , n327195 , n327196 );
buf ( n327198 , n7349 );
buf ( n327199 , n327198 );
nand ( n7352 , n327194 , n327199 );
buf ( n327201 , n7352 );
buf ( n327202 , n327201 );
nand ( n7355 , n7345 , n327202 );
buf ( n327204 , n7355 );
buf ( n327205 , n327204 );
xor ( n7358 , n7340 , n327205 );
buf ( n327207 , n7358 );
buf ( n327208 , n327207 );
xor ( n7361 , n7317 , n327208 );
buf ( n327210 , n7361 );
buf ( n327211 , n327210 );
xor ( n7364 , n7308 , n327211 );
buf ( n327213 , n7364 );
buf ( n327214 , n327213 );
xor ( n7367 , n327104 , n327214 );
xor ( n7368 , n327076 , n327082 );
and ( n7369 , n7368 , n327089 );
and ( n7370 , n327076 , n327082 );
or ( n7371 , n7369 , n7370 );
buf ( n327220 , n7371 );
buf ( n327221 , n327220 );
xor ( n7374 , n7367 , n327221 );
buf ( n327223 , n7374 );
buf ( n327224 , n327223 );
xor ( n7377 , n327023 , n327029 );
and ( n7378 , n7377 , n327092 );
and ( n7379 , n327023 , n327029 );
or ( n7380 , n7378 , n7379 );
buf ( n327229 , n7380 );
buf ( n327230 , n327229 );
xor ( n7383 , n327224 , n327230 );
not ( n7384 , n6860 );
not ( n7385 , n7384 );
not ( n7386 , n326718 );
not ( n7387 , n326727 );
not ( n7388 , n7387 );
or ( n7389 , n7386 , n7388 );
or ( n7390 , n7387 , n326718 );
nand ( n7391 , n7389 , n7390 );
not ( n7392 , n7391 );
or ( n7393 , n7385 , n7392 );
or ( n7394 , n7384 , n7391 );
nand ( n7395 , n7393 , n7394 );
buf ( n327244 , n7395 );
xor ( n7397 , n324990 , n324996 );
and ( n7398 , n7397 , n325003 );
and ( n7399 , n324990 , n324996 );
or ( n7400 , n7398 , n7399 );
buf ( n327249 , n7400 );
buf ( n327250 , n327249 );
xor ( n7403 , n327244 , n327250 );
buf ( n327252 , n326912 );
buf ( n327253 , n326922 );
and ( n7406 , n327252 , n327253 );
not ( n7407 , n327252 );
buf ( n327256 , n326939 );
and ( n7409 , n7407 , n327256 );
or ( n7410 , n7406 , n7409 );
buf ( n327259 , n7410 );
xnor ( n327260 , n327259 , n326932 );
buf ( n327261 , n327260 );
and ( n327262 , n7403 , n327261 );
and ( n7415 , n327244 , n327250 );
or ( n327264 , n327262 , n7415 );
buf ( n327265 , n327264 );
buf ( n327266 , n327265 );
xor ( n7419 , n7383 , n327266 );
buf ( n327268 , n7419 );
xor ( n7421 , n7250 , n327268 );
xor ( n7422 , n327244 , n327250 );
xor ( n7423 , n7422 , n327261 );
buf ( n327272 , n7423 );
xor ( n7425 , n5509 , n325920 );
and ( n7426 , n7425 , n326251 );
and ( n7427 , n5509 , n325920 );
or ( n7428 , n7426 , n7427 );
buf ( n327277 , n7428 );
xor ( n7430 , n327272 , n327277 );
xor ( n7431 , n7106 , n326959 );
xor ( n7432 , n7431 , n327094 );
and ( n7433 , n7430 , n7432 );
and ( n7434 , n327272 , n327277 );
or ( n7435 , n7433 , n7434 );
nor ( n7436 , n7421 , n7435 );
xor ( n7437 , n326258 , n326357 );
xor ( n7438 , n7437 , n326362 );
buf ( n327287 , n7438 );
buf ( n327288 , n327287 );
xor ( n7441 , n326311 , n326323 );
xnor ( n7442 , n7441 , n326345 );
not ( n7443 , n7442 );
not ( n7444 , n7443 );
not ( n7445 , n3086 );
not ( n7446 , n322981 );
or ( n7447 , n7445 , n7446 );
buf ( n327296 , n3086 );
buf ( n327297 , n322981 );
nor ( n7450 , n327296 , n327297 );
buf ( n327299 , n7450 );
or ( n7452 , n327299 , n3043 );
nand ( n7453 , n7447 , n7452 );
not ( n7454 , n7453 );
not ( n7455 , n6486 );
and ( n7456 , n326331 , n7455 );
not ( n7457 , n326331 );
and ( n7458 , n7457 , n6486 );
nor ( n7459 , n7456 , n7458 );
and ( n7460 , n7459 , n326341 );
not ( n7461 , n7459 );
not ( n7462 , n326341 );
and ( n7463 , n7461 , n7462 );
nor ( n7464 , n7460 , n7463 );
not ( n7465 , n7464 );
xor ( n7466 , n3357 , n323229 );
and ( n7467 , n7466 , n3427 );
and ( n7468 , n3357 , n323229 );
or ( n7469 , n7467 , n7468 );
not ( n7470 , n7469 );
nand ( n7471 , n7465 , n7470 );
not ( n7472 , n7471 );
or ( n7473 , n7454 , n7472 );
nand ( n7474 , n7469 , n7464 );
nand ( n7475 , n7473 , n7474 );
not ( n7476 , n7475 );
not ( n7477 , n7476 );
or ( n7478 , n7444 , n7477 );
xor ( n7479 , n326499 , n326503 );
xor ( n7480 , n7479 , n326542 );
buf ( n327329 , n7480 );
nand ( n7482 , n7478 , n327329 );
buf ( n327331 , n7482 );
buf ( n327332 , n7475 );
buf ( n327333 , n7442 );
nand ( n7486 , n327332 , n327333 );
buf ( n327335 , n7486 );
buf ( n327336 , n327335 );
nand ( n7489 , n327331 , n327336 );
buf ( n327338 , n7489 );
buf ( n327339 , n327338 );
xor ( n7492 , n326427 , n326439 );
xor ( n7493 , n7492 , n326459 );
buf ( n327342 , n7493 );
buf ( n327343 , n327342 );
xor ( n7496 , n326443 , n326448 );
xor ( n7497 , n7496 , n326454 );
buf ( n327346 , n7497 );
not ( n7499 , n327346 );
xor ( n7500 , n324212 , n324248 );
and ( n7501 , n7500 , n324255 );
and ( n7502 , n324212 , n324248 );
or ( n7503 , n7501 , n7502 );
buf ( n327352 , n7503 );
not ( n7505 , n327352 );
or ( n7506 , n7499 , n7505 );
not ( n7507 , n327352 );
not ( n7508 , n7507 );
not ( n7509 , n327346 );
not ( n7510 , n7509 );
or ( n7511 , n7508 , n7510 );
or ( n7512 , n4319 , n4255 );
nand ( n7513 , n7512 , n4329 );
nand ( n7514 , n4319 , n4255 );
nand ( n7515 , n7513 , n7514 );
nand ( n7516 , n7511 , n7515 );
nand ( n7517 , n7506 , n7516 );
buf ( n327366 , n7517 );
xor ( n7519 , n327343 , n327366 );
xor ( n7520 , n326574 , n6771 );
xor ( n7521 , n7520 , n326623 );
buf ( n327370 , n7521 );
and ( n7523 , n7519 , n327370 );
and ( n7524 , n327343 , n327366 );
or ( n7525 , n7523 , n7524 );
buf ( n327374 , n7525 );
buf ( n327375 , n327374 );
xor ( n7528 , n327339 , n327375 );
xor ( n7529 , n326571 , n326626 );
xor ( n7530 , n7529 , n326630 );
buf ( n327379 , n7530 );
and ( n7532 , n7528 , n327379 );
and ( n7533 , n327339 , n327375 );
or ( n7534 , n7532 , n7533 );
buf ( n327383 , n7534 );
buf ( n327384 , n327383 );
xor ( n7537 , n327288 , n327384 );
xor ( n7538 , n326568 , n326634 );
xor ( n7539 , n7538 , n326639 );
buf ( n327388 , n7539 );
buf ( n327389 , n327388 );
and ( n7542 , n7537 , n327389 );
and ( n7543 , n327288 , n327384 );
or ( n7544 , n7542 , n7543 );
buf ( n327393 , n7544 );
buf ( n327394 , n327393 );
xor ( n7547 , n6640 , n326644 );
xor ( n7548 , n7547 , n326649 );
buf ( n327397 , n7548 );
buf ( n327398 , n327397 );
nor ( n7551 , n327394 , n327398 );
buf ( n327400 , n7551 );
nor ( n7553 , n7436 , n327400 );
xor ( n7554 , n327272 , n327277 );
xor ( n7555 , n7554 , n7432 );
not ( n7556 , n7555 );
xor ( n327405 , n5166 , n326253 );
and ( n7558 , n327405 , n326483 );
and ( n327407 , n5166 , n326253 );
or ( n327408 , n7558 , n327407 );
buf ( n327409 , n327408 );
not ( n327410 , n327409 );
buf ( n327411 , n327410 );
nand ( n7564 , n7556 , n327411 );
and ( n7565 , n6809 , n7553 , n7564 );
xor ( n327414 , n323191 , n323272 );
and ( n327415 , n327414 , n323390 );
and ( n7568 , n323191 , n323272 );
or ( n327417 , n327415 , n7568 );
buf ( n327418 , n327417 );
buf ( n327419 , n327418 );
buf ( n327420 , n326513 );
buf ( n327421 , n6691 );
xor ( n7574 , n327420 , n327421 );
buf ( n327423 , n326509 );
xnor ( n327424 , n7574 , n327423 );
buf ( n327425 , n327424 );
buf ( n327426 , n327425 );
not ( n7579 , n327426 );
buf ( n327428 , n7579 );
buf ( n327429 , n327428 );
and ( n7582 , n327419 , n327429 );
not ( n7583 , n327419 );
buf ( n327432 , n327425 );
and ( n7585 , n7583 , n327432 );
nor ( n7586 , n7582 , n7585 );
buf ( n327435 , n7586 );
buf ( n327436 , n327435 );
and ( n7589 , n7469 , n7464 );
not ( n7590 , n7469 );
and ( n7591 , n7590 , n7465 );
nor ( n7592 , n7589 , n7591 );
and ( n7593 , n7592 , n7453 );
not ( n327442 , n7592 );
not ( n7595 , n7453 );
and ( n7596 , n327442 , n7595 );
nor ( n327445 , n7593 , n7596 );
buf ( n327446 , n327445 );
buf ( n327447 , n327446 );
buf ( n327448 , n327447 );
buf ( n7601 , n327448 );
xor ( n7602 , n327436 , n7601 );
buf ( n7603 , n7602 );
buf ( n327452 , n7603 );
xor ( n7605 , n324051 , n4214 );
and ( n327454 , n7605 , n324271 );
and ( n327455 , n324051 , n4214 );
or ( n327456 , n327454 , n327455 );
buf ( n327457 , n327456 );
buf ( n7610 , n327457 );
xor ( n7611 , n327452 , n7610 );
xor ( n7612 , n324182 , n324188 );
and ( n327461 , n7612 , n324268 );
and ( n7614 , n324182 , n324188 );
or ( n7615 , n327461 , n7614 );
buf ( n327464 , n7615 );
buf ( n327465 , n327464 );
buf ( n327466 , n322984 );
not ( n327467 , n327466 );
buf ( n327468 , n327467 );
buf ( n327469 , n327468 );
not ( n327470 , n327469 );
buf ( n327471 , n323183 );
not ( n7624 , n327471 );
or ( n327473 , n327470 , n7624 );
buf ( n327474 , n323183 );
buf ( n327475 , n327468 );
or ( n7628 , n327474 , n327475 );
buf ( n327477 , n323392 );
nand ( n7630 , n7628 , n327477 );
buf ( n327479 , n7630 );
buf ( n327480 , n327479 );
nand ( n327481 , n327473 , n327480 );
buf ( n327482 , n327481 );
buf ( n327483 , n327482 );
xor ( n7636 , n327465 , n327483 );
buf ( n327485 , n326583 );
not ( n7638 , n327485 );
xor ( n7639 , n326615 , n6738 );
buf ( n327488 , n7639 );
not ( n7641 , n327488 );
or ( n7642 , n7638 , n7641 );
buf ( n327491 , n7639 );
buf ( n327492 , n326583 );
or ( n7645 , n327491 , n327492 );
nand ( n7646 , n7642 , n7645 );
buf ( n327495 , n7646 );
buf ( n327496 , n327495 );
xor ( n7649 , n324195 , n324258 );
and ( n7650 , n7649 , n324265 );
and ( n7651 , n324195 , n324258 );
or ( n7652 , n7650 , n7651 );
buf ( n327501 , n7652 );
buf ( n327502 , n327501 );
xor ( n327503 , n327496 , n327502 );
xor ( n7656 , n7507 , n7515 );
xnor ( n7657 , n7656 , n327346 );
buf ( n327506 , n7657 );
xor ( n7659 , n327503 , n327506 );
buf ( n327508 , n7659 );
buf ( n327509 , n327508 );
xor ( n327510 , n7636 , n327509 );
buf ( n327511 , n327510 );
buf ( n327512 , n327511 );
and ( n327513 , n7611 , n327512 );
and ( n7666 , n327452 , n7610 );
or ( n327515 , n327513 , n7666 );
buf ( n327516 , n327515 );
not ( n7669 , n327516 );
buf ( n327518 , n7475 );
xor ( n327519 , n7442 , n327518 );
xor ( n7672 , n327519 , n327329 );
xor ( n327521 , n327465 , n327483 );
and ( n327522 , n327521 , n327509 );
and ( n7675 , n327465 , n327483 );
or ( n327524 , n327522 , n7675 );
buf ( n327525 , n327524 );
xor ( n7678 , n7672 , n327525 );
not ( n7679 , n327418 );
nand ( n327528 , n7679 , n327425 );
not ( n327529 , n327528 );
not ( n7682 , n327445 );
or ( n327531 , n327529 , n7682 );
buf ( n327532 , n327418 );
buf ( n327533 , n327428 );
nand ( n327534 , n327532 , n327533 );
buf ( n327535 , n327534 );
nand ( n7688 , n327531 , n327535 );
buf ( n327537 , n7688 );
xor ( n7690 , n327496 , n327502 );
and ( n7691 , n7690 , n327506 );
and ( n7692 , n327496 , n327502 );
or ( n7693 , n7691 , n7692 );
buf ( n327542 , n7693 );
buf ( n327543 , n327542 );
xor ( n7696 , n327537 , n327543 );
xor ( n7697 , n327343 , n327366 );
xor ( n327546 , n7697 , n327370 );
buf ( n327547 , n327546 );
buf ( n327548 , n327547 );
xor ( n327549 , n7696 , n327548 );
buf ( n327550 , n327549 );
xor ( n7703 , n7678 , n327550 );
not ( n327552 , n7703 );
and ( n327553 , n7669 , n327552 );
xor ( n327554 , n327452 , n7610 );
xor ( n327555 , n327554 , n327512 );
buf ( n327556 , n327555 );
xor ( n327557 , n323396 , n324011 );
and ( n327558 , n327557 , n324274 );
and ( n7711 , n323396 , n324011 );
or ( n327560 , n327558 , n7711 );
buf ( n327561 , n327560 );
nor ( n327562 , n327556 , n327561 );
nor ( n7715 , n327553 , n327562 );
buf ( n327564 , n7715 );
buf ( n327565 , n6646 );
not ( n7718 , n327565 );
buf ( n327567 , n326546 );
buf ( n327568 , n326563 );
and ( n327569 , n327567 , n327568 );
not ( n7722 , n327567 );
buf ( n327571 , n326554 );
and ( n327572 , n7722 , n327571 );
or ( n7725 , n327569 , n327572 );
buf ( n7726 , n7725 );
buf ( n327575 , n7726 );
not ( n7728 , n327575 );
or ( n7729 , n7718 , n7728 );
buf ( n327578 , n7726 );
buf ( n327579 , n6646 );
or ( n327580 , n327578 , n327579 );
buf ( n327581 , n327580 );
buf ( n327582 , n327581 );
nand ( n7735 , n7729 , n327582 );
buf ( n327584 , n7735 );
buf ( n327585 , n327584 );
xor ( n327586 , n327537 , n327543 );
and ( n327587 , n327586 , n327548 );
and ( n7740 , n327537 , n327543 );
or ( n327589 , n327587 , n7740 );
buf ( n327590 , n327589 );
buf ( n327591 , n327590 );
xor ( n327592 , n327585 , n327591 );
xor ( n7745 , n327339 , n327375 );
xor ( n327594 , n7745 , n327379 );
buf ( n327595 , n327594 );
buf ( n327596 , n327595 );
xor ( n7749 , n327592 , n327596 );
buf ( n327598 , n7749 );
buf ( n327599 , n327598 );
xor ( n327600 , n7672 , n327525 );
and ( n7753 , n327600 , n327550 );
and ( n327602 , n7672 , n327525 );
or ( n327603 , n7753 , n327602 );
buf ( n327604 , n327603 );
nor ( n327605 , n327599 , n327604 );
buf ( n327606 , n327605 );
buf ( n327607 , n327606 );
not ( n7760 , n327607 );
buf ( n7761 , n7760 );
buf ( n327610 , n7761 );
xor ( n7763 , n327288 , n327384 );
xor ( n327612 , n7763 , n327389 );
buf ( n327613 , n327612 );
buf ( n327614 , n327613 );
xor ( n7767 , n327585 , n327591 );
and ( n327616 , n7767 , n327596 );
and ( n327617 , n327585 , n327591 );
or ( n7770 , n327616 , n327617 );
buf ( n327619 , n7770 );
buf ( n327620 , n327619 );
nor ( n7773 , n327614 , n327620 );
buf ( n7774 , n7773 );
buf ( n327623 , n7774 );
not ( n7776 , n327623 );
buf ( n327625 , n7776 );
buf ( n327626 , n327625 );
and ( n7779 , n327564 , n327610 , n327626 );
buf ( n327628 , n7779 );
nand ( n327629 , n7565 , n327628 );
not ( n7782 , n327629 );
buf ( n327631 , n7782 );
not ( n327632 , n327631 );
or ( n7785 , n4656 , n327632 );
buf ( n327634 , n7564 );
not ( n327635 , n327634 );
buf ( n327636 , n327635 );
nor ( n7789 , n7421 , n7435 );
nor ( n7790 , n327636 , n7789 );
not ( n327639 , n7790 );
buf ( n327640 , n327397 );
buf ( n327641 , n327393 );
nand ( n7794 , n327640 , n327641 );
buf ( n327643 , n7794 );
buf ( n327644 , n327643 );
not ( n7797 , n327644 );
buf ( n327646 , n7797 );
not ( n7799 , n327646 );
not ( n7800 , n6809 );
or ( n7801 , n7799 , n7800 );
buf ( n327650 , n326656 );
not ( n7803 , n327650 );
buf ( n327652 , n6636 );
nand ( n7805 , n7803 , n327652 );
buf ( n327654 , n7805 );
nand ( n327655 , n7801 , n327654 );
not ( n7808 , n327655 );
or ( n327657 , n327639 , n7808 );
not ( n7810 , n327411 );
nand ( n327659 , n7810 , n7555 );
not ( n7812 , n327659 );
not ( n327661 , n7789 );
and ( n7814 , n7812 , n327661 );
and ( n7815 , n7435 , n7421 );
nor ( n327664 , n7814 , n7815 );
nand ( n7817 , n327657 , n327664 );
not ( n327666 , n7817 );
nor ( n7819 , n7774 , n327606 );
not ( n327668 , n7819 );
nor ( n327669 , n327516 , n7703 );
nand ( n327670 , n327561 , n327556 );
or ( n327671 , n327669 , n327670 );
nand ( n7824 , n7703 , n327516 );
nand ( n327673 , n327671 , n7824 );
not ( n7826 , n327673 );
or ( n7827 , n327668 , n7826 );
nand ( n7828 , n327598 , n327603 );
nor ( n7829 , n7774 , n7828 );
buf ( n327678 , n327613 );
buf ( n327679 , n327619 );
and ( n7832 , n327678 , n327679 );
buf ( n327681 , n7832 );
nor ( n7834 , n7829 , n327681 );
nand ( n7835 , n7827 , n7834 );
nand ( n7836 , n7835 , n7565 );
nand ( n7837 , n327666 , n7836 );
buf ( n327686 , n7837 );
not ( n7839 , n327686 );
buf ( n327688 , n7839 );
buf ( n327689 , n327688 );
nand ( n327690 , n7785 , n327689 );
buf ( n327691 , n327690 );
buf ( n327692 , n327691 );
xor ( n7845 , n326837 , n326852 );
and ( n327694 , n7845 , n326897 );
and ( n7847 , n326837 , n326852 );
or ( n327696 , n327694 , n7847 );
buf ( n327697 , n327696 );
buf ( n327698 , n327697 );
xor ( n327699 , n326807 , n326814 );
and ( n327700 , n327699 , n326832 );
and ( n327701 , n326807 , n326814 );
or ( n7854 , n327700 , n327701 );
buf ( n327703 , n7854 );
buf ( n327704 , n327703 );
buf ( n327705 , n326887 );
not ( n327706 , n327705 );
buf ( n327707 , n7031 );
not ( n7860 , n327707 );
or ( n327709 , n327706 , n7860 );
buf ( n7862 , n324855 );
buf ( n327711 , n549 );
buf ( n327712 , n560 );
xor ( n327713 , n327711 , n327712 );
buf ( n327714 , n327713 );
buf ( n327715 , n327714 );
nand ( n7868 , n7862 , n327715 );
buf ( n327717 , n7868 );
buf ( n327718 , n327717 );
nand ( n7871 , n327709 , n327718 );
buf ( n7872 , n7871 );
buf ( n327721 , n551 );
buf ( n327722 , n560 );
nand ( n7875 , n327721 , n327722 );
buf ( n327724 , n7875 );
xor ( n327725 , n7872 , n327724 );
buf ( n327726 , n326825 );
not ( n7879 , n327726 );
buf ( n327728 , n1975 );
not ( n327729 , n327728 );
or ( n7882 , n7879 , n327729 );
buf ( n327731 , n321771 );
buf ( n327732 , n566 );
nand ( n7885 , n327731 , n327732 );
buf ( n7886 , n7885 );
buf ( n327735 , n7886 );
nand ( n7888 , n7882 , n327735 );
buf ( n327737 , n7888 );
xnor ( n327738 , n327725 , n327737 );
buf ( n327739 , n327738 );
xor ( n7892 , n327704 , n327739 );
buf ( n327741 , n326800 );
not ( n327742 , n327741 );
buf ( n327743 , n3157 );
not ( n7896 , n327743 );
or ( n327745 , n327742 , n7896 );
buf ( n327746 , n323009 );
buf ( n327747 , n547 );
buf ( n327748 , n562 );
xor ( n7901 , n327747 , n327748 );
buf ( n327750 , n7901 );
buf ( n327751 , n327750 );
nand ( n327752 , n327746 , n327751 );
buf ( n327753 , n327752 );
buf ( n327754 , n327753 );
nand ( n327755 , n327745 , n327754 );
buf ( n327756 , n327755 );
buf ( n327757 , n327756 );
buf ( n327758 , n326868 );
not ( n7911 , n327758 );
buf ( n327760 , n321592 );
not ( n7913 , n327760 );
or ( n7914 , n7911 , n7913 );
buf ( n327763 , n1857 );
buf ( n327764 , n545 );
buf ( n327765 , n564 );
xor ( n7918 , n327764 , n327765 );
buf ( n327767 , n7918 );
buf ( n327768 , n327767 );
nand ( n7921 , n327763 , n327768 );
buf ( n327770 , n7921 );
buf ( n327771 , n327770 );
nand ( n7924 , n7914 , n327771 );
buf ( n327773 , n7924 );
buf ( n327774 , n327773 );
not ( n327775 , n327774 );
buf ( n327776 , n327775 );
buf ( n327777 , n327776 );
xor ( n327778 , n327757 , n327777 );
xor ( n7931 , n326858 , n326875 );
and ( n327780 , n7931 , n326894 );
and ( n327781 , n326858 , n326875 );
or ( n7934 , n327780 , n327781 );
buf ( n327783 , n7934 );
buf ( n327784 , n327783 );
xor ( n7937 , n327778 , n327784 );
buf ( n327786 , n7937 );
buf ( n327787 , n327786 );
xor ( n327788 , n7892 , n327787 );
buf ( n327789 , n327788 );
buf ( n327790 , n327789 );
xor ( n327791 , n327698 , n327790 );
xor ( n7944 , n326790 , n326835 );
and ( n327793 , n7944 , n326900 );
and ( n327794 , n326790 , n326835 );
or ( n7947 , n327793 , n327794 );
buf ( n327796 , n7947 );
buf ( n327797 , n327796 );
xor ( n327798 , n327791 , n327797 );
buf ( n327799 , n327798 );
buf ( n7952 , n327799 );
xor ( n327801 , n327157 , n327164 );
and ( n7954 , n327801 , n327208 );
and ( n327803 , n327157 , n327164 );
or ( n7956 , n7954 , n327803 );
buf ( n327805 , n7956 );
buf ( n327806 , n327805 );
buf ( n327807 , n551 );
buf ( n327808 , n576 );
and ( n7961 , n327807 , n327808 );
buf ( n327810 , n7961 );
buf ( n327811 , n327810 );
buf ( n327812 , n327180 );
not ( n7965 , n327812 );
buf ( n327814 , n325952 );
not ( n7967 , n327814 );
or ( n327816 , n7965 , n7967 );
buf ( n327817 , n5580 );
buf ( n327818 , n549 );
buf ( n327819 , n576 );
xor ( n7972 , n327818 , n327819 );
buf ( n327821 , n7972 );
buf ( n327822 , n327821 );
nand ( n7975 , n327817 , n327822 );
buf ( n327824 , n7975 );
buf ( n327825 , n327824 );
nand ( n327826 , n327816 , n327825 );
buf ( n327827 , n327826 );
buf ( n327828 , n327827 );
xor ( n327829 , n327811 , n327828 );
buf ( n327830 , n327120 );
not ( n7983 , n327830 );
buf ( n327832 , n322554 );
not ( n327833 , n327832 );
or ( n7986 , n7983 , n327833 );
buf ( n327835 , n323755 );
buf ( n327836 , n582 );
nand ( n327837 , n327835 , n327836 );
buf ( n327838 , n327837 );
buf ( n327839 , n327838 );
nand ( n327840 , n7986 , n327839 );
buf ( n327841 , n327840 );
buf ( n327842 , n327841 );
xor ( n327843 , n327829 , n327842 );
buf ( n327844 , n327843 );
buf ( n327845 , n327844 );
xor ( n327846 , n327127 , n327144 );
and ( n327847 , n327846 , n327152 );
and ( n327848 , n327127 , n327144 );
or ( n327849 , n327847 , n327848 );
buf ( n327850 , n327849 );
buf ( n327851 , n327850 );
xor ( n8004 , n327845 , n327851 );
buf ( n327853 , n327137 );
not ( n327854 , n327853 );
buf ( n327855 , n3865 );
not ( n327856 , n327855 );
or ( n8009 , n327854 , n327856 );
buf ( n327858 , n323715 );
buf ( n327859 , n547 );
buf ( n327860 , n578 );
xor ( n8013 , n327859 , n327860 );
buf ( n8014 , n8013 );
buf ( n327863 , n8014 );
nand ( n8016 , n327858 , n327863 );
buf ( n327865 , n8016 );
buf ( n327866 , n327865 );
nand ( n327867 , n8009 , n327866 );
buf ( n327868 , n327867 );
buf ( n327869 , n327868 );
buf ( n327870 , n327198 );
not ( n327871 , n327870 );
buf ( n327872 , n5650 );
not ( n327873 , n327872 );
or ( n327874 , n327871 , n327873 );
buf ( n327875 , n322474 );
buf ( n327876 , n545 );
buf ( n327877 , n580 );
xor ( n327878 , n327876 , n327877 );
buf ( n327879 , n327878 );
buf ( n327880 , n327879 );
nand ( n327881 , n327875 , n327880 );
buf ( n327882 , n327881 );
buf ( n327883 , n327882 );
nand ( n327884 , n327874 , n327883 );
buf ( n327885 , n327884 );
buf ( n327886 , n327885 );
not ( n8039 , n327886 );
buf ( n8040 , n8039 );
buf ( n8041 , n8040 );
xor ( n8042 , n327869 , n8041 );
xor ( n327891 , n327170 , n327187 );
and ( n8044 , n327891 , n327205 );
and ( n327893 , n327170 , n327187 );
or ( n8046 , n8044 , n327893 );
buf ( n327895 , n8046 );
buf ( n327896 , n327895 );
xor ( n8049 , n8042 , n327896 );
buf ( n327898 , n8049 );
buf ( n327899 , n327898 );
xor ( n8052 , n8004 , n327899 );
buf ( n327901 , n8052 );
buf ( n327902 , n327901 );
xor ( n327903 , n327806 , n327902 );
xor ( n8056 , n327110 , n327155 );
and ( n327905 , n8056 , n327211 );
and ( n8058 , n327110 , n327155 );
or ( n327907 , n327905 , n8058 );
buf ( n327908 , n327907 );
buf ( n327909 , n327908 );
xor ( n327910 , n327903 , n327909 );
buf ( n327911 , n327910 );
xor ( n8064 , n327104 , n327214 );
and ( n327913 , n8064 , n327221 );
and ( n327914 , n327104 , n327214 );
or ( n8067 , n327913 , n327914 );
buf ( n327916 , n8067 );
xor ( n8069 , n327911 , n327916 );
xor ( n327918 , n6883 , n326903 );
and ( n8071 , n327918 , n326946 );
and ( n8072 , n6883 , n326903 );
or ( n327921 , n8071 , n8072 );
buf ( n327922 , n327921 );
xor ( n327923 , n8069 , n327922 );
buf ( n327924 , n327923 );
xor ( n327925 , n7952 , n327924 );
xor ( n327926 , n327224 , n327230 );
and ( n8079 , n327926 , n327266 );
and ( n327928 , n327224 , n327230 );
or ( n327929 , n8079 , n327928 );
buf ( n327930 , n327929 );
buf ( n327931 , n327930 );
xor ( n327932 , n327925 , n327931 );
buf ( n327933 , n327932 );
xor ( n327934 , n326948 , n7249 );
and ( n8087 , n327934 , n327268 );
and ( n327936 , n326948 , n7249 );
or ( n8089 , n8087 , n327936 );
or ( n8090 , n327933 , n8089 );
buf ( n327939 , n8090 );
nand ( n8092 , n327933 , n8089 );
buf ( n8093 , n8092 );
nand ( n8094 , n327939 , n8093 );
buf ( n327943 , n8094 );
buf ( n327944 , n327943 );
xnor ( n327945 , n327692 , n327944 );
buf ( n327946 , n327945 );
not ( n8099 , n327946 );
not ( n327948 , n544 );
or ( n327949 , n570 , n586 );
or ( n8102 , n571 , n587 );
nand ( n327951 , n327949 , n8102 );
not ( n8104 , n327951 );
not ( n327953 , n8104 );
nor ( n327954 , n573 , n589 );
nor ( n8107 , n572 , n588 );
nor ( n327956 , n327954 , n8107 );
not ( n327957 , n327956 );
nand ( n8110 , n575 , n591 );
nor ( n8111 , n574 , n590 );
or ( n8112 , n8110 , n8111 );
nand ( n8113 , n574 , n590 );
nand ( n327962 , n8112 , n8113 );
not ( n327963 , n327962 );
or ( n8116 , n327957 , n327963 );
nor ( n8117 , n572 , n588 );
not ( n8118 , n8117 );
nand ( n8119 , n573 , n589 );
not ( n8120 , n8119 );
and ( n8121 , n8118 , n8120 );
and ( n8122 , n572 , n588 );
nor ( n8123 , n8121 , n8122 );
nand ( n8124 , n8116 , n8123 );
not ( n8125 , n8124 );
or ( n327974 , n327953 , n8125 );
nand ( n8127 , n571 , n587 );
nor ( n327976 , n570 , n586 );
or ( n8129 , n8127 , n327976 );
nand ( n8130 , n570 , n586 );
nand ( n8131 , n8129 , n8130 );
not ( n8132 , n8131 );
nand ( n8133 , n327974 , n8132 );
nand ( n8134 , n569 , n585 );
not ( n8135 , n8134 );
nor ( n327984 , n569 , n585 );
nor ( n8137 , n8135 , n327984 );
and ( n327986 , n8133 , n8137 );
not ( n8139 , n8133 );
not ( n327988 , n327984 );
nand ( n8141 , n327988 , n8134 );
and ( n327990 , n8139 , n8141 );
nor ( n8143 , n327986 , n327990 );
not ( n8144 , n8143 );
not ( n327993 , n8144 );
or ( n327994 , n327948 , n327993 );
not ( n327995 , n8133 );
not ( n8148 , n8141 );
nand ( n327997 , n327995 , n8148 );
not ( n327998 , n8137 );
nand ( n8151 , n327998 , n8133 );
nand ( n328000 , n327997 , n8151 );
not ( n328001 , n544 );
nand ( n8154 , n328000 , n328001 );
nand ( n328003 , n327994 , n8154 );
not ( n8156 , n328003 );
not ( n8157 , n8156 );
xor ( n8158 , n545 , n546 );
not ( n8159 , n8158 );
xor ( n8160 , n544 , n545 );
nand ( n8161 , n8159 , n8160 );
not ( n8162 , n8161 );
and ( n8163 , n8157 , n8162 );
not ( n8164 , n544 );
nor ( n8165 , n569 , n585 );
nor ( n8166 , n327951 , n8165 );
not ( n8167 , n8166 );
not ( n8168 , n8124 );
or ( n8169 , n8167 , n8168 );
and ( n8170 , n8131 , n327988 );
not ( n328019 , n8134 );
nor ( n8172 , n8170 , n328019 );
nand ( n8173 , n8169 , n8172 );
xor ( n8174 , n568 , n584 );
and ( n8175 , n8173 , n8174 );
not ( n8176 , n8173 );
not ( n8177 , n8174 );
and ( n328026 , n8176 , n8177 );
nor ( n328027 , n8175 , n328026 );
buf ( n8180 , n328027 );
not ( n328029 , n8180 );
not ( n8182 , n328029 );
or ( n8183 , n8164 , n8182 );
not ( n328032 , n328027 );
not ( n328033 , n328032 );
nand ( n8186 , n328033 , n328001 );
nand ( n328035 , n8183 , n8186 );
and ( n8188 , n328035 , n8158 );
nor ( n328037 , n8163 , n8188 );
not ( n328038 , n328037 );
nor ( n328039 , n571 , n587 );
not ( n8192 , n328039 );
not ( n328041 , n8192 );
not ( n328042 , n8124 );
or ( n8195 , n328041 , n328042 );
buf ( n328044 , n8127 );
nand ( n8197 , n8195 , n328044 );
not ( n8198 , n8130 );
nor ( n328047 , n8198 , n327976 );
and ( n328048 , n8197 , n328047 );
not ( n328049 , n8197 );
xnor ( n8202 , n570 , n586 );
and ( n328051 , n328049 , n8202 );
nor ( n328052 , n328048 , n328051 );
buf ( n8205 , n328052 );
buf ( n328054 , n8205 );
nand ( n8207 , n328054 , n544 );
xor ( n8208 , n328038 , n8207 );
and ( n8209 , n553 , n554 );
not ( n8210 , n553 );
not ( n8211 , n554 );
and ( n328060 , n8210 , n8211 );
nor ( n328061 , n8209 , n328060 );
not ( n328062 , n328061 );
xor ( n8215 , n552 , n553 );
nand ( n328064 , n328062 , n8215 );
not ( n328065 , n328064 );
not ( n8218 , n328065 );
nor ( n328067 , n563 , n579 );
nor ( n8220 , n562 , n578 );
nor ( n8221 , n328067 , n8220 );
not ( n328070 , n8221 );
or ( n8223 , n564 , n580 );
not ( n328072 , n581 );
nand ( n328073 , n328072 , n3089 );
or ( n8226 , n567 , n583 );
not ( n328075 , n582 );
nand ( n328076 , n328075 , n1842 );
nand ( n8229 , n8223 , n328073 , n8226 , n328076 );
nor ( n8230 , n328070 , n8229 );
not ( n8231 , n8230 );
nor ( n8232 , n568 , n584 );
nor ( n8233 , n569 , n585 );
nor ( n8234 , n8232 , n8233 );
not ( n8235 , n587 );
not ( n8236 , n571 );
nand ( n8237 , n8235 , n8236 );
not ( n8238 , n588 );
not ( n8239 , n572 );
nand ( n328088 , n8238 , n8239 );
not ( n8241 , n570 );
nand ( n8242 , n5703 , n8241 );
nand ( n8243 , n8234 , n8237 , n328088 , n8242 );
not ( n8244 , n8243 );
not ( n8245 , n8244 );
nand ( n8246 , n574 , n590 );
nand ( n8247 , n575 , n591 );
nand ( n8248 , n8246 , n8247 );
not ( n8249 , n8248 );
nor ( n328098 , n574 , n590 );
nor ( n328099 , n573 , n589 );
nor ( n328100 , n328098 , n328099 );
not ( n8253 , n328100 );
or ( n328102 , n8249 , n8253 );
not ( n8255 , n589 );
not ( n328104 , n573 );
or ( n328105 , n8255 , n328104 );
nand ( n328106 , n588 , n572 );
nand ( n328107 , n328105 , n328106 );
not ( n8260 , n328107 );
nand ( n328109 , n328102 , n8260 );
not ( n328110 , n328109 );
or ( n328111 , n8245 , n328110 );
or ( n8264 , n570 , n586 );
nand ( n328113 , n8264 , n571 , n587 );
not ( n328114 , n328113 );
nand ( n328115 , n568 , n584 );
nand ( n8268 , n570 , n586 );
nand ( n328117 , n569 , n585 );
nand ( n8270 , n328115 , n8268 , n328117 );
not ( n8271 , n8270 );
not ( n328120 , n8271 );
or ( n328121 , n328114 , n328120 );
not ( n8274 , n584 );
not ( n328123 , n568 );
nand ( n328124 , n8274 , n328123 );
not ( n328125 , n328124 );
not ( n8278 , n8165 );
not ( n328127 , n8278 );
or ( n328128 , n328125 , n328127 );
nand ( n8281 , n328128 , n328115 );
nand ( n328130 , n328121 , n8281 );
nand ( n328131 , n328111 , n328130 );
not ( n8284 , n328131 );
or ( n328133 , n8231 , n8284 );
nor ( n328134 , n565 , n581 );
nor ( n328135 , n564 , n580 );
nor ( n8288 , n328134 , n328135 );
not ( n328137 , n8288 );
nand ( n8290 , n567 , n583 );
nor ( n8291 , n566 , n582 );
or ( n328140 , n8290 , n8291 );
nand ( n8293 , n566 , n582 );
nand ( n328142 , n328140 , n8293 );
not ( n328143 , n328142 );
or ( n8296 , n328137 , n328143 );
and ( n328145 , n565 , n581 );
not ( n8298 , n564 );
nand ( n328147 , n8298 , n5821 );
and ( n328148 , n328145 , n328147 );
and ( n8301 , n564 , n580 );
nor ( n328150 , n328148 , n8301 );
nand ( n328151 , n8296 , n328150 );
and ( n8304 , n328151 , n8221 );
nand ( n8305 , n563 , n579 );
nor ( n8306 , n562 , n578 );
or ( n8307 , n8305 , n8306 );
nand ( n8308 , n562 , n578 );
nand ( n328157 , n8307 , n8308 );
nor ( n328158 , n8304 , n328157 );
nand ( n8311 , n328133 , n328158 );
nor ( n328160 , n561 , n577 );
not ( n328161 , n328160 );
nand ( n8314 , n561 , n577 );
and ( n8315 , n328161 , n8314 );
and ( n8316 , n8311 , n8315 );
not ( n8317 , n8311 );
not ( n8318 , n8315 );
and ( n328167 , n8317 , n8318 );
nor ( n328168 , n8316 , n328167 );
not ( n8321 , n328168 );
and ( n328170 , n8321 , n552 );
not ( n328171 , n8321 );
not ( n8324 , n552 );
and ( n328173 , n328171 , n8324 );
or ( n328174 , n328170 , n328173 );
not ( n8327 , n328174 );
or ( n328176 , n8218 , n8327 );
not ( n328177 , n552 );
not ( n8330 , n562 );
not ( n328179 , n578 );
and ( n328180 , n8330 , n328179 );
nor ( n8333 , n328180 , n328067 );
not ( n8334 , n8333 );
nor ( n8335 , n8334 , n328160 );
not ( n8336 , n8335 );
nor ( n328185 , n8336 , n8229 );
not ( n328186 , n328185 );
not ( n8339 , n328109 );
not ( n328188 , n8244 );
or ( n8341 , n8339 , n328188 );
nand ( n328190 , n8341 , n328130 );
not ( n8343 , n328190 );
or ( n328192 , n328186 , n8343 );
not ( n328193 , n8335 );
not ( n328194 , n8288 );
not ( n8347 , n328142 );
or ( n328196 , n328194 , n8347 );
nand ( n328197 , n328196 , n328150 );
not ( n8350 , n328197 );
or ( n328199 , n328193 , n8350 );
and ( n8352 , n328157 , n328161 );
not ( n8353 , n8314 );
nor ( n8354 , n8352 , n8353 );
nand ( n8355 , n328199 , n8354 );
not ( n8356 , n8355 );
nand ( n8357 , n328192 , n8356 );
nor ( n8358 , n560 , n576 );
not ( n8359 , n8358 );
nand ( n8360 , n560 , n576 );
nand ( n8361 , n8359 , n8360 );
not ( n8362 , n8361 );
and ( n8363 , n8357 , n8362 );
not ( n8364 , n8357 );
and ( n8365 , n8364 , n8361 );
nor ( n8366 , n8363 , n8365 );
not ( n8367 , n8366 );
not ( n8368 , n8367 );
or ( n8369 , n328177 , n8368 );
nand ( n8370 , n8366 , n8324 );
nand ( n8371 , n8369 , n8370 );
not ( n8372 , n328062 );
nand ( n8373 , n8371 , n8372 );
nand ( n8374 , n328176 , n8373 );
xor ( n8375 , n8208 , n8374 );
xor ( n8376 , n547 , n548 );
not ( n8377 , n8376 );
not ( n8378 , n546 );
not ( n8379 , n8378 );
or ( n8380 , n583 , n567 );
not ( n8381 , n8380 );
not ( n8382 , n328131 );
or ( n8383 , n8381 , n8382 );
buf ( n8384 , n8290 );
nand ( n8385 , n8383 , n8384 );
not ( n8386 , n8293 );
nor ( n8387 , n8386 , n8291 );
and ( n8388 , n8385 , n8387 );
not ( n8389 , n8385 );
not ( n8390 , n1842 );
not ( n8391 , n323949 );
or ( n8392 , n8390 , n8391 );
nand ( n8393 , n8392 , n8293 );
and ( n8394 , n8389 , n8393 );
nor ( n8395 , n8388 , n8394 );
not ( n8396 , n8395 );
buf ( n8397 , n8396 );
not ( n8398 , n8397 );
not ( n8399 , n8398 );
or ( n8400 , n8379 , n8399 );
not ( n8401 , n8395 );
nand ( n8402 , n546 , n8401 );
nand ( n8403 , n8400 , n8402 );
not ( n8404 , n8403 );
or ( n8405 , n8377 , n8404 );
not ( n8406 , n546 );
nand ( n8407 , n567 , n583 );
and ( n8408 , n8380 , n8407 );
xor ( n8409 , n8408 , n328190 );
buf ( n8410 , n8409 );
not ( n8411 , n8410 );
not ( n8412 , n8411 );
or ( n8413 , n8406 , n8412 );
nand ( n8414 , n8410 , n8378 );
nand ( n8415 , n8413 , n8414 );
xnor ( n8416 , n546 , n547 );
nor ( n8417 , n8376 , n8416 );
nand ( n8418 , n8415 , n8417 );
nand ( n8419 , n8405 , n8418 );
not ( n8420 , n8419 );
xor ( n8421 , n550 , n549 );
not ( n8422 , n8421 );
not ( n8423 , n8422 );
not ( n8424 , n8423 );
not ( n8425 , n548 );
and ( n8426 , n8226 , n328073 , n328076 );
not ( n8427 , n8426 );
not ( n8428 , n328190 );
or ( n8429 , n8427 , n8428 );
not ( n8430 , n328073 );
not ( n8431 , n328142 );
or ( n8432 , n8430 , n8431 );
nand ( n8433 , n565 , n581 );
nand ( n8434 , n8432 , n8433 );
not ( n8435 , n8434 );
nand ( n8436 , n8429 , n8435 );
nor ( n8437 , n8301 , n328135 );
and ( n8438 , n8436 , n8437 );
not ( n8439 , n8436 );
xnor ( n8440 , n564 , n580 );
and ( n8441 , n8439 , n8440 );
nor ( n8442 , n8438 , n8441 );
not ( n8443 , n8442 );
not ( n8444 , n8443 );
or ( n8445 , n8425 , n8444 );
buf ( n8446 , n8442 );
not ( n8447 , n548 );
nand ( n8448 , n8446 , n8447 );
nand ( n8449 , n8445 , n8448 );
not ( n8450 , n8449 );
or ( n8451 , n8424 , n8450 );
not ( n8452 , n548 );
and ( n8453 , n8226 , n328076 );
not ( n8454 , n8453 );
not ( n8455 , n328190 );
or ( n8456 , n8454 , n8455 );
not ( n8457 , n328142 );
nand ( n8458 , n8456 , n8457 );
or ( n8459 , n328145 , n328134 );
and ( n8460 , n8458 , n8459 );
not ( n8461 , n8458 );
and ( n8462 , n328073 , n8433 );
and ( n8463 , n8461 , n8462 );
nor ( n8464 , n8460 , n8463 );
not ( n8465 , n8464 );
not ( n8466 , n8465 );
not ( n8467 , n8466 );
or ( n8468 , n8452 , n8467 );
not ( n8469 , n548 );
nand ( n8470 , n8469 , n8465 );
nand ( n8471 , n8468 , n8470 );
xnor ( n8472 , n548 , n549 );
not ( n8473 , n8472 );
and ( n8474 , n8473 , n8422 );
buf ( n8475 , n8474 );
nand ( n8476 , n8471 , n8475 );
nand ( n8477 , n8451 , n8476 );
not ( n8478 , n8477 );
not ( n8479 , n8478 );
and ( n8480 , n8420 , n8479 );
not ( n8481 , n8420 );
and ( n8482 , n8481 , n8478 );
nor ( n8483 , n8480 , n8482 );
xor ( n8484 , n551 , n552 );
buf ( n8485 , n8484 );
not ( n8486 , n8485 );
not ( n8487 , n562 );
not ( n8488 , n578 );
and ( n8489 , n8487 , n8488 );
and ( n8490 , n562 , n578 );
nor ( n8491 , n8489 , n8490 );
not ( n8492 , n8491 );
nor ( n8493 , n563 , n579 );
nor ( n8494 , n8229 , n8493 );
not ( n8495 , n8494 );
not ( n8496 , n328131 );
or ( n8497 , n8495 , n8496 );
not ( n8498 , n328067 );
not ( n8499 , n8498 );
not ( n8500 , n328151 );
or ( n8501 , n8499 , n8500 );
nand ( n8502 , n563 , n579 );
nand ( n8503 , n8501 , n8502 );
not ( n8504 , n8503 );
nand ( n8505 , n8497 , n8504 );
not ( n8506 , n8505 );
not ( n8507 , n8506 );
or ( n8508 , n8492 , n8507 );
not ( n8509 , n8491 );
nand ( n8510 , n8509 , n8505 );
nand ( n8511 , n8508 , n8510 );
buf ( n8512 , n8511 );
not ( n8513 , n8512 );
not ( n8514 , n550 );
not ( n8515 , n8514 );
or ( n8516 , n8513 , n8515 );
not ( n8517 , n8512 );
nand ( n8518 , n8517 , n550 );
nand ( n8519 , n8516 , n8518 );
not ( n8520 , n8519 );
or ( n8521 , n8486 , n8520 );
not ( n8522 , n8229 );
not ( n8523 , n8522 );
not ( n8524 , n328131 );
or ( n8525 , n8523 , n8524 );
not ( n8526 , n328197 );
nand ( n8527 , n8525 , n8526 );
not ( n8528 , n8502 );
nor ( n8529 , n8528 , n8493 );
and ( n8530 , n8527 , n8529 );
not ( n8531 , n8527 );
not ( n8532 , n8502 );
nor ( n8533 , n8532 , n8493 );
not ( n8534 , n8533 );
and ( n8535 , n8531 , n8534 );
nor ( n8536 , n8530 , n8535 );
buf ( n8537 , n8536 );
and ( n8538 , n550 , n8537 );
not ( n8539 , n550 );
not ( n8540 , n8537 );
and ( n8541 , n8539 , n8540 );
nor ( n8542 , n8538 , n8541 );
or ( n8543 , n550 , n551 );
nand ( n8544 , n550 , n551 );
nand ( n8545 , n8543 , n8544 );
nor ( n8546 , n8545 , n8484 );
nand ( n8547 , n8542 , n8546 );
nand ( n8548 , n8521 , n8547 );
buf ( n8549 , n8548 );
and ( n8550 , n8483 , n8549 );
not ( n8551 , n8483 );
not ( n8552 , n8549 );
and ( n8553 , n8551 , n8552 );
nor ( n8554 , n8550 , n8553 );
xor ( n8555 , n8375 , n8554 );
not ( n8556 , n328065 );
not ( n8557 , n552 );
not ( n8558 , n8517 );
or ( n8559 , n8557 , n8558 );
nand ( n328408 , n8512 , n8324 );
nand ( n8561 , n8559 , n328408 );
not ( n8562 , n8561 );
or ( n8563 , n8556 , n8562 );
not ( n8564 , n328062 );
nand ( n8565 , n328174 , n8564 );
nand ( n8566 , n8563 , n8565 );
xnor ( n328415 , n554 , n555 );
xor ( n328416 , n555 , n556 );
or ( n328417 , n328415 , n328416 );
not ( n8570 , n328417 );
not ( n328419 , n8570 );
not ( n328420 , n554 );
not ( n328421 , n8367 );
or ( n8574 , n328420 , n328421 );
not ( n328423 , n8367 );
nand ( n328424 , n328423 , n8211 );
nand ( n8577 , n8574 , n328424 );
not ( n328426 , n8577 );
or ( n328427 , n328419 , n328426 );
not ( n8580 , n8211 );
not ( n328429 , n561 );
not ( n328430 , n577 );
and ( n8583 , n328429 , n328430 );
nor ( n328432 , n8583 , n8358 );
nand ( n328433 , n328432 , n8221 );
nor ( n8586 , n8229 , n328433 );
not ( n328435 , n8586 );
not ( n328436 , n328190 );
or ( n328437 , n328435 , n328436 );
not ( n8590 , n328433 );
not ( n328439 , n8590 );
not ( n8592 , n328151 );
or ( n328441 , n328439 , n8592 );
and ( n8594 , n328157 , n328432 );
or ( n328443 , n8358 , n8314 );
nand ( n328444 , n328443 , n8360 );
nor ( n8597 , n8594 , n328444 );
nand ( n8598 , n328441 , n8597 );
not ( n328447 , n8598 );
nand ( n8600 , n328437 , n328447 );
buf ( n328449 , n8600 );
not ( n8602 , n328449 );
or ( n328451 , n8580 , n8602 );
not ( n328452 , n328449 );
nand ( n8605 , n328452 , n554 );
nand ( n328454 , n328451 , n8605 );
buf ( n328455 , n328416 );
nand ( n8608 , n328454 , n328455 );
nand ( n8609 , n328427 , n8608 );
or ( n328458 , n8566 , n8609 );
not ( n8611 , n8475 );
not ( n328460 , n548 );
not ( n8613 , n8401 );
or ( n8614 , n328460 , n8613 );
not ( n328463 , n8401 );
nand ( n328464 , n328463 , n8447 );
nand ( n8617 , n8614 , n328464 );
not ( n328466 , n8617 );
or ( n328467 , n8611 , n328466 );
nand ( n8620 , n8471 , n8423 );
nand ( n328469 , n328467 , n8620 );
and ( n328470 , n328458 , n328469 );
and ( n328471 , n8609 , n8566 );
nor ( n8624 , n328470 , n328471 );
and ( n328473 , n8555 , n8624 );
and ( n328474 , n8375 , n8554 );
or ( n8627 , n328473 , n328474 );
not ( n328476 , n328065 );
not ( n328477 , n8371 );
or ( n8630 , n328476 , n328477 );
not ( n8631 , n8324 );
not ( n328480 , n328449 );
or ( n328481 , n8631 , n328480 );
nand ( n8634 , n328452 , n552 );
nand ( n328483 , n328481 , n8634 );
nand ( n8636 , n8564 , n328483 );
nand ( n328485 , n8630 , n8636 );
not ( n8638 , n8421 );
not ( n8639 , n548 );
not ( n328488 , n8537 );
not ( n8641 , n328488 );
or ( n8642 , n8639 , n8641 );
nand ( n328491 , n8447 , n8537 );
nand ( n328492 , n8642 , n328491 );
not ( n8645 , n328492 );
or ( n328494 , n8638 , n8645 );
nand ( n328495 , n8449 , n8475 );
nand ( n8648 , n328494 , n328495 );
or ( n328497 , n328485 , n8648 );
nand ( n328498 , n8648 , n328485 );
nand ( n8651 , n328497 , n328498 );
not ( n8652 , n8376 );
not ( n328501 , n546 );
not ( n8654 , n8466 );
not ( n328503 , n8654 );
not ( n8656 , n328503 );
or ( n8657 , n328501 , n8656 );
nand ( n328506 , n8654 , n8378 );
nand ( n328507 , n8657 , n328506 );
not ( n8660 , n328507 );
or ( n328509 , n8652 , n8660 );
nand ( n328510 , n8403 , n8417 );
nand ( n8663 , n328509 , n328510 );
and ( n328512 , n8651 , n8663 );
not ( n328513 , n8651 );
not ( n328514 , n8663 );
and ( n8667 , n328513 , n328514 );
nor ( n328516 , n328512 , n8667 );
not ( n328517 , n328516 );
or ( n8670 , n8548 , n8477 );
nand ( n328519 , n8670 , n8419 );
nand ( n328520 , n8548 , n8477 );
nand ( n8673 , n328519 , n328520 );
not ( n8674 , n8673 );
not ( n8675 , n328455 );
not ( n328524 , n8675 );
not ( n328525 , n8570 );
not ( n328526 , n328525 );
or ( n8679 , n328524 , n328526 );
nand ( n328528 , n8679 , n554 );
not ( n8681 , n328000 );
not ( n328530 , n8681 );
nand ( n8683 , n328530 , n544 );
not ( n328532 , n8683 );
xor ( n328533 , n328528 , n328532 );
not ( n8686 , n8161 );
not ( n8687 , n8686 );
not ( n328536 , n328035 );
or ( n328537 , n8687 , n328536 );
not ( n8690 , n544 );
not ( n328539 , n8410 );
not ( n328540 , n328539 );
or ( n8693 , n8690 , n328540 );
not ( n328542 , n328539 );
nand ( n328543 , n328542 , n328001 );
nand ( n8696 , n8693 , n328543 );
nand ( n8697 , n8696 , n8158 );
nand ( n328546 , n328537 , n8697 );
xnor ( n8699 , n328533 , n328546 );
not ( n328548 , n8699 );
not ( n8701 , n328548 );
or ( n8702 , n8674 , n8701 );
or ( n328551 , n328548 , n8673 );
nand ( n328552 , n8702 , n328551 );
not ( n8705 , n328552 );
not ( n328554 , n8705 );
or ( n328555 , n328517 , n328554 );
not ( n8708 , n328516 );
nand ( n328557 , n328552 , n8708 );
nand ( n328558 , n328555 , n328557 );
not ( n328559 , n328558 );
buf ( n8712 , n8570 );
not ( n328561 , n8712 );
not ( n328562 , n328454 );
or ( n8715 , n328561 , n328562 );
nand ( n328564 , n328455 , n554 );
nand ( n328565 , n8715 , n328564 );
xor ( n8718 , n557 , n558 );
not ( n328567 , n8718 );
not ( n8720 , n328567 );
xor ( n328569 , n556 , n557 );
nand ( n8722 , n328567 , n328569 );
not ( n8723 , n8722 );
or ( n328572 , n8720 , n8723 );
nand ( n328573 , n328572 , n556 );
not ( n8726 , n8248 );
not ( n328575 , n328100 );
or ( n328576 , n8726 , n328575 );
nand ( n8729 , n573 , n589 );
nand ( n328578 , n328576 , n8729 );
not ( n328579 , n328578 );
not ( n328580 , n328579 );
and ( n8733 , n572 , n588 );
not ( n328582 , n572 );
and ( n8735 , n328582 , n320600 );
or ( n8736 , n8733 , n8735 );
not ( n328585 , n8736 );
or ( n328586 , n328580 , n328585 );
not ( n8739 , n8736 );
nand ( n328588 , n8739 , n328578 );
nand ( n328589 , n328586 , n328588 );
not ( n8742 , n328589 );
nand ( n328591 , n8742 , n544 );
not ( n328592 , n328591 );
xor ( n8745 , n328573 , n328592 );
not ( n8746 , n8124 );
and ( n8747 , n571 , n587 );
nor ( n328596 , n8747 , n328039 );
not ( n328597 , n328596 );
and ( n8750 , n8746 , n328597 );
not ( n328599 , n8746 );
and ( n328600 , n328599 , n328596 );
nor ( n8753 , n8750 , n328600 );
buf ( n8754 , n8753 );
and ( n8755 , n8754 , n544 );
and ( n328604 , n8745 , n8755 );
and ( n328605 , n328573 , n328592 );
or ( n8758 , n328604 , n328605 );
not ( n8759 , n8758 );
nand ( n8760 , n328565 , n8759 );
not ( n8761 , n8760 );
not ( n8762 , n8686 );
not ( n328611 , n544 );
not ( n328612 , n8205 );
not ( n8765 , n328612 );
or ( n8766 , n328611 , n8765 );
nand ( n328615 , n328054 , n328001 );
nand ( n328616 , n8766 , n328615 );
not ( n8769 , n328616 );
or ( n328618 , n8762 , n8769 );
nand ( n8771 , n328003 , n8158 );
nand ( n328620 , n328618 , n8771 );
buf ( n8773 , n328620 );
not ( n8774 , n8773 );
not ( n328623 , n8417 );
not ( n328624 , n546 );
not ( n8777 , n328029 );
or ( n328626 , n328624 , n8777 );
nand ( n328627 , n8180 , n8378 );
nand ( n8780 , n328626 , n328627 );
not ( n328629 , n8780 );
or ( n328630 , n328623 , n328629 );
not ( n8783 , n8376 );
not ( n328632 , n8783 );
nand ( n328633 , n328632 , n8415 );
nand ( n8786 , n328630 , n328633 );
buf ( n8787 , n8786 );
not ( n8788 , n8787 );
or ( n328637 , n8774 , n8788 );
or ( n328638 , n8787 , n8773 );
not ( n8791 , n8546 );
not ( n8792 , n8446 );
and ( n8793 , n550 , n8792 );
not ( n8794 , n550 );
and ( n8795 , n8794 , n8446 );
or ( n328644 , n8793 , n8795 );
not ( n328645 , n328644 );
or ( n328646 , n8791 , n328645 );
nand ( n8799 , n8542 , n8485 );
nand ( n8800 , n328646 , n8799 );
nand ( n8801 , n328638 , n8800 );
nand ( n8802 , n328637 , n8801 );
not ( n8803 , n8802 );
or ( n328652 , n8761 , n8803 );
and ( n328653 , n328454 , n8570 );
not ( n328654 , n328564 );
nor ( n8807 , n328653 , n328654 );
nand ( n328656 , n8807 , n8758 );
nand ( n8809 , n328652 , n328656 );
not ( n328658 , n8207 );
not ( n328659 , n328037 );
or ( n8812 , n328658 , n328659 );
nand ( n328661 , n8812 , n8374 );
not ( n8814 , n8207 );
nand ( n8815 , n8814 , n328038 );
nand ( n328664 , n328661 , n8815 );
not ( n328665 , n8519 );
not ( n8818 , n328665 );
not ( n328667 , n8545 );
not ( n8820 , n8484 );
nand ( n328669 , n328667 , n8820 );
not ( n328670 , n328669 );
and ( n8823 , n8818 , n328670 );
not ( n328672 , n550 );
not ( n8825 , n328672 );
not ( n8826 , n8321 );
not ( n328675 , n8826 );
or ( n8828 , n8825 , n328675 );
or ( n328677 , n8826 , n328672 );
nand ( n8830 , n8828 , n328677 );
and ( n8831 , n8830 , n8484 );
nor ( n328680 , n8823 , n8831 );
and ( n8833 , n328680 , n8807 );
not ( n328682 , n328680 );
and ( n8835 , n328682 , n328565 );
nor ( n8836 , n8833 , n8835 );
xor ( n328685 , n328664 , n8836 );
not ( n328686 , n328685 );
and ( n8839 , n8809 , n328686 );
not ( n328688 , n8809 );
and ( n8841 , n328688 , n328685 );
nor ( n8842 , n8839 , n8841 );
not ( n8843 , n8842 );
and ( n328692 , n328559 , n8843 );
and ( n8845 , n328558 , n8842 );
nor ( n8846 , n328692 , n8845 );
xor ( n8847 , n8627 , n8846 );
not ( n8848 , n8158 );
not ( n8849 , n328616 );
or ( n8850 , n8848 , n8849 );
not ( n8851 , n544 );
not ( n8852 , n8754 );
not ( n8853 , n8852 );
or ( n328702 , n8851 , n8853 );
nand ( n8855 , n328001 , n8754 );
nand ( n328704 , n328702 , n8855 );
nand ( n8857 , n328704 , n8686 );
nand ( n8858 , n8850 , n8857 );
not ( n8859 , n8858 );
not ( n8860 , n8376 );
not ( n328709 , n8780 );
or ( n8862 , n8860 , n328709 );
not ( n328711 , n8417 );
not ( n328712 , n328711 );
not ( n8865 , n546 );
not ( n328714 , n8144 );
or ( n328715 , n8865 , n328714 );
nand ( n8868 , n328000 , n8378 );
nand ( n8869 , n328715 , n8868 );
nand ( n328718 , n328712 , n8869 );
nand ( n328719 , n8862 , n328718 );
not ( n8872 , n328719 );
nand ( n328721 , n8859 , n8872 );
not ( n328722 , n328721 );
not ( n328723 , n8485 );
not ( n8876 , n328644 );
or ( n328725 , n328723 , n8876 );
not ( n8878 , n550 );
not ( n8879 , n8466 );
or ( n328728 , n8878 , n8879 );
not ( n8881 , n550 );
nand ( n328730 , n8881 , n8465 );
nand ( n8883 , n328728 , n328730 );
nand ( n8884 , n8883 , n8546 );
nand ( n328733 , n328725 , n8884 );
not ( n8886 , n328733 );
or ( n328735 , n328722 , n8886 );
nand ( n8888 , n8858 , n328719 );
nand ( n8889 , n328735 , n8888 );
not ( n328738 , n8889 );
xor ( n328739 , n8609 , n8566 );
not ( n328740 , n328469 );
and ( n8893 , n328739 , n328740 );
not ( n328742 , n328739 );
and ( n328743 , n328742 , n328469 );
nor ( n8896 , n8893 , n328743 );
nand ( n328745 , n328738 , n8896 );
not ( n328746 , n8423 );
not ( n8899 , n8617 );
or ( n328748 , n328746 , n8899 );
not ( n8901 , n8475 );
not ( n8902 , n8901 );
not ( n8903 , n548 );
not ( n8904 , n8411 );
or ( n8905 , n8903 , n8904 );
nand ( n8906 , n8410 , n8447 );
nand ( n8907 , n8905 , n8906 );
nand ( n8908 , n8902 , n8907 );
nand ( n8909 , n328748 , n8908 );
not ( n8910 , n8909 );
not ( n328759 , n328455 );
not ( n328760 , n8577 );
or ( n328761 , n328759 , n328760 );
not ( n8914 , n554 );
not ( n328763 , n8321 );
or ( n328764 , n8914 , n328763 );
not ( n8917 , n554 );
nand ( n328766 , n8917 , n328168 );
nand ( n8919 , n328764 , n328766 );
nand ( n328768 , n8919 , n8570 );
nand ( n8921 , n328761 , n328768 );
not ( n328770 , n8921 );
nand ( n8923 , n8910 , n328770 );
not ( n8924 , n8923 );
not ( n328773 , n328065 );
and ( n328774 , n552 , n8540 );
not ( n328775 , n552 );
and ( n8928 , n328775 , n8537 );
or ( n328777 , n328774 , n8928 );
not ( n328778 , n328777 );
or ( n8931 , n328773 , n328778 );
nand ( n328780 , n8561 , n8564 );
nand ( n328781 , n8931 , n328780 );
not ( n8934 , n328781 );
or ( n328783 , n8924 , n8934 );
not ( n8936 , n328770 );
nand ( n328785 , n8936 , n8909 );
nand ( n8938 , n328783 , n328785 );
and ( n328787 , n328745 , n8938 );
not ( n8940 , n8889 );
nor ( n8941 , n8940 , n8896 );
nor ( n328790 , n328787 , n8941 );
not ( n328791 , n328790 );
and ( n328792 , n328565 , n8759 );
not ( n8945 , n328565 );
and ( n328794 , n8945 , n8758 );
nor ( n328795 , n328792 , n328794 );
not ( n8948 , n328795 );
and ( n328797 , n8802 , n8948 );
not ( n328798 , n8802 );
and ( n8951 , n328798 , n328795 );
nor ( n328800 , n328797 , n8951 );
not ( n8953 , n328800 );
and ( n328802 , n328791 , n8953 );
nand ( n8955 , n328790 , n328800 );
xor ( n328804 , n328573 , n328592 );
xor ( n8957 , n328804 , n8755 );
not ( n8958 , n8957 );
not ( n328807 , n544 );
not ( n328808 , n589 );
not ( n8961 , n328808 );
not ( n328810 , n573 );
not ( n8963 , n328810 );
or ( n328812 , n8961 , n8963 );
nand ( n8965 , n573 , n589 );
nand ( n8966 , n328812 , n8965 );
not ( n8967 , n8966 );
nand ( n8968 , n575 , n591 );
nor ( n8969 , n574 , n590 );
or ( n8970 , n8968 , n8969 );
nand ( n8971 , n574 , n590 );
nand ( n8972 , n8970 , n8971 );
not ( n8973 , n8972 );
or ( n328822 , n8967 , n8973 );
not ( n8975 , n327962 );
not ( n8976 , n328808 );
not ( n8977 , n328810 );
or ( n8978 , n8976 , n8977 );
nand ( n8979 , n8978 , n8965 );
not ( n8980 , n8979 );
nand ( n8981 , n8975 , n8980 );
nand ( n8982 , n328822 , n8981 );
buf ( n8983 , n8982 );
not ( n328832 , n8983 );
or ( n8985 , n328807 , n328832 );
nand ( n328834 , n8985 , n558 );
not ( n8987 , n328834 );
nand ( n328836 , n328592 , n8987 );
not ( n8989 , n328836 );
not ( n8990 , n328567 );
not ( n328839 , n556 );
not ( n328840 , n328839 );
and ( n328841 , n8990 , n328840 );
and ( n8994 , n556 , n328449 );
not ( n328843 , n556 );
not ( n328844 , n8600 );
and ( n8997 , n328843 , n328844 );
nor ( n328846 , n8994 , n8997 );
not ( n328847 , n8722 );
and ( n9000 , n328846 , n328847 );
nor ( n328849 , n328841 , n9000 );
not ( n328850 , n328849 );
not ( n9003 , n328850 );
or ( n328852 , n8989 , n9003 );
not ( n328853 , n8987 );
nand ( n9006 , n328853 , n328591 );
nand ( n328855 , n328852 , n9006 );
not ( n9008 , n328855 );
nand ( n9009 , n8958 , n9008 );
not ( n9010 , n9009 );
xor ( n9011 , n8786 , n328620 );
and ( n9012 , n328644 , n8546 );
and ( n9013 , n8542 , n8485 );
nor ( n9014 , n9012 , n9013 );
and ( n328863 , n9011 , n9014 );
not ( n9016 , n9011 );
and ( n9017 , n9016 , n8800 );
nor ( n9018 , n328863 , n9017 );
not ( n9019 , n9018 );
not ( n9020 , n9019 );
or ( n9021 , n9010 , n9020 );
not ( n9022 , n9008 );
nand ( n9023 , n9022 , n8957 );
nand ( n9024 , n9021 , n9023 );
and ( n328873 , n8955 , n9024 );
nor ( n328874 , n328802 , n328873 );
xor ( n9027 , n8847 , n328874 );
xor ( n328876 , n8375 , n8554 );
xor ( n328877 , n328876 , n8624 );
not ( n9030 , n328849 );
not ( n328879 , n328591 );
not ( n9032 , n8987 );
or ( n9033 , n328879 , n9032 );
or ( n328882 , n8987 , n328591 );
nand ( n328883 , n9033 , n328882 );
not ( n9036 , n328883 );
and ( n328885 , n9030 , n9036 );
and ( n9038 , n328849 , n328883 );
nor ( n328887 , n328885 , n9038 );
not ( n328888 , n544 );
not ( n9041 , n8736 );
not ( n328890 , n328579 );
or ( n9043 , n9041 , n328890 );
nand ( n328892 , n9043 , n328588 );
not ( n9045 , n328892 );
or ( n328894 , n328888 , n9045 );
not ( n328895 , n328892 );
nand ( n9048 , n328895 , n328001 );
nand ( n328897 , n328894 , n9048 );
buf ( n328898 , n328897 );
nand ( n9051 , n328898 , n8686 );
not ( n9052 , n9051 );
nand ( n328901 , n328704 , n8158 );
not ( n9054 , n328901 );
or ( n328903 , n9052 , n9054 );
not ( n9056 , n558 );
and ( n328905 , n8983 , n9056 , n544 );
not ( n328906 , n328905 );
nand ( n9059 , n328906 , n328834 );
nand ( n328908 , n328903 , n9059 );
nand ( n9061 , n328887 , n328908 );
not ( n9062 , n9061 );
buf ( n9063 , n8546 );
not ( n328912 , n9063 );
not ( n328913 , n328672 );
buf ( n328914 , n8395 );
not ( n9067 , n328914 );
or ( n328916 , n328913 , n9067 );
nand ( n328917 , n550 , n8401 );
nand ( n9070 , n328916 , n328917 );
not ( n328919 , n9070 );
or ( n9072 , n328912 , n328919 );
nand ( n9073 , n8883 , n8484 );
nand ( n9074 , n9072 , n9073 );
not ( n9075 , n8570 );
not ( n9076 , n8211 );
not ( n328925 , n8512 );
or ( n9078 , n9076 , n328925 );
or ( n328927 , n8512 , n8211 );
nand ( n9080 , n9078 , n328927 );
not ( n328929 , n9080 );
or ( n9082 , n9075 , n328929 );
nand ( n9083 , n8919 , n328455 );
nand ( n328932 , n9082 , n9083 );
nor ( n9085 , n9074 , n328932 );
not ( n328934 , n556 );
not ( n9087 , n8367 );
or ( n9088 , n328934 , n9087 );
or ( n328937 , n8367 , n556 );
nand ( n328938 , n9088 , n328937 );
nand ( n9091 , n328847 , n328938 );
buf ( n328940 , n8718 );
nand ( n328941 , n328846 , n328940 );
and ( n9094 , n9091 , n328941 );
or ( n328943 , n9085 , n9094 );
nand ( n328944 , n9074 , n328932 );
nand ( n328945 , n328943 , n328944 );
not ( n9098 , n328945 );
or ( n328947 , n9062 , n9098 );
not ( n9100 , n328908 );
not ( n328949 , n328887 );
nand ( n9102 , n9100 , n328949 );
nand ( n328951 , n328947 , n9102 );
not ( n9104 , n328951 );
not ( n9105 , n9104 );
xor ( n328954 , n328855 , n8957 );
not ( n328955 , n328954 );
not ( n9108 , n328955 );
not ( n328957 , n9019 );
or ( n328958 , n9108 , n328957 );
nand ( n328959 , n9018 , n328954 );
nand ( n9112 , n328958 , n328959 );
not ( n328961 , n9112 );
not ( n328962 , n328961 );
or ( n9115 , n9105 , n328962 );
not ( n328964 , n8376 );
not ( n9117 , n8869 );
or ( n9118 , n328964 , n9117 );
and ( n9119 , n8205 , n8378 );
not ( n328968 , n8205 );
and ( n9121 , n328968 , n546 );
or ( n328970 , n9119 , n9121 );
nand ( n9123 , n328970 , n8417 );
nand ( n9124 , n9118 , n9123 );
not ( n328973 , n9124 );
not ( n328974 , n8475 );
not ( n328975 , n548 );
not ( n9128 , n328032 );
or ( n328977 , n328975 , n9128 );
nand ( n328978 , n8180 , n8447 );
nand ( n9131 , n328977 , n328978 );
not ( n328980 , n9131 );
or ( n328981 , n328974 , n328980 );
not ( n9134 , n8422 );
nand ( n328983 , n8907 , n9134 );
nand ( n328984 , n328981 , n328983 );
not ( n328985 , n328984 );
or ( n9138 , n328973 , n328985 );
not ( n328987 , n328065 );
not ( n9140 , n552 );
not ( n9141 , n8443 );
or ( n328990 , n9140 , n9141 );
nand ( n328991 , n8446 , n8324 );
nand ( n328992 , n328990 , n328991 );
not ( n9145 , n328992 );
or ( n328994 , n328987 , n9145 );
nand ( n328995 , n328777 , n8564 );
nand ( n9148 , n328994 , n328995 );
not ( n328997 , n328984 );
not ( n328998 , n9124 );
nand ( n9151 , n328997 , n328998 );
nand ( n329000 , n9148 , n9151 );
nand ( n329001 , n9138 , n329000 );
not ( n9154 , n328719 );
not ( n329003 , n8859 );
or ( n9156 , n9154 , n329003 );
nand ( n329005 , n8858 , n8872 );
nand ( n9158 , n9156 , n329005 );
and ( n9159 , n9158 , n328733 );
not ( n329008 , n9158 );
not ( n329009 , n328733 );
and ( n329010 , n329008 , n329009 );
nor ( n9163 , n9159 , n329010 );
or ( n329012 , n329001 , n9163 );
xor ( n329013 , n8921 , n8909 );
xor ( n9166 , n329013 , n328781 );
nand ( n329015 , n329012 , n9166 );
nand ( n329016 , n9163 , n329001 );
nand ( n9169 , n329015 , n329016 );
nand ( n329018 , n9115 , n9169 );
not ( n329019 , n328961 );
nand ( n9172 , n329019 , n328951 );
and ( n329021 , n329018 , n9172 );
xor ( n329022 , n328877 , n329021 );
not ( n9175 , n328800 );
and ( n329024 , n9024 , n9175 );
not ( n9177 , n9024 );
and ( n329026 , n9177 , n328800 );
nor ( n9179 , n329024 , n329026 );
xor ( n9180 , n9179 , n328790 );
and ( n9181 , n329022 , n9180 );
and ( n9182 , n328877 , n329021 );
or ( n329031 , n9181 , n9182 );
nand ( n329032 , n9027 , n329031 );
not ( n9185 , n328546 );
nand ( n9186 , n9185 , n8683 );
and ( n9187 , n9186 , n328528 );
and ( n9188 , n328546 , n328532 );
nor ( n9189 , n9187 , n9188 );
not ( n329038 , n328065 );
not ( n329039 , n328483 );
or ( n329040 , n329038 , n329039 );
nand ( n9193 , n8564 , n552 );
nand ( n329042 , n329040 , n9193 );
not ( n9195 , n8423 );
and ( n9196 , n8517 , n548 );
not ( n329045 , n8517 );
and ( n9198 , n329045 , n8447 );
or ( n329047 , n9196 , n9198 );
not ( n329048 , n329047 );
or ( n329049 , n9195 , n329048 );
nand ( n9202 , n328492 , n8475 );
nand ( n329051 , n329049 , n9202 );
xor ( n9204 , n329042 , n329051 );
buf ( n329053 , n8158 );
not ( n329054 , n329053 );
xor ( n9207 , n328463 , n544 );
not ( n329056 , n9207 );
or ( n329057 , n329054 , n329056 );
nand ( n9210 , n8696 , n8686 );
nand ( n9211 , n329057 , n9210 );
xor ( n329060 , n9204 , n9211 );
xor ( n329061 , n9189 , n329060 );
or ( n9214 , n8663 , n328485 );
and ( n9215 , n9214 , n8648 );
and ( n9216 , n8663 , n328485 );
nor ( n9217 , n9215 , n9216 );
xor ( n329066 , n329061 , n9217 );
not ( n9219 , n328516 );
not ( n9220 , n8673 );
not ( n9221 , n9220 );
and ( n9222 , n9219 , n9221 );
nand ( n9223 , n9220 , n328516 );
and ( n9224 , n9223 , n328548 );
nor ( n9225 , n9222 , n9224 );
not ( n329074 , n9225 );
not ( n9227 , n328664 );
nand ( n329076 , n328680 , n8807 );
not ( n329077 , n329076 );
or ( n9230 , n9227 , n329077 );
not ( n329079 , n328680 );
nand ( n329080 , n329079 , n328565 );
nand ( n9233 , n9230 , n329080 );
not ( n329082 , n9233 );
not ( n9235 , n328029 );
nand ( n9236 , n9235 , n544 );
not ( n9237 , n8484 );
and ( n9238 , n550 , n8367 );
not ( n9239 , n550 );
and ( n9240 , n9239 , n328423 );
or ( n9241 , n9238 , n9240 );
not ( n9242 , n9241 );
or ( n9243 , n9237 , n9242 );
nand ( n9244 , n8830 , n8546 );
nand ( n329093 , n9243 , n9244 );
not ( n9246 , n329093 );
xor ( n9247 , n9236 , n9246 );
buf ( n9248 , n8443 );
and ( n9249 , n9248 , n546 );
not ( n9250 , n9248 );
and ( n9251 , n9250 , n8378 );
or ( n329100 , n9249 , n9251 );
not ( n9253 , n329100 );
not ( n329102 , n9253 );
not ( n329103 , n8783 );
and ( n9256 , n329102 , n329103 );
buf ( n329105 , n8417 );
and ( n329106 , n328507 , n329105 );
nor ( n329107 , n9256 , n329106 );
xor ( n9260 , n9247 , n329107 );
not ( n329109 , n9260 );
or ( n329110 , n329082 , n329109 );
or ( n9263 , n9233 , n9260 );
nand ( n9264 , n329110 , n9263 );
not ( n329113 , n9264 );
and ( n329114 , n329074 , n329113 );
and ( n9267 , n9225 , n9264 );
nor ( n329116 , n329114 , n9267 );
xor ( n329117 , n329066 , n329116 );
buf ( n9270 , n328558 );
not ( n329119 , n328685 );
not ( n9272 , n8809 );
nand ( n329121 , n329119 , n9272 );
and ( n329122 , n9270 , n329121 );
not ( n9275 , n328685 );
nor ( n329124 , n9275 , n9272 );
nor ( n329125 , n329122 , n329124 );
xor ( n9278 , n329117 , n329125 );
xor ( n329127 , n8627 , n8846 );
and ( n329128 , n329127 , n328874 );
and ( n329129 , n8627 , n8846 );
or ( n329130 , n329128 , n329129 );
nand ( n9283 , n9278 , n329130 );
and ( n329132 , n329032 , n9283 );
not ( n9285 , n329132 );
not ( n329134 , n9134 );
not ( n329135 , n9131 );
or ( n329136 , n329134 , n329135 );
not ( n329137 , n548 );
not ( n329138 , n8143 );
not ( n9291 , n329138 );
or ( n329140 , n329137 , n9291 );
not ( n329141 , n8151 );
not ( n9294 , n327997 );
or ( n329143 , n329141 , n9294 );
nand ( n329144 , n329143 , n8447 );
nand ( n9297 , n329140 , n329144 );
nand ( n329146 , n9297 , n8475 );
nand ( n329147 , n329136 , n329146 );
not ( n9300 , n329147 );
not ( n329149 , n8376 );
not ( n9302 , n328970 );
or ( n9303 , n329149 , n9302 );
not ( n9304 , n546 );
not ( n9305 , n8753 );
not ( n9306 , n9305 );
or ( n9307 , n9304 , n9306 );
not ( n9308 , n546 );
nand ( n9309 , n9308 , n8753 );
nand ( n9310 , n9307 , n9309 );
nand ( n9311 , n9310 , n8417 );
nand ( n9312 , n9303 , n9311 );
buf ( n9313 , n9312 );
not ( n9314 , n9313 );
or ( n9315 , n9300 , n9314 );
not ( n9316 , n329147 );
not ( n9317 , n9316 );
not ( n9318 , n9313 );
not ( n9319 , n9318 );
or ( n9320 , n9317 , n9319 );
not ( n9321 , n8372 );
not ( n9322 , n328992 );
or ( n9323 , n9321 , n9322 );
not ( n9324 , n552 );
not ( n9325 , n8464 );
or ( n9326 , n9324 , n9325 );
nand ( n9327 , n8465 , n8324 );
nand ( n9328 , n9326 , n9327 );
not ( n9329 , n328064 );
nand ( n9330 , n9328 , n9329 );
nand ( n9331 , n9323 , n9330 );
nand ( n9332 , n9320 , n9331 );
nand ( n9333 , n9315 , n9332 );
not ( n9334 , n328940 );
not ( n9335 , n328938 );
or ( n9336 , n9334 , n9335 );
xor ( n9337 , n8315 , n556 );
xnor ( n9338 , n9337 , n8311 );
not ( n9339 , n9338 );
nand ( n9340 , n9339 , n328847 );
nand ( n9341 , n9336 , n9340 );
not ( n9342 , n9341 );
not ( n9343 , n9342 );
not ( n9344 , n8820 );
not ( n9345 , n9344 );
not ( n9346 , n9070 );
or ( n9347 , n9345 , n9346 );
not ( n9348 , n328669 );
xor ( n9349 , n550 , n8410 );
nand ( n9350 , n9348 , n9349 );
nand ( n9351 , n9347 , n9350 );
not ( n9352 , n9351 );
not ( n9353 , n9352 );
and ( n9354 , n9343 , n9353 );
nand ( n9355 , n9342 , n9352 );
not ( n9356 , n544 );
xor ( n9357 , n574 , n590 );
nand ( n9358 , n575 , n591 );
not ( n9359 , n9358 );
and ( n9360 , n9357 , n9359 );
not ( n9361 , n9357 );
and ( n9362 , n9361 , n9358 );
nor ( n9363 , n9360 , n9362 );
not ( n9364 , n9363 );
not ( n9365 , n9364 );
or ( n9366 , n9356 , n9365 );
nand ( n9367 , n9363 , n328001 );
nand ( n9368 , n9366 , n9367 );
not ( n9369 , n9368 );
not ( n9370 , n8686 );
or ( n9371 , n9369 , n9370 );
not ( n9372 , n544 );
and ( n9373 , n8972 , n8966 );
not ( n9374 , n8972 );
and ( n9375 , n9374 , n8980 );
nor ( n9376 , n9373 , n9375 );
not ( n9377 , n9376 );
or ( n9378 , n9372 , n9377 );
nand ( n9379 , n8982 , n328001 );
nand ( n9380 , n9378 , n9379 );
nand ( n9381 , n9380 , n8158 );
nand ( n9382 , n9371 , n9381 );
not ( n9383 , n9382 );
not ( n9384 , n575 );
not ( n9385 , n591 );
not ( n9386 , n9385 );
or ( n9387 , n9384 , n9386 );
not ( n9388 , n575 );
nand ( n9389 , n9388 , n591 );
nand ( n9390 , n9387 , n9389 );
buf ( n9391 , n9390 );
nand ( n9392 , n9391 , n544 );
nand ( n9393 , n9383 , n9392 );
not ( n9394 , n9393 );
not ( n9395 , n8376 );
not ( n9396 , n9310 );
or ( n9397 , n9395 , n9396 );
not ( n9398 , n328711 );
not ( n9399 , n328895 );
not ( n9400 , n8378 );
or ( n9401 , n9399 , n9400 );
nand ( n9402 , n546 , n328892 );
nand ( n9403 , n9401 , n9402 );
nand ( n9404 , n9398 , n9403 );
nand ( n9405 , n9397 , n9404 );
not ( n9406 , n9405 );
or ( n9407 , n9394 , n9406 );
not ( n9408 , n9392 );
nand ( n9409 , n9408 , n9382 );
nand ( n9410 , n9407 , n9409 );
buf ( n9411 , n9410 );
and ( n9412 , n9355 , n9411 );
nor ( n9413 , n9354 , n9412 );
xor ( n9414 , n9333 , n9413 );
not ( n9415 , n8570 );
not ( n9416 , n9080 );
or ( n9417 , n9415 , n9416 );
nand ( n9418 , n9417 , n9083 );
not ( n9419 , n328847 );
not ( n9420 , n328938 );
or ( n9421 , n9419 , n9420 );
nand ( n9422 , n9421 , n328941 );
not ( n9423 , n9422 );
and ( n9424 , n9418 , n9423 );
not ( n9425 , n9418 );
and ( n9426 , n9425 , n9422 );
nor ( n9427 , n9424 , n9426 );
buf ( n9428 , n9074 );
not ( n9429 , n9428 );
and ( n9430 , n9427 , n9429 );
not ( n9431 , n9427 );
and ( n9432 , n9431 , n9428 );
nor ( n9433 , n9430 , n9432 );
xor ( n9434 , n9414 , n9433 );
buf ( n9435 , n9434 );
not ( n9436 , n9435 );
not ( n9437 , n9316 );
not ( n9438 , n9312 );
or ( n9439 , n9437 , n9438 );
not ( n9440 , n9312 );
nand ( n9441 , n9440 , n329147 );
nand ( n9442 , n9439 , n9441 );
and ( n9443 , n9442 , n9331 );
not ( n9444 , n9442 );
not ( n9445 , n9331 );
and ( n9446 , n9444 , n9445 );
nor ( n9447 , n9443 , n9446 );
not ( n9448 , n9447 );
not ( n9449 , n552 );
not ( n9450 , n8396 );
or ( n9451 , n9449 , n9450 );
nand ( n9452 , n320990 , n8395 );
nand ( n9453 , n9451 , n9452 );
not ( n9454 , n9453 );
not ( n9455 , n9454 );
not ( n9456 , n328064 );
and ( n9457 , n9455 , n9456 );
and ( n9458 , n9328 , n8372 );
nor ( n9459 , n9457 , n9458 );
not ( n9460 , n559 );
nand ( n9461 , n9460 , n558 );
not ( n9462 , n9461 );
not ( n9463 , n9462 );
and ( n9464 , n558 , n8361 );
and ( n9465 , n8362 , n9056 );
nor ( n9466 , n9464 , n9465 );
not ( n9467 , n9466 );
buf ( n9468 , n8357 );
not ( n9469 , n9468 );
or ( n9470 , n9467 , n9469 );
or ( n9471 , n9468 , n9466 );
nand ( n9472 , n9470 , n9471 );
not ( n9473 , n9472 );
or ( n9474 , n9463 , n9473 );
not ( n9475 , n558 );
not ( n9476 , n328844 );
or ( n9477 , n9475 , n9476 );
nand ( n9478 , n8600 , n9056 );
nand ( n9479 , n9477 , n9478 );
nand ( n9480 , n9479 , n559 );
nand ( n9481 , n9474 , n9480 );
not ( n9482 , n9481 );
nand ( n9483 , n9459 , n9482 );
not ( n9484 , n9483 );
not ( n9485 , n328940 );
not ( n9486 , n9338 );
not ( n9487 , n9486 );
or ( n9488 , n9485 , n9487 );
xor ( n9489 , n8491 , n556 );
buf ( n9490 , n8505 );
and ( n9491 , n9489 , n9490 );
not ( n9492 , n9489 );
not ( n9493 , n9490 );
and ( n9494 , n9492 , n9493 );
nor ( n9495 , n9491 , n9494 );
nand ( n9496 , n9495 , n328847 );
nand ( n9497 , n9488 , n9496 );
not ( n9498 , n9497 );
or ( n9499 , n9484 , n9498 );
not ( n9500 , n9482 );
not ( n9501 , n9459 );
nand ( n9502 , n9500 , n9501 );
nand ( n9503 , n9499 , n9502 );
not ( n9504 , n9503 );
nand ( n9505 , n9448 , n9504 );
not ( n9506 , n9505 );
xor ( n9507 , n9341 , n9410 );
and ( n9508 , n9507 , n9351 );
not ( n9509 , n9507 );
and ( n9510 , n9509 , n9352 );
nor ( n9511 , n9508 , n9510 );
not ( n9512 , n9511 );
or ( n9513 , n9506 , n9512 );
nand ( n9514 , n9503 , n9447 );
nand ( n9515 , n9513 , n9514 );
not ( n9516 , n9515 );
not ( n9517 , n328997 );
not ( n9518 , n9124 );
or ( n9519 , n9517 , n9518 );
nand ( n9520 , n328998 , n328984 );
nand ( n9521 , n9519 , n9520 );
and ( n9522 , n9521 , n9148 );
not ( n9523 , n9521 );
not ( n9524 , n9148 );
and ( n9525 , n9523 , n9524 );
nor ( n9526 , n9522 , n9525 );
not ( n9527 , n9526 );
not ( n9528 , n8686 );
not ( n9529 , n328898 );
or ( n329378 , n9528 , n9529 );
nand ( n9531 , n329378 , n328901 );
xor ( n9532 , n9531 , n9059 );
not ( n329381 , n9532 );
and ( n329382 , n9357 , n9359 );
not ( n9535 , n9357 );
and ( n329384 , n9535 , n9358 );
nor ( n329385 , n329382 , n329384 );
buf ( n9538 , n329385 );
nand ( n329387 , n9538 , n544 );
not ( n329388 , n329387 );
not ( n9541 , n9056 );
not ( n329390 , n1768 );
and ( n9543 , n9541 , n329390 );
not ( n329392 , n9461 );
and ( n9545 , n9479 , n329392 );
nor ( n9546 , n9543 , n9545 );
not ( n9547 , n9546 );
or ( n9548 , n329388 , n9547 );
not ( n9549 , n8158 );
not ( n9550 , n328898 );
or ( n9551 , n9549 , n9550 );
nand ( n9552 , n9380 , n8686 );
nand ( n9553 , n9551 , n9552 );
nand ( n9554 , n9548 , n9553 );
not ( n9555 , n9546 );
not ( n9556 , n329387 );
nand ( n9557 , n9555 , n9556 );
and ( n9558 , n9554 , n9557 );
not ( n9559 , n9558 );
and ( n9560 , n329381 , n9559 );
and ( n9561 , n9558 , n9532 );
nor ( n9562 , n9560 , n9561 );
and ( n9563 , n9527 , n9562 );
not ( n9564 , n9527 );
not ( n9565 , n9562 );
and ( n9566 , n9564 , n9565 );
nor ( n9567 , n9563 , n9566 );
not ( n9568 , n9134 );
not ( n9569 , n9297 );
or ( n9570 , n9568 , n9569 );
and ( n9571 , n548 , n8205 );
not ( n9572 , n548 );
not ( n9573 , n8205 );
and ( n9574 , n9572 , n9573 );
nor ( n9575 , n9571 , n9574 );
nand ( n9576 , n8473 , n8422 );
not ( n9577 , n9576 );
nand ( n9578 , n9575 , n9577 );
nand ( n9579 , n9570 , n9578 );
not ( n9580 , n9579 );
not ( n9581 , n9063 );
and ( n9582 , n550 , n328032 );
not ( n9583 , n550 );
and ( n9584 , n9583 , n8180 );
or ( n9585 , n9582 , n9584 );
not ( n9586 , n9585 );
or ( n9587 , n9581 , n9586 );
nand ( n9588 , n9349 , n8484 );
nand ( n9589 , n9587 , n9588 );
not ( n9590 , n9589 );
not ( n9591 , n9590 );
not ( n9592 , n9591 );
or ( n9593 , n9580 , n9592 );
not ( n9594 , n9579 );
not ( n9595 , n9594 );
not ( n9596 , n9590 );
or ( n9597 , n9595 , n9596 );
and ( n9598 , n9390 , n328001 );
not ( n9599 , n9390 );
and ( n9600 , n9599 , n544 );
nor ( n9601 , n9598 , n9600 );
not ( n9602 , n9601 );
not ( n9603 , n8161 );
and ( n9604 , n9602 , n9603 );
and ( n9605 , n9368 , n8158 );
nor ( n9606 , n9604 , n9605 );
not ( n9607 , n9606 );
or ( n9608 , n545 , n546 );
and ( n9609 , n9391 , n9608 );
not ( n9610 , n545 );
not ( n9611 , n546 );
or ( n9612 , n9610 , n9611 );
nand ( n9613 , n9612 , n544 );
nor ( n9614 , n9609 , n9613 );
nand ( n9615 , n9607 , n9614 );
not ( n9616 , n9615 );
nand ( n9617 , n9597 , n9616 );
nand ( n9618 , n9593 , n9617 );
not ( n9619 , n9618 );
not ( n9620 , n8570 );
and ( n9621 , n8211 , n328488 );
not ( n9622 , n8211 );
and ( n9623 , n9622 , n8537 );
nor ( n9624 , n9621 , n9623 );
not ( n9625 , n9624 );
or ( n9626 , n9620 , n9625 );
nand ( n9627 , n9080 , n328455 );
nand ( n9628 , n9626 , n9627 );
not ( n9629 , n9628 );
not ( n9630 , n8158 );
not ( n9631 , n328897 );
or ( n9632 , n9630 , n9631 );
nand ( n9633 , n9632 , n9552 );
and ( n9634 , n9633 , n9556 );
not ( n9635 , n9633 );
and ( n9636 , n9635 , n329387 );
nor ( n9637 , n9634 , n9636 );
and ( n9638 , n9637 , n9555 );
not ( n9639 , n9637 );
and ( n9640 , n9639 , n9546 );
nor ( n9641 , n9638 , n9640 );
not ( n9642 , n9641 );
nand ( n9643 , n9629 , n9642 );
not ( n9644 , n9643 );
or ( n9645 , n9619 , n9644 );
not ( n9646 , n9642 );
nand ( n9647 , n9646 , n9628 );
nand ( n9648 , n9645 , n9647 );
not ( n9649 , n9648 );
and ( n9650 , n9567 , n9649 );
not ( n9651 , n9567 );
and ( n9652 , n9651 , n9648 );
nor ( n9653 , n9650 , n9652 );
not ( n9654 , n9653 );
or ( n9655 , n9516 , n9654 );
not ( n9656 , n9653 );
not ( n9657 , n9515 );
nand ( n9658 , n9656 , n9657 );
nand ( n9659 , n9655 , n9658 );
or ( n9660 , n9436 , n9659 );
xor ( n9661 , n9615 , n9589 );
xnor ( n9662 , n9661 , n9594 );
not ( n9663 , n8484 );
not ( n9664 , n9585 );
or ( n9665 , n9663 , n9664 );
and ( n9666 , n8514 , n8143 );
not ( n9667 , n8514 );
and ( n9668 , n9667 , n329138 );
nor ( n9669 , n9666 , n9668 );
not ( n9670 , n9669 );
nand ( n9671 , n9670 , n8546 );
nand ( n9672 , n9665 , n9671 );
buf ( n9673 , n9462 );
not ( n9674 , n9673 );
not ( n9675 , n558 );
not ( n9676 , n8321 );
or ( n9677 , n9675 , n9676 );
nand ( n9678 , n9056 , n328168 );
nand ( n9679 , n9677 , n9678 );
not ( n9680 , n9679 );
or ( n9681 , n9674 , n9680 );
not ( n9682 , n1768 );
nand ( n9683 , n9682 , n9472 );
nand ( n9684 , n9681 , n9683 );
or ( n9685 , n9672 , n9684 );
not ( n9686 , n328065 );
not ( n9687 , n552 );
not ( n9688 , n8411 );
or ( n329537 , n9687 , n9688 );
nand ( n329538 , n8410 , n8324 );
nand ( n329539 , n329537 , n329538 );
not ( n329540 , n329539 );
or ( n9693 , n9686 , n329540 );
nand ( n329542 , n9453 , n328061 );
nand ( n329543 , n9693 , n329542 );
nand ( n9696 , n9685 , n329543 );
nand ( n9697 , n9672 , n9684 );
nand ( n329546 , n9696 , n9697 );
not ( n329547 , n329546 );
nand ( n9700 , n9662 , n329547 );
not ( n329549 , n9700 );
not ( n9702 , n8712 );
and ( n9703 , n8466 , n554 );
not ( n9704 , n8466 );
and ( n9705 , n9704 , n8211 );
or ( n329554 , n9703 , n9705 );
not ( n9707 , n329554 );
or ( n329556 , n9702 , n9707 );
not ( n329557 , n554 );
not ( n9710 , n8443 );
or ( n329559 , n329557 , n9710 );
not ( n329560 , n554 );
nand ( n9713 , n329560 , n8442 );
nand ( n329562 , n329559 , n9713 );
buf ( n9715 , n329562 );
nand ( n329564 , n9715 , n328455 );
nand ( n9717 , n329556 , n329564 );
not ( n9718 , n9717 );
not ( n329567 , n328847 );
xor ( n329568 , n8537 , n556 );
not ( n329569 , n329568 );
or ( n9722 , n329567 , n329569 );
nand ( n329571 , n9495 , n328940 );
nand ( n329572 , n9722 , n329571 );
not ( n9725 , n329572 );
or ( n329574 , n9718 , n9725 );
not ( n329575 , n329572 );
not ( n9728 , n329575 );
not ( n329577 , n9715 );
not ( n329578 , n329577 );
not ( n9731 , n8675 );
and ( n329580 , n329578 , n9731 );
and ( n9733 , n329554 , n8712 );
nor ( n9734 , n329580 , n9733 );
not ( n329583 , n9734 );
or ( n329584 , n9728 , n329583 );
not ( n329585 , n8376 );
not ( n9738 , n546 );
not ( n329587 , n9376 );
or ( n329588 , n9738 , n329587 );
nand ( n9741 , n8982 , n8378 );
nand ( n329590 , n329588 , n9741 );
not ( n329591 , n329590 );
or ( n9744 , n329585 , n329591 );
not ( n329593 , n546 );
not ( n9746 , n9364 );
or ( n329595 , n329593 , n9746 );
nand ( n9748 , n8378 , n329385 );
nand ( n329597 , n329595 , n9748 );
nor ( n9750 , n8416 , n8376 );
nand ( n9751 , n329597 , n9750 );
nand ( n329600 , n9744 , n9751 );
not ( n9753 , n329600 );
not ( n329602 , n575 );
not ( n9755 , n9385 );
or ( n329604 , n329602 , n9755 );
nand ( n329605 , n9388 , n591 );
nand ( n9758 , n329604 , n329605 );
nand ( n329607 , n9758 , n8158 );
nand ( n9760 , n9753 , n329607 );
not ( n9761 , n9760 );
not ( n9762 , n8376 );
not ( n9763 , n329597 );
or ( n9764 , n9762 , n9763 );
nand ( n329613 , n9390 , n8378 );
not ( n9766 , n329613 );
not ( n9767 , n9390 );
nand ( n9768 , n9767 , n546 );
not ( n9769 , n9768 );
or ( n329618 , n9766 , n9769 );
nand ( n9771 , n329618 , n9750 );
nand ( n329620 , n9764 , n9771 );
not ( n329621 , n329620 );
or ( n9774 , n547 , n548 );
not ( n9775 , n9774 );
not ( n9776 , n9390 );
not ( n9777 , n9776 );
not ( n329626 , n9777 );
or ( n9779 , n9775 , n329626 );
nand ( n329628 , n547 , n548 );
and ( n329629 , n329628 , n546 );
nand ( n9782 , n9779 , n329629 );
nor ( n9783 , n329621 , n9782 );
not ( n329632 , n9783 );
or ( n9785 , n9761 , n329632 );
or ( n9786 , n9753 , n329607 );
nand ( n329635 , n9785 , n9786 );
nand ( n9788 , n329584 , n329635 );
nand ( n9789 , n329574 , n9788 );
not ( n329638 , n9789 );
or ( n9791 , n329549 , n329638 );
not ( n329640 , n9662 );
nand ( n9793 , n329640 , n329546 );
nand ( n9794 , n9791 , n9793 );
not ( n329643 , n9794 );
and ( n9796 , n544 , n9391 );
and ( n9797 , n9382 , n9796 );
not ( n9798 , n9382 );
and ( n329647 , n9798 , n9392 );
nor ( n9800 , n9797 , n329647 );
xor ( n9801 , n9800 , n9405 );
not ( n329650 , n9801 );
not ( n329651 , n329650 );
not ( n329652 , n8570 );
not ( n9805 , n329562 );
or ( n329654 , n329652 , n9805 );
not ( n329655 , n8675 );
nand ( n9808 , n329655 , n9624 );
nand ( n329657 , n329654 , n9808 );
not ( n329658 , n329657 );
not ( n9811 , n329658 );
or ( n329660 , n329651 , n9811 );
not ( n329661 , n8376 );
not ( n9814 , n9403 );
or ( n329663 , n329661 , n9814 );
nand ( n9816 , n8417 , n329590 );
nand ( n9817 , n329663 , n9816 );
buf ( n329666 , n9817 );
not ( n329667 , n329666 );
not ( n329668 , n8422 );
not ( n9821 , n329668 );
not ( n329670 , n9575 );
or ( n329671 , n9821 , n329670 );
not ( n9824 , n548 );
not ( n329673 , n8852 );
or ( n329674 , n9824 , n329673 );
nand ( n9827 , n8754 , n8447 );
nand ( n329676 , n329674 , n9827 );
nand ( n9829 , n329676 , n8474 );
nand ( n329678 , n329671 , n9829 );
not ( n9831 , n329678 );
or ( n329680 , n329667 , n9831 );
not ( n9833 , n329666 );
not ( n9834 , n9833 );
not ( n329683 , n329678 );
not ( n329684 , n329683 );
or ( n329685 , n9834 , n329684 );
not ( n9838 , n9606 );
not ( n329687 , n9614 );
not ( n329688 , n329687 );
or ( n9841 , n9838 , n329688 );
nand ( n329690 , n9841 , n9615 );
not ( n329691 , n329690 );
nand ( n9844 , n329685 , n329691 );
nand ( n329693 , n329680 , n9844 );
nand ( n9846 , n329660 , n329693 );
or ( n329695 , n329658 , n329650 );
nand ( n9848 , n9846 , n329695 );
not ( n329697 , n9618 );
not ( n329698 , n329697 );
and ( n9851 , n9628 , n9642 );
not ( n329700 , n9628 );
and ( n329701 , n329700 , n9641 );
nor ( n9854 , n9851 , n329701 );
not ( n9855 , n9854 );
not ( n329704 , n9855 );
or ( n329705 , n329698 , n329704 );
nand ( n9858 , n9854 , n9618 );
nand ( n329707 , n329705 , n9858 );
or ( n329708 , n9848 , n329707 );
not ( n9861 , n329708 );
or ( n329710 , n329643 , n9861 );
nand ( n329711 , n329707 , n9848 );
nand ( n9864 , n329710 , n329711 );
nand ( n9865 , n9660 , n9864 );
not ( n329714 , n9435 );
nand ( n9867 , n329714 , n9659 );
nand ( n329716 , n9865 , n9867 );
not ( n9869 , n329716 );
not ( n329718 , n9869 );
not ( n329719 , n9515 );
not ( n9872 , n9648 );
not ( n9873 , n9567 );
nand ( n9874 , n9872 , n9873 );
not ( n9875 , n9874 );
or ( n9876 , n329719 , n9875 );
not ( n329725 , n9873 );
nand ( n329726 , n329725 , n9648 );
nand ( n9879 , n9876 , n329726 );
not ( n329728 , n9166 );
xor ( n9881 , n329001 , n9163 );
xnor ( n9882 , n329728 , n9881 );
not ( n9883 , n9532 );
nand ( n9884 , n9883 , n9558 );
not ( n9885 , n9884 );
not ( n9886 , n9526 );
or ( n9887 , n9885 , n9886 );
not ( n9888 , n9558 );
nand ( n9889 , n9888 , n9532 );
nand ( n9890 , n9887 , n9889 );
and ( n329739 , n328908 , n328887 );
not ( n9892 , n328908 );
and ( n329741 , n9892 , n328949 );
nor ( n9894 , n329739 , n329741 );
xnor ( n329743 , n328945 , n9894 );
not ( n329744 , n329743 );
and ( n9897 , n9890 , n329744 );
not ( n329746 , n9890 );
and ( n9899 , n329746 , n329743 );
nor ( n9900 , n9897 , n9899 );
not ( n329749 , n9333 );
not ( n329750 , n9433 );
or ( n9903 , n329749 , n329750 );
or ( n329752 , n9333 , n9433 );
not ( n9905 , n9413 );
nand ( n329754 , n329752 , n9905 );
nand ( n329755 , n9903 , n329754 );
and ( n9908 , n9900 , n329755 );
not ( n329757 , n9900 );
not ( n329758 , n329755 );
and ( n9911 , n329757 , n329758 );
nor ( n329760 , n9908 , n9911 );
xor ( n9913 , n9882 , n329760 );
xor ( n329762 , n9879 , n9913 );
not ( n9915 , n329762 );
not ( n9916 , n9915 );
or ( n329765 , n329718 , n9916 );
xor ( n329766 , n9434 , n9864 );
xnor ( n9919 , n329766 , n9659 );
not ( n329768 , n9919 );
not ( n9921 , n9848 );
and ( n329770 , n329707 , n9921 );
not ( n329771 , n329707 );
and ( n9924 , n329771 , n9848 );
nor ( n329773 , n329770 , n9924 );
not ( n329774 , n9794 );
and ( n9927 , n329773 , n329774 );
not ( n9928 , n329773 );
and ( n9929 , n9928 , n9794 );
nor ( n9930 , n9927 , n9929 );
not ( n329779 , n9930 );
and ( n329780 , n9447 , n9503 );
not ( n9933 , n9447 );
and ( n329782 , n9933 , n9504 );
nor ( n329783 , n329780 , n329782 );
not ( n9936 , n9511 );
and ( n329785 , n329783 , n9936 );
not ( n329786 , n329783 );
and ( n329787 , n329786 , n9511 );
nor ( n9940 , n329785 , n329787 );
buf ( n329789 , n9940 );
or ( n9942 , n329779 , n329789 );
not ( n329791 , n329789 );
not ( n329792 , n329779 );
or ( n9945 , n329791 , n329792 );
not ( n329794 , n329690 );
xor ( n329795 , n9817 , n329794 );
xor ( n9948 , n329678 , n329795 );
not ( n9949 , n9134 );
not ( n329798 , n329676 );
or ( n9951 , n9949 , n329798 );
not ( n329800 , n548 );
not ( n329801 , n8742 );
not ( n9954 , n329801 );
or ( n329803 , n329800 , n9954 );
not ( n9956 , n328895 );
not ( n329805 , n9956 );
nand ( n329806 , n329805 , n8447 );
nand ( n9959 , n329803 , n329806 );
nand ( n329808 , n8474 , n9959 );
nand ( n329809 , n9951 , n329808 );
not ( n9962 , n329809 );
not ( n329811 , n9669 );
not ( n329812 , n8820 );
and ( n329813 , n329811 , n329812 );
and ( n9966 , n8205 , n5763 );
not ( n329815 , n8205 );
and ( n9968 , n329815 , n550 );
or ( n9969 , n9966 , n9968 );
and ( n329818 , n9969 , n9063 );
nor ( n9971 , n329813 , n329818 );
not ( n329820 , n9971 );
not ( n9973 , n329820 );
or ( n329822 , n9962 , n9973 );
not ( n329823 , n329809 );
not ( n9976 , n329823 );
not ( n329825 , n9971 );
or ( n329826 , n9976 , n329825 );
not ( n9979 , n328065 );
not ( n329828 , n552 );
not ( n329829 , n328029 );
or ( n9982 , n329828 , n329829 );
nand ( n329831 , n328033 , n8324 );
nand ( n9984 , n9982 , n329831 );
not ( n9985 , n9984 );
or ( n329834 , n9979 , n9985 );
nand ( n329835 , n329539 , n8372 );
nand ( n329836 , n329834 , n329835 );
nand ( n9989 , n329826 , n329836 );
nand ( n329838 , n329822 , n9989 );
xor ( n329839 , n9948 , n329838 );
not ( n9992 , n558 );
not ( n329841 , n8517 );
or ( n329842 , n9992 , n329841 );
nand ( n9995 , n8512 , n9056 );
nand ( n329844 , n329842 , n9995 );
nand ( n9997 , n329844 , n9673 );
nand ( n9998 , n9679 , n559 );
nand ( n9999 , n9997 , n9998 );
not ( n10000 , n328940 );
not ( n329849 , n329568 );
or ( n329850 , n10000 , n329849 );
not ( n10003 , n556 );
not ( n329852 , n8443 );
or ( n329853 , n10003 , n329852 );
not ( n329854 , n556 );
nand ( n10007 , n329854 , n8442 );
nand ( n329856 , n329853 , n10007 );
nand ( n10009 , n329856 , n328847 );
nand ( n10010 , n329850 , n10009 );
nor ( n10011 , n9999 , n10010 );
not ( n10012 , n9783 );
not ( n10013 , n329607 );
not ( n10014 , n10013 );
not ( n10015 , n9753 );
or ( n329864 , n10014 , n10015 );
not ( n10017 , n8159 );
nand ( n10018 , n10017 , n9777 );
nand ( n10019 , n10018 , n329600 );
nand ( n10020 , n329864 , n10019 );
not ( n10021 , n10020 );
or ( n329870 , n10012 , n10021 );
or ( n329871 , n10020 , n9783 );
nand ( n10024 , n329870 , n329871 );
or ( n329873 , n10011 , n10024 );
not ( n329874 , n9997 );
not ( n10027 , n9998 );
or ( n10028 , n329874 , n10027 );
nand ( n10029 , n10028 , n10010 );
nand ( n10030 , n329873 , n10029 );
and ( n329879 , n329839 , n10030 );
and ( n329880 , n9948 , n329838 );
or ( n10033 , n329879 , n329880 );
not ( n329882 , n10033 );
xor ( n10035 , n9481 , n9497 );
xnor ( n329884 , n10035 , n9459 );
not ( n10037 , n329884 );
and ( n10038 , n329657 , n9801 );
not ( n329887 , n329657 );
and ( n10040 , n329887 , n329650 );
nor ( n329889 , n10038 , n10040 );
and ( n10042 , n329693 , n329889 );
not ( n329891 , n329693 );
not ( n329892 , n329889 );
and ( n10045 , n329891 , n329892 );
or ( n329894 , n10042 , n10045 );
nand ( n329895 , n10037 , n329894 );
not ( n329896 , n329895 );
or ( n10049 , n329882 , n329896 );
not ( n329898 , n329894 );
nand ( n10051 , n329898 , n329884 );
nand ( n10052 , n10049 , n10051 );
nand ( n329901 , n9945 , n10052 );
nand ( n10054 , n9942 , n329901 );
not ( n329903 , n10054 );
nand ( n10056 , n329768 , n329903 );
nand ( n329905 , n329765 , n10056 );
xor ( n329906 , n8889 , n8938 );
xor ( n10059 , n329906 , n8896 );
xor ( n329908 , n9104 , n9112 );
xor ( n329909 , n329908 , n9169 );
xor ( n10062 , n10059 , n329909 );
not ( n329911 , n329758 );
buf ( n10064 , n329743 );
not ( n329913 , n10064 );
and ( n10066 , n329911 , n329913 );
nand ( n10067 , n329758 , n10064 );
buf ( n329916 , n9890 );
and ( n10069 , n10067 , n329916 );
nor ( n329918 , n10066 , n10069 );
xor ( n10071 , n10062 , n329918 );
or ( n329920 , n329760 , n9882 );
and ( n329921 , n329920 , n9879 );
and ( n10074 , n9882 , n329760 );
nor ( n329923 , n329921 , n10074 );
nand ( n329924 , n10071 , n329923 );
xor ( n10077 , n328877 , n329021 );
xor ( n329926 , n10077 , n9180 );
xor ( n329927 , n10059 , n329909 );
and ( n10080 , n329927 , n329918 );
and ( n329929 , n10059 , n329909 );
or ( n329930 , n10080 , n329929 );
nand ( n329931 , n329926 , n329930 );
nand ( n10084 , n329924 , n329931 );
nor ( n329933 , n329905 , n10084 );
not ( n10086 , n329933 );
nand ( n329935 , n9696 , n9697 );
and ( n329936 , n9662 , n329935 );
not ( n10089 , n9662 );
and ( n10090 , n10089 , n329547 );
or ( n10091 , n329936 , n10090 );
not ( n10092 , n9789 );
and ( n329941 , n10091 , n10092 );
not ( n10094 , n10091 );
and ( n329943 , n10094 , n9789 );
nor ( n329944 , n329941 , n329943 );
not ( n10097 , n9497 );
xor ( n329946 , n9481 , n10097 );
xnor ( n10099 , n329946 , n9501 );
and ( n329948 , n329693 , n329889 );
not ( n10101 , n329693 );
and ( n329950 , n10101 , n329892 );
nor ( n10103 , n329948 , n329950 );
xor ( n329952 , n10099 , n10103 );
xnor ( n329953 , n329952 , n10033 );
xor ( n10106 , n329944 , n329953 );
xor ( n10107 , n9948 , n329838 );
xor ( n329956 , n10107 , n10030 );
xor ( n10109 , n9672 , n329543 );
buf ( n329958 , n9684 );
not ( n10111 , n329958 );
and ( n329960 , n10109 , n10111 );
not ( n329961 , n10109 );
and ( n10114 , n329961 , n329958 );
nor ( n329963 , n329960 , n10114 );
not ( n329964 , n329635 );
not ( n329965 , n329575 );
or ( n329966 , n329964 , n329965 );
not ( n10119 , n329635 );
nand ( n329968 , n10119 , n329572 );
nand ( n10121 , n329966 , n329968 );
and ( n329970 , n10121 , n9734 );
not ( n329971 , n10121 );
and ( n329972 , n329971 , n9717 );
nor ( n329973 , n329970 , n329972 );
nand ( n10126 , n329963 , n329973 );
and ( n329975 , n329956 , n10126 );
nor ( n329976 , n329963 , n329973 );
nor ( n10129 , n329975 , n329976 );
and ( n329978 , n10106 , n10129 );
and ( n329979 , n329944 , n329953 );
or ( n10132 , n329978 , n329979 );
not ( n10133 , n10132 );
xor ( n10134 , n9940 , n10052 );
xor ( n10135 , n10134 , n9930 );
not ( n329984 , n10135 );
or ( n329985 , n10133 , n329984 );
xor ( n10138 , n329944 , n329953 );
xor ( n329987 , n10138 , n10129 );
not ( n329988 , n328455 );
not ( n10141 , n329554 );
or ( n329990 , n329988 , n10141 );
not ( n10143 , n554 );
not ( n10144 , n8397 );
or ( n329993 , n10143 , n10144 );
nand ( n10146 , n8398 , n8211 );
nand ( n329995 , n329993 , n10146 );
nand ( n329996 , n329995 , n8570 );
nand ( n10149 , n329990 , n329996 );
not ( n329998 , n10149 );
xor ( n329999 , n329809 , n329836 );
xnor ( n10152 , n329999 , n329820 );
not ( n330001 , n10152 );
not ( n330002 , n330001 );
or ( n10155 , n329998 , n330002 );
not ( n330004 , n10149 );
not ( n330005 , n330004 );
not ( n10158 , n10152 );
or ( n330007 , n330005 , n10158 );
nand ( n10160 , n9969 , n8484 );
not ( n10161 , n548 );
buf ( n10162 , n9376 );
not ( n10163 , n10162 );
or ( n10164 , n10161 , n10163 );
not ( n10165 , n9376 );
nand ( n10166 , n10165 , n8447 );
nand ( n10167 , n10164 , n10166 );
not ( n10168 , n10167 );
not ( n330017 , n10168 );
not ( n330018 , n9576 );
and ( n10171 , n330017 , n330018 );
and ( n330020 , n9959 , n8421 );
nor ( n10173 , n10171 , n330020 );
nand ( n10174 , n10160 , n10173 );
and ( n10175 , n550 , n8852 );
not ( n10176 , n550 );
and ( n10177 , n10176 , n8754 );
or ( n10178 , n10175 , n10177 );
not ( n10179 , n10178 );
nor ( n10180 , n10179 , n328669 );
or ( n10181 , n10174 , n10180 );
not ( n10182 , n9782 );
not ( n10183 , n329620 );
or ( n10184 , n10182 , n10183 );
or ( n10185 , n9782 , n329620 );
nand ( n10186 , n10184 , n10185 );
nand ( n10187 , n10181 , n10186 );
not ( n10188 , n10173 );
not ( n10189 , n328669 );
not ( n10190 , n10189 );
not ( n10191 , n10178 );
or ( n10192 , n10190 , n10191 );
nand ( n10193 , n10192 , n10160 );
nand ( n10194 , n10188 , n10193 );
nand ( n10195 , n10187 , n10194 );
nand ( n10196 , n330007 , n10195 );
nand ( n10197 , n10155 , n10196 );
not ( n10198 , n10197 );
xnor ( n10199 , n329963 , n329973 );
xor ( n10200 , n329956 , n10199 );
nand ( n10201 , n10198 , n10200 );
and ( n10202 , n10024 , n10010 );
not ( n10203 , n10024 );
not ( n10204 , n10010 );
and ( n10205 , n10203 , n10204 );
nor ( n10206 , n10202 , n10205 );
and ( n10207 , n10206 , n9999 );
not ( n10208 , n10206 );
not ( n10209 , n9999 );
and ( n10210 , n10208 , n10209 );
nor ( n10211 , n10207 , n10210 );
not ( n10212 , n10211 );
not ( n10213 , n10212 );
not ( n10214 , n329856 );
not ( n10215 , n10214 );
not ( n10216 , n328940 );
not ( n10217 , n10216 );
and ( n10218 , n10215 , n10217 );
not ( n10219 , n556 );
not ( n10220 , n8466 );
or ( n10221 , n10219 , n10220 );
nand ( n10222 , n8465 , n328839 );
nand ( n10223 , n10221 , n10222 );
and ( n10224 , n10223 , n328847 );
nor ( n10225 , n10218 , n10224 );
not ( n10226 , n10225 );
not ( n10227 , n552 );
not ( n10228 , n8144 );
or ( n10229 , n10227 , n10228 );
not ( n10230 , n8144 );
nand ( n10231 , n10230 , n8324 );
nand ( n10232 , n10229 , n10231 );
not ( n10233 , n10232 );
not ( n10234 , n10233 );
not ( n10235 , n328064 );
and ( n10236 , n10234 , n10235 );
and ( n10237 , n9984 , n8564 );
nor ( n10238 , n10236 , n10237 );
not ( n10239 , n10238 );
and ( n10240 , n10226 , n10239 );
nand ( n10241 , n10225 , n10238 );
nand ( n10242 , n9758 , n8376 );
not ( n10243 , n10242 );
not ( n10244 , n8421 );
not ( n10245 , n10167 );
or ( n10246 , n10244 , n10245 );
and ( n10247 , n9538 , n8447 );
not ( n10248 , n9538 );
and ( n10249 , n10248 , n548 );
or ( n10250 , n10247 , n10249 );
nor ( n10251 , n8472 , n9134 );
nand ( n10252 , n10250 , n10251 );
nand ( n10253 , n10246 , n10252 );
not ( n10254 , n10253 );
not ( n10255 , n10254 );
or ( n10256 , n10243 , n10255 );
or ( n10257 , n549 , n550 );
nand ( n10258 , n10257 , n9391 );
nand ( n10259 , n549 , n550 );
and ( n10260 , n10258 , n10259 , n548 );
not ( n10261 , n8421 );
not ( n10262 , n10250 );
or ( n10263 , n10261 , n10262 );
not ( n10264 , n548 );
not ( n10265 , n9391 );
not ( n10266 , n10265 );
or ( n10267 , n10264 , n10266 );
nand ( n10268 , n8447 , n9758 );
nand ( n10269 , n10267 , n10268 );
nand ( n10270 , n10269 , n10251 );
nand ( n10271 , n10263 , n10270 );
and ( n10272 , n10260 , n10271 );
nand ( n10273 , n10256 , n10272 );
not ( n10274 , n10254 );
not ( n10275 , n10242 );
nand ( n10276 , n10274 , n10275 );
nand ( n10277 , n10273 , n10276 );
buf ( n10278 , n10277 );
and ( n10279 , n10241 , n10278 );
nor ( n10280 , n10240 , n10279 );
not ( n10281 , n10280 );
not ( n10282 , n10281 );
or ( n10283 , n10213 , n10282 );
not ( n10284 , n10280 );
not ( n10285 , n10211 );
or ( n10286 , n10284 , n10285 );
not ( n10287 , n9673 );
not ( n10288 , n558 );
not ( n10289 , n328488 );
or ( n10290 , n10288 , n10289 );
not ( n10291 , n8540 );
nand ( n10292 , n10291 , n9056 );
nand ( n10293 , n10290 , n10292 );
not ( n10294 , n10293 );
or ( n10295 , n10287 , n10294 );
nand ( n10296 , n329844 , n559 );
nand ( n10297 , n10295 , n10296 );
not ( n10298 , n10297 );
not ( n10299 , n10298 );
xnor ( n10300 , n8410 , n554 );
not ( n10301 , n10300 );
not ( n10302 , n328525 );
and ( n10303 , n10301 , n10302 );
and ( n10304 , n329995 , n328455 );
nor ( n10305 , n10303 , n10304 );
not ( n10306 , n10305 );
and ( n10307 , n10299 , n10306 );
not ( n10308 , n10173 );
not ( n10309 , n10186 );
or ( n10310 , n10308 , n10309 );
or ( n10311 , n10186 , n10173 );
nand ( n10312 , n10310 , n10311 );
and ( n10313 , n10193 , n10312 );
not ( n10314 , n10193 );
not ( n10315 , n10312 );
and ( n10316 , n10314 , n10315 );
nor ( n10317 , n10313 , n10316 );
nand ( n10318 , n10298 , n10305 );
and ( n10319 , n10317 , n10318 );
nor ( n10320 , n10307 , n10319 );
not ( n10321 , n10320 );
nand ( n10322 , n10286 , n10321 );
nand ( n10323 , n10283 , n10322 );
not ( n10324 , n10323 );
not ( n10325 , n10324 );
and ( n10326 , n10201 , n10325 );
not ( n10327 , n10197 );
nor ( n10328 , n10327 , n10200 );
nor ( n10329 , n10326 , n10328 );
nand ( n10330 , n329987 , n10329 );
nand ( n10331 , n329985 , n10330 );
not ( n10332 , n10331 );
xor ( n10333 , n10275 , n10254 );
xor ( n330182 , n10333 , n10272 );
not ( n10335 , n330182 );
not ( n330184 , n10335 );
not ( n10337 , n328847 );
and ( n330186 , n556 , n8397 );
not ( n330187 , n556 );
and ( n10340 , n330187 , n328463 );
or ( n330189 , n330186 , n10340 );
not ( n330190 , n330189 );
or ( n330191 , n10337 , n330190 );
nand ( n10344 , n328940 , n10223 );
nand ( n330193 , n330191 , n10344 );
not ( n10346 , n330193 );
not ( n10347 , n10346 );
or ( n330196 , n330184 , n10347 );
nand ( n10349 , n330193 , n330182 );
nand ( n330198 , n330196 , n10349 );
not ( n10351 , n559 );
not ( n330200 , n10293 );
or ( n330201 , n10351 , n330200 );
not ( n10354 , n558 );
not ( n330203 , n8792 );
or ( n330204 , n10354 , n330203 );
nand ( n10357 , n8446 , n9056 );
nand ( n330206 , n330204 , n10357 );
nand ( n10359 , n330206 , n9462 );
nand ( n330208 , n330201 , n10359 );
buf ( n10361 , n330208 );
not ( n10362 , n10361 );
and ( n330211 , n330198 , n10362 );
not ( n330212 , n330198 );
and ( n330213 , n330212 , n10361 );
nor ( n10366 , n330211 , n330213 );
buf ( n330215 , n10366 );
not ( n330216 , n559 );
not ( n10369 , n330206 );
or ( n330218 , n330216 , n10369 );
not ( n330219 , n558 );
not ( n10372 , n8466 );
or ( n330221 , n330219 , n10372 );
nand ( n330222 , n8654 , n9056 );
nand ( n10375 , n330221 , n330222 );
nand ( n330224 , n10375 , n9462 );
nand ( n330225 , n330218 , n330224 );
xor ( n330226 , n10162 , n550 );
not ( n10379 , n330226 );
not ( n10380 , n328669 );
and ( n330229 , n10379 , n10380 );
and ( n10382 , n5763 , n8742 );
not ( n10383 , n5763 );
and ( n330232 , n10383 , n329801 );
nor ( n330233 , n10382 , n330232 );
nor ( n330234 , n330233 , n8820 );
nor ( n10387 , n330229 , n330234 );
not ( n330236 , n10387 );
xor ( n330237 , n10260 , n10271 );
not ( n10390 , n330237 );
and ( n330239 , n330236 , n10390 );
and ( n330240 , n10387 , n330237 );
nor ( n10393 , n330239 , n330240 );
not ( n330242 , n328061 );
not ( n330243 , n8324 );
not ( n330244 , n9573 );
not ( n10397 , n330244 );
or ( n330246 , n330243 , n10397 );
not ( n10399 , n8205 );
nand ( n330248 , n10399 , n552 );
nand ( n10401 , n330246 , n330248 );
not ( n10402 , n10401 );
or ( n330251 , n330242 , n10402 );
not ( n330252 , n552 );
not ( n10405 , n8852 );
or ( n330254 , n330252 , n10405 );
nand ( n330255 , n8754 , n8324 );
nand ( n10408 , n330254 , n330255 );
nand ( n330257 , n10408 , n9329 );
nand ( n330258 , n330251 , n330257 );
not ( n10411 , n330258 );
xor ( n330260 , n10393 , n10411 );
xor ( n330261 , n330225 , n330260 );
and ( n10414 , n556 , n328032 );
not ( n330263 , n556 );
and ( n330264 , n330263 , n8180 );
or ( n10417 , n10414 , n330264 );
not ( n10418 , n10417 );
not ( n10419 , n10418 );
not ( n10420 , n8722 );
and ( n10421 , n10419 , n10420 );
and ( n330270 , n556 , n328539 );
not ( n330271 , n556 );
not ( n10424 , n8411 );
and ( n330273 , n330271 , n10424 );
or ( n330274 , n330270 , n330273 );
and ( n330275 , n330274 , n328940 );
nor ( n10428 , n10421 , n330275 );
not ( n330277 , n10428 );
not ( n10430 , n330277 );
not ( n330279 , n328525 );
not ( n330280 , n320444 );
not ( n10433 , n9573 );
or ( n10434 , n330280 , n10433 );
nand ( n330283 , n8205 , n554 );
nand ( n10436 , n10434 , n330283 );
not ( n330285 , n10436 );
and ( n330286 , n330279 , n330285 );
not ( n330287 , n554 );
not ( n10440 , n8681 );
or ( n330289 , n330287 , n10440 );
nand ( n10442 , n10230 , n8211 );
nand ( n330291 , n330289 , n10442 );
and ( n330292 , n330291 , n328455 );
nor ( n10445 , n330286 , n330292 );
not ( n330294 , n10445 );
not ( n330295 , n330294 );
or ( n10448 , n10430 , n330295 );
not ( n330297 , n10445 );
not ( n330298 , n10428 );
or ( n10451 , n330297 , n330298 );
not ( n330300 , n8485 );
not ( n330301 , n550 );
not ( n330302 , n9538 );
not ( n10455 , n330302 );
or ( n330304 , n330301 , n10455 );
not ( n330305 , n550 );
nand ( n10458 , n330305 , n9538 );
nand ( n330307 , n330304 , n10458 );
not ( n330308 , n330307 );
or ( n10461 , n330300 , n330308 );
and ( n330310 , n550 , n9776 );
not ( n330311 , n550 );
and ( n330312 , n330311 , n9391 );
or ( n330313 , n330310 , n330312 );
nand ( n10466 , n330313 , n8546 );
nand ( n330315 , n10461 , n10466 );
or ( n10468 , n551 , n552 );
nand ( n10469 , n10468 , n9758 );
nand ( n10470 , n551 , n552 );
and ( n10471 , n10469 , n10470 , n550 );
nand ( n10472 , n330315 , n10471 );
not ( n330321 , n10472 );
nand ( n330322 , n10451 , n330321 );
nand ( n10475 , n10448 , n330322 );
and ( n330324 , n330261 , n10475 );
and ( n10477 , n330225 , n330260 );
or ( n10478 , n330324 , n10477 );
buf ( n10479 , n10478 );
not ( n10480 , n10479 );
nor ( n330329 , n330215 , n10480 );
not ( n10482 , n330258 );
not ( n330331 , n10387 );
not ( n330332 , n330331 );
or ( n10485 , n10482 , n330332 );
not ( n330334 , n10387 );
not ( n10487 , n10411 );
or ( n330336 , n330334 , n10487 );
nand ( n10489 , n330336 , n330237 );
nand ( n10490 , n10485 , n10489 );
not ( n10491 , n10490 );
not ( n10492 , n10491 );
not ( n330341 , n8372 );
not ( n10494 , n10232 );
or ( n330343 , n330341 , n10494 );
nand ( n330344 , n328065 , n10401 );
nand ( n330345 , n330343 , n330344 );
not ( n10498 , n330345 );
not ( n330347 , n10498 );
not ( n10500 , n10300 );
not ( n10501 , n8675 );
and ( n330350 , n10500 , n10501 );
not ( n330351 , n554 );
not ( n330352 , n328032 );
or ( n10505 , n330351 , n330352 );
nand ( n330354 , n328033 , n8211 );
nand ( n330355 , n10505 , n330354 );
and ( n10508 , n330355 , n8570 );
nor ( n330357 , n330350 , n10508 );
not ( n330358 , n330233 );
not ( n10511 , n328669 );
and ( n330360 , n330358 , n10511 );
and ( n330361 , n10178 , n8485 );
nor ( n10514 , n330360 , n330361 );
xor ( n330363 , n330357 , n10514 );
not ( n10516 , n330363 );
not ( n330365 , n10516 );
or ( n10518 , n330347 , n330365 );
not ( n10519 , n10498 );
nand ( n330368 , n10519 , n330363 );
nand ( n330369 , n10518 , n330368 );
not ( n330370 , n330369 );
not ( n10523 , n330370 );
or ( n330372 , n10492 , n10523 );
nand ( n330373 , n330369 , n10490 );
nand ( n10526 , n330372 , n330373 );
not ( n330375 , n8570 );
not ( n330376 , n330291 );
or ( n10529 , n330375 , n330376 );
and ( n330378 , n328032 , n554 );
not ( n330379 , n328032 );
and ( n10532 , n330379 , n8211 );
or ( n330381 , n330378 , n10532 );
nand ( n330382 , n330381 , n328455 );
nand ( n10535 , n10529 , n330382 );
not ( n330384 , n10535 );
not ( n330385 , n330384 );
not ( n10538 , n328940 );
not ( n10539 , n330189 );
or ( n10540 , n10538 , n10539 );
nand ( n330389 , n330274 , n328847 );
nand ( n330390 , n10540 , n330389 );
not ( n330391 , n330390 );
not ( n10544 , n330391 );
or ( n330393 , n330385 , n10544 );
not ( n330394 , n8564 );
not ( n10547 , n10408 );
or ( n330396 , n330394 , n10547 );
not ( n330397 , n552 );
not ( n10550 , n329801 );
or ( n330399 , n330397 , n10550 );
nand ( n330400 , n329805 , n8324 );
nand ( n10553 , n330399 , n330400 );
nand ( n330402 , n10553 , n9329 );
nand ( n330403 , n330396 , n330402 );
not ( n10556 , n330403 );
and ( n10557 , n9391 , n8423 );
not ( n10558 , n10557 );
not ( n10559 , n330307 );
not ( n330408 , n10559 );
not ( n330409 , n328669 );
and ( n10562 , n330408 , n330409 );
not ( n10563 , n330226 );
and ( n330412 , n10563 , n9344 );
nor ( n10565 , n10562 , n330412 );
nand ( n330414 , n10558 , n10565 );
not ( n10567 , n330414 );
or ( n10568 , n10556 , n10567 );
not ( n10569 , n10565 );
nand ( n10570 , n10569 , n10557 );
nand ( n10571 , n10568 , n10570 );
nand ( n330420 , n330393 , n10571 );
nand ( n10573 , n330390 , n10535 );
nand ( n10574 , n330420 , n10573 );
buf ( n10575 , n10574 );
and ( n10576 , n10526 , n10575 );
not ( n330425 , n10526 );
not ( n330426 , n10574 );
and ( n10579 , n330425 , n330426 );
nor ( n330428 , n10576 , n10579 );
or ( n10581 , n330329 , n330428 );
nand ( n330430 , n330215 , n10480 );
nand ( n10583 , n10581 , n330430 );
not ( n10584 , n328455 );
not ( n330433 , n329995 );
or ( n330434 , n10584 , n330433 );
not ( n330435 , n10300 );
nand ( n10588 , n330435 , n8712 );
nand ( n330437 , n330434 , n10588 );
xor ( n330438 , n330437 , n10298 );
xnor ( n10591 , n330438 , n10317 );
not ( n330440 , n10591 );
not ( n330441 , n330440 );
not ( n10594 , n330369 );
not ( n330443 , n10491 );
and ( n330444 , n10594 , n330443 );
nand ( n330445 , n330369 , n10491 );
and ( n330446 , n330445 , n10574 );
nor ( n10599 , n330444 , n330446 );
not ( n330448 , n10599 );
not ( n330449 , n330448 );
or ( n10602 , n330441 , n330449 );
nand ( n330451 , n10599 , n10591 );
nand ( n330452 , n10602 , n330451 );
or ( n10605 , n330357 , n10514 );
and ( n10606 , n330357 , n10514 );
not ( n330455 , n10606 );
not ( n10608 , n10498 );
nand ( n10609 , n330455 , n10608 );
nand ( n330458 , n10605 , n10609 );
not ( n330459 , n330208 );
not ( n10612 , n330193 );
or ( n330461 , n330459 , n10612 );
not ( n10614 , n330208 );
not ( n10615 , n10614 );
not ( n330464 , n10346 );
or ( n10617 , n10615 , n330464 );
nand ( n330466 , n10617 , n10335 );
nand ( n10619 , n330461 , n330466 );
xor ( n330468 , n330458 , n10619 );
not ( n330469 , n10277 );
not ( n10622 , n330469 );
not ( n330471 , n8372 );
not ( n10624 , n9984 );
or ( n330473 , n330471 , n10624 );
nand ( n330474 , n10232 , n9329 );
nand ( n10627 , n330473 , n330474 );
not ( n330476 , n10627 );
not ( n10629 , n330476 );
or ( n10630 , n10622 , n10629 );
nand ( n330479 , n10627 , n10277 );
nand ( n330480 , n10630 , n330479 );
and ( n330481 , n330480 , n10225 );
not ( n10634 , n330480 );
not ( n330483 , n10225 );
and ( n330484 , n10634 , n330483 );
nor ( n10637 , n330481 , n330484 );
xor ( n330486 , n330468 , n10637 );
not ( n330487 , n330486 );
and ( n10640 , n330452 , n330487 );
not ( n330489 , n330452 );
and ( n330490 , n330489 , n330486 );
nor ( n330491 , n10640 , n330490 );
nand ( n10644 , n10583 , n330491 );
not ( n330493 , n10478 );
not ( n10646 , n10366 );
and ( n10647 , n330493 , n10646 );
and ( n330496 , n10478 , n10366 );
nor ( n330497 , n10647 , n330496 );
and ( n10650 , n10526 , n10575 );
not ( n330499 , n10526 );
and ( n330500 , n330499 , n330426 );
nor ( n10653 , n10650 , n330500 );
xor ( n330502 , n330497 , n10653 );
xor ( n330503 , n330225 , n330260 );
xor ( n10656 , n330503 , n10475 );
buf ( n330505 , n10656 );
not ( n330506 , n10571 );
not ( n10659 , n330384 );
or ( n330508 , n330506 , n10659 );
nand ( n10661 , n330403 , n330414 );
nand ( n330510 , n10661 , n10535 , n10570 );
nand ( n330511 , n330508 , n330510 );
and ( n10664 , n330511 , n330390 );
not ( n10665 , n330511 );
not ( n10666 , n330390 );
and ( n10667 , n10665 , n10666 );
nor ( n10668 , n10664 , n10667 );
not ( n330517 , n559 );
not ( n330518 , n10375 );
or ( n10671 , n330517 , n330518 );
not ( n330520 , n9461 );
not ( n330521 , n558 );
and ( n10674 , n330521 , n8401 );
not ( n10675 , n330521 );
and ( n10676 , n10675 , n328463 );
nor ( n10677 , n10674 , n10676 );
nand ( n330526 , n330520 , n10677 );
nand ( n330527 , n10671 , n330526 );
not ( n10680 , n330527 );
not ( n10681 , n10680 );
not ( n10682 , n10557 );
not ( n10683 , n10565 );
or ( n10684 , n10682 , n10683 );
not ( n330533 , n10557 );
nand ( n330534 , n330533 , n10569 );
nand ( n10687 , n10684 , n330534 );
not ( n10688 , n330403 );
and ( n10689 , n10687 , n10688 );
not ( n10690 , n10687 );
and ( n330539 , n10690 , n330403 );
nor ( n330540 , n10689 , n330539 );
not ( n330541 , n330540 );
or ( n10694 , n10681 , n330541 );
not ( n330543 , n328061 );
not ( n10696 , n10553 );
or ( n10697 , n330543 , n10696 );
and ( n330546 , n8983 , n8324 );
not ( n10699 , n8983 );
and ( n330548 , n10699 , n552 );
or ( n10701 , n330546 , n330548 );
nand ( n10702 , n10701 , n9329 );
nand ( n330551 , n10697 , n10702 );
not ( n10704 , n328940 );
not ( n330553 , n10417 );
or ( n330554 , n10704 , n330553 );
and ( n10707 , n556 , n8144 );
not ( n330556 , n556 );
and ( n330557 , n330556 , n328000 );
or ( n10710 , n10707 , n330557 );
nand ( n330559 , n10710 , n328847 );
nand ( n330560 , n330554 , n330559 );
or ( n10713 , n330551 , n330560 );
xor ( n330562 , n10471 , n330315 );
nand ( n10715 , n10713 , n330562 );
nand ( n10716 , n330560 , n330551 );
nand ( n10717 , n10715 , n10716 );
nand ( n10718 , n10694 , n10717 );
not ( n10719 , n330540 );
nand ( n330568 , n10719 , n330527 );
nand ( n330569 , n10718 , n330568 );
or ( n10722 , n10668 , n330569 );
and ( n330571 , n330505 , n10722 );
and ( n10724 , n10668 , n330569 );
nor ( n10725 , n330571 , n10724 );
nand ( n330574 , n330502 , n10725 );
and ( n330575 , n10644 , n330574 );
not ( n330576 , n330575 );
and ( n10729 , n558 , n328029 );
not ( n330578 , n558 );
and ( n330579 , n330578 , n8180 );
or ( n10732 , n10729 , n330579 );
and ( n330581 , n10732 , n559 );
not ( n330582 , n558 );
not ( n10735 , n8144 );
or ( n330584 , n330582 , n10735 );
nand ( n330585 , n328000 , n9056 );
nand ( n10738 , n330584 , n330585 );
not ( n330587 , n10738 );
nor ( n10740 , n330587 , n9461 );
nor ( n330589 , n330581 , n10740 );
not ( n10742 , n330589 );
not ( n10743 , n328455 );
not ( n330592 , n554 );
not ( n10745 , n9364 );
or ( n330594 , n330592 , n10745 );
nand ( n10747 , n9538 , n8211 );
nand ( n330596 , n330594 , n10747 );
not ( n330597 , n330596 );
or ( n10750 , n10743 , n330597 );
not ( n330599 , n554 );
not ( n330600 , n9776 );
or ( n10753 , n330599 , n330600 );
nand ( n330602 , n9758 , n8211 );
nand ( n330603 , n10753 , n330602 );
nor ( n10756 , n328415 , n328416 );
nand ( n330605 , n330603 , n10756 );
nand ( n330606 , n10750 , n330605 );
or ( n10759 , n555 , n556 );
nand ( n10760 , n10759 , n9391 );
nand ( n10761 , n555 , n556 );
and ( n10762 , n10760 , n10761 , n554 );
nand ( n10763 , n330606 , n10762 );
not ( n330612 , n10763 );
not ( n330613 , n330612 );
and ( n10766 , n9391 , n328061 );
not ( n330615 , n10766 );
not ( n330616 , n328455 );
not ( n10769 , n554 );
not ( n330618 , n10162 );
or ( n330619 , n10769 , n330618 );
nand ( n10772 , n8211 , n8982 );
nand ( n330621 , n330619 , n10772 );
not ( n330622 , n330621 );
or ( n10775 , n330616 , n330622 );
nand ( n330624 , n330596 , n8570 );
nand ( n10777 , n10775 , n330624 );
not ( n10778 , n10777 );
nand ( n10779 , n330615 , n10778 );
not ( n10780 , n10779 );
or ( n330629 , n330613 , n10780 );
nand ( n10782 , n10777 , n10766 );
nand ( n330631 , n330629 , n10782 );
not ( n330632 , n330631 );
and ( n10785 , n10742 , n330632 );
and ( n330634 , n330589 , n330631 );
nor ( n10787 , n10785 , n330634 );
not ( n10788 , n10787 );
not ( n10789 , n328940 );
not ( n10790 , n328839 );
not ( n10791 , n328054 );
or ( n10792 , n10790 , n10791 );
nand ( n10793 , n9573 , n556 );
nand ( n10794 , n10792 , n10793 );
not ( n10795 , n10794 );
or ( n10796 , n10789 , n10795 );
and ( n10797 , n556 , n8852 );
not ( n10798 , n556 );
and ( n10799 , n10798 , n8754 );
or ( n10800 , n10797 , n10799 );
nand ( n10801 , n10800 , n328847 );
nand ( n10802 , n10796 , n10801 );
not ( n10803 , n10802 );
not ( n10804 , n10803 );
not ( n10805 , n328455 );
not ( n10806 , n554 );
not ( n10807 , n329801 );
or ( n10808 , n10806 , n10807 );
not ( n10809 , n554 );
nand ( n10810 , n10809 , n8742 );
nand ( n10811 , n10808 , n10810 );
not ( n10812 , n10811 );
or ( n10813 , n10805 , n10812 );
not ( n10814 , n328525 );
nand ( n10815 , n10814 , n330621 );
nand ( n10816 , n10813 , n10815 );
not ( n10817 , n10816 );
not ( n10818 , n10817 );
not ( n10819 , n328061 );
not ( n330668 , n8324 );
not ( n10821 , n9364 );
not ( n330670 , n10821 );
or ( n10823 , n330668 , n330670 );
not ( n10824 , n9538 );
nand ( n10825 , n10824 , n552 );
nand ( n10826 , n10823 , n10825 );
not ( n10827 , n10826 );
or ( n10828 , n10819 , n10827 );
not ( n10829 , n575 );
not ( n10830 , n9385 );
or ( n10831 , n10829 , n10830 );
nand ( n330680 , n10831 , n9389 );
and ( n10833 , n330680 , n8324 );
not ( n10834 , n330680 );
and ( n330683 , n10834 , n552 );
nor ( n10836 , n10833 , n330683 );
not ( n330685 , n10836 );
nand ( n10838 , n330685 , n9329 );
nand ( n330687 , n10828 , n10838 );
or ( n330688 , n553 , n554 );
not ( n10841 , n330688 );
not ( n330690 , n9391 );
or ( n330691 , n10841 , n330690 );
nand ( n10844 , n553 , n554 );
and ( n10845 , n10844 , n552 );
nand ( n330694 , n330691 , n10845 );
not ( n10847 , n330694 );
and ( n10848 , n330687 , n10847 );
not ( n10849 , n330687 );
and ( n10850 , n10849 , n330694 );
nor ( n10851 , n10848 , n10850 );
not ( n330700 , n10851 );
and ( n10853 , n10818 , n330700 );
buf ( n330702 , n10851 );
not ( n10855 , n10816 );
and ( n10856 , n330702 , n10855 );
nor ( n10857 , n10853 , n10856 );
or ( n10858 , n10804 , n10857 );
not ( n330707 , n10851 );
nand ( n10860 , n330707 , n10816 );
nand ( n330709 , n330702 , n10855 );
nand ( n330710 , n10802 , n10860 , n330709 );
nand ( n10863 , n10858 , n330710 );
not ( n10864 , n10863 );
not ( n330713 , n10864 );
or ( n330714 , n10788 , n330713 );
not ( n10867 , n10787 );
nand ( n330716 , n10867 , n10863 );
nand ( n330717 , n330714 , n330716 );
not ( n10870 , n9673 );
not ( n330719 , n558 );
not ( n330720 , n328054 );
not ( n330721 , n330720 );
or ( n330722 , n330719 , n330721 );
not ( n10875 , n328612 );
nand ( n330724 , n10875 , n9056 );
nand ( n330725 , n330722 , n330724 );
not ( n10878 , n330725 );
or ( n330727 , n10870 , n10878 );
nand ( n330728 , n10738 , n559 );
nand ( n10881 , n330727 , n330728 );
not ( n330730 , n328940 );
not ( n330731 , n10800 );
or ( n10884 , n330730 , n330731 );
and ( n330733 , n556 , n329801 );
not ( n330734 , n556 );
and ( n10887 , n330734 , n329805 );
or ( n330736 , n330733 , n10887 );
nand ( n330737 , n330736 , n328847 );
nand ( n10890 , n10884 , n330737 );
or ( n330739 , n10881 , n10890 );
xor ( n330740 , n10766 , n10778 );
xnor ( n10893 , n330740 , n10763 );
not ( n330742 , n10893 );
and ( n330743 , n330739 , n330742 );
and ( n10896 , n10890 , n10881 );
nor ( n330745 , n330743 , n10896 );
nand ( n10898 , n330717 , n330745 );
not ( n330747 , n10898 );
xor ( n10900 , n10890 , n10881 );
and ( n10901 , n10900 , n10893 );
not ( n10902 , n10900 );
and ( n10903 , n10902 , n330742 );
nor ( n10904 , n10901 , n10903 );
xor ( n10905 , n556 , n329805 );
and ( n10906 , n10905 , n328940 );
xor ( n330755 , n556 , n8982 );
not ( n330756 , n330755 );
nor ( n10909 , n330756 , n8722 );
nor ( n330758 , n10906 , n10909 );
not ( n330759 , n10762 );
not ( n10912 , n330606 );
or ( n330761 , n330759 , n10912 );
or ( n330762 , n330606 , n10762 );
nand ( n330763 , n330761 , n330762 );
xor ( n10916 , n330758 , n330763 );
not ( n330765 , n8754 );
not ( n10918 , n9056 );
and ( n10919 , n330765 , n10918 );
and ( n330768 , n8754 , n9056 );
nor ( n330769 , n10919 , n330768 );
not ( n10922 , n330769 );
not ( n330771 , n9461 );
and ( n10924 , n10922 , n330771 );
and ( n10925 , n330725 , n559 );
nor ( n330774 , n10924 , n10925 );
and ( n330775 , n10916 , n330774 );
and ( n10928 , n330758 , n330763 );
or ( n330777 , n330775 , n10928 );
nand ( n330778 , n10904 , n330777 );
not ( n10931 , n330778 );
xor ( n330780 , n330758 , n330763 );
xor ( n330781 , n330780 , n330774 );
not ( n10934 , n330781 );
not ( n330783 , n10934 );
and ( n330784 , n9758 , n328455 );
not ( n10937 , n330784 );
not ( n330786 , n8718 );
not ( n330787 , n330755 );
or ( n10940 , n330786 , n330787 );
not ( n10941 , n8722 );
xor ( n330790 , n556 , n10821 );
nand ( n330791 , n10941 , n330790 );
nand ( n10944 , n10940 , n330791 );
not ( n10945 , n10944 );
and ( n330794 , n10937 , n10945 );
not ( n10947 , n8718 );
not ( n330796 , n330790 );
or ( n10949 , n10947 , n330796 );
not ( n10950 , n8722 );
and ( n10951 , n556 , n9391 );
not ( n10952 , n556 );
and ( n10953 , n10952 , n9776 );
nor ( n10954 , n10951 , n10953 );
nand ( n330803 , n10950 , n10954 );
nand ( n330804 , n10949 , n330803 );
or ( n10957 , n557 , n558 );
nand ( n330806 , n10957 , n9758 );
nand ( n330807 , n557 , n558 );
and ( n10960 , n330806 , n330807 , n556 );
nand ( n330809 , n330804 , n10960 );
nor ( n330810 , n330794 , n330809 );
and ( n10963 , n330784 , n10944 );
nor ( n10964 , n330810 , n10963 );
not ( n10965 , n10964 );
not ( n330814 , n10965 );
or ( n330815 , n330783 , n330814 );
xor ( n10968 , n330784 , n10944 );
xor ( n10969 , n10968 , n330809 );
not ( n10970 , n558 );
not ( n330819 , n329801 );
or ( n10972 , n10970 , n330819 );
nand ( n330821 , n329805 , n9056 );
nand ( n10974 , n10972 , n330821 );
not ( n10975 , n10974 );
not ( n330824 , n10975 );
not ( n330825 , n9461 );
and ( n10978 , n330824 , n330825 );
not ( n330827 , n330769 );
and ( n330828 , n330827 , n559 );
nor ( n10981 , n10978 , n330828 );
nand ( n330830 , n10969 , n10981 );
not ( n330831 , n559 );
and ( n330832 , n8982 , n9056 );
not ( n10985 , n8982 );
and ( n330834 , n10985 , n558 );
or ( n10987 , n330832 , n330834 );
not ( n330836 , n10987 );
or ( n10989 , n330831 , n330836 );
not ( n10990 , n558 );
not ( n10991 , n330302 );
or ( n330840 , n10990 , n10991 );
nand ( n330841 , n9538 , n9056 );
nand ( n10994 , n330840 , n330841 );
nand ( n10995 , n10994 , n329392 );
nand ( n10996 , n10989 , n10995 );
and ( n330845 , n9758 , n328940 );
nor ( n330846 , n10996 , n330845 );
not ( n330847 , n9758 );
nand ( n11000 , n330847 , n9462 );
not ( n330849 , n11000 );
nand ( n11002 , n10994 , n559 );
not ( n11003 , n11002 );
or ( n11004 , n330849 , n11003 );
nand ( n11005 , n9758 , n559 );
and ( n11006 , n11005 , n558 );
nand ( n11007 , n11004 , n11006 );
or ( n11008 , n330846 , n11007 );
nand ( n330857 , n10996 , n330845 );
nand ( n11010 , n11008 , n330857 );
not ( n330859 , n11010 );
not ( n11012 , n10987 );
not ( n11013 , n11012 );
not ( n11014 , n9461 );
and ( n11015 , n11013 , n11014 );
and ( n330864 , n10974 , n559 );
nor ( n330865 , n11015 , n330864 );
not ( n11018 , n10960 );
not ( n330867 , n330804 );
or ( n330868 , n11018 , n330867 );
or ( n11021 , n330804 , n10960 );
nand ( n330870 , n330868 , n11021 );
nand ( n330871 , n330865 , n330870 );
not ( n11024 , n330871 );
or ( n11025 , n330859 , n11024 );
or ( n11026 , n330865 , n330870 );
nand ( n330875 , n11025 , n11026 );
nand ( n330876 , n330830 , n330875 );
not ( n11029 , n330876 );
not ( n11030 , n10969 );
not ( n11031 , n10981 );
nand ( n330880 , n11030 , n11031 );
not ( n330881 , n330880 );
or ( n11034 , n11029 , n330881 );
nand ( n11035 , n330781 , n10964 );
nand ( n11036 , n11034 , n11035 );
nand ( n330885 , n330815 , n11036 );
not ( n330886 , n330885 );
or ( n11039 , n10931 , n330886 );
not ( n11040 , n10904 );
not ( n11041 , n330777 );
nand ( n330890 , n11040 , n11041 );
nand ( n330891 , n11039 , n330890 );
not ( n11044 , n330891 );
or ( n330893 , n330747 , n11044 );
not ( n330894 , n330717 );
not ( n11047 , n330745 );
nand ( n330896 , n330894 , n11047 );
nand ( n11049 , n330893 , n330896 );
not ( n330898 , n328847 );
not ( n11051 , n10794 );
or ( n330900 , n330898 , n11051 );
nand ( n11053 , n10710 , n328940 );
nand ( n330902 , n330900 , n11053 );
not ( n11055 , n330902 );
not ( n11056 , n9673 );
not ( n330905 , n10732 );
or ( n330906 , n11056 , n330905 );
not ( n11059 , n9056 );
not ( n330908 , n8411 );
or ( n330909 , n11059 , n330908 );
nor ( n11062 , n328539 , n9056 );
nor ( n330911 , n11062 , n1768 );
nand ( n330912 , n330909 , n330911 );
nand ( n11065 , n330906 , n330912 );
not ( n11066 , n11065 );
or ( n330915 , n11055 , n11066 );
or ( n11068 , n330902 , n11065 );
nand ( n330917 , n330687 , n10847 );
not ( n11070 , n330917 );
nand ( n11071 , n11068 , n11070 );
nand ( n330920 , n330915 , n11071 );
not ( n330921 , n330920 );
not ( n11074 , n330562 );
and ( n330923 , n11074 , n330551 );
not ( n330924 , n11074 );
not ( n11077 , n330551 );
and ( n330926 , n330924 , n11077 );
nor ( n330927 , n330923 , n330926 );
and ( n330928 , n330927 , n330560 );
not ( n11081 , n330927 );
not ( n330930 , n330560 );
and ( n330931 , n11081 , n330930 );
nor ( n11084 , n330928 , n330931 );
xor ( n330933 , n330921 , n11084 );
not ( n330934 , n10436 );
not ( n330935 , n8675 );
and ( n11088 , n330934 , n330935 );
not ( n330937 , n554 );
not ( n11090 , n8852 );
or ( n11091 , n330937 , n11090 );
not ( n330940 , n554 );
nand ( n11093 , n330940 , n8754 );
nand ( n330942 , n11091 , n11093 );
buf ( n11095 , n330942 );
and ( n330944 , n11095 , n8712 );
nor ( n330945 , n11088 , n330944 );
not ( n11098 , n330945 );
and ( n11099 , n9391 , n9344 );
not ( n330948 , n11099 );
not ( n11101 , n328065 );
not ( n330950 , n10826 );
or ( n330951 , n11101 , n330950 );
nand ( n330952 , n10701 , n8372 );
nand ( n11105 , n330951 , n330952 );
not ( n330954 , n11105 );
or ( n330955 , n330948 , n330954 );
or ( n11108 , n11099 , n11105 );
not ( n330957 , n328455 );
not ( n330958 , n330942 );
or ( n330959 , n330957 , n330958 );
nand ( n11112 , n10811 , n8570 );
nand ( n330961 , n330959 , n11112 );
nand ( n330962 , n11108 , n330961 );
nand ( n11115 , n330955 , n330962 );
xor ( n330964 , n11098 , n11115 );
and ( n330965 , n10677 , n559 );
not ( n330966 , n9673 );
and ( n11119 , n558 , n328539 );
not ( n330968 , n558 );
and ( n11121 , n330968 , n10424 );
nor ( n11122 , n11119 , n11121 );
nor ( n330971 , n330966 , n11122 );
nor ( n11124 , n330965 , n330971 );
xor ( n330973 , n330964 , n11124 );
and ( n11126 , n330933 , n330973 );
not ( n11127 , n330933 );
not ( n330976 , n330973 );
and ( n330977 , n11127 , n330976 );
nor ( n11130 , n11126 , n330977 );
and ( n330979 , n9391 , n8485 );
xor ( n330980 , n330979 , n11105 );
xnor ( n11133 , n330980 , n330961 );
not ( n330982 , n10803 );
not ( n330983 , n10855 );
and ( n330984 , n330982 , n330983 );
not ( n11137 , n10802 );
nand ( n330986 , n11137 , n10855 );
and ( n330987 , n330986 , n330702 );
nor ( n11140 , n330984 , n330987 );
xor ( n330989 , n11133 , n11140 );
not ( n330990 , n328847 );
not ( n11143 , n10794 );
or ( n11144 , n330990 , n11143 );
nand ( n330993 , n11144 , n11053 );
xor ( n330994 , n330917 , n330993 );
xor ( n11147 , n330994 , n11065 );
and ( n11148 , n330989 , n11147 );
and ( n11149 , n11133 , n11140 );
or ( n330998 , n11148 , n11149 );
nand ( n330999 , n11130 , n330998 );
xor ( n331000 , n11133 , n11140 );
xor ( n11153 , n331000 , n11147 );
buf ( n331002 , n330589 );
not ( n11155 , n331002 );
not ( n11156 , n330631 );
not ( n331005 , n11156 );
and ( n11158 , n11155 , n331005 );
buf ( n331007 , n10863 );
nand ( n11160 , n11156 , n331002 );
and ( n11161 , n331007 , n11160 );
nor ( n331010 , n11158 , n11161 );
nand ( n331011 , n11153 , n331010 );
nand ( n11164 , n11049 , n330999 , n331011 );
nor ( n331013 , n11153 , n331010 );
nand ( n331014 , n330999 , n331013 );
not ( n11167 , n11130 );
not ( n331016 , n330998 );
nand ( n331017 , n11167 , n331016 );
nand ( n331018 , n11164 , n331014 , n331017 );
not ( n11171 , n330945 );
not ( n331020 , n11124 );
or ( n331021 , n11171 , n331020 );
nand ( n11174 , n331021 , n11115 );
or ( n331023 , n11124 , n330945 );
nand ( n331024 , n11174 , n331023 );
xor ( n11177 , n10472 , n330277 );
xnor ( n331026 , n11177 , n330294 );
or ( n11179 , n331024 , n331026 );
not ( n331028 , n330540 );
not ( n11181 , n331028 );
not ( n11182 , n10680 );
or ( n331031 , n11181 , n11182 );
nand ( n331032 , n330527 , n330540 );
nand ( n11185 , n331031 , n331032 );
and ( n11186 , n11185 , n10717 );
not ( n331035 , n11185 );
not ( n331036 , n10717 );
and ( n331037 , n331035 , n331036 );
nor ( n11190 , n11186 , n331037 );
and ( n331039 , n11179 , n11190 );
and ( n11192 , n331024 , n331026 );
nor ( n11193 , n331039 , n11192 );
xor ( n331042 , n10668 , n330569 );
not ( n11195 , n10656 );
and ( n331044 , n331042 , n11195 );
not ( n11197 , n331042 );
and ( n11198 , n11197 , n10656 );
nor ( n331047 , n331044 , n11198 );
nand ( n331048 , n11193 , n331047 );
xor ( n11201 , n331024 , n331026 );
not ( n331050 , n11190 );
and ( n331051 , n11201 , n331050 );
not ( n11204 , n11201 );
and ( n331053 , n11204 , n11190 );
nor ( n331054 , n331051 , n331053 );
not ( n331055 , n330921 );
buf ( n11208 , n11084 );
not ( n331057 , n11208 );
and ( n331058 , n331055 , n331057 );
nand ( n11211 , n330921 , n11208 );
and ( n331060 , n330976 , n11211 );
nor ( n331061 , n331058 , n331060 );
nand ( n11214 , n331054 , n331061 );
nand ( n331063 , n331018 , n331048 , n11214 );
nor ( n331064 , n331061 , n331054 );
and ( n11217 , n331048 , n331064 );
nor ( n331066 , n331047 , n11193 );
nor ( n331067 , n11217 , n331066 );
nand ( n11220 , n331063 , n331067 );
not ( n331069 , n11220 );
or ( n331070 , n330576 , n331069 );
not ( n11223 , n10644 );
nor ( n11224 , n330502 , n10725 );
not ( n11225 , n11224 );
or ( n11226 , n11223 , n11225 );
not ( n331075 , n330491 );
not ( n331076 , n10583 );
nand ( n11229 , n331075 , n331076 );
nand ( n331078 , n11226 , n11229 );
not ( n11231 , n331078 );
nand ( n11232 , n331070 , n11231 );
and ( n11233 , n10197 , n10324 );
not ( n331082 , n10197 );
and ( n331083 , n331082 , n10323 );
nor ( n11236 , n11233 , n331083 );
not ( n331085 , n10200 );
and ( n331086 , n11236 , n331085 );
not ( n11239 , n11236 );
and ( n331088 , n11239 , n10200 );
nor ( n11241 , n331086 , n331088 );
xor ( n11242 , n330458 , n10619 );
and ( n331091 , n11242 , n10637 );
and ( n331092 , n330458 , n10619 );
or ( n331093 , n331091 , n331092 );
not ( n11246 , n330004 );
not ( n11247 , n10195 );
and ( n331096 , n11246 , n11247 );
and ( n331097 , n10195 , n330004 );
nor ( n11250 , n331096 , n331097 );
buf ( n11251 , n10152 );
and ( n331100 , n11250 , n11251 );
not ( n11253 , n11250 );
and ( n331102 , n11253 , n330001 );
nor ( n331103 , n331100 , n331102 );
or ( n331104 , n331093 , n331103 );
and ( n11257 , n10320 , n10280 );
not ( n331106 , n10320 );
and ( n11259 , n331106 , n10281 );
nor ( n331108 , n11257 , n11259 );
not ( n331109 , n10211 );
and ( n331110 , n331108 , n331109 );
not ( n331111 , n331108 );
not ( n11264 , n331109 );
and ( n331113 , n331111 , n11264 );
nor ( n11266 , n331110 , n331113 );
and ( n331115 , n331104 , n11266 );
and ( n331116 , n331093 , n331103 );
nor ( n11269 , n331115 , n331116 );
nand ( n331118 , n11241 , n11269 );
not ( n331119 , n331118 );
xor ( n11272 , n331093 , n331103 );
xor ( n11273 , n11272 , n11266 );
not ( n331122 , n330448 );
not ( n331123 , n331122 );
not ( n11276 , n330440 );
or ( n331125 , n331123 , n11276 );
nand ( n11278 , n331125 , n330486 );
nand ( n331127 , n330448 , n10591 );
nand ( n11280 , n11278 , n331127 );
nor ( n11281 , n11273 , n11280 );
nor ( n11282 , n331119 , n11281 );
nand ( n331131 , n10332 , n11232 , n11282 );
nor ( n11284 , n329987 , n10329 );
nand ( n331133 , n10135 , n10132 );
and ( n331134 , n11284 , n331133 );
buf ( n11287 , n10135 );
buf ( n331136 , n10132 );
nor ( n11288 , n11287 , n331136 );
nor ( n331138 , n331134 , n11288 );
not ( n331139 , n331118 );
nand ( n11291 , n11273 , n11280 );
not ( n11292 , n11291 );
not ( n11293 , n11292 );
or ( n331143 , n331139 , n11293 );
not ( n331144 , n11269 );
not ( n11296 , n11241 );
nand ( n11297 , n331144 , n11296 );
nand ( n11298 , n331143 , n11297 );
nand ( n331148 , n11298 , n331133 , n10330 );
nand ( n331149 , n331131 , n331138 , n331148 );
not ( n11301 , n331149 );
or ( n331151 , n10086 , n11301 );
not ( n331152 , n9869 );
not ( n11304 , n9915 );
or ( n331154 , n331152 , n11304 );
not ( n11306 , n329716 );
not ( n331156 , n329762 );
or ( n11308 , n11306 , n331156 );
nand ( n331158 , n9919 , n10054 );
nand ( n11310 , n11308 , n331158 );
nand ( n11311 , n331154 , n11310 );
not ( n331161 , n11311 );
not ( n331162 , n329923 );
not ( n11314 , n10071 );
nand ( n331164 , n331162 , n11314 );
not ( n331165 , n329926 );
not ( n11317 , n329930 );
nand ( n331167 , n331165 , n11317 );
nand ( n331168 , n331164 , n331167 );
or ( n11320 , n331161 , n331168 );
nand ( n11321 , n10084 , n331167 );
nand ( n331171 , n11320 , n11321 );
nand ( n11323 , n331151 , n331171 );
not ( n331173 , n11323 );
or ( n11325 , n9285 , n331173 );
not ( n11326 , n9283 );
nor ( n331176 , n9027 , n329031 );
not ( n331177 , n331176 );
or ( n11329 , n11326 , n331177 );
or ( n331179 , n9278 , n329130 );
nand ( n331180 , n11329 , n331179 );
not ( n11332 , n331180 );
nand ( n331182 , n11325 , n11332 );
buf ( n331183 , n331182 );
xor ( n331184 , n9189 , n329060 );
and ( n11336 , n331184 , n9217 );
and ( n331186 , n9189 , n329060 );
or ( n331187 , n11336 , n331186 );
or ( n11339 , n9211 , n329051 );
not ( n331189 , n329042 );
nand ( n331190 , n11339 , n331189 );
nand ( n11342 , n9211 , n329051 );
nand ( n11343 , n331190 , n11342 );
not ( n11344 , n11343 );
not ( n331194 , n11344 );
and ( n331195 , n8826 , n8447 );
not ( n331196 , n8826 );
and ( n11348 , n331196 , n548 );
or ( n331198 , n331195 , n11348 );
not ( n331199 , n331198 );
not ( n11351 , n329668 );
or ( n11352 , n331199 , n11351 );
nand ( n331202 , n8475 , n329047 );
nand ( n11354 , n11352 , n331202 );
not ( n11355 , n11354 );
not ( n331205 , n329105 );
not ( n331206 , n329100 );
or ( n11358 , n331205 , n331206 );
not ( n11359 , n546 );
not ( n11360 , n328488 );
or ( n11361 , n11359 , n11360 );
not ( n331211 , n328488 );
nand ( n11363 , n331211 , n8378 );
nand ( n331213 , n11361 , n11363 );
nand ( n11365 , n331213 , n8376 );
nand ( n11366 , n11358 , n11365 );
not ( n331216 , n11366 );
or ( n331217 , n11355 , n331216 );
or ( n11369 , n11366 , n11354 );
nand ( n331219 , n331217 , n11369 );
not ( n331220 , n8686 );
not ( n11372 , n9207 );
or ( n331222 , n331220 , n11372 );
not ( n331223 , n329053 );
not ( n11375 , n331223 );
not ( n11376 , n328503 );
xor ( n11377 , n544 , n11376 );
nand ( n11378 , n11375 , n11377 );
nand ( n11379 , n331222 , n11378 );
and ( n331229 , n331219 , n11379 );
not ( n331230 , n331219 );
not ( n331231 , n11379 );
and ( n11383 , n331230 , n331231 );
nor ( n331233 , n331229 , n11383 );
not ( n11385 , n331233 );
or ( n11386 , n331194 , n11385 );
or ( n331236 , n11344 , n331233 );
nand ( n331237 , n11386 , n331236 );
not ( n11389 , n331237 );
not ( n331239 , n328062 );
not ( n331240 , n328064 );
or ( n11392 , n331239 , n331240 );
nand ( n331242 , n11392 , n552 );
buf ( n331243 , n328542 );
nand ( n11395 , n331243 , n544 );
and ( n11396 , n331242 , n11395 );
not ( n11397 , n331242 );
not ( n331247 , n11395 );
and ( n331248 , n11397 , n331247 );
nor ( n11400 , n11396 , n331248 );
not ( n331250 , n11400 );
not ( n331251 , n9063 );
not ( n11403 , n9241 );
or ( n11404 , n331251 , n11403 );
not ( n11405 , n8514 );
buf ( n331255 , n328452 );
not ( n331256 , n331255 );
or ( n11408 , n11405 , n331256 );
not ( n11409 , n331255 );
not ( n11410 , n8514 );
and ( n11411 , n11409 , n11410 );
not ( n11412 , n8485 );
nor ( n331262 , n11411 , n11412 );
nand ( n331263 , n11408 , n331262 );
nand ( n11415 , n11404 , n331263 );
not ( n11416 , n11415 );
or ( n331266 , n331250 , n11416 );
or ( n331267 , n11415 , n11400 );
nand ( n11419 , n331266 , n331267 );
xor ( n331269 , n329042 , n11419 );
and ( n11421 , n9236 , n9246 );
or ( n331271 , n11421 , n329107 );
or ( n11423 , n9246 , n9236 );
nand ( n11424 , n331271 , n11423 );
xor ( n331274 , n331269 , n11424 );
not ( n331275 , n331274 );
and ( n11427 , n11389 , n331275 );
and ( n331277 , n331274 , n331237 );
nor ( n331278 , n11427 , n331277 );
xor ( n11430 , n331187 , n331278 );
not ( n331280 , n9233 );
not ( n331281 , n331280 );
not ( n11433 , n9260 );
and ( n331283 , n331281 , n11433 );
not ( n331284 , n9225 );
nand ( n11436 , n331280 , n9260 );
and ( n331286 , n331284 , n11436 );
nor ( n331287 , n331283 , n331286 );
xor ( n331288 , n11430 , n331287 );
not ( n11440 , n331288 );
xor ( n331290 , n329066 , n329116 );
and ( n11442 , n331290 , n329125 );
and ( n11443 , n329066 , n329116 );
or ( n331293 , n11442 , n11443 );
not ( n11445 , n331293 );
nand ( n331295 , n11440 , n11445 );
buf ( n11447 , n331295 );
nand ( n11448 , n331288 , n331293 );
buf ( n331298 , n11448 );
nand ( n331299 , n11447 , n331298 );
not ( n11451 , n331299 );
and ( n331301 , n331183 , n11451 );
not ( n331302 , n331183 );
and ( n11454 , n331302 , n331299 );
nor ( n331304 , n331301 , n11454 );
nor ( n331305 , n8099 , n331304 );
not ( n331306 , n331305 );
buf ( n331307 , n7565 );
buf ( n331308 , n8090 );
and ( n331309 , n331307 , n331308 );
buf ( n331310 , n331309 );
not ( n331311 , n331310 );
not ( n331312 , n327628 );
not ( n11464 , n2971 );
not ( n11465 , n4617 );
or ( n331315 , n11464 , n11465 );
nand ( n331316 , n331315 , n4651 );
not ( n11468 , n331316 );
or ( n331318 , n331312 , n11468 );
buf ( n331319 , n7835 );
not ( n331320 , n331319 );
buf ( n331321 , n331320 );
nand ( n11473 , n331318 , n331321 );
not ( n331323 , n11473 );
or ( n11475 , n331311 , n331323 );
buf ( n331325 , n7817 );
buf ( n331326 , n8090 );
and ( n11478 , n331325 , n331326 );
not ( n331328 , n8092 );
buf ( n331329 , n331328 );
nor ( n11481 , n11478 , n331329 );
buf ( n11482 , n11481 );
nand ( n331332 , n11475 , n11482 );
xor ( n11484 , n7952 , n327924 );
and ( n331334 , n11484 , n327931 );
and ( n331335 , n7952 , n327924 );
or ( n331336 , n331334 , n331335 );
buf ( n331337 , n331336 );
not ( n331338 , n331337 );
xor ( n331339 , n327911 , n327916 );
and ( n11491 , n331339 , n327922 );
and ( n331341 , n327911 , n327916 );
or ( n331342 , n11491 , n331341 );
not ( n11494 , n331342 );
xor ( n11495 , n327698 , n327790 );
and ( n331345 , n11495 , n327797 );
and ( n331346 , n327698 , n327790 );
or ( n11498 , n331345 , n331346 );
buf ( n331348 , n11498 );
buf ( n331349 , n331348 );
not ( n331350 , n331349 );
buf ( n331351 , n331350 );
nand ( n331352 , n11494 , n331351 );
not ( n11504 , n331352 );
nand ( n331354 , n331342 , n331348 );
not ( n11506 , n331354 );
or ( n11507 , n11504 , n11506 );
xor ( n331357 , n327869 , n8041 );
and ( n11509 , n331357 , n327896 );
and ( n331359 , n327869 , n8041 );
or ( n11511 , n11509 , n331359 );
buf ( n331361 , n11511 );
buf ( n11513 , n331361 );
buf ( n331363 , n550 );
buf ( n331364 , n576 );
and ( n331365 , n331363 , n331364 );
buf ( n331366 , n331365 );
buf ( n331367 , n331366 );
buf ( n331368 , n8014 );
not ( n331369 , n331368 );
buf ( n331370 , n3865 );
not ( n11522 , n331370 );
or ( n331372 , n331369 , n11522 );
buf ( n331373 , n323715 );
buf ( n331374 , n546 );
buf ( n331375 , n578 );
xor ( n331376 , n331374 , n331375 );
buf ( n331377 , n331376 );
buf ( n331378 , n331377 );
nand ( n11530 , n331373 , n331378 );
buf ( n331380 , n11530 );
buf ( n331381 , n331380 );
nand ( n11533 , n331372 , n331381 );
buf ( n331383 , n11533 );
buf ( n331384 , n331383 );
xor ( n11536 , n331367 , n331384 );
buf ( n331386 , n327885 );
xor ( n331387 , n11536 , n331386 );
buf ( n331388 , n331387 );
buf ( n11540 , n331388 );
xor ( n331390 , n327811 , n327828 );
and ( n11542 , n331390 , n327842 );
and ( n331392 , n327811 , n327828 );
or ( n331393 , n11542 , n331392 );
buf ( n331394 , n331393 );
buf ( n331395 , n331394 );
xor ( n331396 , n11540 , n331395 );
buf ( n331397 , n327821 );
not ( n11549 , n331397 );
buf ( n331399 , n325952 );
not ( n11551 , n331399 );
or ( n11552 , n11549 , n11551 );
buf ( n331402 , n5580 );
buf ( n331403 , n548 );
buf ( n331404 , n576 );
xor ( n331405 , n331403 , n331404 );
buf ( n331406 , n331405 );
buf ( n331407 , n331406 );
nand ( n11559 , n331402 , n331407 );
buf ( n331409 , n11559 );
buf ( n331410 , n331409 );
nand ( n331411 , n11552 , n331410 );
buf ( n331412 , n331411 );
buf ( n331413 , n331412 );
buf ( n331414 , n327879 );
not ( n331415 , n331414 );
buf ( n331416 , n5650 );
not ( n331417 , n331416 );
or ( n331418 , n331415 , n331417 );
buf ( n331419 , n322474 );
buf ( n331420 , n544 );
buf ( n331421 , n580 );
xor ( n11573 , n331420 , n331421 );
buf ( n331423 , n11573 );
buf ( n331424 , n331423 );
nand ( n11576 , n331419 , n331424 );
buf ( n331426 , n11576 );
buf ( n331427 , n331426 );
nand ( n331428 , n331418 , n331427 );
buf ( n331429 , n331428 );
buf ( n331430 , n331429 );
xor ( n331431 , n331413 , n331430 );
buf ( n331432 , n323755 );
buf ( n331433 , n323550 );
or ( n11585 , n331432 , n331433 );
buf ( n331435 , n582 );
nand ( n331436 , n11585 , n331435 );
buf ( n331437 , n331436 );
buf ( n331438 , n331437 );
xor ( n11590 , n331431 , n331438 );
buf ( n331440 , n11590 );
buf ( n331441 , n331440 );
xor ( n331442 , n331396 , n331441 );
buf ( n331443 , n331442 );
buf ( n331444 , n331443 );
xor ( n331445 , n11513 , n331444 );
xor ( n11597 , n327845 , n327851 );
and ( n331447 , n11597 , n327899 );
and ( n331448 , n327845 , n327851 );
or ( n11600 , n331447 , n331448 );
buf ( n331450 , n11600 );
buf ( n331451 , n331450 );
xor ( n331452 , n331445 , n331451 );
buf ( n331453 , n331452 );
buf ( n331454 , n331453 );
xor ( n11603 , n327806 , n327902 );
and ( n11604 , n11603 , n327909 );
and ( n11605 , n327806 , n327902 );
or ( n11606 , n11604 , n11605 );
buf ( n331459 , n11606 );
buf ( n331460 , n331459 );
xor ( n11608 , n331454 , n331460 );
xor ( n11609 , n327757 , n327777 );
and ( n331463 , n11609 , n327784 );
and ( n331464 , n327757 , n327777 );
or ( n331465 , n331463 , n331464 );
buf ( n331466 , n331465 );
buf ( n331467 , n331466 );
buf ( n331468 , n327737 );
buf ( n331469 , n327724 );
not ( n11614 , n331469 );
buf ( n331471 , n11614 );
buf ( n331472 , n331471 );
or ( n11617 , n331468 , n331472 );
buf ( n331474 , n7872 );
nand ( n331475 , n11617 , n331474 );
buf ( n331476 , n331475 );
buf ( n331477 , n331476 );
buf ( n331478 , n327737 );
buf ( n331479 , n331471 );
nand ( n331480 , n331478 , n331479 );
buf ( n331481 , n331480 );
buf ( n331482 , n331481 );
nand ( n11626 , n331477 , n331482 );
buf ( n331484 , n11626 );
buf ( n331485 , n331484 );
buf ( n331486 , n550 );
buf ( n331487 , n560 );
and ( n331488 , n331486 , n331487 );
buf ( n331489 , n331488 );
buf ( n331490 , n331489 );
buf ( n331491 , n327773 );
xor ( n11635 , n331490 , n331491 );
buf ( n331493 , n327750 );
not ( n11637 , n331493 );
buf ( n331495 , n3157 );
not ( n331496 , n331495 );
or ( n11640 , n11637 , n331496 );
buf ( n331498 , n323009 );
buf ( n331499 , n546 );
buf ( n331500 , n562 );
xor ( n331501 , n331499 , n331500 );
buf ( n331502 , n331501 );
buf ( n331503 , n331502 );
nand ( n11647 , n331498 , n331503 );
buf ( n331505 , n11647 );
buf ( n331506 , n331505 );
nand ( n11650 , n11640 , n331506 );
buf ( n331508 , n11650 );
buf ( n331509 , n331508 );
xor ( n331510 , n11635 , n331509 );
buf ( n331511 , n331510 );
buf ( n331512 , n331511 );
xor ( n11656 , n331485 , n331512 );
buf ( n331514 , n327714 );
not ( n11658 , n331514 );
buf ( n331516 , n7031 );
not ( n331517 , n331516 );
or ( n11661 , n11658 , n331517 );
buf ( n331519 , n324855 );
buf ( n331520 , n548 );
buf ( n331521 , n560 );
xor ( n331522 , n331520 , n331521 );
buf ( n331523 , n331522 );
buf ( n331524 , n331523 );
nand ( n331525 , n331519 , n331524 );
buf ( n331526 , n331525 );
buf ( n331527 , n331526 );
nand ( n331528 , n11661 , n331527 );
buf ( n331529 , n331528 );
buf ( n331530 , n331529 );
buf ( n331531 , n327767 );
not ( n331532 , n331531 );
buf ( n331533 , n321592 );
not ( n11677 , n331533 );
or ( n11678 , n331532 , n11677 );
buf ( n331536 , n3186 );
buf ( n331537 , n544 );
buf ( n331538 , n564 );
xor ( n331539 , n331537 , n331538 );
buf ( n331540 , n331539 );
buf ( n331541 , n331540 );
nand ( n11685 , n331536 , n331541 );
buf ( n331543 , n11685 );
buf ( n331544 , n331543 );
nand ( n11688 , n11678 , n331544 );
buf ( n331546 , n11688 );
buf ( n331547 , n331546 );
xor ( n11691 , n331530 , n331547 );
buf ( n11692 , n321771 );
not ( n331550 , n11692 );
buf ( n331551 , n331550 );
buf ( n331552 , n331551 );
not ( n331553 , n331552 );
buf ( n331554 , n322973 );
not ( n331555 , n331554 );
or ( n331556 , n331553 , n331555 );
buf ( n331557 , n566 );
nand ( n11701 , n331556 , n331557 );
buf ( n11702 , n11701 );
buf ( n331560 , n11702 );
xor ( n11704 , n11691 , n331560 );
buf ( n331562 , n11704 );
buf ( n331563 , n331562 );
xor ( n11707 , n11656 , n331563 );
buf ( n331565 , n11707 );
buf ( n331566 , n331565 );
xor ( n331567 , n331467 , n331566 );
xor ( n331568 , n327704 , n327739 );
and ( n11712 , n331568 , n327787 );
and ( n11713 , n327704 , n327739 );
or ( n11714 , n11712 , n11713 );
buf ( n11715 , n11714 );
buf ( n331573 , n11715 );
xor ( n11717 , n331567 , n331573 );
buf ( n331575 , n11717 );
buf ( n331576 , n331575 );
xor ( n11720 , n11608 , n331576 );
buf ( n331578 , n11720 );
nand ( n11722 , n11507 , n331578 );
not ( n11723 , n331342 );
not ( n11724 , n331348 );
and ( n331582 , n11723 , n11724 );
nor ( n331583 , n331582 , n331578 );
nand ( n331584 , n331583 , n331354 );
nand ( n11728 , n331338 , n11722 , n331584 );
not ( n331586 , n11722 );
not ( n11730 , n331584 );
or ( n11731 , n331586 , n11730 );
nand ( n331589 , n11731 , n331337 );
and ( n11733 , n11728 , n331589 );
xor ( n331591 , n331332 , n11733 );
not ( n11735 , n331591 );
not ( n11736 , n11447 );
nand ( n331594 , n331182 , n331298 );
not ( n331595 , n331594 );
or ( n11739 , n11736 , n331595 );
not ( n331597 , n8517 );
xor ( n331598 , n331597 , n8378 );
not ( n11742 , n331598 );
not ( n331600 , n8783 );
and ( n331601 , n11742 , n331600 );
and ( n331602 , n331213 , n329105 );
nor ( n11746 , n331601 , n331602 );
not ( n331604 , n9063 );
and ( n331605 , n550 , n331255 );
not ( n11749 , n331605 );
or ( n331607 , n331604 , n11749 );
not ( n331608 , n331255 );
and ( n331609 , n8514 , n9063 , n331608 );
and ( n11753 , n8485 , n550 );
nor ( n331611 , n331609 , n11753 );
nand ( n11755 , n331607 , n331611 );
and ( n11756 , n11746 , n11755 );
not ( n331614 , n11746 );
not ( n11758 , n11755 );
and ( n11759 , n331614 , n11758 );
nor ( n331617 , n11756 , n11759 );
not ( n11761 , n331231 );
not ( n11762 , n11354 );
not ( n331620 , n11762 );
and ( n11764 , n11761 , n331620 );
nand ( n331622 , n331231 , n11762 );
buf ( n11766 , n11366 );
and ( n331624 , n331622 , n11766 );
nor ( n331625 , n11764 , n331624 );
not ( n11769 , n331625 );
and ( n331627 , n331617 , n11769 );
not ( n331628 , n331617 );
and ( n331629 , n331628 , n331625 );
nor ( n11773 , n331627 , n331629 );
not ( n331631 , n331242 );
not ( n331632 , n331247 );
or ( n11776 , n331631 , n331632 );
not ( n331634 , n331242 );
nand ( n331635 , n331634 , n11395 );
nand ( n11779 , n11415 , n331635 );
nand ( n11780 , n11776 , n11779 );
not ( n11781 , n11780 );
not ( n331639 , n11781 );
and ( n331640 , n328463 , n544 );
not ( n11784 , n8475 );
not ( n11785 , n331198 );
or ( n11786 , n11784 , n11785 );
not ( n331644 , n548 );
buf ( n331645 , n328423 );
not ( n11789 , n331645 );
not ( n11790 , n11789 );
or ( n331648 , n331644 , n11790 );
nand ( n331649 , n331645 , n8447 );
nand ( n11793 , n331648 , n331649 );
nand ( n331651 , n11793 , n329668 );
nand ( n11795 , n11786 , n331651 );
xor ( n331653 , n331640 , n11795 );
not ( n11797 , n8686 );
not ( n11798 , n11377 );
or ( n11799 , n11797 , n11798 );
not ( n11800 , n544 );
not ( n11801 , n9248 );
or ( n11802 , n11800 , n11801 );
not ( n11803 , n9248 );
nand ( n11804 , n11803 , n328001 );
nand ( n331662 , n11802 , n11804 );
nand ( n331663 , n331662 , n329053 );
nand ( n11807 , n11799 , n331663 );
xnor ( n331665 , n331653 , n11807 );
not ( n331666 , n331665 );
not ( n11810 , n331666 );
or ( n331668 , n331639 , n11810 );
nand ( n331669 , n11780 , n331665 );
nand ( n11813 , n331668 , n331669 );
xor ( n11814 , n329042 , n11419 );
and ( n11815 , n11814 , n11424 );
and ( n331673 , n329042 , n11419 );
or ( n331674 , n11815 , n331673 );
xor ( n11818 , n11813 , n331674 );
xor ( n331676 , n11773 , n11818 );
not ( n11820 , n331274 );
not ( n11821 , n331233 );
not ( n331679 , n11821 );
nand ( n11823 , n331679 , n11344 );
not ( n331681 , n11823 );
or ( n11825 , n11820 , n331681 );
nand ( n331683 , n11821 , n11343 );
nand ( n11827 , n11825 , n331683 );
xnor ( n11828 , n331676 , n11827 );
not ( n331686 , n11828 );
xor ( n331687 , n331187 , n331278 );
and ( n11831 , n331687 , n331287 );
and ( n331689 , n331187 , n331278 );
or ( n331690 , n11831 , n331689 );
not ( n11834 , n331690 );
nand ( n331692 , n331686 , n11834 );
nand ( n331693 , n11828 , n331690 );
buf ( n11837 , n331693 );
nand ( n11838 , n331692 , n11837 );
nand ( n331696 , n11739 , n11838 );
not ( n11840 , n11447 );
nor ( n331698 , n11840 , n11838 );
nand ( n11842 , n331594 , n331698 );
nand ( n11843 , n331696 , n11842 );
nand ( n331701 , n11735 , n11843 );
not ( n331702 , n331701 );
or ( n11846 , n331306 , n331702 );
not ( n331704 , n11843 );
buf ( n331705 , n331591 );
nand ( n11849 , n331704 , n331705 );
nand ( n331707 , n11846 , n11849 );
not ( n331708 , n331707 );
buf ( n331709 , n11728 );
buf ( n331710 , n8090 );
nand ( n331711 , n331709 , n331710 );
buf ( n331712 , n331711 );
buf ( n331713 , n331712 );
buf ( n331714 , n331578 );
not ( n331715 , n331714 );
buf ( n331716 , n331715 );
buf ( n331717 , n331716 );
buf ( n331718 , n331351 );
nand ( n331719 , n331717 , n331718 );
buf ( n331720 , n331719 );
not ( n11864 , n331720 );
not ( n11865 , n331342 );
or ( n331723 , n11864 , n11865 );
or ( n331724 , n331716 , n331351 );
nand ( n331725 , n331723 , n331724 );
buf ( n331726 , n331725 );
xor ( n331727 , n331467 , n331566 );
and ( n11871 , n331727 , n331573 );
and ( n11872 , n331467 , n331566 );
or ( n331730 , n11871 , n11872 );
buf ( n331731 , n331730 );
not ( n331732 , n331731 );
xor ( n11876 , n331454 , n331460 );
and ( n11877 , n11876 , n331576 );
and ( n11878 , n331454 , n331460 );
or ( n11879 , n11877 , n11878 );
buf ( n331737 , n11879 );
xor ( n11881 , n331732 , n331737 );
xor ( n331739 , n331490 , n331491 );
and ( n331740 , n331739 , n331509 );
and ( n331741 , n331490 , n331491 );
or ( n11885 , n331740 , n331741 );
buf ( n331743 , n11885 );
buf ( n331744 , n331743 );
buf ( n331745 , n331540 );
not ( n331746 , n331745 );
buf ( n331747 , n321592 );
not ( n11891 , n331747 );
or ( n331749 , n331746 , n11891 );
buf ( n331750 , n3186 );
buf ( n331751 , n564 );
nand ( n11895 , n331750 , n331751 );
buf ( n331753 , n11895 );
buf ( n11897 , n331753 );
nand ( n331755 , n331749 , n11897 );
buf ( n331756 , n331755 );
buf ( n331757 , n331756 );
not ( n331758 , n331757 );
buf ( n331759 , n331758 );
buf ( n11903 , n331759 );
buf ( n331761 , n549 );
buf ( n331762 , n560 );
and ( n331763 , n331761 , n331762 );
buf ( n331764 , n331763 );
buf ( n331765 , n331764 );
not ( n331766 , n324728 );
not ( n11910 , n331523 );
or ( n11911 , n331766 , n11910 );
buf ( n11912 , n324855 );
buf ( n331770 , n560 );
buf ( n331771 , n547 );
xor ( n331772 , n331770 , n331771 );
buf ( n331773 , n331772 );
buf ( n331774 , n331773 );
nand ( n11918 , n11912 , n331774 );
buf ( n331776 , n11918 );
nand ( n331777 , n11911 , n331776 );
buf ( n11921 , n331777 );
xor ( n11922 , n331765 , n11921 );
buf ( n331780 , n331502 );
not ( n331781 , n331780 );
buf ( n331782 , n3157 );
not ( n331783 , n331782 );
or ( n331784 , n331781 , n331783 );
buf ( n331785 , n323009 );
buf ( n331786 , n545 );
buf ( n331787 , n562 );
xor ( n331788 , n331786 , n331787 );
buf ( n331789 , n331788 );
buf ( n331790 , n331789 );
nand ( n331791 , n331785 , n331790 );
buf ( n331792 , n331791 );
buf ( n331793 , n331792 );
nand ( n331794 , n331784 , n331793 );
buf ( n331795 , n331794 );
buf ( n331796 , n331795 );
xor ( n331797 , n11922 , n331796 );
buf ( n331798 , n331797 );
buf ( n331799 , n331798 );
xor ( n331800 , n11903 , n331799 );
xor ( n11944 , n331530 , n331547 );
and ( n331802 , n11944 , n331560 );
and ( n331803 , n331530 , n331547 );
or ( n331804 , n331802 , n331803 );
buf ( n331805 , n331804 );
buf ( n331806 , n331805 );
xor ( n331807 , n331800 , n331806 );
buf ( n331808 , n331807 );
buf ( n331809 , n331808 );
xor ( n331810 , n331744 , n331809 );
xor ( n331811 , n331485 , n331512 );
and ( n11955 , n331811 , n331563 );
and ( n11956 , n331485 , n331512 );
or ( n11957 , n11955 , n11956 );
buf ( n331815 , n11957 );
buf ( n331816 , n331815 );
xor ( n11960 , n331810 , n331816 );
buf ( n331818 , n11960 );
buf ( n331819 , n331818 );
xor ( n11963 , n11513 , n331444 );
and ( n331821 , n11963 , n331451 );
and ( n11965 , n11513 , n331444 );
or ( n331823 , n331821 , n11965 );
buf ( n331824 , n331823 );
buf ( n331825 , n331824 );
xor ( n331826 , n331819 , n331825 );
xor ( n11969 , n331367 , n331384 );
and ( n331828 , n11969 , n331386 );
and ( n11971 , n331367 , n331384 );
or ( n331830 , n331828 , n11971 );
buf ( n331831 , n331830 );
buf ( n331832 , n331831 );
xor ( n11975 , n11540 , n331395 );
and ( n11976 , n11975 , n331441 );
and ( n331835 , n11540 , n331395 );
or ( n11978 , n11976 , n331835 );
buf ( n331837 , n11978 );
buf ( n331838 , n331837 );
xor ( n11981 , n331832 , n331838 );
buf ( n331840 , n331423 );
not ( n11983 , n331840 );
buf ( n331842 , n5650 );
not ( n331843 , n331842 );
or ( n11986 , n11983 , n331843 );
buf ( n331845 , n322474 );
buf ( n331846 , n580 );
nand ( n331847 , n331845 , n331846 );
buf ( n331848 , n331847 );
buf ( n331849 , n331848 );
nand ( n11992 , n11986 , n331849 );
buf ( n331851 , n11992 );
buf ( n331852 , n331851 );
not ( n331853 , n331852 );
buf ( n331854 , n331853 );
buf ( n331855 , n331854 );
buf ( n331856 , n549 );
buf ( n11999 , n576 );
and ( n12000 , n331856 , n11999 );
buf ( n331859 , n12000 );
buf ( n12002 , n331859 );
buf ( n331861 , n331406 );
not ( n12004 , n331861 );
buf ( n331863 , n325952 );
not ( n331864 , n331863 );
or ( n12007 , n12004 , n331864 );
buf ( n331866 , n5580 );
buf ( n331867 , n576 );
buf ( n331868 , n547 );
xor ( n331869 , n331867 , n331868 );
buf ( n331870 , n331869 );
buf ( n331871 , n331870 );
nand ( n331872 , n331866 , n331871 );
buf ( n331873 , n331872 );
buf ( n331874 , n331873 );
nand ( n331875 , n12007 , n331874 );
buf ( n331876 , n331875 );
buf ( n331877 , n331876 );
xor ( n331878 , n12002 , n331877 );
buf ( n331879 , n331377 );
not ( n331880 , n331879 );
buf ( n331881 , n3865 );
not ( n331882 , n331881 );
or ( n331883 , n331880 , n331882 );
buf ( n331884 , n323715 );
buf ( n331885 , n545 );
buf ( n12028 , n578 );
xor ( n12029 , n331885 , n12028 );
buf ( n331888 , n12029 );
buf ( n331889 , n331888 );
nand ( n331890 , n331884 , n331889 );
buf ( n331891 , n331890 );
buf ( n331892 , n331891 );
nand ( n12035 , n331883 , n331892 );
buf ( n331894 , n12035 );
buf ( n331895 , n331894 );
xor ( n331896 , n331878 , n331895 );
buf ( n331897 , n331896 );
buf ( n331898 , n331897 );
xor ( n331899 , n331855 , n331898 );
xor ( n12042 , n331413 , n331430 );
and ( n331901 , n12042 , n331438 );
and ( n331902 , n331413 , n331430 );
or ( n12045 , n331901 , n331902 );
buf ( n331904 , n12045 );
buf ( n331905 , n331904 );
xor ( n331906 , n331899 , n331905 );
buf ( n331907 , n331906 );
buf ( n331908 , n331907 );
xor ( n331909 , n11981 , n331908 );
buf ( n331910 , n331909 );
buf ( n331911 , n331910 );
xor ( n331912 , n331826 , n331911 );
buf ( n331913 , n331912 );
xnor ( n12056 , n11881 , n331913 );
buf ( n331915 , n12056 );
nor ( n331916 , n331726 , n331915 );
buf ( n331917 , n331916 );
buf ( n331918 , n331917 );
nor ( n12061 , n331713 , n331918 );
buf ( n331920 , n12061 );
buf ( n331921 , n331920 );
not ( n331922 , n331921 );
buf ( n331923 , n7837 );
not ( n12066 , n331923 );
or ( n331925 , n331922 , n12066 );
buf ( n12068 , n331316 );
nand ( n331927 , n12068 , n331920 );
not ( n12070 , n331927 );
and ( n331929 , n12070 , n7782 );
buf ( n331930 , n331725 );
buf ( n331931 , n12056 );
or ( n331932 , n331930 , n331931 );
buf ( n331933 , n331932 );
buf ( n331934 , n331933 );
not ( n12077 , n331934 );
buf ( n331936 , n11728 );
not ( n12079 , n331936 );
buf ( n331938 , n12079 );
buf ( n331939 , n331938 );
buf ( n331940 , n8092 );
or ( n331941 , n331939 , n331940 );
buf ( n331942 , n331589 );
nand ( n331943 , n331941 , n331942 );
buf ( n331944 , n331943 );
buf ( n331945 , n331944 );
not ( n331946 , n331945 );
or ( n12089 , n12077 , n331946 );
buf ( n331948 , n331725 );
buf ( n331949 , n12056 );
nand ( n12092 , n331948 , n331949 );
buf ( n12093 , n12092 );
buf ( n331952 , n12093 );
nand ( n12095 , n12089 , n331952 );
buf ( n331954 , n12095 );
nor ( n331955 , n331929 , n331954 );
buf ( n331956 , n331955 );
nand ( n331957 , n331925 , n331956 );
buf ( n331958 , n331957 );
not ( n12101 , n331913 );
not ( n12102 , n331737 );
nand ( n12103 , n12102 , n331732 );
not ( n12104 , n12103 );
or ( n12105 , n12101 , n12104 );
nand ( n12106 , n331737 , n331731 );
nand ( n12107 , n12105 , n12106 );
buf ( n12108 , n12107 );
xor ( n12109 , n331744 , n331809 );
and ( n12110 , n12109 , n331816 );
and ( n331969 , n331744 , n331809 );
or ( n331970 , n12110 , n331969 );
buf ( n331971 , n331970 );
buf ( n331972 , n548 );
buf ( n331973 , n560 );
and ( n331974 , n331972 , n331973 );
buf ( n331975 , n331974 );
buf ( n331976 , n331975 );
buf ( n331977 , n3186 );
buf ( n331978 , n321592 );
or ( n331979 , n331977 , n331978 );
buf ( n331980 , n564 );
nand ( n12123 , n331979 , n331980 );
buf ( n331982 , n12123 );
buf ( n331983 , n331982 );
xor ( n331984 , n331976 , n331983 );
buf ( n331985 , n331789 );
not ( n331986 , n331985 );
buf ( n331987 , n3157 );
not ( n331988 , n331987 );
or ( n12131 , n331986 , n331988 );
buf ( n331990 , n323009 );
buf ( n331991 , n544 );
buf ( n331992 , n562 );
xor ( n331993 , n331991 , n331992 );
buf ( n331994 , n331993 );
buf ( n331995 , n331994 );
nand ( n12138 , n331990 , n331995 );
buf ( n331997 , n12138 );
buf ( n331998 , n331997 );
nand ( n331999 , n12131 , n331998 );
buf ( n332000 , n331999 );
buf ( n332001 , n332000 );
xor ( n332002 , n331984 , n332001 );
buf ( n332003 , n332002 );
buf ( n332004 , n332003 );
buf ( n332005 , n331756 );
buf ( n12148 , n331773 );
not ( n12149 , n12148 );
buf ( n12150 , n7031 );
not ( n12151 , n12150 );
or ( n12152 , n12149 , n12151 );
buf ( n332011 , n324855 );
buf ( n332012 , n560 );
buf ( n332013 , n546 );
xor ( n12156 , n332012 , n332013 );
buf ( n332015 , n12156 );
buf ( n332016 , n332015 );
nand ( n332017 , n332011 , n332016 );
buf ( n332018 , n332017 );
buf ( n332019 , n332018 );
nand ( n332020 , n12152 , n332019 );
buf ( n332021 , n332020 );
buf ( n332022 , n332021 );
xor ( n332023 , n332005 , n332022 );
xor ( n12166 , n331765 , n11921 );
and ( n12167 , n12166 , n331796 );
and ( n332026 , n331765 , n11921 );
or ( n332027 , n12167 , n332026 );
buf ( n332028 , n332027 );
buf ( n332029 , n332028 );
xor ( n12172 , n332023 , n332029 );
buf ( n332031 , n12172 );
buf ( n332032 , n332031 );
xor ( n12175 , n332004 , n332032 );
xor ( n332034 , n11903 , n331799 );
and ( n332035 , n332034 , n331806 );
and ( n12178 , n11903 , n331799 );
or ( n332037 , n332035 , n12178 );
buf ( n332038 , n332037 );
buf ( n332039 , n332038 );
xor ( n12182 , n12175 , n332039 );
buf ( n332041 , n12182 );
buf ( n332042 , n332041 );
buf ( n332043 , n548 );
buf ( n332044 , n576 );
and ( n332045 , n332043 , n332044 );
buf ( n332046 , n332045 );
buf ( n332047 , n332046 );
buf ( n332048 , n322474 );
buf ( n332049 , n322468 );
or ( n12192 , n332048 , n332049 );
buf ( n332051 , n580 );
nand ( n332052 , n12192 , n332051 );
buf ( n332053 , n332052 );
buf ( n332054 , n332053 );
xor ( n12197 , n332047 , n332054 );
buf ( n332056 , n331888 );
not ( n12199 , n332056 );
buf ( n332058 , n3865 );
not ( n332059 , n332058 );
or ( n12202 , n12199 , n332059 );
buf ( n332061 , n323715 );
buf ( n332062 , n544 );
buf ( n332063 , n578 );
xor ( n332064 , n332062 , n332063 );
buf ( n332065 , n332064 );
buf ( n12208 , n332065 );
nand ( n12209 , n332061 , n12208 );
buf ( n12210 , n12209 );
buf ( n12211 , n12210 );
nand ( n12212 , n12202 , n12211 );
buf ( n12213 , n12212 );
buf ( n332072 , n12213 );
xor ( n332073 , n12197 , n332072 );
buf ( n332074 , n332073 );
buf ( n332075 , n332074 );
buf ( n332076 , n331851 );
buf ( n332077 , n331870 );
not ( n332078 , n332077 );
buf ( n332079 , n325952 );
not ( n12222 , n332079 );
or ( n12223 , n332078 , n12222 );
buf ( n332082 , n5580 );
buf ( n332083 , n576 );
buf ( n332084 , n546 );
xor ( n12227 , n332083 , n332084 );
buf ( n332086 , n12227 );
buf ( n332087 , n332086 );
nand ( n332088 , n332082 , n332087 );
buf ( n332089 , n332088 );
buf ( n332090 , n332089 );
nand ( n332091 , n12223 , n332090 );
buf ( n332092 , n332091 );
buf ( n332093 , n332092 );
xor ( n12236 , n332076 , n332093 );
xor ( n12237 , n12002 , n331877 );
and ( n12238 , n12237 , n331895 );
and ( n12239 , n12002 , n331877 );
or ( n12240 , n12238 , n12239 );
buf ( n332099 , n12240 );
buf ( n332100 , n332099 );
xor ( n12243 , n12236 , n332100 );
buf ( n332102 , n12243 );
buf ( n332103 , n332102 );
xor ( n12246 , n332075 , n332103 );
xor ( n332105 , n331855 , n331898 );
and ( n332106 , n332105 , n331905 );
and ( n12249 , n331855 , n331898 );
or ( n332108 , n332106 , n12249 );
buf ( n332109 , n332108 );
buf ( n332110 , n332109 );
xor ( n12253 , n12246 , n332110 );
buf ( n332112 , n12253 );
buf ( n332113 , n332112 );
xor ( n332114 , n332042 , n332113 );
xor ( n12257 , n331832 , n331838 );
and ( n12258 , n12257 , n331908 );
and ( n332117 , n331832 , n331838 );
or ( n332118 , n12258 , n332117 );
buf ( n332119 , n332118 );
buf ( n332120 , n332119 );
xor ( n332121 , n332114 , n332120 );
buf ( n332122 , n332121 );
xor ( n12265 , n331971 , n332122 );
xor ( n12266 , n331819 , n331825 );
and ( n12267 , n12266 , n331911 );
and ( n12268 , n331819 , n331825 );
or ( n12269 , n12267 , n12268 );
buf ( n332128 , n12269 );
xor ( n332129 , n12265 , n332128 );
buf ( n332130 , n332129 );
nor ( n332131 , n12108 , n332130 );
buf ( n332132 , n332131 );
buf ( n332133 , n332132 );
not ( n332134 , n332133 );
buf ( n332135 , n12107 );
buf ( n332136 , n332129 );
nand ( n332137 , n332135 , n332136 );
buf ( n332138 , n332137 );
buf ( n332139 , n332138 );
nand ( n332140 , n332134 , n332139 );
buf ( n332141 , n332140 );
xor ( n332142 , n331958 , n332141 );
and ( n12285 , n11448 , n331693 );
nand ( n332144 , n12285 , n329132 );
nand ( n12287 , n11746 , n11755 );
not ( n332146 , n12287 );
not ( n12289 , n11769 );
or ( n12290 , n332146 , n12289 );
not ( n332149 , n11746 );
nand ( n12292 , n332149 , n11758 );
nand ( n332151 , n12290 , n12292 );
not ( n12294 , n8820 );
not ( n332153 , n328669 );
or ( n332154 , n12294 , n332153 );
nand ( n12297 , n332154 , n550 );
not ( n332156 , n329053 );
not ( n332157 , n544 );
not ( n12300 , n328488 );
or ( n12301 , n332157 , n12300 );
nand ( n332160 , n331211 , n328001 );
nand ( n332161 , n12301 , n332160 );
not ( n12304 , n332161 );
or ( n12305 , n332156 , n12304 );
nand ( n332164 , n331662 , n8686 );
nand ( n12307 , n12305 , n332164 );
xor ( n12308 , n12297 , n12307 );
not ( n332167 , n8475 );
not ( n332168 , n11793 );
or ( n332169 , n332167 , n332168 );
not ( n12312 , n548 );
not ( n332171 , n331255 );
or ( n332172 , n12312 , n332171 );
nand ( n12315 , n331608 , n8447 );
nand ( n332174 , n332172 , n12315 );
nand ( n332175 , n332174 , n329668 );
nand ( n12318 , n332169 , n332175 );
xor ( n332177 , n12308 , n12318 );
and ( n332178 , n544 , n11376 );
xor ( n12321 , n332178 , n11755 );
not ( n332180 , n8376 );
and ( n12323 , n8826 , n8378 );
not ( n332182 , n8826 );
and ( n332183 , n332182 , n546 );
or ( n332184 , n12323 , n332183 );
not ( n332185 , n332184 );
or ( n12328 , n332180 , n332185 );
not ( n12329 , n331598 );
nand ( n332188 , n12329 , n329105 );
nand ( n12331 , n12328 , n332188 );
xor ( n332190 , n12321 , n12331 );
xor ( n332191 , n332177 , n332190 );
buf ( n12334 , n11807 );
or ( n332193 , n12334 , n331640 );
nand ( n332194 , n332193 , n11795 );
nand ( n12337 , n12334 , n331640 );
nand ( n332196 , n332194 , n12337 );
xor ( n332197 , n332191 , n332196 );
xor ( n12340 , n332151 , n332197 );
not ( n332199 , n11780 );
buf ( n12342 , n331665 );
nand ( n332201 , n332199 , n12342 );
not ( n12344 , n332201 );
not ( n12345 , n331674 );
or ( n332204 , n12344 , n12345 );
not ( n332205 , n12342 );
nand ( n12348 , n332205 , n11780 );
nand ( n332207 , n332204 , n12348 );
xor ( n332208 , n12340 , n332207 );
or ( n12351 , n11773 , n11818 );
nand ( n332210 , n12351 , n11827 );
nand ( n332211 , n11818 , n11773 );
nand ( n12354 , n332210 , n332211 );
nor ( n332213 , n332208 , n12354 );
nor ( n12355 , n332144 , n332213 );
nand ( n332215 , n11323 , n12355 );
not ( n332216 , n332213 );
nand ( n12358 , n331180 , n11837 , n11448 );
not ( n12359 , n331295 );
nand ( n12360 , n11837 , n12359 );
nand ( n332220 , n12358 , n12360 , n331692 );
nand ( n332221 , n332216 , n332220 );
nand ( n12363 , n332208 , n12354 );
nand ( n12364 , n332215 , n332221 , n12363 );
xor ( n12365 , n332151 , n332197 );
and ( n332225 , n12365 , n332207 );
and ( n332226 , n332151 , n332197 );
or ( n12368 , n332225 , n332226 );
nand ( n12369 , n11803 , n544 );
not ( n12370 , n331597 );
not ( n332230 , n328001 );
and ( n12372 , n12370 , n332230 );
and ( n12373 , n331597 , n328001 );
nor ( n332233 , n12372 , n12373 );
not ( n12375 , n332233 );
not ( n12376 , n331223 );
and ( n12377 , n12375 , n12376 );
and ( n332237 , n332161 , n8686 );
nor ( n12379 , n12377 , n332237 );
not ( n332239 , n12379 );
xor ( n12381 , n12369 , n332239 );
not ( n332241 , n329105 );
not ( n332242 , n332184 );
or ( n12384 , n332241 , n332242 );
not ( n12385 , n546 );
not ( n332245 , n11789 );
or ( n12387 , n12385 , n332245 );
nand ( n12388 , n331645 , n8378 );
nand ( n332248 , n12387 , n12388 );
nand ( n332249 , n332248 , n8376 );
nand ( n12391 , n12384 , n332249 );
xnor ( n12392 , n12381 , n12391 );
not ( n12393 , n8422 );
not ( n12394 , n8447 );
and ( n12395 , n12393 , n12394 );
and ( n332255 , n332174 , n8475 );
nor ( n332256 , n12395 , n332255 );
xor ( n12398 , n12297 , n12307 );
and ( n332258 , n12398 , n12318 );
and ( n12400 , n12297 , n12307 );
or ( n332260 , n332258 , n12400 );
xor ( n332261 , n332256 , n332260 );
xor ( n12403 , n332178 , n11755 );
and ( n332263 , n12403 , n12331 );
and ( n332264 , n332178 , n11755 );
or ( n12406 , n332263 , n332264 );
xor ( n332266 , n332261 , n12406 );
xor ( n12408 , n12392 , n332266 );
xor ( n12409 , n332177 , n332190 );
and ( n12410 , n12409 , n332196 );
and ( n12411 , n332177 , n332190 );
or ( n12412 , n12410 , n12411 );
xor ( n12413 , n12408 , n12412 );
or ( n12414 , n12368 , n12413 );
nand ( n12415 , n12368 , n12413 );
nand ( n12416 , n12414 , n12415 );
not ( n12417 , n12416 );
and ( n12418 , n12364 , n12417 );
not ( n12419 , n12364 );
and ( n12420 , n12419 , n12416 );
nor ( n12421 , n12418 , n12420 );
nand ( n12422 , n332142 , n12421 );
not ( n332282 , n12422 );
and ( n12424 , n331933 , n12093 );
buf ( n332284 , n331712 );
not ( n332285 , n332284 );
buf ( n332286 , n332285 );
not ( n12428 , n332286 );
not ( n332288 , n7837 );
or ( n12430 , n12428 , n332288 );
buf ( n332290 , n7782 );
buf ( n332291 , n4654 );
buf ( n332292 , n332286 );
and ( n332293 , n332290 , n332291 , n332292 );
not ( n332294 , n11728 );
not ( n12436 , n331328 );
or ( n12437 , n332294 , n12436 );
nand ( n332297 , n12437 , n331589 );
buf ( n332298 , n332297 );
nor ( n332299 , n332293 , n332298 );
buf ( n332300 , n332299 );
nand ( n12442 , n12430 , n332300 );
xor ( n332302 , n12424 , n12442 );
not ( n332303 , n332144 );
not ( n12445 , n332303 );
buf ( n332305 , n11323 );
not ( n332306 , n332305 );
or ( n332307 , n12445 , n332306 );
not ( n12449 , n332220 );
nand ( n332309 , n332307 , n12449 );
not ( n12451 , n332213 );
nand ( n12452 , n12451 , n12363 );
and ( n332312 , n332309 , n12452 );
not ( n332313 , n332309 );
not ( n12455 , n12452 );
and ( n332315 , n332313 , n12455 );
nor ( n332316 , n332312 , n332315 );
nor ( n12458 , n332302 , n332316 );
nor ( n332318 , n332282 , n12458 );
not ( n332319 , n332318 );
or ( n332320 , n331708 , n332319 );
buf ( n12462 , n12422 );
not ( n332322 , n332302 );
not ( n12464 , n332316 );
nor ( n332324 , n332322 , n12464 );
and ( n12466 , n12462 , n332324 );
nor ( n332326 , n332142 , n12421 );
nor ( n332327 , n12466 , n332326 );
nand ( n12469 , n332320 , n332327 );
not ( n332329 , n12469 );
not ( n332330 , n332329 );
not ( n332331 , n332330 );
not ( n332332 , n332129 );
not ( n12474 , n12107 );
and ( n332334 , n332332 , n12474 );
nor ( n332335 , n332334 , n331917 );
nand ( n12477 , n332335 , n332286 );
buf ( n332337 , n12477 );
xor ( n332338 , n331971 , n332122 );
and ( n12480 , n332338 , n332128 );
and ( n332340 , n331971 , n332122 );
or ( n332341 , n12480 , n332340 );
buf ( n332342 , n332341 );
not ( n12484 , n332342 );
xor ( n332344 , n332004 , n332032 );
and ( n332345 , n332344 , n332039 );
and ( n12487 , n332004 , n332032 );
or ( n332347 , n332345 , n12487 );
buf ( n332348 , n332347 );
xor ( n12490 , n332042 , n332113 );
and ( n12491 , n12490 , n332120 );
and ( n332351 , n332042 , n332113 );
or ( n332352 , n12491 , n332351 );
buf ( n332353 , n332352 );
xor ( n332354 , n332348 , n332353 );
and ( n332355 , n331867 , n331868 );
buf ( n332356 , n332355 );
buf ( n332357 , n332356 );
buf ( n332358 , n332086 );
not ( n12500 , n332358 );
buf ( n332360 , n325952 );
not ( n332361 , n332360 );
or ( n12503 , n12500 , n332361 );
buf ( n332363 , n5580 );
buf ( n332364 , n545 );
buf ( n332365 , n576 );
xor ( n332366 , n332364 , n332365 );
buf ( n332367 , n332366 );
buf ( n332368 , n332367 );
nand ( n12509 , n332363 , n332368 );
buf ( n332370 , n12509 );
buf ( n332371 , n332370 );
nand ( n12512 , n12503 , n332371 );
buf ( n332373 , n12512 );
buf ( n332374 , n332373 );
xor ( n12515 , n332357 , n332374 );
buf ( n332376 , n332065 );
not ( n12517 , n332376 );
buf ( n332378 , n3865 );
not ( n12519 , n332378 );
or ( n332380 , n12517 , n12519 );
buf ( n332381 , n323715 );
buf ( n332382 , n578 );
nand ( n332383 , n332381 , n332382 );
buf ( n332384 , n332383 );
buf ( n332385 , n332384 );
nand ( n12526 , n332380 , n332385 );
buf ( n332387 , n12526 );
buf ( n332388 , n332387 );
not ( n12529 , n332388 );
buf ( n332390 , n12529 );
buf ( n332391 , n332390 );
xor ( n332392 , n12515 , n332391 );
buf ( n332393 , n332392 );
buf ( n332394 , n332393 );
xor ( n332395 , n332047 , n332054 );
and ( n12536 , n332395 , n332072 );
and ( n332397 , n332047 , n332054 );
or ( n12538 , n12536 , n332397 );
buf ( n332399 , n12538 );
buf ( n332400 , n332399 );
xor ( n12541 , n332394 , n332400 );
xor ( n332402 , n332076 , n332093 );
and ( n12543 , n332402 , n332100 );
and ( n12544 , n332076 , n332093 );
or ( n332405 , n12543 , n12544 );
buf ( n332406 , n332405 );
buf ( n332407 , n332406 );
xor ( n12548 , n12541 , n332407 );
buf ( n332409 , n12548 );
buf ( n332410 , n332409 );
xor ( n12551 , n331976 , n331983 );
and ( n12552 , n12551 , n332001 );
and ( n12553 , n331976 , n331983 );
or ( n332414 , n12552 , n12553 );
buf ( n332415 , n332414 );
buf ( n332416 , n332415 );
and ( n12557 , n331770 , n331771 );
buf ( n332418 , n12557 );
buf ( n332419 , n332418 );
buf ( n332420 , n332015 );
not ( n332421 , n332420 );
buf ( n332422 , n7031 );
not ( n12563 , n332422 );
or ( n12564 , n332421 , n12563 );
buf ( n332425 , n324855 );
buf ( n12566 , n545 );
buf ( n332427 , n560 );
xor ( n332428 , n12566 , n332427 );
buf ( n332429 , n332428 );
buf ( n332430 , n332429 );
nand ( n332431 , n332425 , n332430 );
buf ( n332432 , n332431 );
buf ( n332433 , n332432 );
nand ( n332434 , n12564 , n332433 );
buf ( n332435 , n332434 );
buf ( n332436 , n332435 );
xor ( n332437 , n332419 , n332436 );
buf ( n332438 , n3157 );
not ( n332439 , n332438 );
buf ( n332440 , n332439 );
buf ( n332441 , n332440 );
not ( n332442 , n332441 );
buf ( n332443 , n331994 );
not ( n12584 , n332443 );
buf ( n332445 , n12584 );
buf ( n332446 , n332445 );
not ( n12587 , n332446 );
and ( n12588 , n332442 , n12587 );
buf ( n332449 , n562 );
not ( n12590 , n332449 );
buf ( n12591 , n323009 );
not ( n332452 , n12591 );
buf ( n332453 , n332452 );
buf ( n332454 , n332453 );
nor ( n12595 , n12590 , n332454 );
buf ( n332456 , n12595 );
buf ( n332457 , n332456 );
nor ( n12598 , n12588 , n332457 );
buf ( n332459 , n12598 );
buf ( n332460 , n332459 );
xor ( n12601 , n332437 , n332460 );
buf ( n332462 , n12601 );
buf ( n332463 , n332462 );
xor ( n332464 , n332416 , n332463 );
xor ( n12605 , n332005 , n332022 );
and ( n12606 , n12605 , n332029 );
and ( n12607 , n332005 , n332022 );
or ( n12608 , n12606 , n12607 );
buf ( n332469 , n12608 );
buf ( n332470 , n332469 );
xor ( n12611 , n332464 , n332470 );
buf ( n332472 , n12611 );
buf ( n332473 , n332472 );
xor ( n332474 , n332410 , n332473 );
xor ( n12615 , n332075 , n332103 );
and ( n332476 , n12615 , n332110 );
and ( n332477 , n332075 , n332103 );
or ( n12618 , n332476 , n332477 );
buf ( n332479 , n12618 );
buf ( n332480 , n332479 );
xor ( n12621 , n332474 , n332480 );
buf ( n332482 , n12621 );
xnor ( n12623 , n332354 , n332482 );
buf ( n332484 , n12623 );
nand ( n332485 , n12484 , n332484 );
buf ( n332486 , n332485 );
buf ( n332487 , n332486 );
xor ( n332488 , n332416 , n332463 );
and ( n12629 , n332488 , n332470 );
and ( n332490 , n332416 , n332463 );
or ( n12631 , n12629 , n332490 );
buf ( n332492 , n12631 );
buf ( n12633 , n332492 );
buf ( n332494 , n332459 );
not ( n12635 , n332494 );
buf ( n12636 , n12635 );
buf ( n332497 , n12636 );
xor ( n12638 , n332419 , n332436 );
and ( n332499 , n12638 , n332460 );
and ( n332500 , n332419 , n332436 );
or ( n12641 , n332499 , n332500 );
buf ( n332502 , n12641 );
buf ( n332503 , n332502 );
xor ( n332504 , n332497 , n332503 );
and ( n12645 , n332012 , n332013 );
buf ( n332506 , n12645 );
buf ( n332507 , n332506 );
buf ( n332508 , n332453 );
not ( n12649 , n332508 );
buf ( n332510 , n332440 );
not ( n332511 , n332510 );
or ( n12652 , n12649 , n332511 );
buf ( n332513 , n562 );
nand ( n332514 , n12652 , n332513 );
buf ( n332515 , n332514 );
buf ( n332516 , n332515 );
xor ( n332517 , n332507 , n332516 );
buf ( n332518 , n332429 );
not ( n12659 , n332518 );
buf ( n332520 , n7031 );
not ( n332521 , n332520 );
or ( n12662 , n12659 , n332521 );
buf ( n332523 , n324855 );
buf ( n332524 , n560 );
buf ( n332525 , n544 );
xor ( n332526 , n332524 , n332525 );
buf ( n332527 , n332526 );
buf ( n332528 , n332527 );
nand ( n332529 , n332523 , n332528 );
buf ( n332530 , n332529 );
buf ( n332531 , n332530 );
nand ( n12672 , n12662 , n332531 );
buf ( n332533 , n12672 );
buf ( n332534 , n332533 );
xor ( n12675 , n332517 , n332534 );
buf ( n332536 , n12675 );
buf ( n332537 , n332536 );
xor ( n332538 , n332504 , n332537 );
buf ( n332539 , n332538 );
buf ( n332540 , n332539 );
buf ( n332541 , n332387 );
and ( n332542 , n332083 , n332084 );
buf ( n332543 , n332542 );
buf ( n332544 , n332543 );
buf ( n332545 , n332367 );
not ( n12686 , n332545 );
buf ( n332547 , n325952 );
not ( n332548 , n332547 );
or ( n332549 , n12686 , n332548 );
buf ( n332550 , n544 );
buf ( n332551 , n576 );
xnor ( n332552 , n332550 , n332551 );
buf ( n332553 , n332552 );
buf ( n332554 , n332553 );
not ( n332555 , n332554 );
buf ( n332556 , n5580 );
nand ( n332557 , n332555 , n332556 );
buf ( n332558 , n332557 );
buf ( n332559 , n332558 );
nand ( n332560 , n332549 , n332559 );
buf ( n332561 , n332560 );
buf ( n332562 , n332561 );
xor ( n332563 , n332544 , n332562 );
buf ( n332564 , n3865 );
buf ( n332565 , n323715 );
or ( n332566 , n332564 , n332565 );
buf ( n332567 , n578 );
nand ( n12708 , n332566 , n332567 );
buf ( n332569 , n12708 );
buf ( n332570 , n332569 );
xor ( n12711 , n332563 , n332570 );
buf ( n332572 , n12711 );
buf ( n332573 , n332572 );
xor ( n12714 , n332541 , n332573 );
xor ( n332575 , n332357 , n332374 );
and ( n332576 , n332575 , n332391 );
and ( n12717 , n332357 , n332374 );
or ( n332578 , n332576 , n12717 );
buf ( n332579 , n332578 );
buf ( n332580 , n332579 );
xor ( n332581 , n12714 , n332580 );
buf ( n332582 , n332581 );
buf ( n332583 , n332582 );
xor ( n12724 , n332540 , n332583 );
xor ( n332585 , n332394 , n332400 );
and ( n332586 , n332585 , n332407 );
and ( n12727 , n332394 , n332400 );
or ( n332588 , n332586 , n12727 );
buf ( n332589 , n332588 );
buf ( n332590 , n332589 );
xor ( n332591 , n12724 , n332590 );
buf ( n332592 , n332591 );
buf ( n332593 , n332592 );
xor ( n12734 , n12633 , n332593 );
xor ( n332595 , n332410 , n332473 );
and ( n332596 , n332595 , n332480 );
and ( n12737 , n332410 , n332473 );
or ( n12738 , n332596 , n12737 );
buf ( n332599 , n12738 );
buf ( n332600 , n332599 );
xor ( n12741 , n12734 , n332600 );
buf ( n332602 , n12741 );
buf ( n12743 , n332602 );
not ( n12744 , n12743 );
buf ( n12745 , n12744 );
xor ( n332606 , n332482 , n332348 );
and ( n12747 , n332606 , n332353 );
and ( n332608 , n332482 , n332348 );
nor ( n12749 , n12747 , n332608 );
nand ( n12750 , n12745 , n12749 );
buf ( n332611 , n12750 );
and ( n332612 , n332487 , n332611 );
buf ( n332613 , n332612 );
buf ( n332614 , n332613 );
xor ( n12755 , n12633 , n332593 );
and ( n12756 , n12755 , n332600 );
and ( n12757 , n12633 , n332593 );
or ( n12758 , n12756 , n12757 );
buf ( n332619 , n12758 );
buf ( n332620 , n332619 );
xor ( n12761 , n332497 , n332503 );
and ( n332622 , n12761 , n332537 );
and ( n332623 , n332497 , n332503 );
or ( n12764 , n332622 , n332623 );
buf ( n332625 , n12764 );
buf ( n332626 , n332625 );
buf ( n12767 , n545 );
buf ( n332628 , n560 );
nand ( n332629 , n12767 , n332628 );
buf ( n332630 , n332629 );
buf ( n332631 , n332630 );
buf ( n332632 , n332527 );
not ( n12773 , n332632 );
buf ( n332634 , n7031 );
not ( n332635 , n332634 );
or ( n12776 , n12773 , n332635 );
buf ( n332637 , n324855 );
buf ( n332638 , n560 );
nand ( n12779 , n332637 , n332638 );
buf ( n332640 , n12779 );
buf ( n332641 , n332640 );
nand ( n12782 , n12776 , n332641 );
buf ( n332643 , n12782 );
buf ( n332644 , n332643 );
xor ( n332645 , n332631 , n332644 );
xor ( n332646 , n332507 , n332516 );
and ( n12787 , n332646 , n332534 );
and ( n332648 , n332507 , n332516 );
or ( n332649 , n12787 , n332648 );
buf ( n332650 , n332649 );
buf ( n332651 , n332650 );
xor ( n12792 , n332645 , n332651 );
buf ( n332653 , n12792 );
buf ( n332654 , n332653 );
buf ( n332655 , n545 );
buf ( n332656 , n576 );
nand ( n332657 , n332655 , n332656 );
buf ( n332658 , n332657 );
buf ( n12799 , n332658 );
buf ( n332660 , n325952 );
not ( n12801 , n332660 );
buf ( n12802 , n12801 );
buf ( n332663 , n12802 );
buf ( n332664 , n332553 );
or ( n12805 , n332663 , n332664 );
buf ( n332666 , n5580 );
not ( n332667 , n332666 );
buf ( n332668 , n332667 );
buf ( n332669 , n332668 );
buf ( n332670 , n576 );
not ( n12811 , n332670 );
buf ( n332672 , n12811 );
buf ( n332673 , n332672 );
or ( n332674 , n332669 , n332673 );
nand ( n332675 , n12805 , n332674 );
buf ( n332676 , n332675 );
buf ( n332677 , n332676 );
xor ( n332678 , n12799 , n332677 );
xor ( n12819 , n332544 , n332562 );
and ( n332680 , n12819 , n332570 );
and ( n12821 , n332544 , n332562 );
or ( n12822 , n332680 , n12821 );
buf ( n332683 , n12822 );
buf ( n332684 , n332683 );
xor ( n12825 , n332678 , n332684 );
buf ( n332686 , n12825 );
buf ( n332687 , n332686 );
xor ( n12828 , n332654 , n332687 );
xor ( n12829 , n332541 , n332573 );
and ( n12830 , n12829 , n332580 );
and ( n12831 , n332541 , n332573 );
or ( n12832 , n12830 , n12831 );
buf ( n332693 , n12832 );
buf ( n332694 , n332693 );
xor ( n12835 , n12828 , n332694 );
buf ( n332696 , n12835 );
buf ( n332697 , n332696 );
xor ( n332698 , n332626 , n332697 );
xor ( n332699 , n332540 , n332583 );
and ( n12840 , n332699 , n332590 );
and ( n332701 , n332540 , n332583 );
or ( n12842 , n12840 , n332701 );
buf ( n332703 , n12842 );
buf ( n332704 , n332703 );
xor ( n12845 , n332698 , n332704 );
buf ( n332706 , n12845 );
buf ( n12847 , n332706 );
or ( n12848 , n332620 , n12847 );
buf ( n12849 , n12848 );
buf ( n332710 , n12849 );
nand ( n12851 , n332614 , n332710 );
buf ( n12852 , n12851 );
buf ( n332713 , n12852 );
nor ( n12854 , n332337 , n332713 );
buf ( n332715 , n12854 );
not ( n332716 , n332715 );
buf ( n332717 , n7837 );
buf ( n12858 , n332717 );
buf ( n12859 , n12858 );
not ( n332720 , n12859 );
or ( n12861 , n332716 , n332720 );
not ( n332722 , n327629 );
and ( n332723 , n332715 , n4654 , n332722 );
buf ( n332724 , n332297 );
buf ( n332725 , n332335 );
and ( n12866 , n332724 , n332725 );
buf ( n332727 , n332132 );
buf ( n332728 , n12093 );
or ( n332729 , n332727 , n332728 );
buf ( n332730 , n332138 );
nand ( n332731 , n332729 , n332730 );
buf ( n332732 , n332731 );
buf ( n332733 , n332732 );
nor ( n12874 , n12866 , n332733 );
buf ( n332735 , n12874 );
buf ( n332736 , n332735 );
buf ( n12877 , n332736 );
buf ( n332738 , n12877 );
or ( n332739 , n12852 , n332738 );
buf ( n332740 , n12623 );
not ( n332741 , n332740 );
buf ( n332742 , n332341 );
nand ( n12883 , n332741 , n332742 );
buf ( n12884 , n12883 );
not ( n332745 , n12750 );
or ( n12886 , n12884 , n332745 );
buf ( n332747 , n12749 );
buf ( n332748 , n12745 );
or ( n332749 , n332747 , n332748 );
buf ( n332750 , n332749 );
nand ( n332751 , n12886 , n332750 );
buf ( n332752 , n332751 );
buf ( n332753 , n12849 );
and ( n12894 , n332752 , n332753 );
buf ( n332755 , n332619 );
buf ( n332756 , n332706 );
nand ( n12897 , n332755 , n332756 );
buf ( n332758 , n12897 );
buf ( n12899 , n332758 );
not ( n12900 , n12899 );
buf ( n332761 , n12900 );
buf ( n332762 , n332761 );
nor ( n12903 , n12894 , n332762 );
buf ( n332764 , n12903 );
nand ( n332765 , n332739 , n332764 );
nor ( n12906 , n332723 , n332765 );
nand ( n332767 , n12861 , n12906 );
and ( n12908 , n332524 , n332525 );
buf ( n332769 , n12908 );
buf ( n332770 , n332769 );
buf ( n332771 , n332630 );
xor ( n12912 , n332770 , n332771 );
buf ( n332773 , n324855 );
buf ( n332774 , n7031 );
or ( n12915 , n332773 , n332774 );
buf ( n332776 , n560 );
nand ( n12917 , n12915 , n332776 );
buf ( n332778 , n12917 );
buf ( n332779 , n332778 );
xnor ( n12920 , n12912 , n332779 );
buf ( n332781 , n12920 );
buf ( n332782 , n332781 );
buf ( n12923 , n544 );
buf ( n12924 , n576 );
nand ( n12925 , n12923 , n12924 );
buf ( n12926 , n12925 );
xor ( n12927 , n332658 , n12926 );
buf ( n332788 , n325952 );
buf ( n332789 , n5580 );
or ( n332790 , n332788 , n332789 );
buf ( n332791 , n576 );
nand ( n332792 , n332790 , n332791 );
buf ( n332793 , n332792 );
xor ( n332794 , n12927 , n332793 );
buf ( n332795 , n332794 );
xor ( n332796 , n332782 , n332795 );
xor ( n12937 , n12799 , n332677 );
and ( n332798 , n12937 , n332684 );
and ( n12939 , n12799 , n332677 );
or ( n332800 , n332798 , n12939 );
buf ( n332801 , n332800 );
buf ( n332802 , n332801 );
xor ( n12943 , n332796 , n332802 );
buf ( n332804 , n12943 );
buf ( n332805 , n332804 );
xor ( n12946 , n332654 , n332687 );
and ( n332807 , n12946 , n332694 );
and ( n332808 , n332654 , n332687 );
or ( n12949 , n332807 , n332808 );
buf ( n332810 , n12949 );
buf ( n332811 , n332810 );
xor ( n12952 , n332631 , n332644 );
and ( n12953 , n12952 , n332651 );
and ( n12954 , n332631 , n332644 );
or ( n12955 , n12953 , n12954 );
buf ( n332816 , n12955 );
buf ( n332817 , n332816 );
xnor ( n332818 , n332811 , n332817 );
buf ( n332819 , n332818 );
buf ( n332820 , n332819 );
xnor ( n332821 , n332805 , n332820 );
buf ( n332822 , n332821 );
buf ( n12963 , n332822 );
not ( n12964 , n12963 );
xor ( n332825 , n332626 , n332697 );
and ( n12966 , n332825 , n332704 );
and ( n332827 , n332626 , n332697 );
or ( n12968 , n12966 , n332827 );
buf ( n332829 , n12968 );
buf ( n332830 , n332829 );
not ( n332831 , n332830 );
or ( n12972 , n12964 , n332831 );
buf ( n332833 , n332829 );
buf ( n332834 , n332822 );
or ( n12975 , n332833 , n332834 );
nand ( n332836 , n12972 , n12975 );
buf ( n332837 , n332836 );
not ( n12978 , n332837 );
and ( n12979 , n332767 , n12978 );
not ( n332840 , n332767 );
and ( n332841 , n332840 , n332837 );
nor ( n12982 , n12979 , n332841 );
not ( n332843 , n12982 );
not ( n332844 , n8422 );
not ( n12985 , n8901 );
or ( n332846 , n332844 , n12985 );
nand ( n332847 , n332846 , n548 );
and ( n12988 , n331211 , n544 );
xor ( n332849 , n332847 , n12988 );
not ( n332850 , n329105 );
not ( n12991 , n332248 );
or ( n332852 , n332850 , n12991 );
not ( n332853 , n546 );
not ( n12994 , n331255 );
or ( n332855 , n332853 , n12994 );
nand ( n332856 , n331608 , n8378 );
nand ( n12997 , n332855 , n332856 );
nand ( n332858 , n12997 , n8376 );
nand ( n332859 , n332852 , n332858 );
and ( n13000 , n332849 , n332859 );
and ( n13001 , n332847 , n12988 );
or ( n13002 , n13000 , n13001 );
and ( n13003 , n331597 , n544 );
and ( n332864 , n12997 , n329105 );
and ( n332865 , n8376 , n546 );
nor ( n13006 , n332864 , n332865 );
xor ( n13007 , n13003 , n13006 );
not ( n13008 , n8686 );
and ( n13009 , n8826 , n328001 );
not ( n13010 , n8826 );
and ( n332871 , n13010 , n544 );
or ( n332872 , n13009 , n332871 );
not ( n332873 , n332872 );
or ( n13014 , n13008 , n332873 );
not ( n13015 , n544 );
not ( n13016 , n11789 );
or ( n13017 , n13015 , n13016 );
nand ( n13018 , n331645 , n328001 );
nand ( n332879 , n13017 , n13018 );
nand ( n13020 , n332879 , n329053 );
nand ( n13021 , n13014 , n13020 );
xor ( n332882 , n13007 , n13021 );
xor ( n332883 , n13002 , n332882 );
not ( n13024 , n332872 );
not ( n332885 , n329053 );
or ( n332886 , n13024 , n332885 );
not ( n13027 , n332233 );
nand ( n332888 , n13027 , n8686 );
nand ( n332889 , n332886 , n332888 );
not ( n13030 , n332889 );
nand ( n332891 , n13030 , n332256 );
not ( n13032 , n332891 );
not ( n332893 , n12369 );
not ( n13034 , n12379 );
or ( n13035 , n332893 , n13034 );
nand ( n13036 , n13035 , n12391 );
not ( n13037 , n12369 );
nand ( n13038 , n13037 , n332239 );
nand ( n13039 , n13036 , n13038 );
not ( n13040 , n13039 );
or ( n13041 , n13032 , n13040 );
not ( n13042 , n332256 );
nand ( n13043 , n13042 , n332889 );
nand ( n13044 , n13041 , n13043 );
and ( n13045 , n332883 , n13044 );
and ( n13046 , n13002 , n332882 );
or ( n13047 , n13045 , n13046 );
not ( n13048 , n13006 );
or ( n13049 , n329105 , n8376 );
nand ( n13050 , n13049 , n546 );
and ( n332911 , n8826 , n544 );
xor ( n332912 , n13050 , n332911 );
not ( n332913 , n8686 );
not ( n332914 , n332879 );
or ( n13055 , n332913 , n332914 );
and ( n332916 , n544 , n331608 );
not ( n332917 , n544 );
and ( n332918 , n332917 , n331255 );
nor ( n13059 , n332916 , n332918 );
nand ( n332920 , n13059 , n329053 );
nand ( n13061 , n13055 , n332920 );
xor ( n13062 , n332912 , n13061 );
xor ( n332923 , n13048 , n13062 );
xor ( n332924 , n13003 , n13006 );
and ( n332925 , n332924 , n13021 );
and ( n13066 , n13003 , n13006 );
or ( n332927 , n332925 , n13066 );
xor ( n332928 , n332923 , n332927 );
nor ( n13069 , n13047 , n332928 );
not ( n332930 , n13069 );
not ( n332931 , n332930 );
xor ( n13072 , n332847 , n12988 );
xor ( n332933 , n13072 , n332859 );
xor ( n332934 , n332256 , n332889 );
xnor ( n13075 , n332934 , n13039 );
xor ( n332936 , n332933 , n13075 );
xor ( n13077 , n332256 , n332260 );
and ( n332938 , n13077 , n12406 );
and ( n13079 , n332256 , n332260 );
or ( n13080 , n332938 , n13079 );
and ( n332941 , n332936 , n13080 );
and ( n13082 , n332933 , n13075 );
or ( n332943 , n332941 , n13082 );
xor ( n13084 , n13002 , n332882 );
xor ( n332945 , n13084 , n13044 );
nor ( n332946 , n332943 , n332945 );
not ( n13087 , n332946 );
not ( n332948 , n13087 );
not ( n332949 , n12414 );
xor ( n13090 , n12392 , n332266 );
and ( n332951 , n13090 , n12412 );
and ( n332952 , n12392 , n332266 );
or ( n13093 , n332951 , n332952 );
xor ( n13094 , n332933 , n13075 );
xor ( n13095 , n13094 , n13080 );
nor ( n13096 , n13093 , n13095 );
nor ( n332957 , n332949 , n13096 );
not ( n332958 , n332957 );
buf ( n332959 , n12363 );
nand ( n13100 , n332215 , n332221 , n332959 );
not ( n332961 , n13100 );
or ( n332962 , n332958 , n332961 );
and ( n13103 , n12368 , n12413 );
not ( n332964 , n13096 );
and ( n13105 , n13103 , n332964 );
and ( n13106 , n13093 , n13095 );
nor ( n332967 , n13105 , n13106 );
nand ( n13108 , n332962 , n332967 );
not ( n332969 , n13108 );
or ( n13110 , n332948 , n332969 );
nand ( n13111 , n332943 , n332945 );
nand ( n332972 , n13110 , n13111 );
not ( n332973 , n332972 );
or ( n332974 , n332931 , n332973 );
nand ( n13115 , n13047 , n332928 );
nand ( n332976 , n332974 , n13115 );
not ( n332977 , n332976 );
and ( n13118 , n13059 , n8686 );
and ( n332979 , n329053 , n544 );
nor ( n332980 , n13118 , n332979 );
nand ( n13121 , n331645 , n544 );
and ( n332982 , n332980 , n13121 );
nor ( n13123 , n332980 , n13121 );
nor ( n13124 , n332982 , n13123 );
not ( n13125 , n13124 );
xor ( n13126 , n13050 , n332911 );
and ( n13127 , n13126 , n13061 );
and ( n13128 , n13050 , n332911 );
or ( n13129 , n13127 , n13128 );
not ( n13130 , n13129 );
or ( n13131 , n13125 , n13130 );
or ( n332992 , n13129 , n13124 );
nand ( n13133 , n13131 , n332992 );
not ( n332994 , n13133 );
xor ( n332995 , n13048 , n13062 );
and ( n13136 , n332995 , n332927 );
and ( n13137 , n13048 , n13062 );
or ( n13138 , n13136 , n13137 );
not ( n13139 , n13138 );
or ( n333000 , n332994 , n13139 );
or ( n333001 , n13138 , n13133 );
nand ( n13142 , n333000 , n333001 );
not ( n13143 , n13142 );
or ( n13144 , n332977 , n13143 );
not ( n13145 , n332930 );
not ( n13146 , n332972 );
or ( n333007 , n13145 , n13146 );
not ( n333008 , n13115 );
nor ( n13149 , n333008 , n13142 );
nand ( n13150 , n333007 , n13149 );
nand ( n13151 , n13144 , n13150 );
nand ( n13152 , n332843 , n13151 );
buf ( n333013 , n12477 );
buf ( n13154 , n332613 );
not ( n13155 , n13154 );
buf ( n333016 , n13155 );
buf ( n333017 , n333016 );
nor ( n13158 , n333013 , n333017 );
buf ( n333019 , n13158 );
not ( n333020 , n333019 );
not ( n13161 , n12859 );
or ( n333022 , n333020 , n13161 );
buf ( n333023 , n332722 );
buf ( n333024 , n333019 );
buf ( n333025 , n4654 );
and ( n13166 , n333023 , n333024 , n333025 );
buf ( n333027 , n332738 );
buf ( n333028 , n333016 );
or ( n333029 , n333027 , n333028 );
buf ( n333030 , n332751 );
not ( n333031 , n333030 );
buf ( n333032 , n333031 );
buf ( n333033 , n333032 );
nand ( n333034 , n333029 , n333033 );
buf ( n333035 , n333034 );
buf ( n333036 , n333035 );
nor ( n333037 , n13166 , n333036 );
buf ( n333038 , n333037 );
nand ( n13179 , n333022 , n333038 );
nand ( n13180 , n12849 , n332758 );
not ( n333041 , n13180 );
and ( n13182 , n13179 , n333041 );
not ( n333043 , n13179 );
and ( n13184 , n333043 , n13180 );
nor ( n333045 , n13182 , n13184 );
not ( n13186 , n333045 );
not ( n13187 , n13069 );
nand ( n333048 , n13187 , n13115 );
not ( n333049 , n333048 );
not ( n333050 , n332972 );
or ( n13191 , n333049 , n333050 );
or ( n333052 , n333048 , n332972 );
nand ( n333053 , n13191 , n333052 );
nand ( n13194 , n13186 , n333053 );
buf ( n333055 , n13108 );
not ( n333056 , n332946 );
nand ( n13197 , n333056 , n13111 );
not ( n333058 , n13197 );
and ( n333059 , n333055 , n333058 );
not ( n13200 , n333055 );
and ( n333061 , n13200 , n13197 );
nor ( n333062 , n333059 , n333061 );
not ( n13203 , n332286 );
nand ( n333064 , n332486 , n332335 );
nor ( n333065 , n13203 , n333064 );
not ( n13206 , n333065 );
not ( n13207 , n12859 );
or ( n13208 , n13206 , n13207 );
buf ( n333069 , n332722 );
buf ( n333070 , n333065 );
buf ( n333071 , n4654 );
and ( n333072 , n333069 , n333070 , n333071 );
buf ( n333073 , n332735 );
buf ( n333074 , n332486 );
not ( n333075 , n333074 );
buf ( n333076 , n333075 );
buf ( n333077 , n333076 );
or ( n333078 , n333073 , n333077 );
buf ( n333079 , n12884 );
nand ( n13220 , n333078 , n333079 );
buf ( n333081 , n13220 );
buf ( n333082 , n333081 );
nor ( n333083 , n333072 , n333082 );
buf ( n333084 , n333083 );
nand ( n13225 , n13208 , n333084 );
nand ( n13226 , n332750 , n12750 );
xor ( n13227 , n13225 , n13226 );
nand ( n13228 , n333062 , n13227 );
not ( n13229 , n12414 );
not ( n333090 , n13100 );
or ( n333091 , n13229 , n333090 );
nand ( n13232 , n333091 , n12415 );
not ( n13233 , n332964 );
nor ( n13234 , n13233 , n13106 );
and ( n13235 , n13232 , n13234 );
not ( n333096 , n13232 );
or ( n333097 , n13096 , n13106 );
and ( n13238 , n333096 , n333097 );
nor ( n13239 , n13235 , n13238 );
and ( n13240 , n332486 , n12884 );
not ( n13241 , n13240 );
buf ( n333102 , n332335 );
not ( n333103 , n333102 );
buf ( n333104 , n331712 );
nor ( n333105 , n333103 , n333104 );
buf ( n333106 , n333105 );
nand ( n13247 , n4654 , n333106 , n332722 );
nand ( n333108 , n12859 , n333106 );
nand ( n333109 , n13247 , n333108 , n332738 );
not ( n13250 , n333109 );
or ( n13251 , n13241 , n13250 );
not ( n13252 , n332738 );
nor ( n13253 , n13252 , n13240 );
nand ( n13254 , n13247 , n333108 , n13253 );
nand ( n13255 , n13251 , n13254 );
nand ( n13256 , n13239 , n13255 );
and ( n13257 , n13228 , n13256 );
not ( n13258 , n13257 );
not ( n13259 , n13258 );
nand ( n13260 , n13152 , n13194 , n13259 );
nor ( n333121 , n332331 , n13260 );
buf ( n13262 , n13228 );
not ( n333123 , n13262 );
not ( n13264 , n13255 );
not ( n333125 , n13239 );
nand ( n13266 , n13264 , n333125 );
not ( n13267 , n13266 );
not ( n333128 , n13267 );
or ( n13269 , n333123 , n333128 );
or ( n333130 , n333062 , n13227 );
nand ( n13271 , n13269 , n333130 );
not ( n333132 , n13271 );
and ( n333133 , n13152 , n13194 );
not ( n13274 , n333133 );
or ( n333135 , n333132 , n13274 );
buf ( n333136 , n13152 );
nor ( n13277 , n13186 , n333053 );
and ( n333138 , n333136 , n13277 );
not ( n333139 , n12982 );
nor ( n13280 , n333139 , n13151 );
nor ( n333141 , n333138 , n13280 );
nand ( n13282 , n333135 , n333141 );
nor ( n333143 , n333121 , n13282 );
buf ( n13284 , n10056 );
not ( n13285 , n13284 );
not ( n333146 , n331149 );
or ( n333147 , n13285 , n333146 );
buf ( n333148 , n331158 );
nand ( n13289 , n333147 , n333148 );
nor ( n333150 , n9915 , n9869 );
not ( n333151 , n333150 );
nand ( n13292 , n9869 , n9915 );
nand ( n333153 , n333151 , n13292 );
xnor ( n333154 , n13289 , n333153 );
buf ( n333155 , n7715 );
buf ( n333156 , n7761 );
and ( n333157 , n333155 , n333156 );
buf ( n333158 , n333157 );
not ( n13299 , n333158 );
not ( n333160 , n331316 );
or ( n13301 , n13299 , n333160 );
and ( n13302 , n327673 , n7761 );
not ( n333163 , n7828 );
nor ( n13304 , n13302 , n333163 );
nand ( n333165 , n13301 , n13304 );
buf ( n333166 , n327625 );
not ( n333167 , n333166 );
buf ( n333168 , n327681 );
nor ( n13309 , n333167 , n333168 );
buf ( n13310 , n13309 );
and ( n333171 , n333165 , n13310 );
not ( n13312 , n333165 );
buf ( n333173 , n13310 );
not ( n333174 , n333173 );
buf ( n333175 , n333174 );
and ( n13316 , n13312 , n333175 );
nor ( n333177 , n333171 , n13316 );
not ( n333178 , n333177 );
and ( n13319 , n333154 , n333178 );
buf ( n333180 , n331149 );
nand ( n333181 , n13284 , n333148 );
xnor ( n13322 , n333180 , n333181 );
not ( n13323 , n7715 );
not ( n13324 , n2971 );
not ( n13325 , n4617 );
or ( n333186 , n13324 , n13325 );
nand ( n333187 , n333186 , n4651 );
not ( n13328 , n333187 );
or ( n13329 , n13323 , n13328 );
not ( n13330 , n327673 );
nand ( n13331 , n13329 , n13330 );
nand ( n13332 , n7761 , n7828 );
not ( n333193 , n13332 );
and ( n333194 , n13331 , n333193 );
not ( n333195 , n13331 );
and ( n333196 , n333195 , n13332 );
nor ( n13337 , n333194 , n333196 );
not ( n333198 , n13337 );
nand ( n13339 , n13322 , n333198 );
not ( n333200 , n13339 );
nor ( n333201 , n13319 , n333200 );
not ( n333202 , n333201 );
not ( n333203 , n327561 );
buf ( n13344 , n327556 );
not ( n333205 , n13344 );
or ( n333206 , n333203 , n333205 );
or ( n13347 , n13344 , n327561 );
nand ( n333208 , n333206 , n13347 );
buf ( n333209 , n333208 );
not ( n13350 , n333209 );
buf ( n333211 , n4652 );
not ( n13352 , n333211 );
or ( n13353 , n13350 , n13352 );
buf ( n333214 , n12068 );
buf ( n333215 , n333208 );
or ( n13356 , n333214 , n333215 );
nand ( n333217 , n13353 , n13356 );
buf ( n333218 , n333217 );
not ( n333219 , n333218 );
not ( n13360 , n11282 );
not ( n13361 , n11220 );
not ( n333222 , n330575 );
or ( n333223 , n13361 , n333222 );
nand ( n333224 , n333223 , n11231 );
not ( n13365 , n333224 );
or ( n333226 , n13360 , n13365 );
buf ( n333227 , n11297 );
buf ( n13368 , n11291 );
nand ( n333229 , n333227 , n13368 );
buf ( n333230 , n331118 );
nand ( n13371 , n333229 , n333230 );
nand ( n333232 , n333226 , n13371 );
not ( n333233 , n11284 );
buf ( n13374 , n10330 );
nand ( n333235 , n333233 , n13374 );
xnor ( n13376 , n333232 , n333235 );
nand ( n13377 , n333219 , n13376 );
not ( n333238 , n13374 );
not ( n333239 , n333232 );
or ( n333240 , n333238 , n333239 );
nand ( n13381 , n333240 , n333233 );
buf ( n333242 , n331133 );
or ( n333243 , n11287 , n331136 );
nand ( n13384 , n333242 , n333243 );
not ( n333245 , n13384 );
and ( n333246 , n13381 , n333245 );
not ( n13387 , n13381 );
and ( n333248 , n13387 , n13384 );
nor ( n13389 , n333246 , n333248 );
or ( n13390 , n13344 , n327561 );
nand ( n333251 , n13390 , n331316 );
not ( n13392 , n333251 );
buf ( n333253 , n327670 );
not ( n13394 , n333253 );
buf ( n333255 , n327669 );
not ( n333256 , n333255 );
buf ( n333257 , n7824 );
nand ( n333258 , n333256 , n333257 );
buf ( n333259 , n333258 );
buf ( n333260 , n333259 );
nor ( n13401 , n13394 , n333260 );
buf ( n333262 , n13401 );
not ( n333263 , n333262 );
or ( n13404 , n13392 , n333263 );
not ( n13405 , n333187 );
nand ( n13406 , n13405 , n327670 );
nand ( n13407 , n13406 , n333259 , n13390 );
nand ( n13408 , n13404 , n13407 );
not ( n333269 , n13408 );
nand ( n333270 , n13389 , n333269 );
nand ( n13411 , n13377 , n333270 );
nor ( n333272 , n333202 , n13411 );
buf ( n333273 , n329032 );
not ( n13414 , n333273 );
not ( n333275 , n11323 );
or ( n333276 , n13414 , n333275 );
not ( n13417 , n331176 );
buf ( n333278 , n13417 );
nand ( n333279 , n333276 , n333278 );
nand ( n13420 , n331179 , n9283 );
not ( n333281 , n13420 );
and ( n13422 , n333279 , n333281 );
not ( n13423 , n333279 );
and ( n13424 , n13423 , n13420 );
nor ( n13425 , n13422 , n13424 );
nor ( n333286 , n7815 , n7436 );
not ( n13427 , n333286 );
buf ( n13428 , n327655 );
buf ( n333289 , n7564 );
and ( n333290 , n13428 , n333289 );
not ( n13431 , n327659 );
nor ( n333292 , n333290 , n13431 );
buf ( n13433 , n333187 );
and ( n13434 , n326656 , n326485 );
nor ( n13435 , n13434 , n327400 );
buf ( n333296 , n13435 );
buf ( n333297 , n7564 );
and ( n333298 , n333296 , n333297 );
buf ( n333299 , n333298 );
nand ( n13440 , n327628 , n13433 , n333299 );
buf ( n333301 , n7835 );
buf ( n333302 , n333299 );
nand ( n333303 , n333301 , n333302 );
buf ( n333304 , n333303 );
nand ( n13445 , n333292 , n13440 , n333304 );
not ( n333306 , n13445 );
or ( n13447 , n13427 , n333306 );
not ( n13448 , n333286 );
nand ( n13449 , n13448 , n333292 , n13440 , n333304 );
nand ( n13450 , n13447 , n13449 );
nand ( n13451 , n13425 , n13450 );
buf ( n13452 , n13451 );
buf ( n333313 , n6809 );
buf ( n333314 , n327654 );
nand ( n13455 , n333313 , n333314 );
buf ( n333316 , n13455 );
not ( n13457 , n333316 );
buf ( n333318 , n327400 );
not ( n13459 , n333318 );
buf ( n333320 , n13459 );
nand ( n13461 , n327628 , n333187 , n333320 );
buf ( n333322 , n7835 );
buf ( n333323 , n333320 );
nand ( n13464 , n333322 , n333323 );
buf ( n333325 , n13464 );
buf ( n333326 , n327643 );
buf ( n13467 , n333326 );
buf ( n333328 , n13467 );
nand ( n13469 , n13461 , n333325 , n333328 );
not ( n13470 , n13469 );
or ( n13471 , n13457 , n13470 );
not ( n13472 , n333328 );
nor ( n13473 , n13472 , n333316 );
nand ( n13474 , n333325 , n13473 , n13461 );
nand ( n13475 , n13471 , n13474 );
not ( n13476 , n13475 );
not ( n13477 , n13476 );
nand ( n13478 , n329931 , n331167 );
not ( n13479 , n13478 );
not ( n13480 , n10056 );
nor ( n13481 , n329716 , n329762 );
nor ( n13482 , n13480 , n13481 );
not ( n13483 , n13482 );
not ( n13484 , n331149 );
or ( n13485 , n13483 , n13484 );
not ( n13486 , n331161 );
nand ( n13487 , n13485 , n13486 );
buf ( n13488 , n329924 );
nand ( n13489 , n13487 , n13488 );
not ( n13490 , n331164 );
not ( n13491 , n13490 );
nand ( n13492 , n13489 , n13491 );
not ( n13493 , n13492 );
or ( n13494 , n13479 , n13493 );
not ( n13495 , n13478 );
nand ( n13496 , n13495 , n13489 , n13491 );
nand ( n13497 , n13494 , n13496 );
not ( n13498 , n13497 );
or ( n13499 , n13477 , n13498 );
buf ( n333360 , n333320 );
buf ( n333361 , n333328 );
nand ( n13502 , n333360 , n333361 );
buf ( n333363 , n13502 );
xor ( n13504 , n333363 , n11473 );
not ( n13505 , n13487 );
not ( n13506 , n13505 );
nand ( n13507 , n13491 , n13488 );
not ( n13508 , n13507 );
not ( n13509 , n13508 );
or ( n13510 , n13506 , n13509 );
or ( n13511 , n13508 , n13505 );
nand ( n13512 , n13510 , n13511 );
nand ( n13513 , n13504 , n13512 );
nand ( n13514 , n13499 , n13513 );
not ( n13515 , n13514 );
nand ( n13516 , n13417 , n333273 );
not ( n13517 , n13516 );
and ( n13518 , n332305 , n13517 );
not ( n13519 , n332305 );
and ( n13520 , n13519 , n13516 );
nor ( n13521 , n13518 , n13520 );
not ( n13522 , n13428 );
buf ( n333383 , n331316 );
buf ( n333384 , n327628 );
buf ( n13525 , n13435 );
buf ( n333386 , n13525 );
nand ( n13527 , n333383 , n333384 , n333386 );
buf ( n333388 , n13527 );
buf ( n333389 , n7835 );
buf ( n333390 , n13525 );
nand ( n13531 , n333389 , n333390 );
buf ( n333392 , n13531 );
nand ( n13533 , n13522 , n333388 , n333392 );
nand ( n13534 , n333289 , n327659 );
and ( n13535 , n13533 , n13534 );
not ( n13536 , n13533 );
not ( n13537 , n13534 );
and ( n13538 , n13536 , n13537 );
nor ( n13539 , n13535 , n13538 );
nand ( n13540 , n13521 , n13539 );
buf ( n13541 , n13540 );
nand ( n13542 , n333272 , n13452 , n13515 , n13541 );
not ( n13543 , n13542 );
buf ( n13544 , n13543 );
not ( n13545 , n331017 );
not ( n13546 , n13545 );
buf ( n13547 , n330999 );
nand ( n13548 , n13546 , n13547 );
not ( n13549 , n13548 );
not ( n13550 , n13549 );
buf ( n13551 , n11049 );
buf ( n13552 , n331011 );
nand ( n13553 , n13551 , n13552 );
not ( n13554 , n331013 );
nand ( n13555 , n13553 , n13554 );
not ( n13556 , n13555 );
not ( n13557 , n13556 );
or ( n13558 , n13550 , n13557 );
nand ( n13559 , n13555 , n13548 );
nand ( n13560 , n13558 , n13559 );
buf ( n333421 , n322776 );
not ( n13562 , n333421 );
buf ( n333423 , n13562 );
not ( n13564 , n333423 );
not ( n13565 , n1832 );
or ( n13566 , n13564 , n13565 );
nand ( n13567 , n13566 , n322789 );
not ( n13568 , n13567 );
buf ( n333429 , n322731 );
not ( n13570 , n333429 );
buf ( n333431 , n322759 );
not ( n13572 , n333431 );
buf ( n333433 , n13572 );
buf ( n333434 , n333433 );
nand ( n13575 , n13570 , n333434 );
buf ( n333436 , n13575 );
buf ( n333437 , n333436 );
buf ( n333438 , n322794 );
nand ( n13579 , n333437 , n333438 );
buf ( n333440 , n13579 );
not ( n13581 , n333440 );
nand ( n13582 , n13568 , n13581 );
nand ( n13583 , n333440 , n13567 );
nand ( n13584 , n13560 , n13582 , n13583 );
not ( n13585 , n13584 );
nand ( n13586 , n13554 , n13552 );
not ( n13587 , n13551 );
and ( n13588 , n13586 , n13587 );
not ( n13589 , n13586 );
and ( n333450 , n13589 , n13551 );
nor ( n13591 , n13588 , n333450 );
not ( n333452 , n13591 );
buf ( n333453 , n333423 );
buf ( n333454 , n322789 );
nand ( n13595 , n333453 , n333454 );
buf ( n333456 , n13595 );
not ( n13597 , n333456 );
not ( n13598 , n1832 );
or ( n13599 , n13597 , n13598 );
not ( n13600 , n333456 );
nand ( n13601 , n13600 , n1833 );
nand ( n13602 , n13599 , n13601 );
nand ( n333463 , n333452 , n13602 );
not ( n13604 , n333463 );
not ( n333465 , n13604 );
or ( n333466 , n13585 , n333465 );
nand ( n13607 , n13582 , n13583 );
not ( n13608 , n13560 );
nand ( n333469 , n13607 , n13608 );
nand ( n13610 , n333466 , n333469 );
not ( n333471 , n13610 );
and ( n333472 , n333436 , n333423 );
not ( n333473 , n333472 );
not ( n13614 , n2882 );
and ( n333475 , n1832 , n13614 );
not ( n333476 , n333475 );
or ( n13617 , n333473 , n333476 );
or ( n333478 , n322675 , n322721 );
and ( n333479 , n333478 , n2952 );
nor ( n13620 , n333479 , n322806 );
nand ( n13621 , n13617 , n13620 );
not ( n333482 , n2965 );
nand ( n333483 , n2955 , n322801 );
nand ( n13624 , n333482 , n333483 );
and ( n333485 , n13621 , n13624 );
not ( n333486 , n13621 );
not ( n13627 , n13624 );
and ( n333488 , n333486 , n13627 );
nor ( n333489 , n333485 , n333488 );
not ( n13630 , n331066 );
buf ( n333491 , n331048 );
nand ( n333492 , n13630 , n333491 );
not ( n13633 , n333492 );
not ( n333494 , n11214 );
not ( n13635 , n331018 );
or ( n13636 , n333494 , n13635 );
not ( n13637 , n331064 );
nand ( n13638 , n13636 , n13637 );
not ( n333499 , n13638 );
or ( n13640 , n13633 , n333499 );
or ( n333501 , n13638 , n333492 );
nand ( n333502 , n13640 , n333501 );
nand ( n333503 , n333489 , n333502 );
buf ( n333504 , n322806 );
not ( n333505 , n333504 );
buf ( n333506 , n333478 );
nand ( n13647 , n333505 , n333506 );
buf ( n13648 , n13647 );
not ( n333509 , n13648 );
not ( n13650 , n322779 );
not ( n333511 , n1832 );
or ( n13652 , n13650 , n333511 );
not ( n13653 , n2952 );
nand ( n13654 , n13652 , n13653 );
not ( n13655 , n13654 );
not ( n13656 , n13655 );
or ( n13657 , n333509 , n13656 );
buf ( n13658 , n13648 );
not ( n13659 , n13658 );
buf ( n13660 , n13659 );
nand ( n13661 , n13660 , n13654 );
nand ( n13662 , n13657 , n13661 );
not ( n13663 , n331018 );
nand ( n13664 , n13637 , n11214 );
and ( n13665 , n13663 , n13664 );
not ( n13666 , n13663 );
not ( n13667 , n13664 );
and ( n13668 , n13666 , n13667 );
nor ( n13669 , n13665 , n13668 );
nand ( n13670 , n13662 , n13669 );
and ( n13671 , n333503 , n13670 );
not ( n13672 , n13671 );
or ( n13673 , n333471 , n13672 );
buf ( n13674 , n333503 );
not ( n13675 , n13669 );
not ( n13676 , n13662 );
nand ( n13677 , n13675 , n13676 );
not ( n13678 , n13677 );
and ( n13679 , n13674 , n13678 );
nor ( n13680 , n333489 , n333502 );
nor ( n13681 , n13679 , n13680 );
nand ( n13682 , n13673 , n13681 );
not ( n13683 , n13682 );
not ( n13684 , n13683 );
buf ( n13685 , n324364 );
and ( n13686 , n324276 , n324361 );
nor ( n13687 , n13685 , n13686 );
not ( n13688 , n13687 );
buf ( n333549 , n324459 );
buf ( n13690 , n333549 );
buf ( n333551 , n13690 );
buf ( n333552 , n324402 );
not ( n13693 , n333552 );
buf ( n333554 , n13693 );
nand ( n13695 , n333551 , n333554 );
buf ( n333556 , n2967 );
buf ( n13697 , n333556 );
buf ( n333558 , n13697 );
buf ( n333559 , n322782 );
buf ( n333560 , n1834 );
and ( n13701 , n333559 , n333560 );
buf ( n333562 , n13701 );
nor ( n13703 , n333558 , n333562 );
or ( n13704 , n13695 , n13703 );
and ( n13705 , n324478 , n324486 );
nand ( n13706 , n13704 , n13705 );
not ( n13707 , n13706 );
or ( n13708 , n13688 , n13707 );
or ( n13709 , n13687 , n13706 );
nand ( n13710 , n13708 , n13709 );
not ( n13711 , n13710 );
or ( n13712 , n11273 , n11280 );
not ( n13713 , n13712 );
not ( n13714 , n333224 );
or ( n13715 , n13713 , n13714 );
nand ( n13716 , n13715 , n13368 );
nand ( n13717 , n333227 , n333230 );
not ( n13718 , n13717 );
and ( n13719 , n13716 , n13718 );
not ( n13720 , n13716 );
and ( n13721 , n13720 , n13717 );
nor ( n13722 , n13719 , n13721 );
not ( n13723 , n13722 );
or ( n13724 , n13711 , n13723 );
nand ( n13725 , n13368 , n13712 );
xnor ( n13726 , n333224 , n13725 );
and ( n13727 , n322782 , n1834 );
and ( n13728 , n333551 , n13727 );
and ( n13729 , n324475 , n324468 );
nor ( n13730 , n13728 , n13729 );
buf ( n333591 , n333551 );
buf ( n333592 , n333558 );
nand ( n13733 , n333591 , n333592 );
buf ( n333594 , n13733 );
nand ( n13735 , n13730 , n333594 );
and ( n13736 , n324486 , n333554 );
xnor ( n13737 , n13735 , n13736 );
nand ( n13738 , n13726 , n13737 );
nand ( n13739 , n13724 , n13738 );
not ( n13740 , n13739 );
buf ( n333601 , n2967 );
buf ( n333602 , n324453 );
buf ( n333603 , n324445 );
nand ( n13744 , n333602 , n333603 );
buf ( n333605 , n13744 );
buf ( n333606 , n333605 );
nand ( n13747 , n333601 , n333606 );
buf ( n333608 , n13747 );
buf ( n333609 , n322782 );
buf ( n333610 , n1834 );
buf ( n333611 , n333605 );
nand ( n13752 , n333609 , n333610 , n333611 );
buf ( n333613 , n13752 );
nand ( n13754 , n333608 , n333613 , n324474 );
buf ( n13755 , n4627 );
nand ( n13756 , n324468 , n13755 );
xor ( n13757 , n13754 , n13756 );
not ( n13758 , n13757 );
buf ( n13759 , n10644 );
nand ( n13760 , n11229 , n13759 );
not ( n13761 , n13760 );
not ( n13762 , n330574 );
buf ( n13763 , n11220 );
not ( n13764 , n13763 );
or ( n13765 , n13762 , n13764 );
not ( n13766 , n11224 );
nand ( n13767 , n13765 , n13766 );
not ( n13768 , n13767 );
or ( n13769 , n13761 , n13768 );
not ( n13770 , n330574 );
not ( n13771 , n13763 );
or ( n13772 , n13770 , n13771 );
nand ( n13773 , n13772 , n13766 );
or ( n13774 , n13773 , n13760 );
nand ( n13775 , n13769 , n13774 );
not ( n13776 , n13775 );
or ( n13777 , n13758 , n13776 );
buf ( n333638 , n324456 );
buf ( n333639 , n324474 );
nand ( n13780 , n333638 , n333639 );
buf ( n333641 , n13780 );
xnor ( n13782 , n2971 , n333641 );
not ( n13783 , n13782 );
nand ( n13784 , n330574 , n13766 );
not ( n13785 , n13763 );
and ( n13786 , n13784 , n13785 );
not ( n13787 , n13784 );
and ( n13788 , n13787 , n13763 );
nor ( n13789 , n13786 , n13788 );
nand ( n13790 , n13783 , n13789 );
nand ( n13791 , n13777 , n13790 );
not ( n13792 , n13791 );
nand ( n13793 , n13684 , n13740 , n13792 );
not ( n13794 , n13789 );
nand ( n13795 , n13794 , n13782 );
not ( n13796 , n13795 );
not ( n13797 , n13796 );
nand ( n13798 , n13775 , n13757 );
not ( n13799 , n13798 );
or ( n13800 , n13797 , n13799 );
not ( n13801 , n13775 );
not ( n13802 , n13757 );
nand ( n13803 , n13801 , n13802 );
nand ( n13804 , n13800 , n13803 );
and ( n13805 , n13740 , n13804 );
nand ( n13806 , n13722 , n13710 );
not ( n13807 , n13806 );
nor ( n13808 , n13737 , n13726 );
not ( n13809 , n13808 );
or ( n13810 , n13807 , n13809 );
not ( n13811 , n13710 );
not ( n13812 , n13722 );
nand ( n13813 , n13811 , n13812 );
nand ( n13814 , n13810 , n13813 );
nor ( n13815 , n13805 , n13814 );
nor ( n13816 , n13608 , n13607 );
nor ( n13817 , n333452 , n13602 );
nor ( n13818 , n13816 , n13817 );
nand ( n13819 , n13669 , n13662 );
nand ( n13820 , n1656 , n320972 );
nand ( n13821 , n1489 , n320978 );
nand ( n13822 , n1826 , n13820 , n13821 );
or ( n13823 , n320978 , n1489 );
buf ( n333684 , n321556 );
not ( n13825 , n333684 );
buf ( n333686 , n321545 );
nor ( n13827 , n13825 , n333686 );
buf ( n333688 , n13827 );
nand ( n13829 , n320972 , n333688 , n321541 );
nand ( n13830 , n13823 , n13829 );
or ( n13831 , n13822 , n13830 );
not ( n13832 , n13821 );
not ( n13833 , n13823 );
or ( n333694 , n13832 , n13833 );
nand ( n333695 , n13829 , n13820 , n1826 );
nand ( n13836 , n333694 , n333695 );
nand ( n13837 , n13831 , n13836 );
not ( n13838 , n13837 );
not ( n13839 , n330778 );
not ( n333700 , n330885 );
or ( n333701 , n13839 , n333700 );
nand ( n13842 , n333701 , n330890 );
not ( n13843 , n13842 );
not ( n13844 , n330745 );
not ( n13845 , n330717 );
or ( n13846 , n13844 , n13845 );
nand ( n333707 , n13846 , n330896 );
not ( n333708 , n333707 );
or ( n333709 , n13843 , n333708 );
or ( n13850 , n13842 , n333707 );
nand ( n333711 , n333709 , n13850 );
buf ( n13852 , n333711 );
and ( n13853 , n13838 , n13852 );
buf ( n333714 , n330885 );
not ( n333715 , n333714 );
nand ( n13856 , n330890 , n330778 );
not ( n333717 , n13856 );
or ( n333718 , n333715 , n333717 );
not ( n13859 , n13856 );
not ( n333720 , n333714 );
nand ( n333721 , n13859 , n333720 );
nand ( n13862 , n333718 , n333721 );
not ( n333723 , n13862 );
nand ( n333724 , n1826 , n320972 );
not ( n13865 , n333724 );
and ( n13866 , n1819 , n13865 );
not ( n13867 , n1819 );
and ( n13868 , n13867 , n333724 );
nor ( n333729 , n13866 , n13868 );
nor ( n333730 , n333723 , n333729 );
nor ( n13871 , n13853 , n333730 );
not ( n13872 , n13871 );
not ( n13873 , n1558 );
not ( n13874 , n321304 );
or ( n13875 , n13873 , n13874 );
nand ( n333736 , n13875 , n321394 );
buf ( n333737 , n333736 );
not ( n13878 , n333737 );
buf ( n333739 , n1799 );
not ( n333740 , n333739 );
buf ( n333741 , n321549 );
buf ( n333742 , n321553 );
nand ( n13883 , n333741 , n333742 );
buf ( n333744 , n13883 );
buf ( n333745 , n333744 );
not ( n13886 , n333745 );
or ( n333747 , n333740 , n13886 );
buf ( n333748 , n1649 );
nand ( n333749 , n333747 , n333748 );
buf ( n333750 , n333749 );
buf ( n333751 , n333750 );
not ( n333752 , n333751 );
or ( n13893 , n13878 , n333752 );
buf ( n333754 , n333736 );
buf ( n333755 , n333750 );
or ( n13896 , n333754 , n333755 );
nand ( n333757 , n13893 , n13896 );
buf ( n333758 , n333757 );
not ( n333759 , n333758 );
or ( n333760 , n330781 , n10964 );
buf ( n13901 , n11035 );
nand ( n333762 , n333760 , n13901 );
nand ( n333763 , n330876 , n330880 );
and ( n333764 , n333762 , n333763 );
not ( n13905 , n333762 );
not ( n333766 , n333763 );
and ( n13907 , n13905 , n333766 );
nor ( n13908 , n333764 , n13907 );
not ( n333769 , n13908 );
nand ( n333770 , n333759 , n333769 );
buf ( n333771 , n333770 );
buf ( n333772 , n321541 );
not ( n333773 , n333772 );
buf ( n333774 , n333773 );
not ( n13915 , n333774 );
buf ( n333776 , n1649 );
buf ( n333777 , n321556 );
nand ( n13918 , n333776 , n333777 );
buf ( n13919 , n13918 );
not ( n333780 , n13919 );
not ( n13921 , n333780 );
or ( n333782 , n13915 , n13921 );
buf ( n333783 , n321541 );
buf ( n333784 , n13919 );
nand ( n13925 , n333783 , n333784 );
buf ( n13926 , n13925 );
nand ( n333787 , n333782 , n13926 );
not ( n13928 , n333787 );
buf ( n13929 , n330875 );
nand ( n333790 , n330880 , n330830 );
xnor ( n333791 , n13929 , n333790 );
nand ( n333792 , n13928 , n333791 );
not ( n13933 , n333792 );
not ( n333794 , n321535 );
not ( n333795 , n321532 );
or ( n13936 , n333794 , n333795 );
nand ( n333797 , n13936 , n1707 );
not ( n333798 , n321528 );
nand ( n13939 , n333798 , n1748 );
or ( n333800 , n333797 , n13939 );
not ( n333801 , n1797 );
not ( n13942 , n1707 );
or ( n333803 , n333801 , n13942 );
not ( n333804 , n321528 );
nand ( n13945 , n333804 , n1748 );
nand ( n333806 , n333803 , n13945 );
nand ( n13947 , n333800 , n333806 );
not ( n333808 , n13947 );
and ( n13949 , n11026 , n330871 );
buf ( n13950 , n11010 );
xor ( n333811 , n13949 , n13950 );
nand ( n333812 , n333808 , n333811 );
not ( n333813 , n333812 );
not ( n13954 , n11007 );
not ( n333815 , n330857 );
nor ( n333816 , n333815 , n330846 );
not ( n13957 , n333816 );
not ( n333818 , n13957 );
or ( n333819 , n13954 , n333818 );
not ( n13960 , n11007 );
nand ( n333821 , n13960 , n333816 );
nand ( n333822 , n333819 , n333821 );
not ( n333823 , n333822 );
xor ( n13964 , n1745 , n1780 );
xor ( n333825 , n13964 , n1747 );
not ( n13966 , n333825 );
and ( n13967 , n333823 , n13966 );
not ( n333828 , n11006 );
nand ( n333829 , n333828 , n11002 , n11000 );
and ( n333830 , n333829 , n11007 );
and ( n13971 , n321502 , n1771 );
not ( n333832 , n321502 );
and ( n333833 , n333832 , n1772 );
nor ( n13974 , n13971 , n333833 );
xor ( n333835 , n13974 , n1776 );
not ( n333836 , n333835 );
nand ( n13977 , n333830 , n333836 );
not ( n333838 , n11005 );
buf ( n333839 , n321499 );
buf ( n333840 , n321494 );
xor ( n333841 , n333839 , n333840 );
buf ( n333842 , n333841 );
not ( n333843 , n333842 );
and ( n13984 , n333838 , n333843 );
not ( n13985 , n13984 );
and ( n333846 , n13977 , n13985 );
nor ( n333847 , n333836 , n333830 );
nor ( n333848 , n333846 , n333847 );
nor ( n13989 , n13967 , n333848 );
not ( n333850 , n13989 );
or ( n333851 , n333813 , n333850 );
nand ( n13992 , n333825 , n333822 );
not ( n333853 , n13992 );
not ( n333854 , n13947 );
nand ( n13995 , n333854 , n333811 );
and ( n333856 , n333853 , n13995 );
not ( n333857 , n13947 );
nor ( n13998 , n333857 , n333811 );
nor ( n333859 , n333856 , n13998 );
nand ( n333860 , n333851 , n333859 );
not ( n14001 , n333860 );
nor ( n333862 , n13933 , n14001 );
and ( n333863 , n333771 , n333862 );
not ( n14004 , n333863 );
or ( n333865 , n13872 , n14004 );
not ( n333866 , n333791 );
nand ( n14007 , n333866 , n333787 );
not ( n333868 , n14007 );
not ( n333869 , n333868 );
not ( n14010 , n333770 );
or ( n14011 , n333869 , n14010 );
nand ( n14012 , n13908 , n333758 );
nand ( n14013 , n14011 , n14012 );
buf ( n333874 , n14013 );
and ( n333875 , n333874 , n13871 );
not ( n14016 , n333711 );
nor ( n14017 , n14016 , n13837 );
not ( n14018 , n13862 );
nand ( n14019 , n14018 , n333729 );
or ( n14020 , n14017 , n14019 );
nand ( n333881 , n13837 , n14016 );
nand ( n333882 , n14020 , n333881 );
nor ( n14023 , n333875 , n333882 );
nand ( n14024 , n333865 , n14023 );
buf ( n14025 , n14024 );
nand ( n14026 , n13674 , n13818 , n13819 , n14025 );
not ( n333887 , n14026 );
nand ( n333888 , n13740 , n13792 , n333887 );
nand ( n14029 , n13793 , n13815 , n333888 );
buf ( n14030 , n14029 );
not ( n14031 , n14030 );
not ( n14032 , n14031 );
and ( n14033 , n13544 , n14032 );
nand ( n333894 , n13451 , n13540 );
nor ( n333895 , n333894 , n13514 );
not ( n333896 , n333895 );
not ( n14037 , n333201 );
not ( n333898 , n333218 );
nor ( n14039 , n333898 , n13376 );
not ( n14040 , n14039 );
nand ( n333901 , n13389 , n333269 );
not ( n333902 , n333901 );
or ( n14043 , n14040 , n333902 );
not ( n333904 , n13389 );
nand ( n333905 , n333904 , n13408 );
nand ( n14046 , n14043 , n333905 );
not ( n333907 , n14046 );
or ( n333908 , n14037 , n333907 );
not ( n14049 , n333177 );
nand ( n333910 , n14049 , n333154 );
not ( n333911 , n13337 );
nor ( n14052 , n333911 , n13322 );
and ( n14053 , n333910 , n14052 );
nor ( n14054 , n333154 , n333178 );
nor ( n14055 , n14053 , n14054 );
nand ( n333916 , n333908 , n14055 );
not ( n333917 , n333916 );
or ( n14058 , n333896 , n333917 );
nand ( n333919 , n13476 , n13497 );
not ( n333920 , n333919 );
nor ( n14061 , n333920 , n333894 );
not ( n333922 , n13497 );
not ( n14063 , n13476 );
nand ( n333924 , n333922 , n14063 );
nand ( n333925 , n333363 , n11473 );
not ( n333926 , n333925 );
or ( n333927 , n333363 , n11473 );
not ( n14068 , n333927 );
or ( n333929 , n333926 , n14068 );
and ( n333930 , n13505 , n13508 );
not ( n14071 , n13505 );
and ( n333932 , n14071 , n13507 );
nor ( n333933 , n333930 , n333932 );
nand ( n14074 , n333929 , n333933 );
nand ( n333935 , n333924 , n14074 );
and ( n333936 , n14061 , n333935 );
not ( n14077 , n13451 );
nor ( n14078 , n13539 , n13521 );
not ( n14079 , n14078 );
or ( n14080 , n14077 , n14079 );
not ( n333941 , n13425 );
not ( n333942 , n13450 );
nand ( n14083 , n333941 , n333942 );
nand ( n333944 , n14080 , n14083 );
nor ( n14085 , n333936 , n333944 );
nand ( n333946 , n14058 , n14085 );
buf ( n14087 , n333946 );
nor ( n14088 , n14033 , n14087 );
not ( n333949 , n14088 );
not ( n333950 , n327946 );
nand ( n14091 , n333950 , n331304 );
and ( n333952 , n331701 , n14091 );
and ( n14093 , n333952 , n332318 );
buf ( n333954 , n14093 );
not ( n333955 , n333954 );
nor ( n14096 , n333955 , n13260 );
nand ( n333957 , n333949 , n14096 );
nand ( n333958 , n333143 , n333957 );
not ( n14099 , n333958 );
buf ( n14100 , n14099 );
nand ( n14101 , n13543 , n14032 );
not ( n14102 , n14101 );
not ( n333963 , n333895 );
not ( n333964 , n333916 );
or ( n333965 , n333963 , n333964 );
nand ( n14106 , n333965 , n14085 );
not ( n333967 , n14106 );
not ( n333968 , n333967 );
or ( n14109 , n14102 , n333968 );
buf ( n333970 , n14091 );
not ( n14111 , n333970 );
buf ( n14112 , n331305 );
nor ( n14113 , n14111 , n14112 );
not ( n14114 , n14113 );
nand ( n14115 , n14109 , n14114 );
nand ( n333976 , n14101 , n333967 , n14113 );
nand ( n333977 , n14115 , n333976 );
buf ( n333978 , n333977 );
nand ( n14119 , n13683 , n14026 );
not ( n333980 , n13782 );
buf ( n333981 , n13789 );
nand ( n14122 , n333980 , n333981 );
nand ( n333983 , n14122 , n13795 );
not ( n14124 , n333983 );
and ( n14125 , n14119 , n14124 );
not ( n333986 , n14119 );
and ( n14127 , n333986 , n333983 );
nor ( n14128 , n14125 , n14127 );
buf ( n14129 , n14128 );
and ( n14130 , n13670 , n13677 );
not ( n333991 , n14024 );
not ( n333992 , n13584 );
nor ( n333993 , n333992 , n13817 );
not ( n14134 , n333993 );
or ( n333995 , n333991 , n14134 );
not ( n333996 , n13610 );
nand ( n14137 , n333995 , n333996 );
xor ( n333998 , n14130 , n14137 );
buf ( n14139 , n333998 );
xor ( n334000 , n13984 , n333836 );
xnor ( n14141 , n334000 , n333830 );
buf ( n334002 , n14141 );
buf ( n14143 , n321273 );
buf ( n14144 , n320864 );
buf ( n334005 , n324348 );
buf ( n14146 , n322653 );
buf ( n334007 , n322408 );
buf ( n14148 , n327922 );
buf ( n334009 , n322071 );
buf ( n334010 , n327547 );
buf ( n14151 , n331453 );
buf ( n334012 , n322433 );
buf ( n14153 , n4574 );
buf ( n334014 , n324270 );
buf ( n334015 , n322581 );
buf ( n14156 , n321222 );
buf ( n334017 , n321100 );
buf ( n14158 , n320550 );
buf ( n14159 , n322706 );
not ( n14160 , n13280 );
nand ( n14161 , n14160 , n333136 );
not ( n14162 , n14161 );
not ( n14163 , n332330 );
not ( n334024 , n333045 );
nand ( n14165 , n334024 , n333053 );
and ( n334026 , n13257 , n14165 );
not ( n334027 , n334026 );
or ( n14168 , n14163 , n334027 );
and ( n334029 , n13271 , n13194 );
nor ( n334030 , n334029 , n13277 );
nand ( n14171 , n14168 , n334030 );
not ( n14172 , n14171 );
nand ( n14173 , n333954 , n334026 , n13544 , n14032 );
not ( n14174 , n14173 );
not ( n14175 , n14174 );
nand ( n334036 , n333954 , n334026 , n14087 );
nand ( n334037 , n14162 , n14172 , n14175 , n334036 );
not ( n14178 , n334037 );
not ( n334039 , n14174 );
not ( n334040 , n14171 );
nand ( n14181 , n334039 , n334040 , n334036 );
buf ( n334042 , n14161 );
nand ( n334043 , n14181 , n334042 );
not ( n14184 , n334043 );
or ( n334045 , n14178 , n14184 );
and ( n334046 , n333952 , n332318 );
buf ( n14187 , n13256 );
nand ( n334048 , n334046 , n13543 , n14032 , n14187 );
nand ( n334049 , n14106 , n14093 , n14187 );
and ( n14190 , n14187 , n12469 );
nor ( n14191 , n14190 , n13267 );
nand ( n14192 , n334048 , n334049 , n14191 );
nand ( n14193 , n333130 , n13262 );
not ( n334054 , n14193 );
and ( n334055 , n14192 , n334054 );
not ( n14196 , n14192 );
and ( n334057 , n14196 , n14193 );
nor ( n334058 , n334055 , n334057 );
buf ( n14199 , n334058 );
nand ( n334060 , n334045 , n14199 );
not ( n334061 , n334060 );
nand ( n14202 , n11849 , n331701 );
not ( n334063 , n14202 );
nand ( n14204 , n14106 , n333970 );
not ( n14205 , n14031 );
nand ( n14206 , n14205 , n333970 , n13543 );
not ( n14207 , n14112 );
nand ( n14208 , n14204 , n14206 , n14207 );
not ( n14209 , n14208 );
or ( n334070 , n334063 , n14209 );
nor ( n14211 , n14202 , n14112 );
nand ( n334072 , n14204 , n14206 , n14211 );
nand ( n14213 , n334070 , n334072 );
and ( n14214 , n14213 , n333977 );
nand ( n14215 , n13452 , n14083 );
not ( n14216 , n14215 );
nand ( n14217 , n13539 , n13521 );
and ( n14218 , n13515 , n14217 );
not ( n14219 , n13411 );
and ( n14220 , n333201 , n14219 );
nand ( n14221 , n14218 , n14220 , n14030 );
nand ( n14222 , n14218 , n333916 );
buf ( n334083 , n14217 );
and ( n14224 , n14074 , n333924 );
nor ( n334085 , n14224 , n333920 );
and ( n14226 , n334083 , n334085 );
nor ( n14227 , n14226 , n14078 );
nand ( n334088 , n14221 , n14222 , n14227 );
not ( n14229 , n334088 );
or ( n334090 , n14216 , n14229 );
not ( n14231 , n14215 );
nand ( n334092 , n14221 , n14222 , n14227 , n14231 );
nand ( n14233 , n334090 , n334092 );
not ( n334094 , n13377 );
buf ( n14235 , n14029 );
not ( n14236 , n14235 );
or ( n14237 , n334094 , n14236 );
not ( n14238 , n14039 );
nand ( n14239 , n14237 , n14238 );
and ( n14240 , n333905 , n333270 );
not ( n14241 , n14240 );
nand ( n14242 , n14239 , n14241 );
not ( n14243 , n14242 );
not ( n14244 , n14239 );
nand ( n14245 , n14244 , n14240 );
not ( n14246 , n14245 );
or ( n14247 , n14243 , n14246 );
nand ( n14248 , n13377 , n14238 );
not ( n14249 , n14248 );
not ( n14250 , n14030 );
or ( n14251 , n14249 , n14250 );
or ( n14252 , n14030 , n14248 );
nand ( n14253 , n14251 , n14252 );
buf ( n14254 , n14253 );
nand ( n14255 , n14247 , n14254 );
not ( n14256 , n14255 );
nand ( n14257 , n333924 , n333919 );
not ( n14258 , n14257 );
buf ( n14259 , n13513 );
nand ( n14260 , n333916 , n14259 );
nand ( n14261 , n14235 , n333272 , n14259 );
not ( n14262 , n333925 );
not ( n14263 , n333927 );
or ( n14264 , n14262 , n14263 );
nand ( n14265 , n14264 , n333933 );
nand ( n14266 , n14260 , n14261 , n14265 );
not ( n14267 , n14266 );
or ( n14268 , n14258 , n14267 );
not ( n14269 , n14257 );
nand ( n14270 , n14269 , n14260 , n14265 , n14261 );
nand ( n14271 , n14268 , n14270 );
nand ( n14272 , n14233 , n14256 , n14271 );
nand ( n14273 , n333916 , n13515 );
nand ( n14274 , n14220 , n14030 , n13515 );
not ( n14275 , n334085 );
nand ( n14276 , n14273 , n14274 , n14275 );
not ( n14277 , n14078 );
nand ( n14278 , n14277 , n334083 );
not ( n14279 , n14278 );
and ( n14280 , n14276 , n14279 );
not ( n14281 , n14276 );
and ( n14282 , n14281 , n14278 );
nor ( n14283 , n14280 , n14282 );
not ( n14284 , n14235 );
not ( n14285 , n14220 );
or ( n14286 , n14284 , n14285 );
not ( n14287 , n333916 );
nand ( n14288 , n14286 , n14287 );
nand ( n14289 , n14265 , n14259 );
not ( n14290 , n14289 );
and ( n14291 , n14288 , n14290 );
not ( n14292 , n14288 );
and ( n14293 , n14292 , n14289 );
nor ( n14294 , n14291 , n14293 );
and ( n14295 , n14283 , n14294 );
buf ( n14296 , n333200 );
nor ( n14297 , n14296 , n13411 );
not ( n14298 , n14297 );
not ( n14299 , n14235 );
or ( n14300 , n14298 , n14299 );
not ( n14301 , n14296 );
buf ( n14302 , n14046 );
and ( n14303 , n14301 , n14302 );
buf ( n14304 , n14052 );
nor ( n14305 , n14303 , n14304 );
nand ( n14306 , n14300 , n14305 );
not ( n14307 , n14054 );
nand ( n14308 , n14307 , n333910 );
not ( n14309 , n14308 );
and ( n14310 , n14306 , n14309 );
not ( n14311 , n14306 );
and ( n14312 , n14311 , n14308 );
nor ( n14313 , n14310 , n14312 );
not ( n14314 , n14219 );
not ( n14315 , n14235 );
or ( n14316 , n14314 , n14315 );
not ( n14317 , n14302 );
nand ( n14318 , n14316 , n14317 );
not ( n14319 , n14301 );
nor ( n14320 , n14319 , n14304 );
and ( n14321 , n14318 , n14320 );
not ( n14322 , n14318 );
not ( n14323 , n14320 );
and ( n14324 , n14322 , n14323 );
nor ( n14325 , n14321 , n14324 );
nand ( n14326 , n14313 , n14325 );
not ( n14327 , n14326 );
nand ( n14328 , n14295 , n14327 );
nor ( n14329 , n14272 , n14328 );
and ( n14330 , n14214 , n14329 );
not ( n14331 , n13277 );
nand ( n14332 , n14331 , n13194 );
not ( n14333 , n14332 );
nand ( n14334 , n13259 , n333954 );
and ( n14335 , n13544 , n14032 );
nor ( n14336 , n14335 , n14087 );
or ( n14337 , n14334 , n14336 );
buf ( n14338 , n12469 );
not ( n14339 , n13258 );
and ( n14340 , n14338 , n14339 );
nor ( n14341 , n14340 , n13271 );
nand ( n14342 , n14337 , n14341 );
not ( n14343 , n14342 );
or ( n14344 , n14333 , n14343 );
or ( n14345 , n14334 , n14336 );
nand ( n14346 , n14345 , n14341 );
or ( n14347 , n14346 , n14332 );
nand ( n14348 , n14344 , n14347 );
not ( n14349 , n14348 );
not ( n14350 , n333952 );
buf ( n14351 , n12458 );
nor ( n14352 , n14350 , n14351 );
nand ( n14353 , n14352 , n13543 , n14032 );
not ( n14354 , n14351 );
buf ( n14355 , n331707 );
and ( n14356 , n14354 , n14355 );
buf ( n14357 , n332324 );
nor ( n14358 , n14356 , n14357 );
not ( n14359 , n332326 );
nand ( n14360 , n14359 , n12462 );
not ( n14361 , n14360 );
nand ( n14362 , n14353 , n14358 , n14361 );
not ( n14363 , n14362 );
not ( n14364 , n14363 );
nand ( n14365 , n14352 , n14106 );
not ( n14366 , n14365 );
or ( n14367 , n14364 , n14366 );
not ( n14368 , n14365 );
nand ( n14369 , n14353 , n14358 );
or ( n14370 , n14368 , n14369 );
nand ( n14371 , n14370 , n14360 );
nand ( n334232 , n14367 , n14371 );
nand ( n14373 , n331701 , n14091 );
not ( n334234 , n14373 );
not ( n14375 , n334234 );
not ( n334236 , n14106 );
or ( n14377 , n14375 , n334236 );
nor ( n334238 , n14373 , n14031 );
and ( n334239 , n334238 , n13543 );
nor ( n14380 , n334239 , n14355 );
nand ( n14381 , n14377 , n14380 );
nor ( n14382 , n14357 , n14351 );
and ( n14383 , n14381 , n14382 );
not ( n14384 , n14381 );
not ( n14385 , n14382 );
and ( n334246 , n14384 , n14385 );
nor ( n14387 , n14383 , n334246 );
nand ( n334248 , n334232 , n14387 );
nor ( n334249 , n14349 , n334248 );
nand ( n14390 , n14093 , n13543 , n14032 );
nand ( n334251 , n14106 , n334046 );
nand ( n14392 , n14390 , n334251 , n332329 );
nand ( n14393 , n14187 , n13266 );
nand ( n14394 , n14392 , n14393 );
not ( n14395 , n14394 );
not ( n334256 , n14392 );
not ( n334257 , n14393 );
nand ( n334258 , n334256 , n334257 );
not ( n14399 , n334258 );
or ( n334260 , n14395 , n14399 );
buf ( n14401 , n13738 );
and ( n14402 , n13804 , n14401 );
not ( n334263 , n13808 );
not ( n334264 , n334263 );
nor ( n334265 , n14402 , n334264 );
nand ( n14406 , n13792 , n333887 , n14401 );
nand ( n334267 , n13684 , n14401 , n13792 );
nand ( n334268 , n334265 , n14406 , n334267 );
nand ( n14409 , n13813 , n13806 );
not ( n334270 , n14409 );
and ( n334271 , n334268 , n334270 );
not ( n14412 , n334268 );
and ( n334273 , n14412 , n14409 );
nor ( n334274 , n334271 , n334273 );
not ( n334275 , n334274 );
not ( n14416 , n576 );
and ( n334277 , n334275 , n14416 );
and ( n14418 , n333503 , n13818 , n13819 );
and ( n334279 , n14418 , n14025 );
nand ( n334280 , n13792 , n334279 );
not ( n14421 , n13791 );
nand ( n14422 , n14421 , n13682 );
not ( n334283 , n13804 );
nand ( n334284 , n334280 , n14422 , n334283 );
nand ( n334285 , n334263 , n14401 );
nand ( n14426 , n334284 , n334285 );
not ( n334287 , n334285 );
nand ( n334288 , n334287 , n14422 , n334283 , n334280 );
not ( n14429 , n577 );
and ( n334290 , n14426 , n334288 , n14429 );
nor ( n334291 , n334277 , n334290 );
not ( n14432 , n334291 );
nand ( n334293 , n13801 , n13802 );
and ( n334294 , n334293 , n13798 );
nand ( n14435 , n13682 , n14122 );
nand ( n334296 , n14122 , n14418 , n14025 );
buf ( n334297 , n13795 );
nand ( n14438 , n14435 , n334296 , n334297 );
xor ( n334299 , n334294 , n14438 );
not ( n14440 , n334299 );
not ( n334301 , n578 );
nand ( n334302 , n14440 , n334301 );
not ( n14443 , n334302 );
and ( n334304 , n14128 , n579 );
not ( n334305 , n334304 );
or ( n14446 , n14443 , n334305 );
not ( n334307 , n334301 );
buf ( n14448 , n334299 );
nand ( n334309 , n334307 , n14448 );
nand ( n14450 , n14446 , n334309 );
not ( n14451 , n14450 );
nor ( n334312 , n579 , n14128 );
not ( n334313 , n334312 );
and ( n334314 , n334302 , n334313 );
not ( n14455 , n581 );
not ( n334316 , n14455 );
not ( n334317 , n333998 );
not ( n14458 , n334317 );
or ( n334319 , n334316 , n14458 );
nand ( n334320 , n13610 , n13819 );
nand ( n14461 , n333993 , n13670 , n14024 );
nand ( n334322 , n334320 , n14461 , n13677 );
not ( n334323 , n333502 );
not ( n334324 , n334323 );
not ( n14465 , n333489 );
not ( n334326 , n14465 );
or ( n14467 , n334324 , n334326 );
nand ( n14468 , n14467 , n13674 );
not ( n334329 , n14468 );
and ( n334330 , n334322 , n334329 );
not ( n334331 , n334322 );
and ( n14472 , n334331 , n14468 );
nor ( n334333 , n334330 , n14472 );
not ( n334334 , n334333 );
not ( n14475 , n580 );
nand ( n334336 , n334334 , n14475 );
nand ( n334337 , n334319 , n334336 );
not ( n14478 , n13602 );
nand ( n334339 , n14478 , n13591 );
not ( n334340 , n334339 );
not ( n14481 , n13871 );
not ( n334342 , n333863 );
or ( n14483 , n14481 , n334342 );
nand ( n334344 , n14483 , n14023 );
not ( n14485 , n334344 );
or ( n14486 , n334340 , n14485 );
buf ( n334347 , n333463 );
nand ( n334348 , n14486 , n334347 );
or ( n334349 , n13608 , n13607 );
not ( n14490 , n334349 );
not ( n334351 , n333469 );
nor ( n334352 , n14490 , n334351 );
and ( n14493 , n334348 , n334352 );
not ( n334354 , n334348 );
nand ( n334355 , n334349 , n333469 );
and ( n14496 , n334354 , n334355 );
nor ( n334357 , n14493 , n14496 );
nor ( n334358 , n334357 , n582 );
and ( n14499 , n334339 , n333463 );
not ( n334360 , n14499 );
not ( n334361 , n334344 );
not ( n14502 , n334361 );
or ( n334363 , n334360 , n14502 );
not ( n334364 , n333463 );
not ( n14505 , n334339 );
or ( n14506 , n334364 , n14505 );
nand ( n14507 , n14506 , n334344 );
nand ( n14508 , n334363 , n14507 );
nand ( n334369 , n583 , n14508 );
or ( n334370 , n334358 , n334369 );
nand ( n14511 , n582 , n334357 );
nand ( n334372 , n334370 , n14511 );
not ( n334373 , n334372 );
nor ( n14514 , n334337 , n334373 );
nand ( n334375 , n333998 , n581 );
not ( n334376 , n334375 );
not ( n334377 , n334376 );
not ( n14518 , n334336 );
or ( n14519 , n334377 , n14518 );
not ( n14520 , n334334 );
nand ( n14521 , n14520 , n580 );
nand ( n14522 , n14519 , n14521 );
nor ( n334383 , n14514 , n14522 );
not ( n334384 , n333729 );
nand ( n14525 , n334384 , n13862 );
nand ( n334386 , n14525 , n14019 );
not ( n334387 , n14013 );
nand ( n14528 , n333770 , n333860 , n333792 );
nand ( n14529 , n334387 , n14528 );
nor ( n14530 , n334386 , n14529 );
not ( n14531 , n14530 );
nand ( n334392 , n14529 , n334386 );
not ( n334393 , n585 );
nand ( n14534 , n14531 , n334392 , n334393 );
buf ( n14535 , n14534 );
not ( n14536 , n14017 );
nand ( n14537 , n14536 , n333881 );
not ( n14538 , n14537 );
nand ( n334399 , n14525 , n333771 , n333862 );
nand ( n334400 , n14525 , n14013 );
nand ( n14541 , n334399 , n334400 , n14019 );
not ( n334402 , n14541 );
not ( n334403 , n334402 );
or ( n14544 , n14538 , n334403 );
nand ( n334405 , n14541 , n14536 , n333881 );
nand ( n14546 , n14544 , n334405 );
nand ( n14547 , n321199 , n14546 );
not ( n14548 , n333860 );
nand ( n14549 , n13928 , n333791 );
not ( n14550 , n14549 );
or ( n14551 , n14548 , n14550 );
nand ( n14552 , n14551 , n14007 );
not ( n14553 , n14552 );
and ( n334414 , n333770 , n14012 );
not ( n334415 , n334414 );
not ( n334416 , n334415 );
or ( n14557 , n14553 , n334416 );
not ( n334418 , n14552 );
nand ( n14559 , n334414 , n334418 );
nand ( n334420 , n14557 , n14559 );
nor ( n334421 , n334420 , n586 );
not ( n334422 , n334421 );
not ( n14563 , n333791 );
not ( n334424 , n13928 );
or ( n14565 , n14563 , n334424 );
nand ( n14566 , n14565 , n14007 );
not ( n14567 , n14566 );
nand ( n14568 , n14567 , n14001 );
nand ( n334429 , n333860 , n14566 );
nand ( n14570 , n14568 , n334429 );
not ( n334431 , n14570 );
not ( n334432 , n587 );
nand ( n14573 , n334431 , n334432 );
not ( n334434 , n588 );
not ( n14575 , n13998 );
nand ( n334436 , n14575 , n13995 );
not ( n14577 , n13989 );
not ( n14578 , n14577 );
nor ( n334439 , n14578 , n333853 );
and ( n334440 , n334436 , n334439 );
not ( n334441 , n334436 );
nand ( n14582 , n14577 , n13992 );
and ( n334443 , n334441 , n14582 );
nor ( n334444 , n334440 , n334443 );
not ( n14585 , n334444 );
nand ( n334446 , n334434 , n14585 );
xnor ( n334447 , n333825 , n333822 );
and ( n14588 , n334447 , n333848 );
not ( n334449 , n334447 );
not ( n334450 , n333848 );
and ( n14591 , n334449 , n334450 );
nor ( n334452 , n14588 , n14591 );
not ( n334453 , n334452 );
nand ( n14594 , n334453 , n328808 );
not ( n334455 , n333838 );
not ( n14596 , n334455 );
not ( n334457 , n333842 );
or ( n14598 , n14596 , n334457 );
nand ( n14599 , n14598 , n13985 );
and ( n334460 , n14599 , n591 );
xor ( n334461 , n590 , n334460 );
and ( n334462 , n334461 , n14141 );
and ( n14603 , n590 , n334460 );
or ( n334464 , n334462 , n14603 );
and ( n334465 , n14594 , n334464 );
nand ( n14606 , n334446 , n334465 );
nand ( n334467 , n334452 , n589 );
not ( n334468 , n334467 );
nand ( n14609 , n334446 , n334468 );
not ( n334470 , n14585 );
nand ( n334471 , n334470 , n588 );
nand ( n334472 , n14606 , n14609 , n334471 );
and ( n14613 , n334422 , n14573 , n334472 );
nand ( n334474 , n14535 , n14547 , n14613 );
not ( n14615 , n14534 );
not ( n334476 , n334429 );
not ( n334477 , n14568 );
or ( n14618 , n334476 , n334477 );
nand ( n14619 , n14618 , n587 );
or ( n334480 , n334421 , n14619 );
nand ( n334481 , n334420 , n586 );
nand ( n334482 , n334480 , n334481 );
not ( n14623 , n334482 );
or ( n334484 , n14615 , n14623 );
and ( n334485 , n14019 , n14525 );
and ( n14626 , n14529 , n334485 );
not ( n334487 , n14529 );
and ( n334488 , n334487 , n334386 );
nor ( n14629 , n14626 , n334488 );
nand ( n334490 , n14629 , n585 );
nand ( n334491 , n334484 , n334490 );
nand ( n14632 , n334491 , n14547 );
not ( n334493 , n14546 );
nand ( n14634 , n334493 , n584 );
nand ( n334495 , n334474 , n14632 , n14634 );
not ( n14636 , n334495 );
not ( n334497 , n14636 );
not ( n334498 , n333998 );
nand ( n14639 , n334498 , n14455 );
and ( n14640 , n334336 , n334497 , n14639 );
not ( n334501 , n334357 );
not ( n334502 , n582 );
and ( n334503 , n334501 , n334502 );
not ( n14644 , n14508 );
nand ( n334505 , n14644 , n323556 );
not ( n334506 , n334505 );
nor ( n14647 , n334503 , n334506 );
buf ( n334508 , n14647 );
nand ( n334509 , n14640 , n334508 );
nand ( n14650 , n334383 , n334509 );
nand ( n334511 , n334314 , n14650 );
nand ( n334512 , n14451 , n334511 );
not ( n14653 , n334512 );
or ( n334514 , n14432 , n14653 );
not ( n334515 , n334274 );
nand ( n14656 , n334515 , n332672 );
nand ( n334517 , n14426 , n334288 );
nand ( n334518 , n334517 , n577 );
not ( n334519 , n334518 );
and ( n334520 , n14656 , n334519 );
nor ( n14661 , n334515 , n332672 );
nor ( n334522 , n334520 , n14661 );
nand ( n14663 , n334514 , n334522 );
not ( n14664 , n14663 );
buf ( n14665 , n14664 );
not ( n14666 , n14665 );
nand ( n14667 , n334260 , n14666 );
not ( n14668 , n14667 );
nand ( n14669 , n334061 , n14330 , n334249 , n14668 );
nand ( n14670 , n14669 , n14100 );
not ( n334531 , n14670 );
not ( n14672 , n14100 );
not ( n14673 , n14672 );
not ( n14674 , n14669 );
not ( n14675 , n14674 );
or ( n334536 , n14673 , n14675 );
nand ( n334537 , n334536 , n14670 );
not ( n14678 , n14665 );
nand ( n14679 , n14271 , n14294 );
not ( n14680 , n14679 );
nand ( n14681 , n14325 , n14313 );
not ( n14682 , n14242 );
not ( n334543 , n14245 );
or ( n334544 , n14682 , n334543 );
nand ( n14685 , n334544 , n14254 );
nor ( n334546 , n14681 , n14685 );
nand ( n334547 , n14678 , n14680 , n334546 );
buf ( n14688 , n14283 );
buf ( n14689 , n14688 );
not ( n14690 , n14689 );
and ( n14691 , n334547 , n14690 );
not ( n14692 , n334547 );
and ( n334553 , n14692 , n14689 );
nor ( n334554 , n14691 , n334553 );
buf ( n14695 , n334554 );
not ( n334556 , n14664 );
not ( n14697 , n14685 );
buf ( n14698 , n14325 );
nand ( n14699 , n334556 , n14697 , n14698 );
not ( n14700 , n14699 );
buf ( n334561 , n14313 );
buf ( n334562 , n334561 );
not ( n14703 , n334562 );
buf ( n334564 , n14703 );
nand ( n14705 , n14700 , n334564 );
buf ( n14706 , n333977 );
nand ( n334567 , n14706 , n14678 );
not ( n14708 , n334567 );
nand ( n14709 , n14708 , n14329 );
nand ( n14710 , n334232 , n14666 );
nor ( n14711 , n14665 , n14328 );
and ( n14712 , n14381 , n14382 );
not ( n14713 , n14381 );
and ( n334574 , n14713 , n14385 );
nor ( n14715 , n14712 , n334574 );
not ( n334576 , n14715 );
not ( n14717 , n14666 );
nor ( n334578 , n334576 , n14717 );
not ( n334579 , n14665 );
not ( n14720 , n14717 );
not ( n14721 , n334312 );
nand ( n14722 , n14129 , n579 );
and ( n14723 , n14721 , n14722 );
and ( n334584 , n14650 , n14723 );
not ( n334585 , n14650 );
not ( n14726 , n14723 );
and ( n334587 , n334585 , n14726 );
nor ( n334588 , n334584 , n334587 );
nand ( n14729 , n14647 , n14639 , n334497 );
nand ( n334590 , n334422 , n334481 );
not ( n334591 , n334472 );
not ( n14732 , n14573 );
or ( n334593 , n334591 , n14732 );
nand ( n14734 , n334593 , n14619 );
nand ( n14735 , n334590 , n14734 );
nand ( n334596 , n14573 , n14619 );
nand ( n14737 , n334472 , n334596 );
nor ( n334598 , n334465 , n334468 );
nand ( n14739 , n334471 , n334446 , n334598 );
not ( n14740 , n334598 );
nand ( n14741 , n14594 , n334467 );
not ( n14742 , n334464 );
and ( n14743 , n14741 , n14742 );
not ( n14744 , n14741 );
and ( n14745 , n14744 , n334464 );
nor ( n14746 , n14743 , n14745 );
xor ( n14747 , n590 , n334460 );
xor ( n14748 , n14747 , n14141 );
buf ( n14749 , n14748 );
nor ( n334610 , n14514 , n14522 );
not ( n14751 , n334610 );
buf ( n334612 , n14751 );
not ( n14753 , n334491 );
nand ( n334614 , n334372 , n14639 );
nor ( n334615 , n14706 , n14272 );
nor ( n14756 , n14681 , n14255 );
and ( n334617 , n333977 , n14756 );
buf ( n334618 , n334617 );
nand ( n14759 , n14688 , n14233 );
not ( n334620 , n14759 );
nand ( n14761 , n334620 , n14680 );
nor ( n14762 , n14761 , n334576 );
not ( n334623 , n14272 );
buf ( n14764 , n334302 );
nand ( n334625 , n14764 , n334309 );
not ( n14766 , n334625 );
not ( n14767 , n334290 );
and ( n14768 , n14767 , n334518 );
not ( n334629 , n14768 );
nand ( n334630 , n334471 , n334446 );
nor ( n14771 , n14759 , n14679 );
nor ( n334632 , n14681 , n14685 );
buf ( n334633 , n14214 );
not ( n14774 , n334376 );
or ( n334635 , n334472 , n334596 );
nand ( n14776 , n334635 , n14737 );
buf ( n334637 , n332492 );
buf ( n334638 , n332539 );
and ( n14779 , n581 , n582 );
not ( n14780 , n581 );
and ( n14781 , n14780 , n323949 );
nor ( n14782 , n14779 , n14781 );
buf ( n334643 , n14782 );
buf ( n334644 , n334643 );
not ( n14785 , n334644 );
not ( n334646 , n14294 );
not ( n334647 , n334646 );
buf ( n334648 , n580 );
not ( n14789 , n334648 );
buf ( n334650 , n14789 );
and ( n14791 , n334647 , n334650 );
not ( n14792 , n334647 );
and ( n334653 , n14792 , n580 );
or ( n334654 , n14791 , n334653 );
buf ( n334655 , n334654 );
not ( n14796 , n334655 );
or ( n334657 , n14785 , n14796 );
buf ( n334658 , n580 );
not ( n14799 , n334658 );
buf ( n334660 , n334561 );
not ( n334661 , n334660 );
buf ( n334662 , n334661 );
buf ( n334663 , n334662 );
not ( n334664 , n334663 );
or ( n14805 , n14799 , n334664 );
buf ( n334666 , n334561 );
buf ( n334667 , n334650 );
nand ( n14808 , n334666 , n334667 );
buf ( n334669 , n14808 );
buf ( n334670 , n334669 );
nand ( n334671 , n14805 , n334670 );
buf ( n334672 , n334671 );
buf ( n334673 , n334672 );
buf ( n334674 , n580 );
buf ( n334675 , n581 );
nor ( n14816 , n334674 , n334675 );
buf ( n14817 , n14816 );
not ( n334678 , n14817 );
and ( n14819 , n580 , n581 );
nor ( n334680 , n14819 , n14782 );
nand ( n334681 , n334678 , n334680 );
not ( n14822 , n334681 );
buf ( n334683 , n14822 );
nand ( n14824 , n334673 , n334683 );
buf ( n334685 , n14824 );
buf ( n334686 , n334685 );
nand ( n334687 , n334657 , n334686 );
buf ( n334688 , n334687 );
buf ( n334689 , n334688 );
buf ( n334690 , n583 );
buf ( n334691 , n584 );
xor ( n14832 , n334690 , n334691 );
buf ( n334693 , n14832 );
buf ( n334694 , n334693 );
buf ( n334695 , n334694 );
not ( n334696 , n334695 );
not ( n14837 , n14688 );
and ( n14838 , n14837 , n582 );
not ( n14839 , n14837 );
buf ( n334700 , n582 );
not ( n334701 , n334700 );
buf ( n334702 , n334701 );
and ( n334703 , n14839 , n334702 );
or ( n14844 , n14838 , n334703 );
buf ( n14845 , n14844 );
not ( n14846 , n14845 );
or ( n14847 , n334696 , n14846 );
buf ( n334708 , n582 );
buf ( n334709 , n14271 );
buf ( n334710 , n334709 );
and ( n334711 , n334708 , n334710 );
not ( n334712 , n334708 );
buf ( n334713 , n334709 );
not ( n334714 , n334713 );
buf ( n334715 , n334714 );
buf ( n334716 , n334715 );
and ( n334717 , n334712 , n334716 );
nor ( n14858 , n334711 , n334717 );
buf ( n334719 , n14858 );
buf ( n14860 , n334719 );
and ( n14861 , n582 , n583 );
buf ( n334722 , n582 );
buf ( n334723 , n583 );
nor ( n334724 , n334722 , n334723 );
buf ( n334725 , n334724 );
nor ( n14866 , n14861 , n334725 , n334694 );
buf ( n334727 , n14866 );
buf ( n334728 , n334727 );
nand ( n334729 , n14860 , n334728 );
buf ( n334730 , n334729 );
buf ( n334731 , n334730 );
nand ( n14872 , n14847 , n334731 );
buf ( n334733 , n14872 );
buf ( n334734 , n334733 );
xor ( n334735 , n334689 , n334734 );
buf ( n334736 , n334517 );
not ( n14877 , n334736 );
not ( n334738 , n14877 );
buf ( n334739 , n334738 );
buf ( n334740 , n576 );
and ( n334741 , n334739 , n334740 );
buf ( n334742 , n334741 );
buf ( n334743 , n334742 );
and ( n334744 , n577 , n578 );
not ( n14885 , n577 );
buf ( n334746 , n578 );
not ( n14887 , n334746 );
buf ( n334748 , n14887 );
and ( n14889 , n14885 , n334748 );
or ( n14890 , n334744 , n14889 );
not ( n14891 , n14890 );
buf ( n334752 , n14891 );
not ( n334753 , n334752 );
buf ( n334754 , n576 );
not ( n334755 , n334754 );
not ( n14896 , n14253 );
not ( n14897 , n14896 );
not ( n14898 , n14897 );
buf ( n334759 , n14898 );
not ( n14900 , n334759 );
or ( n334761 , n334755 , n14900 );
buf ( n334762 , n14254 );
buf ( n334763 , n332672 );
nand ( n14904 , n334762 , n334763 );
buf ( n334765 , n14904 );
buf ( n334766 , n334765 );
nand ( n14907 , n334761 , n334766 );
buf ( n334768 , n14907 );
buf ( n334769 , n334768 );
not ( n14910 , n334769 );
or ( n14911 , n334753 , n14910 );
buf ( n334772 , n576 );
not ( n14913 , n334515 );
buf ( n334774 , n14913 );
xor ( n14915 , n334772 , n334774 );
buf ( n334776 , n14915 );
buf ( n334777 , n334776 );
buf ( n334778 , n577 );
buf ( n334779 , n576 );
and ( n334780 , n334778 , n334779 );
not ( n14921 , n334778 );
buf ( n334782 , n332672 );
and ( n14923 , n14921 , n334782 );
nor ( n14924 , n334780 , n14923 );
buf ( n334785 , n14924 );
and ( n334786 , n14890 , n334785 );
buf ( n334787 , n334786 );
nand ( n14928 , n334777 , n334787 );
buf ( n334789 , n14928 );
buf ( n334790 , n334789 );
nand ( n334791 , n14911 , n334790 );
buf ( n334792 , n334791 );
buf ( n334793 , n334792 );
xor ( n14934 , n334743 , n334793 );
buf ( n334795 , n578 );
buf ( n334796 , n579 );
and ( n14937 , n334795 , n334796 );
and ( n14938 , n579 , n580 );
not ( n14939 , n579 );
and ( n334800 , n14939 , n5821 );
nor ( n14941 , n14938 , n334800 );
buf ( n334802 , n14941 );
buf ( n334803 , n578 );
buf ( n334804 , n579 );
nor ( n334805 , n334803 , n334804 );
buf ( n334806 , n334805 );
buf ( n334807 , n334806 );
nor ( n14948 , n14937 , n334802 , n334807 );
buf ( n14949 , n14948 );
buf ( n334810 , n14949 );
not ( n14951 , n334810 );
buf ( n334812 , n578 );
not ( n334813 , n334812 );
and ( n14954 , n14239 , n14241 );
not ( n334815 , n14239 );
and ( n14956 , n334815 , n14240 );
nor ( n14957 , n14954 , n14956 );
not ( n14958 , n14957 );
buf ( n334819 , n14958 );
not ( n14960 , n334819 );
buf ( n334821 , n14960 );
buf ( n334822 , n334821 );
not ( n14963 , n334822 );
or ( n334824 , n334813 , n14963 );
buf ( n334825 , n14958 );
buf ( n334826 , n334748 );
nand ( n334827 , n334825 , n334826 );
buf ( n334828 , n334827 );
buf ( n334829 , n334828 );
nand ( n14970 , n334824 , n334829 );
buf ( n14971 , n14970 );
buf ( n334832 , n14971 );
not ( n14973 , n334832 );
or ( n334834 , n14951 , n14973 );
buf ( n334835 , n578 );
not ( n14976 , n334835 );
not ( n334837 , n14698 );
buf ( n334838 , n334837 );
not ( n14979 , n334838 );
or ( n14980 , n14976 , n14979 );
buf ( n334841 , n14698 );
buf ( n334842 , n334748 );
nand ( n334843 , n334841 , n334842 );
buf ( n334844 , n334843 );
buf ( n334845 , n334844 );
nand ( n334846 , n14980 , n334845 );
buf ( n334847 , n334846 );
buf ( n334848 , n334847 );
not ( n14989 , n14941 );
not ( n334850 , n14989 );
buf ( n334851 , n334850 );
nand ( n334852 , n334848 , n334851 );
buf ( n334853 , n334852 );
buf ( n334854 , n334853 );
nand ( n14995 , n334834 , n334854 );
buf ( n334856 , n14995 );
buf ( n334857 , n334856 );
xor ( n334858 , n14934 , n334857 );
buf ( n334859 , n334858 );
buf ( n334860 , n334859 );
xor ( n334861 , n334735 , n334860 );
buf ( n334862 , n334861 );
buf ( n334863 , n334862 );
and ( n334864 , n585 , n586 );
not ( n334865 , n585 );
and ( n15006 , n334865 , n325557 );
nor ( n334867 , n334864 , n15006 );
buf ( n334868 , n334867 );
not ( n15009 , n334868 );
buf ( n334870 , n584 );
not ( n15011 , n334870 );
buf ( n15012 , n14233 );
not ( n334873 , n15012 );
buf ( n334874 , n334873 );
not ( n334875 , n334874 );
or ( n15016 , n15011 , n334875 );
buf ( n334877 , n584 );
not ( n334878 , n334877 );
buf ( n334879 , n334878 );
nand ( n334880 , n15012 , n334879 );
buf ( n334881 , n334880 );
nand ( n334882 , n15016 , n334881 );
buf ( n334883 , n334882 );
not ( n334884 , n334883 );
or ( n334885 , n15009 , n334884 );
buf ( n334886 , n584 );
not ( n334887 , n334886 );
buf ( n15028 , n14688 );
not ( n334889 , n15028 );
buf ( n334890 , n334889 );
buf ( n334891 , n334890 );
not ( n334892 , n334891 );
or ( n334893 , n334887 , n334892 );
buf ( n334894 , n334890 );
not ( n334895 , n334894 );
buf ( n334896 , n334895 );
buf ( n334897 , n334896 );
buf ( n334898 , n334879 );
nand ( n15039 , n334897 , n334898 );
buf ( n334900 , n15039 );
buf ( n334901 , n334900 );
nand ( n334902 , n334893 , n334901 );
buf ( n334903 , n334902 );
buf ( n334904 , n584 );
buf ( n334905 , n585 );
and ( n334906 , n334904 , n334905 );
buf ( n334907 , n334867 );
buf ( n334908 , n584 );
buf ( n334909 , n585 );
nor ( n15050 , n334908 , n334909 );
buf ( n334911 , n15050 );
buf ( n334912 , n334911 );
nor ( n334913 , n334906 , n334907 , n334912 );
buf ( n334914 , n334913 );
buf ( n334915 , n334914 );
buf ( n334916 , n334915 );
buf ( n334917 , n334916 );
nand ( n15058 , n334903 , n334917 );
nand ( n15059 , n334885 , n15058 );
buf ( n334920 , n15059 );
not ( n15061 , n14822 );
buf ( n334922 , n580 );
not ( n334923 , n334922 );
buf ( n334924 , n334837 );
not ( n334925 , n334924 );
or ( n15066 , n334923 , n334925 );
buf ( n334927 , n14698 );
buf ( n334928 , n334650 );
nand ( n15069 , n334927 , n334928 );
buf ( n334930 , n15069 );
buf ( n334931 , n334930 );
nand ( n15072 , n15066 , n334931 );
buf ( n334933 , n15072 );
not ( n15074 , n334933 );
or ( n334935 , n15061 , n15074 );
buf ( n334936 , n334672 );
buf ( n334937 , n334643 );
nand ( n15078 , n334936 , n334937 );
buf ( n334939 , n15078 );
nand ( n15080 , n334935 , n334939 );
not ( n15081 , n15080 );
not ( n15082 , n14891 );
not ( n15083 , n334776 );
or ( n15084 , n15082 , n15083 );
and ( n15085 , n334736 , n332672 );
not ( n15086 , n334736 );
and ( n15087 , n15086 , n576 );
or ( n15088 , n15085 , n15087 );
buf ( n334949 , n15088 );
buf ( n334950 , n334786 );
nand ( n15091 , n334949 , n334950 );
buf ( n334952 , n15091 );
nand ( n15093 , n15084 , n334952 );
not ( n15094 , n15093 );
not ( n15095 , n14448 );
not ( n15096 , n15095 );
nand ( n15097 , n15096 , n576 );
not ( n15098 , n15097 );
and ( n15099 , n15094 , n15098 );
and ( n15100 , n15093 , n15097 );
nor ( n15101 , n15099 , n15100 );
not ( n15102 , n15101 );
or ( n15103 , n15081 , n15102 );
or ( n15104 , n15101 , n15080 );
nand ( n15105 , n15103 , n15104 );
buf ( n334966 , n15105 );
xor ( n15107 , n334920 , n334966 );
and ( n15108 , n587 , n588 );
not ( n15109 , n587 );
buf ( n334970 , n588 );
not ( n15111 , n334970 );
buf ( n334972 , n15111 );
and ( n15113 , n15109 , n334972 );
nor ( n15114 , n15108 , n15113 );
buf ( n15115 , n15114 );
buf ( n334976 , n15115 );
buf ( n15117 , n334976 );
buf ( n334978 , n15117 );
not ( n15119 , n334978 );
buf ( n334980 , n586 );
not ( n15121 , n334980 );
buf ( n334982 , n15121 );
not ( n15123 , n334982 );
not ( n15124 , n14202 );
not ( n15125 , n14208 );
or ( n15126 , n15124 , n15125 );
nand ( n15127 , n15126 , n334072 );
not ( n15128 , n15127 );
buf ( n15129 , n15128 );
buf ( n334990 , n15129 );
not ( n15131 , n334990 );
buf ( n334992 , n15131 );
not ( n15133 , n334992 );
or ( n15134 , n15123 , n15133 );
nand ( n15135 , n15129 , n586 );
nand ( n15136 , n15134 , n15135 );
not ( n15137 , n15136 );
or ( n15138 , n15119 , n15137 );
buf ( n334999 , n586 );
not ( n15140 , n334999 );
buf ( n335001 , n333978 );
not ( n15142 , n335001 );
buf ( n335003 , n15142 );
buf ( n335004 , n335003 );
not ( n15145 , n335004 );
or ( n15146 , n15140 , n15145 );
buf ( n335007 , n333978 );
buf ( n335008 , n334982 );
nand ( n15149 , n335007 , n335008 );
buf ( n335010 , n15149 );
buf ( n335011 , n335010 );
nand ( n15152 , n15146 , n335011 );
buf ( n335013 , n15152 );
buf ( n335014 , n335013 );
not ( n15155 , n15114 );
and ( n15156 , n586 , n587 );
buf ( n335017 , n586 );
buf ( n335018 , n587 );
nor ( n15159 , n335017 , n335018 );
buf ( n335020 , n15159 );
nor ( n15161 , n15156 , n335020 );
and ( n15162 , n15155 , n15161 );
buf ( n15163 , n15162 );
buf ( n15164 , n15163 );
buf ( n335025 , n15164 );
nand ( n15166 , n335014 , n335025 );
buf ( n335027 , n15166 );
nand ( n15168 , n15138 , n335027 );
buf ( n335029 , n15168 );
and ( n15170 , n15107 , n335029 );
and ( n15171 , n334920 , n334966 );
or ( n15172 , n15170 , n15171 );
buf ( n335033 , n15172 );
buf ( n335034 , n335033 );
buf ( n15175 , n335034 );
buf ( n335036 , n15175 );
buf ( n335037 , n335036 );
xor ( n15178 , n334863 , n335037 );
not ( n15179 , n15093 );
nand ( n15180 , n15179 , n15097 );
not ( n15181 , n15180 );
not ( n15182 , n15080 );
or ( n15183 , n15181 , n15182 );
not ( n15184 , n15097 );
nand ( n15185 , n15184 , n15093 );
nand ( n15186 , n15183 , n15185 );
buf ( n335047 , n15186 );
buf ( n335048 , n334868 );
not ( n15189 , n335048 );
buf ( n335050 , n584 );
not ( n15191 , n335050 );
buf ( n335052 , n335003 );
not ( n15193 , n335052 );
or ( n15194 , n15191 , n15193 );
buf ( n335055 , n333978 );
buf ( n335056 , n334879 );
nand ( n15197 , n335055 , n335056 );
buf ( n335058 , n15197 );
buf ( n335059 , n335058 );
nand ( n15200 , n15194 , n335059 );
buf ( n335061 , n15200 );
buf ( n335062 , n335061 );
not ( n15203 , n335062 );
or ( n15204 , n15189 , n15203 );
buf ( n335065 , n334883 );
buf ( n335066 , n334917 );
nand ( n15207 , n335065 , n335066 );
buf ( n335068 , n15207 );
buf ( n335069 , n335068 );
nand ( n15210 , n15204 , n335069 );
buf ( n335071 , n15210 );
buf ( n335072 , n335071 );
xor ( n15213 , n335047 , n335072 );
not ( n15214 , n15164 );
not ( n15215 , n15136 );
or ( n15216 , n15214 , n15215 );
buf ( n15217 , n14715 );
and ( n15218 , n15217 , n334982 );
not ( n15219 , n15217 );
and ( n15220 , n15219 , n586 );
or ( n15221 , n15218 , n15220 );
nand ( n15222 , n15221 , n334978 );
nand ( n15223 , n15216 , n15222 );
buf ( n335084 , n15223 );
xor ( n15225 , n15213 , n335084 );
buf ( n335086 , n15225 );
buf ( n335087 , n335086 );
buf ( n15228 , n335087 );
buf ( n335089 , n15228 );
buf ( n335090 , n335089 );
xor ( n15231 , n15178 , n335090 );
buf ( n335092 , n15231 );
and ( n15233 , n589 , n590 );
not ( n15234 , n589 );
buf ( n335095 , n590 );
not ( n15236 , n335095 );
buf ( n335097 , n15236 );
and ( n15238 , n15234 , n335097 );
or ( n15239 , n15233 , n15238 );
buf ( n335100 , n15239 );
buf ( n335101 , n589 );
buf ( n335102 , n588 );
and ( n15243 , n335101 , n335102 );
not ( n15244 , n335101 );
buf ( n335105 , n334972 );
and ( n15246 , n15244 , n335105 );
nor ( n15247 , n15243 , n15246 );
buf ( n335108 , n15247 );
buf ( n335109 , n335108 );
nand ( n15250 , n335100 , n335109 );
buf ( n335111 , n15250 );
buf ( n335112 , n335111 );
not ( n15253 , n335112 );
buf ( n335114 , n15253 );
buf ( n335115 , n335114 );
not ( n15256 , n335115 );
not ( n15257 , n334972 );
buf ( n15258 , n15127 );
buf ( n335119 , n15258 );
buf ( n15260 , n335119 );
buf ( n335121 , n15260 );
not ( n15262 , n335121 );
or ( n15263 , n15257 , n15262 );
not ( n15264 , n15258 );
buf ( n335125 , n15264 );
buf ( n335126 , n588 );
nand ( n15267 , n335125 , n335126 );
buf ( n335128 , n15267 );
nand ( n15269 , n15263 , n335128 );
buf ( n335130 , n15269 );
not ( n15271 , n335130 );
or ( n15272 , n15256 , n15271 );
xor ( n15273 , n588 , n15217 );
buf ( n335134 , n15273 );
not ( n15275 , n15239 );
buf ( n335136 , n15275 );
nand ( n15277 , n335134 , n335136 );
buf ( n335138 , n15277 );
buf ( n335139 , n335138 );
nand ( n15280 , n15272 , n335139 );
buf ( n335141 , n15280 );
buf ( n335142 , n335141 );
not ( n15283 , n335142 );
buf ( n335144 , n591 );
not ( n15285 , n335144 );
not ( n15286 , n334257 );
not ( n15287 , n334256 );
or ( n15288 , n15286 , n15287 );
nand ( n15289 , n15288 , n14394 );
buf ( n15290 , n15289 );
and ( n15291 , n15290 , n335097 );
not ( n15292 , n15290 );
and ( n15293 , n15292 , n590 );
or ( n15294 , n15291 , n15293 );
buf ( n335155 , n15294 );
not ( n15296 , n335155 );
or ( n15297 , n15285 , n15296 );
buf ( n335158 , n590 );
not ( n15299 , n335158 );
buf ( n15300 , n334232 );
buf ( n335161 , n15300 );
not ( n15302 , n335161 );
buf ( n335163 , n15302 );
buf ( n335164 , n335163 );
not ( n15305 , n335164 );
or ( n15306 , n15299 , n15305 );
buf ( n335167 , n15300 );
buf ( n335168 , n335097 );
nand ( n15309 , n335167 , n335168 );
buf ( n335170 , n15309 );
buf ( n335171 , n335170 );
nand ( n15312 , n15306 , n335171 );
buf ( n335173 , n15312 );
buf ( n335174 , n335173 );
buf ( n335175 , n591 );
not ( n15316 , n335175 );
buf ( n335177 , n15316 );
buf ( n335178 , n335177 );
buf ( n335179 , n590 );
and ( n15320 , n335178 , n335179 );
buf ( n335181 , n15320 );
buf ( n15322 , n335181 );
nand ( n15323 , n335174 , n15322 );
buf ( n15324 , n15323 );
buf ( n335185 , n15324 );
nand ( n15326 , n15297 , n335185 );
buf ( n335187 , n15326 );
buf ( n335188 , n335187 );
not ( n15329 , n335188 );
or ( n15330 , n15283 , n15329 );
buf ( n335191 , n335141 );
buf ( n335192 , n335187 );
or ( n15333 , n335191 , n335192 );
buf ( n335194 , n334978 );
not ( n15335 , n335194 );
buf ( n335196 , n335013 );
not ( n15337 , n335196 );
or ( n335198 , n15335 , n15337 );
buf ( n335199 , n15164 );
not ( n15340 , n334982 );
buf ( n15341 , n15012 );
not ( n15342 , n15341 );
or ( n335203 , n15340 , n15342 );
nand ( n335204 , n334873 , n586 );
nand ( n335205 , n335203 , n335204 );
buf ( n335206 , n335205 );
nand ( n335207 , n335199 , n335206 );
buf ( n335208 , n335207 );
buf ( n335209 , n335208 );
nand ( n15350 , n335198 , n335209 );
buf ( n335211 , n15350 );
buf ( n335212 , n335211 );
nand ( n15353 , n15333 , n335212 );
buf ( n335214 , n15353 );
buf ( n335215 , n335214 );
nand ( n15356 , n15330 , n335215 );
buf ( n335217 , n15356 );
buf ( n335218 , n334868 );
not ( n335219 , n335218 );
buf ( n335220 , n584 );
not ( n15361 , n335220 );
buf ( n335222 , n334715 );
not ( n335223 , n335222 );
or ( n15364 , n15361 , n335223 );
buf ( n15365 , n334709 );
buf ( n15366 , n334879 );
nand ( n15367 , n15365 , n15366 );
buf ( n15368 , n15367 );
buf ( n335229 , n15368 );
nand ( n335230 , n15364 , n335229 );
buf ( n335231 , n335230 );
buf ( n15372 , n335231 );
not ( n15373 , n15372 );
or ( n15374 , n335219 , n15373 );
buf ( n335235 , n584 );
not ( n335236 , n335235 );
buf ( n335237 , n334646 );
buf ( n335238 , n335237 );
not ( n335239 , n335238 );
or ( n335240 , n335236 , n335239 );
not ( n15381 , n334646 );
buf ( n335242 , n15381 );
buf ( n335243 , n334879 );
nand ( n15384 , n335242 , n335243 );
buf ( n15385 , n15384 );
buf ( n335246 , n15385 );
nand ( n15387 , n335240 , n335246 );
buf ( n335248 , n15387 );
buf ( n335249 , n335248 );
buf ( n335250 , n334917 );
nand ( n15391 , n335249 , n335250 );
buf ( n335252 , n15391 );
buf ( n335253 , n335252 );
nand ( n335254 , n15374 , n335253 );
buf ( n335255 , n335254 );
buf ( n335256 , n335255 );
buf ( n335257 , n334727 );
not ( n335258 , n335257 );
buf ( n335259 , n582 );
not ( n335260 , n335259 );
not ( n335261 , n14698 );
buf ( n335262 , n335261 );
not ( n335263 , n335262 );
or ( n335264 , n335260 , n335263 );
buf ( n335265 , n14698 );
buf ( n335266 , n334702 );
nand ( n335267 , n335265 , n335266 );
buf ( n335268 , n335267 );
buf ( n335269 , n335268 );
nand ( n335270 , n335264 , n335269 );
buf ( n335271 , n335270 );
buf ( n15412 , n335271 );
not ( n15413 , n15412 );
or ( n15414 , n335258 , n15413 );
buf ( n335275 , n582 );
not ( n335276 , n335275 );
buf ( n335277 , n334564 );
not ( n15418 , n335277 );
or ( n335279 , n335276 , n15418 );
buf ( n335280 , n334662 );
not ( n15421 , n335280 );
buf ( n335282 , n334702 );
nand ( n335283 , n15421 , n335282 );
buf ( n335284 , n335283 );
buf ( n335285 , n335284 );
nand ( n335286 , n335279 , n335285 );
buf ( n335287 , n335286 );
buf ( n335288 , n335287 );
buf ( n335289 , n334694 );
nand ( n15430 , n335288 , n335289 );
buf ( n335291 , n15430 );
buf ( n335292 , n335291 );
nand ( n335293 , n15414 , n335292 );
buf ( n335294 , n335293 );
buf ( n335295 , n335294 );
or ( n335296 , n335256 , n335295 );
buf ( n335297 , n335296 );
not ( n15438 , n14891 );
not ( n15439 , n576 );
buf ( n335300 , n334333 );
not ( n335301 , n335300 );
not ( n15442 , n335301 );
or ( n15443 , n15439 , n15442 );
or ( n335304 , n335301 , n576 );
nand ( n335305 , n15443 , n335304 );
not ( n335306 , n335305 );
or ( n335307 , n15438 , n335306 );
buf ( n335308 , n14139 );
not ( n335309 , n335308 );
buf ( n335310 , n335309 );
buf ( n335311 , n335310 );
not ( n15452 , n335311 );
buf ( n335313 , n15452 );
xor ( n335314 , n576 , n335313 );
nand ( n15455 , n335314 , n334786 );
nand ( n15456 , n335307 , n15455 );
not ( n15457 , n15456 );
not ( n15458 , n15457 );
and ( n15459 , n334348 , n334352 );
not ( n15460 , n334348 );
and ( n335321 , n15460 , n334355 );
nor ( n15462 , n15459 , n335321 );
buf ( n15463 , n15462 );
buf ( n335324 , n15463 );
not ( n335325 , n335324 );
buf ( n335326 , n335325 );
buf ( n335327 , n335326 );
buf ( n15468 , n335327 );
buf ( n335329 , n15468 );
or ( n15470 , n335329 , n332672 );
not ( n15471 , n15470 );
and ( n335332 , n15458 , n15471 );
not ( n335333 , n15456 );
nand ( n15474 , n335333 , n15470 );
not ( n335335 , n14941 );
buf ( n335336 , n578 );
not ( n15477 , n335336 );
buf ( n335338 , n15095 );
not ( n15479 , n335338 );
or ( n15480 , n15477 , n15479 );
buf ( n15481 , n14448 );
buf ( n335342 , n15481 );
buf ( n335343 , n334748 );
nand ( n335344 , n335342 , n335343 );
buf ( n335345 , n335344 );
buf ( n335346 , n335345 );
nand ( n335347 , n15480 , n335346 );
buf ( n335348 , n335347 );
not ( n15489 , n335348 );
or ( n15490 , n335335 , n15489 );
buf ( n335351 , n578 );
not ( n15492 , n335351 );
buf ( n335353 , n14129 );
not ( n15494 , n335353 );
buf ( n335355 , n15494 );
buf ( n335356 , n335355 );
not ( n15497 , n335356 );
or ( n15498 , n15492 , n15497 );
buf ( n335359 , n14129 );
buf ( n335360 , n335359 );
buf ( n335361 , n335360 );
buf ( n335362 , n335361 );
buf ( n335363 , n334748 );
nand ( n15504 , n335362 , n335363 );
buf ( n335365 , n15504 );
buf ( n335366 , n335365 );
nand ( n15507 , n15498 , n335366 );
buf ( n335368 , n15507 );
buf ( n335369 , n335368 );
buf ( n335370 , n14949 );
nand ( n335371 , n335369 , n335370 );
buf ( n335372 , n335371 );
nand ( n15513 , n15490 , n335372 );
and ( n15514 , n15474 , n15513 );
nor ( n15515 , n335332 , n15514 );
buf ( n335376 , n580 );
not ( n15517 , n335376 );
buf ( n335378 , n14898 );
not ( n335379 , n335378 );
or ( n335380 , n15517 , n335379 );
buf ( n335381 , n14897 );
buf ( n335382 , n334650 );
nand ( n15523 , n335381 , n335382 );
buf ( n335384 , n15523 );
buf ( n335385 , n335384 );
nand ( n335386 , n335380 , n335385 );
buf ( n335387 , n335386 );
buf ( n15528 , n334643 );
and ( n335389 , n335387 , n15528 );
buf ( n335390 , n580 );
not ( n15531 , n335390 );
buf ( n335392 , n334515 );
buf ( n335393 , n335392 );
not ( n15534 , n335393 );
or ( n335395 , n15531 , n15534 );
buf ( n15536 , n14913 );
buf ( n335397 , n334650 );
nand ( n15538 , n15536 , n335397 );
buf ( n335399 , n15538 );
buf ( n335400 , n335399 );
nand ( n335401 , n335395 , n335400 );
buf ( n335402 , n335401 );
not ( n335403 , n335402 );
buf ( n335404 , n14822 );
not ( n335405 , n335404 );
buf ( n335406 , n335405 );
nor ( n15547 , n335403 , n335406 );
nor ( n335408 , n335389 , n15547 );
xor ( n335409 , n15515 , n335408 );
not ( n335410 , n14891 );
buf ( n335411 , n576 );
not ( n335412 , n335411 );
buf ( n335413 , n335355 );
not ( n15554 , n335413 );
or ( n335415 , n335412 , n15554 );
buf ( n335416 , n14129 );
buf ( n335417 , n332672 );
nand ( n335418 , n335416 , n335417 );
buf ( n335419 , n335418 );
buf ( n335420 , n335419 );
nand ( n335421 , n335415 , n335420 );
buf ( n335422 , n335421 );
not ( n15563 , n335422 );
or ( n15564 , n335410 , n15563 );
nand ( n15565 , n335305 , n334786 );
nand ( n15566 , n15564 , n15565 );
and ( n15567 , n576 , n335313 );
nor ( n15568 , n15566 , n15567 );
not ( n15569 , n15568 );
nand ( n15570 , n15566 , n15567 );
nand ( n335431 , n15569 , n15570 );
buf ( n335432 , n14941 );
not ( n15573 , n335432 );
not ( n335434 , n334517 );
not ( n335435 , n335434 );
xor ( n15576 , n578 , n335435 );
not ( n335437 , n15576 );
or ( n15578 , n15573 , n335437 );
buf ( n335439 , n14949 );
not ( n335440 , n335439 );
buf ( n335441 , n335440 );
not ( n335442 , n335441 );
nand ( n15583 , n335442 , n335348 );
nand ( n335444 , n15578 , n15583 );
xor ( n335445 , n335431 , n335444 );
and ( n15586 , n335409 , n335445 );
and ( n335447 , n15515 , n335408 );
or ( n335448 , n15586 , n335447 );
buf ( n335449 , n335448 );
not ( n335450 , n335449 );
buf ( n335451 , n335450 );
and ( n335452 , n335297 , n335451 );
and ( n15593 , n335255 , n335294 );
nor ( n335454 , n335452 , n15593 );
buf ( n335455 , n335454 );
not ( n15596 , n335455 );
buf ( n335457 , n15596 );
not ( n335458 , n335457 );
buf ( n335459 , n335300 );
buf ( n335460 , n335459 );
not ( n335461 , n335460 );
buf ( n15602 , n332672 );
nor ( n15603 , n335461 , n15602 );
buf ( n15604 , n15603 );
buf ( n335465 , n15604 );
not ( n15606 , n335465 );
xor ( n335467 , n576 , n14448 );
and ( n15608 , n14891 , n335467 );
and ( n15609 , n335422 , n334786 );
nor ( n335470 , n15608 , n15609 );
buf ( n335471 , n335470 );
nand ( n335472 , n15606 , n335471 );
buf ( n335473 , n335472 );
buf ( n335474 , n335473 );
not ( n335475 , n335474 );
not ( n335476 , n15576 );
not ( n15617 , n335476 );
not ( n15618 , n335441 );
and ( n15619 , n15617 , n15618 );
not ( n15620 , n578 );
not ( n15621 , n334515 );
not ( n15622 , n15621 );
not ( n15623 , n15622 );
or ( n335484 , n15620 , n15623 );
buf ( n335485 , n15621 );
buf ( n335486 , n334748 );
nand ( n335487 , n335485 , n335486 );
buf ( n335488 , n335487 );
nand ( n335489 , n335484 , n335488 );
and ( n335490 , n335489 , n334850 );
nor ( n15631 , n15619 , n335490 );
not ( n335492 , n15631 );
buf ( n335493 , n335492 );
not ( n15634 , n335493 );
or ( n335495 , n335475 , n15634 );
buf ( n335496 , n335470 );
not ( n335497 , n335496 );
buf ( n15638 , n15604 );
nand ( n15639 , n335497 , n15638 );
buf ( n15640 , n15639 );
buf ( n335501 , n15640 );
nand ( n15642 , n335495 , n335501 );
buf ( n335503 , n15642 );
buf ( n335504 , n335503 );
buf ( n335505 , n14822 );
not ( n15646 , n335505 );
buf ( n335507 , n580 );
not ( n15648 , n335507 );
buf ( n335509 , n334821 );
not ( n15650 , n335509 );
or ( n15651 , n15648 , n15650 );
buf ( n335512 , n14958 );
not ( n15653 , n335512 );
buf ( n335514 , n15653 );
buf ( n335515 , n335514 );
not ( n15656 , n335515 );
buf ( n335517 , n334650 );
nand ( n15658 , n15656 , n335517 );
buf ( n335519 , n15658 );
buf ( n335520 , n335519 );
nand ( n15661 , n15651 , n335520 );
buf ( n335522 , n15661 );
buf ( n335523 , n335522 );
not ( n15664 , n335523 );
or ( n15665 , n15646 , n15664 );
buf ( n335526 , n334933 );
buf ( n335527 , n15528 );
nand ( n15668 , n335526 , n335527 );
buf ( n335529 , n15668 );
buf ( n335530 , n335529 );
nand ( n15671 , n15665 , n335530 );
buf ( n335532 , n15671 );
buf ( n335533 , n335532 );
xor ( n15674 , n335504 , n335533 );
buf ( n335535 , n334694 );
not ( n15676 , n335535 );
and ( n15677 , n334647 , n334702 );
not ( n15678 , n334647 );
and ( n15679 , n15678 , n582 );
or ( n15680 , n15677 , n15679 );
buf ( n335541 , n15680 );
not ( n15682 , n335541 );
or ( n15683 , n15676 , n15682 );
buf ( n335544 , n335287 );
buf ( n335545 , n334727 );
nand ( n15686 , n335544 , n335545 );
buf ( n335547 , n15686 );
buf ( n335548 , n335547 );
nand ( n15689 , n15683 , n335548 );
buf ( n335550 , n15689 );
buf ( n335551 , n335550 );
xnor ( n15692 , n15674 , n335551 );
buf ( n335553 , n15692 );
buf ( n335554 , n335553 );
not ( n15695 , n335554 );
buf ( n335556 , n15695 );
not ( n15697 , n335556 );
or ( n15698 , n335458 , n15697 );
not ( n15699 , n335553 );
not ( n15700 , n335454 );
or ( n15701 , n15699 , n15700 );
buf ( n335562 , n335361 );
buf ( n335563 , n576 );
nand ( n15704 , n335562 , n335563 );
buf ( n335565 , n15704 );
buf ( n335566 , n335467 );
not ( n15707 , n335566 );
buf ( n335568 , n15707 );
buf ( n335569 , n335568 );
not ( n15710 , n335569 );
not ( n15711 , n334786 );
buf ( n335572 , n15711 );
not ( n15713 , n335572 );
and ( n15714 , n15710 , n15713 );
buf ( n335575 , n15088 );
buf ( n335576 , n14891 );
and ( n15717 , n335575 , n335576 );
nor ( n15718 , n15714 , n15717 );
buf ( n335579 , n15718 );
xor ( n15720 , n335565 , n335579 );
buf ( n335581 , n335489 );
not ( n15722 , n335581 );
buf ( n335583 , n15722 );
buf ( n335584 , n335583 );
not ( n15725 , n335584 );
buf ( n335586 , n335441 );
not ( n15727 , n335586 );
and ( n15728 , n15725 , n15727 );
buf ( n335589 , n334748 );
not ( n15730 , n335589 );
buf ( n335591 , n14254 );
not ( n15732 , n335591 );
or ( n15733 , n15730 , n15732 );
buf ( n335594 , n14897 );
buf ( n335595 , n334748 );
or ( n15736 , n335594 , n335595 );
nand ( n15737 , n15733 , n15736 );
buf ( n335598 , n15737 );
buf ( n335599 , n335598 );
buf ( n335600 , n335432 );
and ( n15741 , n335599 , n335600 );
nor ( n15742 , n15728 , n15741 );
buf ( n335603 , n15742 );
xnor ( n15744 , n15720 , n335603 );
buf ( n335605 , n15744 );
buf ( n335606 , n334868 );
not ( n15747 , n335606 );
buf ( n335608 , n334903 );
not ( n15749 , n335608 );
or ( n15750 , n15747 , n15749 );
buf ( n335611 , n335231 );
buf ( n335612 , n334917 );
nand ( n15753 , n335611 , n335612 );
buf ( n335614 , n15753 );
buf ( n335615 , n335614 );
nand ( n15756 , n15750 , n335615 );
buf ( n335617 , n15756 );
buf ( n335618 , n335617 );
xor ( n15759 , n335605 , n335618 );
not ( n15760 , n15568 );
not ( n15761 , n15760 );
not ( n15762 , n335444 );
or ( n15763 , n15761 , n15762 );
nand ( n15764 , n15763 , n15570 );
not ( n15765 , n15528 );
not ( n15766 , n335522 );
or ( n15767 , n15765 , n15766 );
buf ( n335628 , n335387 );
buf ( n335629 , n14822 );
nand ( n15770 , n335628 , n335629 );
buf ( n335631 , n15770 );
nand ( n15772 , n15767 , n335631 );
or ( n15773 , n15764 , n15772 );
not ( n15774 , n15604 );
not ( n15775 , n335470 );
or ( n15776 , n15774 , n15775 );
or ( n15777 , n335470 , n15604 );
nand ( n15778 , n15776 , n15777 );
not ( n15779 , n15778 );
not ( n15780 , n15779 );
not ( n15781 , n335492 );
or ( n15782 , n15780 , n15781 );
nand ( n15783 , n15778 , n15631 );
nand ( n15784 , n15782 , n15783 );
nand ( n15785 , n15773 , n15784 );
buf ( n335646 , n15785 );
nand ( n15787 , n15772 , n15764 );
buf ( n335648 , n15787 );
nand ( n15789 , n335646 , n335648 );
buf ( n335650 , n15789 );
buf ( n335651 , n335650 );
xor ( n15792 , n15759 , n335651 );
buf ( n335653 , n15792 );
nand ( n15794 , n15701 , n335653 );
nand ( n15795 , n15698 , n15794 );
xor ( n15796 , n335217 , n15795 );
buf ( n335657 , n15275 );
not ( n15798 , n335657 );
buf ( n335659 , n588 );
not ( n15800 , n335659 );
buf ( n335661 , n335163 );
not ( n15802 , n335661 );
or ( n15803 , n15800 , n15802 );
buf ( n335664 , n15300 );
buf ( n335665 , n334972 );
nand ( n15806 , n335664 , n335665 );
buf ( n335667 , n15806 );
buf ( n335668 , n335667 );
nand ( n15809 , n15803 , n335668 );
buf ( n335670 , n15809 );
buf ( n335671 , n335670 );
not ( n15812 , n335671 );
or ( n15813 , n15798 , n15812 );
buf ( n335674 , n15273 );
buf ( n335675 , n335114 );
nand ( n335676 , n335674 , n335675 );
buf ( n335677 , n335676 );
buf ( n335678 , n335677 );
nand ( n15819 , n15813 , n335678 );
buf ( n335680 , n15819 );
buf ( n15821 , n335680 );
not ( n335682 , n15821 );
buf ( n335683 , n335682 );
buf ( n335684 , n335683 );
buf ( n335685 , n335532 );
not ( n15826 , n335685 );
buf ( n335687 , n335550 );
not ( n15828 , n335687 );
or ( n335689 , n15826 , n15828 );
buf ( n335690 , n335550 );
buf ( n335691 , n335532 );
or ( n335692 , n335690 , n335691 );
buf ( n335693 , n335503 );
nand ( n15834 , n335692 , n335693 );
buf ( n335695 , n15834 );
buf ( n335696 , n335695 );
nand ( n335697 , n335689 , n335696 );
buf ( n335698 , n335697 );
buf ( n335699 , n335698 );
not ( n335700 , n335699 );
buf ( n335701 , n335700 );
buf ( n15842 , n335701 );
and ( n15843 , n335684 , n15842 );
not ( n335704 , n335684 );
buf ( n335705 , n335698 );
and ( n15846 , n335704 , n335705 );
nor ( n335707 , n15843 , n15846 );
buf ( n335708 , n335707 );
buf ( n335709 , n335708 );
buf ( n335710 , n335432 );
not ( n15851 , n335710 );
buf ( n335712 , n14971 );
not ( n15853 , n335712 );
or ( n15854 , n15851 , n15853 );
buf ( n335715 , n14949 );
buf ( n335716 , n335598 );
nand ( n335717 , n335715 , n335716 );
buf ( n335718 , n335717 );
buf ( n335719 , n335718 );
nand ( n335720 , n15854 , n335719 );
buf ( n335721 , n335720 );
buf ( n335722 , n335721 );
buf ( n335723 , n334694 );
not ( n15864 , n335723 );
buf ( n335725 , n334719 );
not ( n335726 , n335725 );
or ( n335727 , n15864 , n335726 );
buf ( n335728 , n15680 );
buf ( n335729 , n334727 );
nand ( n335730 , n335728 , n335729 );
buf ( n335731 , n335730 );
buf ( n335732 , n335731 );
nand ( n335733 , n335727 , n335732 );
buf ( n335734 , n335733 );
buf ( n335735 , n335734 );
xor ( n335736 , n335722 , n335735 );
buf ( n335737 , n335579 );
buf ( n335738 , n335565 );
nand ( n335739 , n335737 , n335738 );
buf ( n335740 , n335739 );
buf ( n335741 , n335740 );
not ( n335742 , n335741 );
buf ( n335743 , n335603 );
not ( n15884 , n335743 );
buf ( n335745 , n15884 );
buf ( n335746 , n335745 );
not ( n335747 , n335746 );
or ( n15888 , n335742 , n335747 );
or ( n335749 , n335579 , n335565 );
buf ( n335750 , n335749 );
nand ( n15891 , n15888 , n335750 );
buf ( n15892 , n15891 );
buf ( n335753 , n15892 );
xnor ( n15894 , n335736 , n335753 );
buf ( n15895 , n15894 );
buf ( n15896 , n15895 );
not ( n15897 , n15896 );
buf ( n15898 , n15897 );
buf ( n15899 , n15898 );
and ( n15900 , n335709 , n15899 );
not ( n15901 , n335709 );
buf ( n335762 , n15895 );
and ( n15903 , n15901 , n335762 );
nor ( n15904 , n15900 , n15903 );
buf ( n335765 , n15904 );
and ( n15906 , n15796 , n335765 );
and ( n335767 , n335217 , n15795 );
or ( n15908 , n15906 , n335767 );
xor ( n335769 , n335092 , n15908 );
buf ( n335770 , n335680 );
not ( n15911 , n335770 );
buf ( n335772 , n15898 );
not ( n335773 , n335772 );
or ( n15914 , n15911 , n335773 );
buf ( n335775 , n335683 );
not ( n15916 , n335775 );
buf ( n335777 , n15895 );
not ( n15918 , n335777 );
or ( n335779 , n15916 , n15918 );
buf ( n335780 , n335698 );
nand ( n15921 , n335779 , n335780 );
buf ( n335782 , n15921 );
buf ( n335783 , n335782 );
nand ( n15924 , n15914 , n335783 );
buf ( n15925 , n15924 );
buf ( n335786 , n15925 );
buf ( n335787 , n335734 );
buf ( n335788 , n335721 );
or ( n335789 , n335787 , n335788 );
buf ( n335790 , n15892 );
nand ( n15931 , n335789 , n335790 );
buf ( n15932 , n15931 );
buf ( n335793 , n15932 );
buf ( n335794 , n335734 );
buf ( n335795 , n335721 );
nand ( n15936 , n335794 , n335795 );
buf ( n335797 , n15936 );
buf ( n335798 , n335797 );
nand ( n15939 , n335793 , n335798 );
buf ( n335800 , n15939 );
buf ( n335801 , n335800 );
buf ( n335802 , n15275 );
not ( n15943 , n335802 );
buf ( n335804 , n588 );
not ( n15945 , n335804 );
buf ( n335806 , n15290 );
not ( n15947 , n335806 );
buf ( n335808 , n15947 );
buf ( n335809 , n335808 );
not ( n15950 , n335809 );
or ( n15951 , n15945 , n15950 );
buf ( n335812 , n15290 );
buf ( n335813 , n334972 );
nand ( n335814 , n335812 , n335813 );
buf ( n335815 , n335814 );
buf ( n335816 , n335815 );
nand ( n335817 , n15951 , n335816 );
buf ( n335818 , n335817 );
buf ( n335819 , n335818 );
not ( n335820 , n335819 );
or ( n335821 , n15943 , n335820 );
buf ( n335822 , n335114 );
buf ( n335823 , n335670 );
nand ( n15964 , n335822 , n335823 );
buf ( n335825 , n15964 );
buf ( n335826 , n335825 );
nand ( n335827 , n335821 , n335826 );
buf ( n335828 , n335827 );
buf ( n335829 , n335828 );
xor ( n335830 , n335801 , n335829 );
buf ( n335831 , n335181 );
not ( n15972 , n335831 );
buf ( n335833 , n590 );
not ( n335834 , n335833 );
not ( n15975 , n14199 );
buf ( n335836 , n15975 );
not ( n335837 , n335836 );
or ( n15978 , n335834 , n335837 );
buf ( n335839 , n14199 );
buf ( n335840 , n335097 );
nand ( n335841 , n335839 , n335840 );
buf ( n335842 , n335841 );
buf ( n335843 , n335842 );
nand ( n335844 , n15978 , n335843 );
buf ( n335845 , n335844 );
buf ( n335846 , n335845 );
not ( n335847 , n335846 );
or ( n335848 , n15972 , n335847 );
buf ( n335849 , n590 );
not ( n335850 , n335849 );
not ( n335851 , n14349 );
not ( n15992 , n335851 );
buf ( n335853 , n15992 );
not ( n335854 , n335853 );
or ( n335855 , n335850 , n335854 );
buf ( n335856 , n335851 );
buf ( n335857 , n335097 );
nand ( n15998 , n335856 , n335857 );
buf ( n335859 , n15998 );
buf ( n16000 , n335859 );
nand ( n16001 , n335855 , n16000 );
buf ( n16002 , n16001 );
buf ( n16003 , n16002 );
buf ( n335864 , n591 );
nand ( n335865 , n16003 , n335864 );
buf ( n335866 , n335865 );
buf ( n335867 , n335866 );
nand ( n335868 , n335848 , n335867 );
buf ( n335869 , n335868 );
buf ( n335870 , n335869 );
xor ( n335871 , n335830 , n335870 );
buf ( n335872 , n335871 );
buf ( n335873 , n335872 );
xor ( n16014 , n335786 , n335873 );
buf ( n335875 , n591 );
not ( n16016 , n335875 );
buf ( n335877 , n335845 );
not ( n335878 , n335877 );
or ( n335879 , n16016 , n335878 );
buf ( n335880 , n15294 );
buf ( n335881 , n335181 );
nand ( n335882 , n335880 , n335881 );
buf ( n335883 , n335882 );
buf ( n335884 , n335883 );
nand ( n335885 , n335879 , n335884 );
buf ( n335886 , n335885 );
buf ( n335887 , n335886 );
not ( n335888 , n335887 );
xor ( n335889 , n334920 , n334966 );
xor ( n335890 , n335889 , n335029 );
buf ( n335891 , n335890 );
buf ( n16032 , n335891 );
not ( n16033 , n16032 );
or ( n16034 , n335888 , n16033 );
buf ( n335895 , n335886 );
buf ( n335896 , n335891 );
or ( n335897 , n335895 , n335896 );
xor ( n16038 , n335605 , n335618 );
and ( n335899 , n16038 , n335651 );
and ( n335900 , n335605 , n335618 );
or ( n16041 , n335899 , n335900 );
buf ( n335902 , n16041 );
buf ( n16043 , n335902 );
nand ( n16044 , n335897 , n16043 );
buf ( n16045 , n16044 );
buf ( n335906 , n16045 );
nand ( n16047 , n16034 , n335906 );
buf ( n16048 , n16047 );
buf ( n335909 , n16048 );
xnor ( n16050 , n16014 , n335909 );
buf ( n335911 , n16050 );
buf ( n335912 , n335911 );
not ( n16053 , n335912 );
buf ( n335914 , n16053 );
and ( n335915 , n335769 , n335914 );
not ( n335916 , n335769 );
and ( n16057 , n335916 , n335911 );
nor ( n335918 , n335915 , n16057 );
not ( n335919 , n335918 );
xor ( n16060 , n335217 , n15795 );
xor ( n335921 , n16060 , n335765 );
buf ( n335922 , n335921 );
not ( n16063 , n335922 );
buf ( n335924 , n16063 );
buf ( n335925 , n335924 );
buf ( n335926 , n335902 );
buf ( n335927 , n335886 );
xor ( n335928 , n335926 , n335927 );
buf ( n335929 , n335891 );
xnor ( n335930 , n335928 , n335929 );
buf ( n335931 , n335930 );
buf ( n335932 , n335931 );
not ( n335933 , n334978 );
not ( n335934 , n335205 );
or ( n16075 , n335933 , n335934 );
nand ( n335936 , n14837 , n586 );
not ( n335937 , n335936 );
buf ( n335938 , n334896 );
buf ( n335939 , n334982 );
nand ( n335940 , n335938 , n335939 );
buf ( n335941 , n335940 );
not ( n335942 , n335941 );
or ( n335943 , n335937 , n335942 );
nand ( n16084 , n335943 , n15164 );
nand ( n335945 , n16075 , n16084 );
not ( n16086 , n335945 );
not ( n16087 , n16086 );
not ( n16088 , n15275 );
not ( n16089 , n15269 );
or ( n16090 , n16088 , n16089 );
and ( n16091 , n335003 , n588 );
not ( n16092 , n335003 );
and ( n16093 , n16092 , n334972 );
or ( n16094 , n16091 , n16093 );
buf ( n16095 , n16094 );
buf ( n335956 , n335114 );
nand ( n16097 , n16095 , n335956 );
buf ( n335958 , n16097 );
nand ( n16099 , n16090 , n335958 );
not ( n335960 , n16099 );
not ( n335961 , n335960 );
or ( n16102 , n16087 , n335961 );
xor ( n335963 , n15764 , n15784 );
xor ( n335964 , n335963 , n15772 );
buf ( n16105 , n335964 );
nand ( n335966 , n16102 , n16105 );
buf ( n16107 , n16099 );
buf ( n335968 , n335945 );
nand ( n335969 , n16107 , n335968 );
buf ( n335970 , n335969 );
nand ( n335971 , n335966 , n335970 );
not ( n335972 , n335971 );
buf ( n335973 , n335211 );
buf ( n335974 , n335141 );
xor ( n16115 , n335973 , n335974 );
buf ( n335976 , n335187 );
xnor ( n16117 , n16115 , n335976 );
buf ( n16118 , n16117 );
buf ( n335979 , n16118 );
not ( n335980 , n335979 );
buf ( n335981 , n335980 );
not ( n335982 , n335981 );
or ( n16123 , n335972 , n335982 );
buf ( n335984 , n335971 );
not ( n335985 , n335984 );
buf ( n335986 , n335985 );
not ( n335987 , n335986 );
not ( n16128 , n16118 );
or ( n16129 , n335987 , n16128 );
buf ( n335990 , n334694 );
not ( n16131 , n335990 );
buf ( n335992 , n335271 );
not ( n16133 , n335992 );
or ( n16134 , n16131 , n16133 );
buf ( n335995 , n582 );
not ( n16136 , n335995 );
buf ( n335997 , n335514 );
not ( n16138 , n335997 );
or ( n335999 , n16136 , n16138 );
buf ( n336000 , n334821 );
not ( n336001 , n336000 );
buf ( n336002 , n334702 );
nand ( n16143 , n336001 , n336002 );
buf ( n336004 , n16143 );
buf ( n336005 , n336004 );
nand ( n16146 , n335999 , n336005 );
buf ( n336007 , n16146 );
buf ( n336008 , n336007 );
buf ( n336009 , n334727 );
nand ( n16150 , n336008 , n336009 );
buf ( n16151 , n16150 );
buf ( n336012 , n16151 );
nand ( n16153 , n16134 , n336012 );
buf ( n336014 , n16153 );
buf ( n336015 , n336014 );
not ( n16156 , n336015 );
not ( n16157 , n334868 );
not ( n336018 , n335248 );
or ( n336019 , n16157 , n336018 );
buf ( n336020 , n584 );
not ( n336021 , n336020 );
buf ( n336022 , n334662 );
buf ( n16163 , n336022 );
buf ( n336024 , n16163 );
buf ( n336025 , n336024 );
not ( n16166 , n336025 );
or ( n16167 , n336021 , n16166 );
buf ( n336028 , n334564 );
not ( n16169 , n336028 );
buf ( n336030 , n16169 );
buf ( n336031 , n336030 );
buf ( n336032 , n334879 );
nand ( n16173 , n336031 , n336032 );
buf ( n336034 , n16173 );
buf ( n336035 , n336034 );
nand ( n336036 , n16167 , n336035 );
buf ( n336037 , n336036 );
buf ( n336038 , n336037 );
buf ( n336039 , n334917 );
nand ( n336040 , n336038 , n336039 );
buf ( n336041 , n336040 );
nand ( n336042 , n336019 , n336041 );
buf ( n336043 , n336042 );
not ( n16184 , n336043 );
or ( n336045 , n16156 , n16184 );
or ( n16186 , n336042 , n336014 );
not ( n336047 , n14891 );
not ( n336048 , n335314 );
or ( n16189 , n336047 , n336048 );
buf ( n336050 , n334786 );
xnor ( n336051 , n332672 , n15463 );
buf ( n336052 , n336051 );
nand ( n336053 , n336050 , n336052 );
buf ( n336054 , n336053 );
nand ( n16195 , n16189 , n336054 );
buf ( n336056 , n16195 );
not ( n336057 , n336056 );
not ( n16198 , n14499 );
not ( n16199 , n334361 );
or ( n16200 , n16198 , n16199 );
nand ( n16201 , n16200 , n14507 );
buf ( n336062 , n16201 );
not ( n336063 , n336062 );
buf ( n336064 , n336063 );
buf ( n336065 , n336064 );
not ( n16206 , n336065 );
buf ( n336067 , n16206 );
buf ( n336068 , n336067 );
buf ( n336069 , n576 );
nand ( n16210 , n336068 , n336069 );
buf ( n336071 , n16210 );
buf ( n336072 , n336071 );
nand ( n16213 , n336057 , n336072 );
buf ( n336074 , n16213 );
buf ( n336075 , n336074 );
not ( n336076 , n336075 );
buf ( n336077 , n335432 );
not ( n336078 , n336077 );
buf ( n336079 , n335368 );
not ( n336080 , n336079 );
or ( n16221 , n336078 , n336080 );
buf ( n16222 , n578 );
not ( n16223 , n16222 );
buf ( n16224 , n335301 );
not ( n16225 , n16224 );
or ( n16226 , n16223 , n16225 );
buf ( n16227 , n335300 );
buf ( n336088 , n334748 );
nand ( n336089 , n16227 , n336088 );
buf ( n336090 , n336089 );
buf ( n336091 , n336090 );
nand ( n336092 , n16226 , n336091 );
buf ( n336093 , n336092 );
buf ( n336094 , n336093 );
buf ( n336095 , n14949 );
nand ( n16236 , n336094 , n336095 );
buf ( n16237 , n16236 );
buf ( n336098 , n16237 );
nand ( n16239 , n16221 , n336098 );
buf ( n336100 , n16239 );
buf ( n336101 , n336100 );
not ( n16242 , n336101 );
or ( n16243 , n336076 , n16242 );
buf ( n336104 , n336071 );
not ( n16245 , n336104 );
buf ( n336106 , n16195 );
nand ( n336107 , n16245 , n336106 );
buf ( n336108 , n336107 );
buf ( n336109 , n336108 );
nand ( n336110 , n16243 , n336109 );
buf ( n336111 , n336110 );
not ( n336112 , n336111 );
not ( n16253 , n15528 );
not ( n16254 , n335402 );
or ( n336115 , n16253 , n16254 );
not ( n16256 , n335406 );
not ( n336117 , n580 );
not ( n336118 , n14877 );
or ( n16259 , n336117 , n336118 );
buf ( n336120 , n334736 );
buf ( n336121 , n334650 );
nand ( n16262 , n336120 , n336121 );
buf ( n336123 , n16262 );
nand ( n336124 , n16259 , n336123 );
nand ( n336125 , n16256 , n336124 );
nand ( n16266 , n336115 , n336125 );
not ( n336127 , n16266 );
nand ( n336128 , n336112 , n336127 );
not ( n16269 , n336128 );
or ( n336130 , n335326 , n332672 );
or ( n336131 , n15457 , n336130 );
nand ( n16272 , n336131 , n15474 );
buf ( n336133 , n16272 );
not ( n16274 , n336133 );
buf ( n336135 , n16274 );
buf ( n336136 , n336135 );
not ( n16277 , n336136 );
not ( n16278 , n15513 );
buf ( n336139 , n16278 );
not ( n336140 , n336139 );
or ( n16281 , n16277 , n336140 );
nand ( n336142 , n16272 , n15513 );
buf ( n336143 , n336142 );
nand ( n16284 , n16281 , n336143 );
buf ( n336145 , n16284 );
not ( n336146 , n336145 );
or ( n336147 , n16269 , n336146 );
buf ( n336148 , n16266 );
buf ( n336149 , n336111 );
nand ( n336150 , n336148 , n336149 );
buf ( n336151 , n336150 );
nand ( n336152 , n336147 , n336151 );
nand ( n336153 , n16186 , n336152 );
buf ( n336154 , n336153 );
nand ( n336155 , n336045 , n336154 );
buf ( n336156 , n336155 );
buf ( n336157 , n336156 );
buf ( n336158 , n591 );
not ( n16299 , n336158 );
buf ( n336160 , n335173 );
not ( n16301 , n336160 );
or ( n16302 , n16299 , n16301 );
buf ( n336163 , n590 );
not ( n336164 , n336163 );
buf ( n336165 , n15217 );
not ( n16306 , n336165 );
buf ( n336167 , n16306 );
buf ( n336168 , n336167 );
not ( n16309 , n336168 );
or ( n336170 , n336164 , n16309 );
buf ( n336171 , n15217 );
buf ( n336172 , n335097 );
nand ( n336173 , n336171 , n336172 );
buf ( n336174 , n336173 );
buf ( n336175 , n336174 );
nand ( n16316 , n336170 , n336175 );
buf ( n336177 , n16316 );
buf ( n336178 , n336177 );
buf ( n336179 , n335181 );
nand ( n336180 , n336178 , n336179 );
buf ( n336181 , n336180 );
buf ( n336182 , n336181 );
nand ( n16323 , n16302 , n336182 );
buf ( n336184 , n16323 );
buf ( n336185 , n336184 );
xor ( n336186 , n336157 , n336185 );
buf ( n16327 , n335294 );
buf ( n336188 , n335255 );
xor ( n16329 , n16327 , n336188 );
buf ( n336190 , n335448 );
not ( n16331 , n336190 );
xor ( n336192 , n16329 , n16331 );
buf ( n336193 , n336192 );
buf ( n336194 , n336193 );
and ( n336195 , n336186 , n336194 );
and ( n16336 , n336157 , n336185 );
or ( n336197 , n336195 , n16336 );
buf ( n336198 , n336197 );
nand ( n336199 , n16129 , n336198 );
nand ( n16340 , n16123 , n336199 );
buf ( n336201 , n16340 );
not ( n16342 , n336201 );
buf ( n336203 , n16342 );
buf ( n336204 , n336203 );
and ( n16345 , n335932 , n336204 );
buf ( n336206 , n16345 );
buf ( n336207 , n336206 );
or ( n336208 , n335925 , n336207 );
buf ( n336209 , n335931 );
not ( n336210 , n336209 );
buf ( n16351 , n16340 );
nand ( n16352 , n336210 , n16351 );
buf ( n16353 , n16352 );
buf ( n16354 , n16353 );
nand ( n16355 , n336208 , n16354 );
buf ( n16356 , n16355 );
not ( n336217 , n16356 );
nand ( n16358 , n335919 , n336217 );
buf ( n336219 , n16358 );
buf ( n336220 , n336219 );
nand ( n16361 , n335918 , n16356 );
buf ( n336222 , n16361 );
buf ( n16363 , n336222 );
buf ( n336224 , n16363 );
buf ( n336225 , n336224 );
nand ( n16366 , n336220 , n336225 );
buf ( n336227 , n16366 );
not ( n336228 , n336227 );
not ( n336229 , n336228 );
buf ( n336230 , n15528 );
not ( n336231 , n336230 );
and ( n336232 , n335300 , n334650 );
not ( n16373 , n335300 );
and ( n336234 , n16373 , n580 );
or ( n336235 , n336232 , n336234 );
buf ( n336236 , n336235 );
not ( n336237 , n336236 );
or ( n336238 , n336231 , n336237 );
buf ( n336239 , n14822 );
not ( n16380 , n580 );
not ( n336241 , n335310 );
or ( n16382 , n16380 , n336241 );
buf ( n336243 , n14139 );
buf ( n336244 , n334650 );
nand ( n16385 , n336243 , n336244 );
buf ( n336246 , n16385 );
nand ( n16387 , n16382 , n336246 );
buf ( n336248 , n16387 );
nand ( n336249 , n336239 , n336248 );
buf ( n336250 , n336249 );
buf ( n336251 , n336250 );
nand ( n336252 , n336238 , n336251 );
buf ( n336253 , n336252 );
buf ( n336254 , n336253 );
not ( n336255 , n336254 );
buf ( n336256 , n336255 );
not ( n336257 , n336256 );
buf ( n336258 , n576 );
buf ( n336259 , n334420 );
buf ( n336260 , n336259 );
not ( n16401 , n336260 );
xor ( n336262 , n336258 , n16401 );
buf ( n336263 , n336262 );
buf ( n336264 , n336263 );
not ( n336265 , n336264 );
buf ( n336266 , n15711 );
not ( n16407 , n336266 );
and ( n16408 , n336265 , n16407 );
buf ( n336269 , n576 );
not ( n16410 , n336269 );
not ( n16411 , n14629 );
buf ( n336272 , n16411 );
not ( n336273 , n336272 );
or ( n16414 , n16410 , n336273 );
not ( n336275 , n16411 );
buf ( n336276 , n336275 );
buf ( n336277 , n332672 );
nand ( n336278 , n336276 , n336277 );
buf ( n336279 , n336278 );
buf ( n336280 , n336279 );
nand ( n336281 , n16414 , n336280 );
buf ( n336282 , n336281 );
buf ( n336283 , n336282 );
buf ( n336284 , n14891 );
and ( n16425 , n336283 , n336284 );
nor ( n336286 , n16408 , n16425 );
buf ( n336287 , n336286 );
buf ( n336288 , n336287 );
not ( n336289 , n336288 );
buf ( n16430 , n14570 );
buf ( n336291 , n16430 );
not ( n336292 , n336291 );
buf ( n336293 , n336292 );
buf ( n336294 , n336293 );
buf ( n336295 , n336294 );
buf ( n336296 , n336295 );
buf ( n336297 , n336296 );
not ( n336298 , n336297 );
buf ( n336299 , n576 );
nand ( n336300 , n336298 , n336299 );
buf ( n336301 , n336300 );
buf ( n336302 , n336301 );
not ( n336303 , n336302 );
and ( n16444 , n336289 , n336303 );
buf ( n336305 , n335432 );
not ( n16446 , n336305 );
and ( n16447 , n16201 , n334748 );
not ( n16448 , n16201 );
and ( n16449 , n16448 , n578 );
or ( n16450 , n16447 , n16449 );
buf ( n336311 , n16450 );
not ( n16452 , n336311 );
or ( n16453 , n16446 , n16452 );
buf ( n336314 , n578 );
not ( n16455 , n336314 );
not ( n16456 , n14546 );
buf ( n336317 , n16456 );
not ( n16458 , n336317 );
buf ( n336319 , n16458 );
buf ( n336320 , n336319 );
not ( n16461 , n336320 );
or ( n16462 , n16455 , n16461 );
buf ( n336323 , n16456 );
buf ( n336324 , n334748 );
nand ( n16465 , n336323 , n336324 );
buf ( n336326 , n16465 );
buf ( n336327 , n336326 );
nand ( n16468 , n16462 , n336327 );
buf ( n336329 , n16468 );
buf ( n336330 , n336329 );
buf ( n336331 , n14949 );
nand ( n16472 , n336330 , n336331 );
buf ( n336333 , n16472 );
buf ( n336334 , n336333 );
nand ( n16475 , n16453 , n336334 );
buf ( n336336 , n16475 );
buf ( n336337 , n336336 );
buf ( n336338 , n336287 );
buf ( n336339 , n336301 );
nand ( n16480 , n336338 , n336339 );
buf ( n336341 , n16480 );
buf ( n336342 , n336341 );
and ( n16483 , n336337 , n336342 );
nor ( n16484 , n16444 , n16483 );
buf ( n336345 , n16484 );
not ( n16486 , n336345 );
and ( n16487 , n336257 , n16486 );
buf ( n336348 , n336256 );
buf ( n336349 , n336345 );
nand ( n16490 , n336348 , n336349 );
buf ( n336351 , n16490 );
buf ( n336352 , n336259 );
not ( n16493 , n336352 );
buf ( n336354 , n16493 );
buf ( n336355 , n336354 );
not ( n16496 , n336355 );
buf ( n336357 , n16496 );
buf ( n336358 , n336357 );
buf ( n336359 , n576 );
and ( n16500 , n336358 , n336359 );
buf ( n336361 , n16500 );
buf ( n336362 , n14891 );
not ( n16503 , n336362 );
and ( n16504 , n16456 , n332672 );
not ( n16505 , n16456 );
and ( n16506 , n16505 , n576 );
or ( n16507 , n16504 , n16506 );
buf ( n336368 , n16507 );
not ( n16509 , n336368 );
or ( n16510 , n16503 , n16509 );
buf ( n336371 , n336282 );
buf ( n336372 , n334786 );
nand ( n16513 , n336371 , n336372 );
buf ( n336374 , n16513 );
buf ( n336375 , n336374 );
nand ( n16516 , n16510 , n336375 );
buf ( n336377 , n16516 );
buf ( n336378 , n336377 );
not ( n16519 , n336378 );
buf ( n336380 , n16519 );
xor ( n16521 , n336361 , n336380 );
buf ( n336382 , n335432 );
not ( n16523 , n336382 );
and ( n16524 , n15463 , n334748 );
not ( n16525 , n15463 );
and ( n16526 , n16525 , n578 );
or ( n16527 , n16524 , n16526 );
buf ( n336388 , n16527 );
not ( n16529 , n336388 );
or ( n16530 , n16523 , n16529 );
buf ( n336391 , n16450 );
buf ( n336392 , n14949 );
nand ( n16533 , n336391 , n336392 );
buf ( n336394 , n16533 );
buf ( n336395 , n336394 );
nand ( n16536 , n16530 , n336395 );
buf ( n336397 , n16536 );
xnor ( n16538 , n16521 , n336397 );
and ( n16539 , n336351 , n16538 );
nor ( n16540 , n16487 , n16539 );
buf ( n336401 , n16540 );
buf ( n16542 , n336401 );
buf ( n336403 , n16542 );
not ( n336404 , n334694 );
not ( n16545 , n582 );
nand ( n16546 , n14426 , n334288 );
not ( n16547 , n16546 );
or ( n16548 , n16545 , n16547 );
or ( n336409 , n16546 , n582 );
nand ( n336410 , n16548 , n336409 );
not ( n16551 , n336410 );
not ( n16552 , n16551 );
or ( n16553 , n336404 , n16552 );
and ( n16554 , n14448 , n334702 );
not ( n16555 , n14448 );
and ( n336416 , n16555 , n582 );
or ( n336417 , n16554 , n336416 );
buf ( n336418 , n336417 );
buf ( n336419 , n334727 );
nand ( n336420 , n336418 , n336419 );
buf ( n336421 , n336420 );
nand ( n16562 , n16553 , n336421 );
not ( n336423 , n16562 );
nand ( n336424 , n336403 , n336423 );
buf ( n336425 , n336424 );
not ( n336426 , n336425 );
buf ( n336427 , n336361 );
not ( n16568 , n336427 );
buf ( n336429 , n336380 );
nand ( n336430 , n16568 , n336429 );
buf ( n336431 , n336430 );
buf ( n336432 , n336431 );
not ( n336433 , n336432 );
buf ( n336434 , n336397 );
not ( n16575 , n336434 );
or ( n16576 , n336433 , n16575 );
buf ( n336437 , n336377 );
buf ( n336438 , n336361 );
nand ( n336439 , n336437 , n336438 );
buf ( n336440 , n336439 );
buf ( n336441 , n336440 );
nand ( n336442 , n16576 , n336441 );
buf ( n336443 , n336442 );
buf ( n336444 , n336443 );
buf ( n336445 , n14891 );
not ( n336446 , n336445 );
and ( n16587 , n16201 , n332672 );
not ( n336448 , n16201 );
and ( n16589 , n336448 , n576 );
or ( n16590 , n16587 , n16589 );
buf ( n336451 , n16590 );
not ( n16592 , n336451 );
or ( n336453 , n336446 , n16592 );
buf ( n336454 , n16507 );
buf ( n336455 , n334786 );
nand ( n336456 , n336454 , n336455 );
buf ( n336457 , n336456 );
buf ( n336458 , n336457 );
nand ( n336459 , n336453 , n336458 );
buf ( n336460 , n336459 );
buf ( n16601 , n336460 );
not ( n16602 , n16601 );
not ( n336463 , n16411 );
buf ( n336464 , n336463 );
buf ( n336465 , n576 );
nand ( n336466 , n336464 , n336465 );
buf ( n336467 , n336466 );
buf ( n336468 , n336467 );
not ( n16609 , n336468 );
and ( n336470 , n16602 , n16609 );
buf ( n336471 , n336460 );
buf ( n336472 , n336467 );
and ( n336473 , n336471 , n336472 );
nor ( n336474 , n336470 , n336473 );
buf ( n336475 , n336474 );
buf ( n336476 , n336475 );
buf ( n336477 , n335432 );
not ( n16618 , n336477 );
and ( n336479 , n14139 , n334748 );
not ( n336480 , n14139 );
and ( n16621 , n336480 , n578 );
or ( n336482 , n336479 , n16621 );
buf ( n336483 , n336482 );
not ( n16624 , n336483 );
or ( n16625 , n16618 , n16624 );
buf ( n336486 , n16527 );
buf ( n336487 , n14949 );
nand ( n16628 , n336486 , n336487 );
buf ( n336489 , n16628 );
buf ( n336490 , n336489 );
nand ( n16631 , n16625 , n336490 );
buf ( n336492 , n16631 );
buf ( n336493 , n336492 );
or ( n16634 , n336476 , n336493 );
buf ( n336495 , n336492 );
buf ( n336496 , n336475 );
nand ( n16637 , n336495 , n336496 );
buf ( n336498 , n16637 );
buf ( n336499 , n336498 );
nand ( n16640 , n16634 , n336499 );
buf ( n336501 , n16640 );
buf ( n336502 , n336501 );
xor ( n16643 , n336444 , n336502 );
buf ( n336504 , n15528 );
not ( n16645 , n336504 );
buf ( n336506 , n580 );
not ( n16647 , n336506 );
buf ( n336508 , n335355 );
not ( n16649 , n336508 );
or ( n336510 , n16647 , n16649 );
buf ( n336511 , n14129 );
buf ( n336512 , n334650 );
nand ( n336513 , n336511 , n336512 );
buf ( n336514 , n336513 );
buf ( n336515 , n336514 );
nand ( n16656 , n336510 , n336515 );
buf ( n336517 , n16656 );
buf ( n336518 , n336517 );
not ( n16659 , n336518 );
or ( n16660 , n16645 , n16659 );
buf ( n336521 , n336235 );
buf ( n336522 , n14822 );
nand ( n16663 , n336521 , n336522 );
buf ( n336524 , n16663 );
buf ( n336525 , n336524 );
nand ( n16666 , n16660 , n336525 );
buf ( n16667 , n16666 );
buf ( n336528 , n16667 );
xor ( n16669 , n16643 , n336528 );
buf ( n336530 , n16669 );
buf ( n336531 , n336530 );
not ( n16672 , n336531 );
or ( n336533 , n336426 , n16672 );
or ( n336534 , n336403 , n336423 );
buf ( n336535 , n336534 );
nand ( n16676 , n336533 , n336535 );
buf ( n16677 , n16676 );
buf ( n336538 , n16677 );
buf ( n336539 , n334868 );
not ( n336540 , n336539 );
buf ( n336541 , n584 );
not ( n16682 , n336541 );
buf ( n336543 , n335514 );
not ( n16684 , n336543 );
or ( n336545 , n16682 , n16684 );
buf ( n16686 , n14957 );
not ( n336547 , n16686 );
nand ( n16688 , n336547 , n334879 );
buf ( n336549 , n16688 );
nand ( n336550 , n336545 , n336549 );
buf ( n336551 , n336550 );
buf ( n336552 , n336551 );
not ( n16693 , n336552 );
or ( n336554 , n336540 , n16693 );
buf ( n336555 , n334879 );
not ( n16696 , n336555 );
buf ( n336557 , n14897 );
not ( n336558 , n336557 );
or ( n16699 , n16696 , n336558 );
buf ( n336560 , n14897 );
buf ( n336561 , n334879 );
or ( n16702 , n336560 , n336561 );
nand ( n16703 , n16699 , n16702 );
buf ( n336564 , n16703 );
buf ( n336565 , n336564 );
buf ( n336566 , n334917 );
nand ( n16707 , n336565 , n336566 );
buf ( n336568 , n16707 );
buf ( n336569 , n336568 );
nand ( n336570 , n336554 , n336569 );
buf ( n336571 , n336570 );
buf ( n336572 , n336571 );
xor ( n336573 , n336538 , n336572 );
not ( n336574 , n15115 );
not ( n16715 , n336030 );
not ( n336576 , n334982 );
or ( n336577 , n16715 , n336576 );
nand ( n16718 , n334662 , n586 );
nand ( n16719 , n336577 , n16718 );
not ( n16720 , n16719 );
or ( n16721 , n336574 , n16720 );
buf ( n336582 , n586 );
not ( n336583 , n336582 );
not ( n16724 , n14698 );
buf ( n336585 , n16724 );
not ( n336586 , n336585 );
or ( n16727 , n336583 , n336586 );
buf ( n336588 , n334837 );
not ( n336589 , n336588 );
buf ( n16730 , n334982 );
nand ( n16731 , n336589 , n16730 );
buf ( n16732 , n16731 );
buf ( n336593 , n16732 );
nand ( n16734 , n16727 , n336593 );
buf ( n16735 , n16734 );
buf ( n336596 , n16735 );
buf ( n336597 , n15164 );
nand ( n16738 , n336596 , n336597 );
buf ( n336599 , n16738 );
nand ( n336600 , n16721 , n336599 );
buf ( n336601 , n336600 );
xnor ( n336602 , n336573 , n336601 );
buf ( n336603 , n336602 );
not ( n16744 , n334694 );
not ( n336605 , n336417 );
or ( n16746 , n16744 , n336605 );
buf ( n336607 , n582 );
not ( n336608 , n336607 );
buf ( n336609 , n335355 );
not ( n16750 , n336609 );
or ( n336611 , n336608 , n16750 );
buf ( n336612 , n335361 );
buf ( n336613 , n334702 );
nand ( n16754 , n336612 , n336613 );
buf ( n336615 , n16754 );
buf ( n336616 , n336615 );
nand ( n16757 , n336611 , n336616 );
buf ( n336618 , n16757 );
buf ( n336619 , n336618 );
buf ( n336620 , n334727 );
nand ( n16761 , n336619 , n336620 );
buf ( n336622 , n16761 );
nand ( n16763 , n16746 , n336622 );
not ( n16764 , n16763 );
not ( n16765 , n334868 );
not ( n16766 , n584 );
not ( n16767 , n335392 );
or ( n16768 , n16766 , n16767 );
buf ( n336629 , n14913 );
buf ( n336630 , n334879 );
nand ( n16771 , n336629 , n336630 );
buf ( n336632 , n16771 );
nand ( n16773 , n16768 , n336632 );
not ( n16774 , n16773 );
or ( n16775 , n16765 , n16774 );
buf ( n336636 , n584 );
not ( n16777 , n336636 );
buf ( n336638 , n335434 );
not ( n16779 , n336638 );
or ( n16780 , n16777 , n16779 );
buf ( n336641 , n334736 );
buf ( n336642 , n334879 );
nand ( n16783 , n336641 , n336642 );
buf ( n336644 , n16783 );
buf ( n336645 , n336644 );
nand ( n16786 , n16780 , n336645 );
buf ( n336647 , n16786 );
nand ( n16788 , n336647 , n334917 );
nand ( n16789 , n16775 , n16788 );
not ( n16790 , n16789 );
or ( n16791 , n16764 , n16790 );
not ( n16792 , n16763 );
buf ( n336653 , n16792 );
not ( n16794 , n336653 );
not ( n16795 , n16789 );
buf ( n336656 , n16795 );
not ( n16797 , n336656 );
or ( n16798 , n16794 , n16797 );
buf ( n16799 , n334444 );
buf ( n336660 , n16799 );
not ( n16801 , n336660 );
buf ( n336662 , n16801 );
buf ( n336663 , n336662 );
not ( n16804 , n336663 );
buf ( n336665 , n16804 );
buf ( n336666 , n336665 );
not ( n16807 , n336666 );
buf ( n336668 , n332672 );
nor ( n16809 , n16807 , n336668 );
buf ( n336670 , n16809 );
buf ( n336671 , n336670 );
not ( n16812 , n336671 );
buf ( n336673 , n336263 );
not ( n16814 , n336673 );
buf ( n336675 , n16814 );
buf ( n336676 , n336675 );
buf ( n336677 , n14891 );
and ( n16818 , n336676 , n336677 );
buf ( n336679 , n16430 );
not ( n16820 , n336679 );
buf ( n336681 , n16820 );
and ( n16822 , n336681 , n576 );
not ( n16823 , n336681 );
and ( n16824 , n16823 , n332672 );
or ( n16825 , n16822 , n16824 );
buf ( n336686 , n16825 );
buf ( n336687 , n334786 );
and ( n16828 , n336686 , n336687 );
buf ( n336689 , n16828 );
buf ( n336690 , n336689 );
nor ( n16831 , n16818 , n336690 );
buf ( n336692 , n16831 );
buf ( n336693 , n336692 );
nand ( n16834 , n16812 , n336693 );
buf ( n336695 , n16834 );
buf ( n336696 , n336695 );
not ( n16837 , n336696 );
not ( n16838 , n335432 );
not ( n16839 , n336329 );
or ( n16840 , n16838 , n16839 );
buf ( n336701 , n578 );
not ( n16842 , n336701 );
not ( n16843 , n336275 );
buf ( n336704 , n16843 );
not ( n16845 , n336704 );
or ( n16846 , n16842 , n16845 );
buf ( n336707 , n336463 );
buf ( n336708 , n334748 );
nand ( n16849 , n336707 , n336708 );
buf ( n336710 , n16849 );
buf ( n336711 , n336710 );
nand ( n16852 , n16846 , n336711 );
buf ( n336713 , n16852 );
buf ( n336714 , n336713 );
buf ( n336715 , n14949 );
nand ( n16856 , n336714 , n336715 );
buf ( n336717 , n16856 );
nand ( n16858 , n16840 , n336717 );
buf ( n336719 , n16858 );
not ( n16860 , n336719 );
or ( n16861 , n16837 , n16860 );
buf ( n336722 , n336692 );
not ( n16863 , n336722 );
buf ( n336724 , n336670 );
nand ( n16865 , n16863 , n336724 );
buf ( n336726 , n16865 );
buf ( n336727 , n336726 );
nand ( n16868 , n16861 , n336727 );
buf ( n336729 , n16868 );
buf ( n336730 , n336729 );
not ( n16871 , n336730 );
not ( n16872 , n334643 );
not ( n16873 , n16387 );
or ( n16874 , n16872 , n16873 );
buf ( n336735 , n580 );
not ( n16876 , n336735 );
buf ( n336737 , n335326 );
not ( n16878 , n336737 );
or ( n16879 , n16876 , n16878 );
buf ( n336740 , n15463 );
buf ( n336741 , n334650 );
nand ( n16882 , n336740 , n336741 );
buf ( n336743 , n16882 );
buf ( n336744 , n336743 );
nand ( n16885 , n16879 , n336744 );
buf ( n336746 , n16885 );
buf ( n336747 , n336746 );
buf ( n336748 , n14822 );
nand ( n16889 , n336747 , n336748 );
buf ( n336750 , n16889 );
nand ( n16891 , n16874 , n336750 );
not ( n16892 , n16891 );
buf ( n336753 , n16892 );
nand ( n16894 , n16871 , n336753 );
buf ( n336755 , n16894 );
buf ( n336756 , n336336 );
buf ( n336757 , n336287 );
buf ( n336758 , n336301 );
xor ( n16899 , n336757 , n336758 );
buf ( n336760 , n16899 );
buf ( n336761 , n336760 );
xor ( n16902 , n336756 , n336761 );
buf ( n336763 , n16902 );
and ( n16904 , n336755 , n336763 );
buf ( n336765 , n16891 );
buf ( n336766 , n336729 );
and ( n16907 , n336765 , n336766 );
buf ( n336768 , n16907 );
nor ( n16909 , n16904 , n336768 );
not ( n16910 , n16909 );
buf ( n336771 , n16910 );
nand ( n336772 , n16798 , n336771 );
buf ( n336773 , n336772 );
nand ( n16914 , n16791 , n336773 );
buf ( n336775 , n16914 );
not ( n16916 , n336775 );
buf ( n336777 , n16916 );
not ( n336778 , n336777 );
buf ( n16919 , n16773 );
not ( n336780 , n16919 );
buf ( n336781 , n336780 );
buf ( n336782 , n336781 );
not ( n336783 , n336782 );
buf ( n336784 , n334917 );
not ( n16925 , n336784 );
buf ( n336786 , n16925 );
buf ( n336787 , n336786 );
not ( n16928 , n336787 );
and ( n336789 , n336783 , n16928 );
buf ( n336790 , n336564 );
buf ( n336791 , n334868 );
and ( n16932 , n336790 , n336791 );
nor ( n16933 , n336789 , n16932 );
buf ( n336794 , n16933 );
not ( n16935 , n336794 );
and ( n336796 , n336778 , n16935 );
buf ( n336797 , n336777 );
buf ( n336798 , n336794 );
nand ( n336799 , n336797 , n336798 );
buf ( n336800 , n336799 );
and ( n16941 , n336423 , n16540 );
not ( n336802 , n336423 );
not ( n336803 , n16540 );
and ( n16944 , n336802 , n336803 );
nor ( n336805 , n16941 , n16944 );
and ( n16946 , n336805 , n336530 );
not ( n336807 , n336805 );
not ( n336808 , n336530 );
and ( n16949 , n336807 , n336808 );
nor ( n336810 , n16946 , n16949 );
buf ( n16951 , n336810 );
buf ( n336812 , n16951 );
buf ( n336813 , n336812 );
and ( n16954 , n336800 , n336813 );
nor ( n336815 , n336796 , n16954 );
or ( n16956 , n336603 , n336815 );
not ( n16957 , n334978 );
not ( n336818 , n16735 );
or ( n336819 , n16957 , n336818 );
buf ( n336820 , n586 );
not ( n16961 , n336820 );
buf ( n336822 , n334821 );
not ( n336823 , n336822 );
or ( n16964 , n16961 , n336823 );
buf ( n336825 , n335514 );
not ( n336826 , n336825 );
buf ( n336827 , n334982 );
nand ( n336828 , n336826 , n336827 );
buf ( n336829 , n336828 );
buf ( n336830 , n336829 );
nand ( n16971 , n16964 , n336830 );
buf ( n336832 , n16971 );
nand ( n16973 , n336832 , n15164 );
nand ( n16974 , n336819 , n16973 );
not ( n336835 , n16974 );
not ( n336836 , n336835 );
buf ( n336837 , n588 );
buf ( n336838 , n336024 );
xor ( n336839 , n336837 , n336838 );
buf ( n336840 , n336839 );
not ( n16981 , n336840 );
not ( n16982 , n335111 );
and ( n16983 , n16981 , n16982 );
not ( n16984 , n588 );
not ( n336845 , n334647 );
not ( n336846 , n336845 );
or ( n16987 , n16984 , n336846 );
buf ( n336848 , n15381 );
buf ( n336849 , n334972 );
nand ( n16990 , n336848 , n336849 );
buf ( n336851 , n16990 );
nand ( n16992 , n16987 , n336851 );
and ( n16993 , n16992 , n15275 );
nor ( n336854 , n16983 , n16993 );
not ( n16995 , n336854 );
or ( n336856 , n336836 , n16995 );
not ( n16997 , n16974 );
not ( n16998 , n336854 );
not ( n336859 , n16998 );
or ( n336860 , n16997 , n336859 );
buf ( n336861 , n590 );
not ( n17002 , n336861 );
buf ( n336863 , n334709 );
buf ( n336864 , n336863 );
buf ( n336865 , n336864 );
buf ( n336866 , n336865 );
not ( n336867 , n336866 );
buf ( n336868 , n336867 );
buf ( n336869 , n336868 );
not ( n17010 , n336869 );
or ( n17011 , n17002 , n17010 );
buf ( n336872 , n336865 );
buf ( n336873 , n335097 );
nand ( n17014 , n336872 , n336873 );
buf ( n336875 , n17014 );
buf ( n336876 , n336875 );
nand ( n17017 , n17011 , n336876 );
buf ( n336878 , n17017 );
buf ( n336879 , n336878 );
buf ( n336880 , n335181 );
and ( n336881 , n336879 , n336880 );
buf ( n336882 , n590 );
not ( n17023 , n336882 );
buf ( n336884 , n14689 );
not ( n336885 , n336884 );
buf ( n336886 , n336885 );
buf ( n336887 , n336886 );
not ( n336888 , n336887 );
or ( n17029 , n17023 , n336888 );
buf ( n336890 , n14689 );
buf ( n336891 , n335097 );
nand ( n336892 , n336890 , n336891 );
buf ( n336893 , n336892 );
buf ( n336894 , n336893 );
nand ( n336895 , n17029 , n336894 );
buf ( n336896 , n336895 );
buf ( n336897 , n336896 );
buf ( n336898 , n591 );
and ( n336899 , n336897 , n336898 );
nor ( n17040 , n336881 , n336899 );
buf ( n17041 , n17040 );
nand ( n336902 , n336860 , n17041 );
nand ( n17043 , n336856 , n336902 );
nand ( n336904 , n16956 , n17043 );
nand ( n336905 , n336603 , n336815 );
nand ( n17046 , n336904 , n336905 );
not ( n336907 , n336410 );
buf ( n336908 , n334727 );
not ( n336909 , n336908 );
buf ( n336910 , n336909 );
not ( n17051 , n336910 );
and ( n336912 , n336907 , n17051 );
buf ( n336913 , n334702 );
not ( n336914 , n336913 );
not ( n17055 , n335392 );
buf ( n336916 , n17055 );
not ( n17057 , n336916 );
or ( n17058 , n336914 , n17057 );
not ( n17059 , n14913 );
nand ( n336920 , n17059 , n582 );
buf ( n336921 , n336920 );
nand ( n336922 , n17058 , n336921 );
buf ( n336923 , n336922 );
and ( n17064 , n336923 , n334694 );
nor ( n17065 , n336912 , n17064 );
xor ( n17066 , n336444 , n336502 );
and ( n17067 , n17066 , n336528 );
and ( n17068 , n336444 , n336502 );
or ( n336929 , n17067 , n17068 );
buf ( n336930 , n336929 );
buf ( n336931 , n336930 );
not ( n336932 , n336931 );
buf ( n336933 , n336932 );
or ( n17074 , n17065 , n336933 );
not ( n336935 , n17074 );
buf ( n336936 , n336460 );
not ( n336937 , n336936 );
buf ( n336938 , n336467 );
nand ( n336939 , n336937 , n336938 );
buf ( n336940 , n336939 );
buf ( n336941 , n336940 );
not ( n17082 , n336941 );
buf ( n336943 , n336492 );
not ( n17084 , n336943 );
or ( n336945 , n17082 , n17084 );
buf ( n336946 , n336467 );
not ( n336947 , n336946 );
buf ( n336948 , n336460 );
nand ( n17089 , n336947 , n336948 );
buf ( n336950 , n17089 );
buf ( n336951 , n336950 );
nand ( n336952 , n336945 , n336951 );
buf ( n336953 , n336952 );
buf ( n336954 , n336953 );
buf ( n336955 , n334643 );
not ( n17096 , n336955 );
buf ( n336957 , n580 );
not ( n336958 , n336957 );
buf ( n336959 , n15095 );
not ( n336960 , n336959 );
or ( n17101 , n336958 , n336960 );
buf ( n336962 , n15481 );
buf ( n336963 , n334650 );
nand ( n17104 , n336962 , n336963 );
buf ( n336965 , n17104 );
buf ( n336966 , n336965 );
nand ( n17107 , n17101 , n336966 );
buf ( n336968 , n17107 );
buf ( n336969 , n336968 );
not ( n17110 , n336969 );
or ( n17111 , n17096 , n17110 );
buf ( n336972 , n336517 );
buf ( n336973 , n14822 );
nand ( n17114 , n336972 , n336973 );
buf ( n336975 , n17114 );
buf ( n336976 , n336975 );
nand ( n17117 , n17111 , n336976 );
buf ( n336978 , n17117 );
buf ( n336979 , n336978 );
xor ( n17120 , n336954 , n336979 );
buf ( n336981 , n336319 );
not ( n17122 , n336981 );
buf ( n336983 , n17122 );
nand ( n17124 , n336983 , n576 );
and ( n17125 , n336051 , n14891 );
buf ( n336986 , n16590 );
not ( n17127 , n336986 );
buf ( n336988 , n15711 );
nor ( n17129 , n17127 , n336988 );
buf ( n336990 , n17129 );
nor ( n17131 , n17125 , n336990 );
xor ( n17132 , n17124 , n17131 );
buf ( n336993 , n14941 );
not ( n17134 , n336993 );
buf ( n336995 , n336093 );
not ( n17136 , n336995 );
or ( n17137 , n17134 , n17136 );
buf ( n336998 , n336482 );
buf ( n336999 , n14949 );
nand ( n17140 , n336998 , n336999 );
buf ( n337001 , n17140 );
buf ( n337002 , n337001 );
nand ( n17143 , n17137 , n337002 );
buf ( n337004 , n17143 );
buf ( n337005 , n337004 );
not ( n17146 , n337005 );
buf ( n337007 , n17146 );
xor ( n17148 , n17132 , n337007 );
buf ( n337009 , n17148 );
xor ( n17150 , n17120 , n337009 );
buf ( n337011 , n17150 );
not ( n17152 , n337011 );
or ( n17153 , n336935 , n17152 );
nand ( n17154 , n17065 , n336933 );
nand ( n17155 , n17153 , n17154 );
buf ( n337016 , n17155 );
not ( n17157 , n336953 );
not ( n17158 , n336978 );
or ( n17159 , n17157 , n17158 );
not ( n17160 , n336953 );
not ( n17161 , n17160 );
not ( n17162 , n336978 );
not ( n17163 , n17162 );
or ( n17164 , n17161 , n17163 );
not ( n17165 , n17148 );
nand ( n17166 , n17164 , n17165 );
nand ( n17167 , n17159 , n17166 );
not ( n337028 , n14897 );
not ( n337029 , n334702 );
or ( n17170 , n337028 , n337029 );
not ( n337031 , n14254 );
nand ( n337032 , n337031 , n582 );
nand ( n17173 , n17170 , n337032 );
not ( n337034 , n17173 );
not ( n17175 , n334694 );
or ( n17176 , n337034 , n17175 );
nand ( n337037 , n336923 , n334727 );
nand ( n337038 , n17176 , n337037 );
xor ( n17179 , n17167 , n337038 );
buf ( n337040 , n334917 );
not ( n17181 , n337040 );
buf ( n337042 , n336551 );
not ( n337043 , n337042 );
or ( n17184 , n17181 , n337043 );
buf ( n337045 , n584 );
not ( n17186 , n337045 );
buf ( n337047 , n16724 );
not ( n337048 , n337047 );
or ( n17189 , n17186 , n337048 );
buf ( n337050 , n14698 );
buf ( n337051 , n334879 );
nand ( n337052 , n337050 , n337051 );
buf ( n337053 , n337052 );
buf ( n337054 , n337053 );
nand ( n337055 , n17189 , n337054 );
buf ( n337056 , n337055 );
buf ( n337057 , n337056 );
buf ( n337058 , n334868 );
nand ( n337059 , n337057 , n337058 );
buf ( n337060 , n337059 );
buf ( n337061 , n337060 );
nand ( n17202 , n17184 , n337061 );
buf ( n337063 , n17202 );
xor ( n17204 , n17179 , n337063 );
buf ( n337065 , n17204 );
xor ( n337066 , n337016 , n337065 );
buf ( n337067 , n336600 );
not ( n17208 , n337067 );
buf ( n337069 , n336571 );
not ( n17210 , n337069 );
or ( n17211 , n17208 , n17210 );
or ( n337072 , n336600 , n336571 );
nand ( n337073 , n337072 , n16677 );
buf ( n337074 , n337073 );
nand ( n17215 , n17211 , n337074 );
buf ( n337076 , n17215 );
buf ( n337077 , n337076 );
xor ( n337078 , n337066 , n337077 );
buf ( n337079 , n337078 );
xor ( n17220 , n17046 , n337079 );
not ( n337081 , n591 );
not ( n337082 , n590 );
buf ( n337083 , n333978 );
buf ( n17224 , n337083 );
buf ( n337085 , n17224 );
buf ( n337086 , n337085 );
not ( n17227 , n337086 );
buf ( n337088 , n17227 );
not ( n337089 , n337088 );
or ( n337090 , n337082 , n337089 );
nand ( n17231 , n337085 , n335097 );
nand ( n337092 , n337090 , n17231 );
not ( n337093 , n337092 );
or ( n17234 , n337081 , n337093 );
buf ( n337095 , n590 );
not ( n337096 , n337095 );
buf ( n337097 , n334873 );
not ( n337098 , n337097 );
or ( n337099 , n337096 , n337098 );
not ( n17240 , n334873 );
buf ( n337101 , n17240 );
buf ( n337102 , n335097 );
nand ( n337103 , n337101 , n337102 );
buf ( n337104 , n337103 );
buf ( n337105 , n337104 );
nand ( n337106 , n337099 , n337105 );
buf ( n337107 , n337106 );
buf ( n337108 , n337107 );
buf ( n337109 , n335181 );
nand ( n337110 , n337108 , n337109 );
buf ( n337111 , n337110 );
nand ( n337112 , n17234 , n337111 );
buf ( n17253 , n337112 );
xor ( n17254 , n17124 , n17131 );
and ( n337115 , n17254 , n337007 );
and ( n337116 , n17124 , n17131 );
nor ( n17257 , n337115 , n337116 );
buf ( n337118 , n17257 );
buf ( n337119 , n334643 );
not ( n17260 , n337119 );
buf ( n337121 , n336124 );
not ( n17262 , n337121 );
or ( n17263 , n17260 , n17262 );
buf ( n337124 , n336968 );
buf ( n337125 , n14822 );
nand ( n17266 , n337124 , n337125 );
buf ( n337127 , n17266 );
buf ( n337128 , n337127 );
nand ( n337129 , n17263 , n337128 );
buf ( n337130 , n337129 );
buf ( n337131 , n337130 );
xor ( n17272 , n337118 , n337131 );
buf ( n337133 , n336100 );
xor ( n17274 , n336071 , n16195 );
buf ( n337135 , n17274 );
xnor ( n337136 , n337133 , n337135 );
buf ( n337137 , n337136 );
buf ( n337138 , n337137 );
xor ( n17279 , n17272 , n337138 );
buf ( n337140 , n17279 );
buf ( n17281 , n337140 );
buf ( n337142 , n15275 );
not ( n17283 , n337142 );
buf ( n337144 , n588 );
not ( n337145 , n337144 );
buf ( n337146 , n14837 );
not ( n337147 , n337146 );
or ( n17288 , n337145 , n337147 );
buf ( n337149 , n334896 );
buf ( n337150 , n334972 );
nand ( n17291 , n337149 , n337150 );
buf ( n337152 , n17291 );
buf ( n337153 , n337152 );
nand ( n17294 , n17288 , n337153 );
buf ( n337155 , n17294 );
buf ( n337156 , n337155 );
not ( n17297 , n337156 );
or ( n17298 , n17283 , n17297 );
and ( n17299 , n588 , n334715 );
not ( n17300 , n588 );
buf ( n337161 , n334715 );
not ( n17302 , n337161 );
buf ( n337163 , n17302 );
and ( n17304 , n17300 , n337163 );
or ( n337165 , n17299 , n17304 );
buf ( n337166 , n337165 );
buf ( n337167 , n335114 );
nand ( n17308 , n337166 , n337167 );
buf ( n337169 , n17308 );
buf ( n337170 , n337169 );
nand ( n337171 , n17298 , n337170 );
buf ( n337172 , n337171 );
buf ( n337173 , n337172 );
xor ( n337174 , n17281 , n337173 );
buf ( n337175 , n15115 );
not ( n17316 , n337175 );
buf ( n337177 , n586 );
not ( n17318 , n337177 );
not ( n17319 , n15381 );
buf ( n337180 , n17319 );
not ( n337181 , n337180 );
or ( n17322 , n17318 , n337181 );
not ( n337183 , n335237 );
buf ( n337184 , n337183 );
buf ( n337185 , n334982 );
nand ( n17326 , n337184 , n337185 );
buf ( n337187 , n17326 );
buf ( n337188 , n337187 );
nand ( n17329 , n17322 , n337188 );
buf ( n337190 , n17329 );
buf ( n337191 , n337190 );
not ( n17332 , n337191 );
or ( n337193 , n17316 , n17332 );
buf ( n17334 , n16719 );
buf ( n337195 , n15164 );
nand ( n337196 , n17334 , n337195 );
buf ( n337197 , n337196 );
buf ( n337198 , n337197 );
nand ( n337199 , n337193 , n337198 );
buf ( n337200 , n337199 );
buf ( n337201 , n337200 );
xnor ( n337202 , n337174 , n337201 );
buf ( n337203 , n337202 );
buf ( n337204 , n337203 );
not ( n17345 , n337204 );
buf ( n337206 , n17345 );
buf ( n337207 , n337206 );
xor ( n17348 , n17253 , n337207 );
buf ( n337209 , n15275 );
not ( n17350 , n337209 );
buf ( n337211 , n337165 );
not ( n17352 , n337211 );
or ( n17353 , n17350 , n17352 );
nand ( n17354 , n16992 , n335114 );
buf ( n337215 , n17354 );
nand ( n17356 , n17353 , n337215 );
buf ( n337217 , n17356 );
not ( n17358 , n337217 );
not ( n17359 , n17358 );
buf ( n337220 , n591 );
not ( n17361 , n337220 );
buf ( n337222 , n337107 );
not ( n17363 , n337222 );
or ( n17364 , n17361 , n17363 );
buf ( n337225 , n336896 );
buf ( n337226 , n335181 );
nand ( n17367 , n337225 , n337226 );
buf ( n337228 , n17367 );
buf ( n337229 , n337228 );
nand ( n17370 , n17364 , n337229 );
buf ( n337231 , n17370 );
not ( n17372 , n337231 );
not ( n17373 , n17372 );
or ( n17374 , n17359 , n17373 );
not ( n17375 , n336930 );
not ( n17376 , n17065 );
and ( n17377 , n17375 , n17376 );
and ( n17378 , n17065 , n336930 );
nor ( n17379 , n17377 , n17378 );
and ( n17380 , n17379 , n337011 );
not ( n17381 , n17379 );
not ( n17382 , n337011 );
and ( n17383 , n17381 , n17382 );
nor ( n17384 , n17380 , n17383 );
not ( n17385 , n17384 );
not ( n17386 , n17385 );
nand ( n17387 , n17374 , n17386 );
nand ( n17388 , n337217 , n337231 );
nand ( n17389 , n17387 , n17388 );
buf ( n337250 , n17389 );
xnor ( n17391 , n17348 , n337250 );
buf ( n337252 , n17391 );
xor ( n17393 , n17220 , n337252 );
xor ( n17394 , n336815 , n17043 );
xnor ( n17395 , n17394 , n336603 );
xor ( n17396 , n17384 , n337217 );
xnor ( n17397 , n17396 , n337231 );
not ( n17398 , n17397 );
or ( n17399 , n17395 , n17398 );
not ( n17400 , n336777 );
buf ( n337261 , n336810 );
buf ( n337262 , n336794 );
nand ( n17403 , n337261 , n337262 );
buf ( n337264 , n17403 );
not ( n17405 , n336810 );
buf ( n337266 , n336794 );
not ( n17407 , n337266 );
buf ( n337268 , n17407 );
nand ( n17409 , n17405 , n337268 );
nand ( n17410 , n337264 , n17409 );
not ( n17411 , n17410 );
or ( n17412 , n17400 , n17411 );
nand ( n17413 , n16914 , n17409 , n337264 );
nand ( n17414 , n17412 , n17413 );
not ( n17415 , n17414 );
xor ( n17416 , n336253 , n336345 );
xnor ( n337277 , n17416 , n16538 );
buf ( n337278 , n334452 );
buf ( n337279 , n337278 );
buf ( n337280 , n576 );
and ( n17421 , n337279 , n337280 );
buf ( n337282 , n17421 );
buf ( n337283 , n337282 );
buf ( n337284 , n14891 );
not ( n337285 , n337284 );
buf ( n337286 , n16825 );
not ( n17427 , n337286 );
or ( n17428 , n337285 , n17427 );
buf ( n337289 , n332672 );
not ( n17430 , n337289 );
buf ( n337291 , n16799 );
not ( n17432 , n337291 );
or ( n17433 , n17430 , n17432 );
buf ( n337294 , n336665 );
not ( n17435 , n337294 );
buf ( n337296 , n576 );
nand ( n337297 , n17435 , n337296 );
buf ( n337298 , n337297 );
buf ( n337299 , n337298 );
nand ( n17440 , n17433 , n337299 );
buf ( n337301 , n17440 );
buf ( n337302 , n337301 );
buf ( n337303 , n334786 );
nand ( n17444 , n337302 , n337303 );
buf ( n337305 , n17444 );
buf ( n337306 , n337305 );
nand ( n17447 , n17428 , n337306 );
buf ( n337308 , n17447 );
buf ( n17449 , n337308 );
xor ( n17450 , n337283 , n17449 );
buf ( n337311 , n334002 );
not ( n337312 , n337311 );
buf ( n337313 , n337312 );
buf ( n337314 , n337313 );
not ( n17455 , n337314 );
buf ( n17456 , n17455 );
buf ( n337317 , n17456 );
buf ( n337318 , n576 );
nand ( n337319 , n337317 , n337318 );
buf ( n337320 , n337319 );
buf ( n337321 , n337320 );
not ( n337322 , n337321 );
buf ( n337323 , n337322 );
buf ( n337324 , n337323 );
not ( n337325 , n337324 );
buf ( n337326 , n337301 );
buf ( n337327 , n14891 );
and ( n17468 , n337326 , n337327 );
not ( n17469 , n576 );
buf ( n337330 , n337278 );
not ( n17471 , n337330 );
buf ( n337332 , n17471 );
not ( n337333 , n337332 );
or ( n17474 , n17469 , n337333 );
buf ( n337335 , n337278 );
buf ( n337336 , n332672 );
nand ( n337337 , n337335 , n337336 );
buf ( n337338 , n337337 );
nand ( n17479 , n17474 , n337338 );
buf ( n337340 , n17479 );
not ( n17481 , n337340 );
buf ( n337342 , n15711 );
nor ( n337343 , n17481 , n337342 );
buf ( n337344 , n337343 );
buf ( n337345 , n337344 );
nor ( n337346 , n17468 , n337345 );
buf ( n337347 , n337346 );
buf ( n337348 , n337347 );
not ( n337349 , n337348 );
buf ( n337350 , n337349 );
buf ( n337351 , n337350 );
not ( n337352 , n337351 );
or ( n17493 , n337325 , n337352 );
buf ( n337354 , n337320 );
not ( n337355 , n337354 );
buf ( n337356 , n337347 );
not ( n337357 , n337356 );
or ( n337358 , n337355 , n337357 );
buf ( n337359 , n14599 );
not ( n337360 , n337359 );
buf ( n337361 , n337360 );
buf ( n337362 , n337361 );
not ( n337363 , n337362 );
buf ( n337364 , n337363 );
buf ( n337365 , n337364 );
buf ( n337366 , n576 );
and ( n17507 , n337365 , n337366 );
buf ( n337368 , n17507 );
buf ( n337369 , n337368 );
buf ( n337370 , n337361 );
buf ( n337371 , n576 );
and ( n17512 , n337370 , n337371 );
buf ( n337373 , n337364 );
buf ( n337374 , n332672 );
and ( n337375 , n337373 , n337374 );
nor ( n337376 , n17512 , n337375 );
buf ( n337377 , n337376 );
not ( n337378 , n337377 );
not ( n337379 , n15711 );
and ( n17520 , n337378 , n337379 );
not ( n17521 , n576 );
buf ( n337382 , n334002 );
not ( n17523 , n337382 );
buf ( n337384 , n17523 );
not ( n337385 , n337384 );
or ( n337386 , n17521 , n337385 );
buf ( n337387 , n17456 );
buf ( n337388 , n332672 );
nand ( n337389 , n337387 , n337388 );
buf ( n337390 , n337389 );
nand ( n337391 , n337386 , n337390 );
and ( n337392 , n337391 , n14891 );
nor ( n17533 , n17520 , n337392 );
buf ( n337394 , n17533 );
buf ( n337395 , n577 );
buf ( n337396 , n578 );
or ( n17537 , n337395 , n337396 );
buf ( n337398 , n337364 );
nand ( n17539 , n17537 , n337398 );
buf ( n17540 , n17539 );
buf ( n337401 , n17540 );
buf ( n337402 , n577 );
buf ( n337403 , n578 );
and ( n17544 , n337402 , n337403 );
buf ( n337405 , n332672 );
nor ( n17546 , n17544 , n337405 );
buf ( n337407 , n17546 );
buf ( n337408 , n337407 );
nand ( n337409 , n337401 , n337408 );
buf ( n337410 , n337409 );
buf ( n337411 , n337410 );
nor ( n337412 , n337394 , n337411 );
buf ( n337413 , n337412 );
buf ( n337414 , n337413 );
xor ( n17555 , n337369 , n337414 );
buf ( n337416 , n14891 );
not ( n337417 , n337416 );
buf ( n337418 , n17479 );
not ( n337419 , n337418 );
or ( n17560 , n337417 , n337419 );
buf ( n337421 , n337391 );
buf ( n337422 , n334786 );
nand ( n17563 , n337421 , n337422 );
buf ( n337424 , n17563 );
buf ( n337425 , n337424 );
nand ( n17566 , n17560 , n337425 );
buf ( n17567 , n17566 );
buf ( n337428 , n17567 );
and ( n17569 , n17555 , n337428 );
and ( n337430 , n337369 , n337414 );
or ( n337431 , n17569 , n337430 );
buf ( n337432 , n337431 );
buf ( n337433 , n337432 );
nand ( n337434 , n337358 , n337433 );
buf ( n337435 , n337434 );
buf ( n337436 , n337435 );
nand ( n337437 , n17493 , n337436 );
buf ( n337438 , n337437 );
buf ( n337439 , n337438 );
and ( n337440 , n17450 , n337439 );
and ( n337441 , n337283 , n17449 );
or ( n17582 , n337440 , n337441 );
buf ( n337443 , n17582 );
buf ( n337444 , n337443 );
buf ( n337445 , n336675 );
buf ( n337446 , n14891 );
and ( n337447 , n337445 , n337446 );
buf ( n337448 , n336689 );
nor ( n337449 , n337447 , n337448 );
buf ( n337450 , n337449 );
buf ( n337451 , n337450 );
not ( n337452 , n337451 );
buf ( n337453 , n336670 );
not ( n17594 , n337453 );
and ( n17595 , n337452 , n17594 );
buf ( n337456 , n336692 );
buf ( n337457 , n336670 );
and ( n337458 , n337456 , n337457 );
nor ( n17599 , n17595 , n337458 );
buf ( n337460 , n17599 );
or ( n17601 , n337460 , n16858 );
nand ( n17602 , n16858 , n337460 );
nand ( n337463 , n17601 , n17602 );
buf ( n337464 , n337463 );
xor ( n337465 , n337444 , n337464 );
buf ( n337466 , n15528 );
not ( n17607 , n337466 );
buf ( n337468 , n336746 );
not ( n337469 , n337468 );
or ( n337470 , n17607 , n337469 );
buf ( n337471 , n580 );
not ( n337472 , n337471 );
buf ( n337473 , n14644 );
not ( n337474 , n337473 );
or ( n17615 , n337472 , n337474 );
buf ( n17616 , n16201 );
buf ( n337477 , n334650 );
nand ( n337478 , n17616 , n337477 );
buf ( n337479 , n337478 );
buf ( n337480 , n337479 );
nand ( n17621 , n17615 , n337480 );
buf ( n337482 , n17621 );
buf ( n337483 , n337482 );
buf ( n17624 , n14822 );
nand ( n17625 , n337483 , n17624 );
buf ( n337486 , n17625 );
buf ( n337487 , n337486 );
nand ( n17628 , n337470 , n337487 );
buf ( n337489 , n17628 );
buf ( n337490 , n337489 );
and ( n337491 , n337465 , n337490 );
and ( n17632 , n337444 , n337464 );
or ( n337493 , n337491 , n17632 );
buf ( n337494 , n337493 );
xor ( n337495 , n336729 , n336763 );
xnor ( n337496 , n337495 , n16892 );
xor ( n17637 , n337494 , n337496 );
buf ( n337498 , n334694 );
not ( n337499 , n337498 );
buf ( n337500 , n336618 );
not ( n17641 , n337500 );
or ( n337502 , n337499 , n17641 );
buf ( n337503 , n582 );
not ( n337504 , n337503 );
buf ( n337505 , n335301 );
not ( n337506 , n337505 );
or ( n17647 , n337504 , n337506 );
buf ( n337508 , n335300 );
buf ( n337509 , n334702 );
nand ( n337510 , n337508 , n337509 );
buf ( n337511 , n337510 );
buf ( n337512 , n337511 );
nand ( n337513 , n17647 , n337512 );
buf ( n337514 , n337513 );
buf ( n337515 , n337514 );
buf ( n337516 , n334727 );
nand ( n17657 , n337515 , n337516 );
buf ( n337518 , n17657 );
buf ( n337519 , n337518 );
nand ( n337520 , n337502 , n337519 );
buf ( n337521 , n337520 );
and ( n17662 , n17637 , n337521 );
and ( n337523 , n337494 , n337496 );
or ( n337524 , n17662 , n337523 );
xor ( n17665 , n337277 , n337524 );
not ( n17666 , n16910 );
not ( n17667 , n16763 );
and ( n17668 , n17666 , n17667 );
and ( n17669 , n16763 , n16910 );
nor ( n337530 , n17668 , n17669 );
and ( n337531 , n337530 , n16789 );
not ( n17672 , n337530 );
and ( n337533 , n17672 , n16795 );
nor ( n337534 , n337531 , n337533 );
and ( n17675 , n17665 , n337534 );
and ( n17676 , n337277 , n337524 );
or ( n17677 , n17675 , n17676 );
buf ( n337538 , n17677 );
not ( n17679 , n337538 );
buf ( n337540 , n17679 );
nand ( n337541 , n17415 , n337540 );
not ( n17682 , n337541 );
buf ( n337543 , n15275 );
not ( n337544 , n337543 );
buf ( n337545 , n336840 );
not ( n337546 , n337545 );
buf ( n337547 , n337546 );
buf ( n337548 , n337547 );
not ( n337549 , n337548 );
or ( n17690 , n337544 , n337549 );
buf ( n337551 , n588 );
not ( n337552 , n16724 );
buf ( n337553 , n337552 );
and ( n337554 , n337551 , n337553 );
not ( n17695 , n337551 );
buf ( n337556 , n335261 );
and ( n17697 , n17695 , n337556 );
nor ( n17698 , n337554 , n17697 );
buf ( n337559 , n17698 );
buf ( n337560 , n337559 );
buf ( n337561 , n335114 );
nand ( n17702 , n337560 , n337561 );
buf ( n337563 , n17702 );
buf ( n337564 , n337563 );
nand ( n17705 , n17690 , n337564 );
buf ( n337566 , n17705 );
buf ( n337567 , n337566 );
not ( n17708 , n337567 );
buf ( n337569 , n15115 );
not ( n17710 , n337569 );
buf ( n337571 , n336832 );
not ( n17712 , n337571 );
or ( n17713 , n17710 , n17712 );
buf ( n337574 , n586 );
not ( n17715 , n337574 );
buf ( n337576 , n14898 );
not ( n17717 , n337576 );
or ( n17718 , n17715 , n17717 );
buf ( n337579 , n14254 );
buf ( n337580 , n334982 );
nand ( n17721 , n337579 , n337580 );
buf ( n337582 , n17721 );
buf ( n337583 , n337582 );
nand ( n17724 , n17718 , n337583 );
buf ( n337585 , n17724 );
buf ( n337586 , n337585 );
buf ( n337587 , n15164 );
nand ( n17728 , n337586 , n337587 );
buf ( n337589 , n17728 );
buf ( n337590 , n337589 );
nand ( n17731 , n17713 , n337590 );
buf ( n337592 , n17731 );
buf ( n337593 , n337592 );
not ( n17734 , n337593 );
or ( n17735 , n17708 , n17734 );
buf ( n337596 , n337566 );
buf ( n337597 , n337592 );
or ( n17738 , n337596 , n337597 );
xor ( n17739 , n337494 , n337496 );
xor ( n17740 , n17739 , n337521 );
not ( n17741 , n17740 );
not ( n17742 , n584 );
not ( n17743 , n15095 );
or ( n17744 , n17742 , n17743 );
or ( n17745 , n15095 , n584 );
nand ( n17746 , n17744 , n17745 );
not ( n17747 , n17746 );
not ( n17748 , n17747 );
not ( n17749 , n336786 );
and ( n17750 , n17748 , n17749 );
and ( n17751 , n336647 , n334868 );
nor ( n17752 , n17750 , n17751 );
buf ( n337613 , n17752 );
buf ( n337614 , n14941 );
not ( n17755 , n337614 );
buf ( n337616 , n336713 );
not ( n17757 , n337616 );
or ( n17758 , n17755 , n17757 );
not ( n17759 , n334415 );
not ( n17760 , n14552 );
or ( n17761 , n17759 , n17760 );
nand ( n17762 , n17761 , n14559 );
not ( n17763 , n17762 );
buf ( n337624 , n17763 );
not ( n17765 , n337624 );
buf ( n337626 , n17765 );
not ( n17767 , n337626 );
not ( n17768 , n334748 );
or ( n17769 , n17767 , n17768 );
nand ( n17770 , n336354 , n578 );
nand ( n17771 , n17769 , n17770 );
buf ( n337632 , n17771 );
buf ( n337633 , n14949 );
nand ( n17774 , n337632 , n337633 );
buf ( n337635 , n17774 );
buf ( n337636 , n337635 );
nand ( n17777 , n17758 , n337636 );
buf ( n337638 , n17777 );
buf ( n337639 , n337638 );
xor ( n17780 , n337283 , n17449 );
xor ( n17781 , n17780 , n337439 );
buf ( n337642 , n17781 );
buf ( n337643 , n337642 );
xor ( n17784 , n337639 , n337643 );
buf ( n337645 , n334643 );
not ( n17786 , n337645 );
buf ( n337647 , n337482 );
not ( n17788 , n337647 );
or ( n17789 , n17786 , n17788 );
not ( n17790 , n580 );
not ( n17791 , n336319 );
or ( n17792 , n17790 , n17791 );
buf ( n337653 , n14546 );
not ( n17794 , n337653 );
buf ( n337655 , n334650 );
nand ( n17796 , n17794 , n337655 );
buf ( n337657 , n17796 );
nand ( n17798 , n17792 , n337657 );
buf ( n337659 , n17798 );
buf ( n337660 , n14822 );
nand ( n17801 , n337659 , n337660 );
buf ( n337662 , n17801 );
buf ( n337663 , n337662 );
nand ( n17804 , n17789 , n337663 );
buf ( n337665 , n17804 );
buf ( n337666 , n337665 );
and ( n17807 , n17784 , n337666 );
and ( n17808 , n337639 , n337643 );
or ( n17809 , n17807 , n17808 );
buf ( n337670 , n17809 );
buf ( n337671 , n337670 );
buf ( n337672 , n334694 );
not ( n17813 , n337672 );
buf ( n337674 , n337514 );
not ( n17815 , n337674 );
or ( n17816 , n17813 , n17815 );
buf ( n337677 , n334727 );
buf ( n337678 , n14139 );
buf ( n17819 , n337678 );
buf ( n337680 , n17819 );
and ( n17821 , n337680 , n334702 );
not ( n17822 , n337680 );
and ( n17823 , n17822 , n582 );
or ( n17824 , n17821 , n17823 );
buf ( n337685 , n17824 );
nand ( n17826 , n337677 , n337685 );
buf ( n337687 , n17826 );
buf ( n337688 , n337687 );
nand ( n17829 , n17816 , n337688 );
buf ( n337690 , n17829 );
buf ( n337691 , n337690 );
xor ( n17832 , n337671 , n337691 );
xor ( n337693 , n337444 , n337464 );
xor ( n17834 , n337693 , n337490 );
buf ( n337695 , n17834 );
buf ( n337696 , n337695 );
and ( n337697 , n17832 , n337696 );
and ( n337698 , n337671 , n337691 );
or ( n17839 , n337697 , n337698 );
buf ( n337700 , n17839 );
buf ( n337701 , n337700 );
not ( n17842 , n337701 );
buf ( n337703 , n17842 );
buf ( n337704 , n337703 );
nand ( n337705 , n337613 , n337704 );
buf ( n337706 , n337705 );
not ( n17847 , n337706 );
or ( n337708 , n17741 , n17847 );
buf ( n337709 , n17752 );
not ( n337710 , n337709 );
buf ( n337711 , n337700 );
nand ( n17852 , n337710 , n337711 );
buf ( n17853 , n17852 );
nand ( n337714 , n337708 , n17853 );
buf ( n337715 , n337714 );
buf ( n337716 , n337715 );
buf ( n337717 , n337716 );
buf ( n337718 , n337717 );
nand ( n17859 , n17738 , n337718 );
buf ( n17860 , n17859 );
buf ( n337721 , n17860 );
nand ( n17862 , n17735 , n337721 );
buf ( n17863 , n17862 );
not ( n337724 , n17863 );
or ( n337725 , n17682 , n337724 );
not ( n337726 , n337540 );
nand ( n337727 , n337726 , n17414 );
nand ( n17868 , n337725 , n337727 );
buf ( n337729 , n17868 );
nand ( n337730 , n17399 , n337729 );
buf ( n337731 , n337730 );
buf ( n337732 , n17398 );
buf ( n337733 , n17395 );
nand ( n337734 , n337732 , n337733 );
buf ( n337735 , n337734 );
buf ( n337736 , n337735 );
and ( n337737 , n337731 , n337736 );
buf ( n337738 , n337737 );
nand ( n337739 , n17393 , n337738 );
buf ( n337740 , n337200 );
not ( n17881 , n337740 );
buf ( n337742 , n15275 );
not ( n17883 , n337742 );
buf ( n337744 , n337155 );
not ( n337745 , n337744 );
or ( n17886 , n17883 , n337745 );
buf ( n337747 , n337169 );
nand ( n337748 , n17886 , n337747 );
buf ( n337749 , n337748 );
buf ( n337750 , n337749 );
not ( n17891 , n337750 );
or ( n337752 , n17881 , n17891 );
buf ( n337753 , n337749 );
buf ( n337754 , n337200 );
or ( n17895 , n337753 , n337754 );
buf ( n337756 , n337140 );
nand ( n337757 , n17895 , n337756 );
buf ( n337758 , n337757 );
buf ( n337759 , n337758 );
nand ( n17900 , n337752 , n337759 );
buf ( n337761 , n17900 );
buf ( n337762 , n336111 );
buf ( n337763 , n336145 );
xor ( n337764 , n337762 , n337763 );
buf ( n337765 , n336127 );
xnor ( n337766 , n337764 , n337765 );
buf ( n337767 , n337766 );
buf ( n337768 , n334978 );
not ( n337769 , n337768 );
buf ( n337770 , n586 );
not ( n337771 , n337770 );
buf ( n337772 , n336868 );
not ( n17913 , n337772 );
or ( n337774 , n337771 , n17913 );
buf ( n337775 , n336865 );
buf ( n337776 , n334982 );
nand ( n337777 , n337775 , n337776 );
buf ( n337778 , n337777 );
buf ( n337779 , n337778 );
nand ( n337780 , n337774 , n337779 );
buf ( n337781 , n337780 );
buf ( n337782 , n337781 );
not ( n17923 , n337782 );
or ( n337784 , n337769 , n17923 );
buf ( n17925 , n15164 );
buf ( n17926 , n337190 );
nand ( n17927 , n17925 , n17926 );
buf ( n17928 , n17927 );
buf ( n337789 , n17928 );
nand ( n17930 , n337784 , n337789 );
buf ( n17931 , n17930 );
xor ( n337792 , n337767 , n17931 );
not ( n17933 , n15275 );
not ( n17934 , n17240 );
not ( n337795 , n334972 );
or ( n337796 , n17934 , n337795 );
not ( n17937 , n15341 );
nand ( n17938 , n17937 , n588 );
nand ( n337799 , n337796 , n17938 );
not ( n337800 , n337799 );
or ( n17941 , n17933 , n337800 );
buf ( n337802 , n337155 );
buf ( n337803 , n335114 );
nand ( n17944 , n337802 , n337803 );
buf ( n337805 , n17944 );
nand ( n337806 , n17941 , n337805 );
xor ( n17947 , n337792 , n337806 );
xor ( n17948 , n337761 , n17947 );
buf ( n337809 , n17155 );
not ( n17950 , n337809 );
buf ( n337811 , n17950 );
buf ( n337812 , n337811 );
not ( n17953 , n337812 );
buf ( n337814 , n17204 );
not ( n337815 , n337814 );
or ( n17956 , n17953 , n337815 );
buf ( n337817 , n17155 );
not ( n337818 , n337817 );
buf ( n337819 , n17204 );
not ( n17960 , n337819 );
buf ( n337821 , n17960 );
buf ( n337822 , n337821 );
not ( n17963 , n337822 );
or ( n337824 , n337818 , n17963 );
buf ( n337825 , n337076 );
nand ( n17966 , n337824 , n337825 );
buf ( n337827 , n17966 );
buf ( n17968 , n337827 );
nand ( n337829 , n17956 , n17968 );
buf ( n337830 , n337829 );
xnor ( n17971 , n17948 , n337830 );
not ( n337832 , n17971 );
buf ( n337833 , n337112 );
not ( n17974 , n337833 );
buf ( n337835 , n17974 );
buf ( n337836 , n337835 );
not ( n17977 , n337836 );
buf ( n337838 , n337203 );
not ( n17979 , n337838 );
or ( n17980 , n17977 , n17979 );
buf ( n337841 , n17389 );
nand ( n17982 , n17980 , n337841 );
buf ( n337843 , n17982 );
buf ( n337844 , n337206 );
buf ( n337845 , n337112 );
nand ( n17986 , n337844 , n337845 );
buf ( n337847 , n17986 );
nand ( n17988 , n337843 , n337847 );
not ( n17989 , n17988 );
xor ( n17990 , n17167 , n337038 );
and ( n17991 , n17990 , n337063 );
and ( n17992 , n17167 , n337038 );
or ( n17993 , n17991 , n17992 );
buf ( n337854 , n17993 );
xor ( n17995 , n337118 , n337131 );
and ( n17996 , n17995 , n337138 );
and ( n17997 , n337118 , n337131 );
or ( n17998 , n17996 , n17997 );
buf ( n337859 , n17998 );
buf ( n337860 , n337859 );
buf ( n337861 , n334694 );
not ( n18002 , n337861 );
buf ( n337863 , n336007 );
not ( n18004 , n337863 );
or ( n18005 , n18002 , n18004 );
buf ( n337866 , n17173 );
buf ( n337867 , n334727 );
nand ( n18008 , n337866 , n337867 );
buf ( n337869 , n18008 );
buf ( n337870 , n337869 );
nand ( n18011 , n18005 , n337870 );
buf ( n337872 , n18011 );
buf ( n337873 , n337872 );
xor ( n18014 , n337860 , n337873 );
buf ( n337875 , n334868 );
not ( n18016 , n337875 );
buf ( n337877 , n336037 );
not ( n18018 , n337877 );
or ( n18019 , n18016 , n18018 );
buf ( n337880 , n337056 );
buf ( n337881 , n334917 );
nand ( n18022 , n337880 , n337881 );
buf ( n337883 , n18022 );
buf ( n337884 , n337883 );
nand ( n18025 , n18019 , n337884 );
buf ( n337886 , n18025 );
buf ( n337887 , n337886 );
xor ( n18028 , n18014 , n337887 );
buf ( n337889 , n18028 );
buf ( n337890 , n337889 );
xor ( n18031 , n337854 , n337890 );
buf ( n337892 , n15264 );
not ( n18033 , n337892 );
buf ( n337894 , n18033 );
buf ( n337895 , n337894 );
not ( n18036 , n337895 );
buf ( n337897 , n335097 );
not ( n18038 , n337897 );
and ( n18039 , n18036 , n18038 );
buf ( n337900 , n15264 );
not ( n18041 , n337900 );
buf ( n337902 , n18041 );
buf ( n337903 , n337902 );
buf ( n337904 , n335097 );
and ( n18045 , n337903 , n337904 );
nor ( n18046 , n18039 , n18045 );
buf ( n337907 , n18046 );
buf ( n337908 , n337907 );
not ( n18049 , n337908 );
buf ( n337910 , n335177 );
not ( n18051 , n337910 );
and ( n18052 , n18049 , n18051 );
buf ( n337913 , n337092 );
buf ( n337914 , n335181 );
and ( n18055 , n337913 , n337914 );
nor ( n18056 , n18052 , n18055 );
buf ( n337917 , n18056 );
buf ( n337918 , n337917 );
xor ( n18059 , n18031 , n337918 );
buf ( n337920 , n18059 );
not ( n18061 , n337920 );
not ( n18062 , n18061 );
or ( n18063 , n17989 , n18062 );
not ( n18064 , n17988 );
nand ( n18065 , n18064 , n337920 );
nand ( n18066 , n18063 , n18065 );
not ( n18067 , n18066 );
or ( n18068 , n337832 , n18067 );
or ( n18069 , n18066 , n17971 );
nand ( n18070 , n18068 , n18069 );
xor ( n18071 , n17046 , n337079 );
and ( n18072 , n18071 , n337252 );
and ( n18073 , n17046 , n337079 );
or ( n18074 , n18072 , n18073 );
nand ( n18075 , n18070 , n18074 );
and ( n18076 , n337739 , n18075 );
not ( n18077 , n18076 );
buf ( n337938 , n334643 );
not ( n18079 , n337938 );
and ( n18080 , n336463 , n334650 );
not ( n18081 , n336463 );
and ( n18082 , n18081 , n580 );
or ( n18083 , n18080 , n18082 );
buf ( n337944 , n18083 );
not ( n18085 , n337944 );
or ( n18086 , n18079 , n18085 );
buf ( n337947 , n580 );
not ( n18088 , n337947 );
buf ( n337949 , n336354 );
not ( n18090 , n337949 );
or ( n18091 , n18088 , n18090 );
buf ( n337952 , n336357 );
buf ( n337953 , n334650 );
nand ( n18094 , n337952 , n337953 );
buf ( n337955 , n18094 );
buf ( n337956 , n337955 );
nand ( n18097 , n18091 , n337956 );
buf ( n337958 , n18097 );
buf ( n337959 , n337958 );
buf ( n337960 , n14822 );
nand ( n18101 , n337959 , n337960 );
buf ( n337962 , n18101 );
buf ( n337963 , n337962 );
nand ( n18104 , n18086 , n337963 );
buf ( n337965 , n18104 );
buf ( n337966 , n337965 );
xor ( n18107 , n337369 , n337414 );
xor ( n18108 , n18107 , n337428 );
buf ( n337969 , n18108 );
buf ( n337970 , n337969 );
buf ( n337971 , n335432 );
not ( n18112 , n337971 );
buf ( n337973 , n578 );
not ( n18114 , n337973 );
buf ( n337975 , n336681 );
not ( n18116 , n337975 );
or ( n18117 , n18114 , n18116 );
buf ( n337978 , n16430 );
buf ( n337979 , n334748 );
nand ( n18120 , n337978 , n337979 );
buf ( n337981 , n18120 );
buf ( n337982 , n337981 );
nand ( n18123 , n18117 , n337982 );
buf ( n337984 , n18123 );
buf ( n337985 , n337984 );
not ( n18126 , n337985 );
or ( n18127 , n18112 , n18126 );
buf ( n337988 , n16799 );
buf ( n18129 , n337988 );
buf ( n337990 , n18129 );
nand ( n18131 , n337990 , n578 );
not ( n18132 , n337990 );
nand ( n18133 , n18132 , n334748 );
nand ( n18134 , n14949 , n18131 , n18133 );
buf ( n337995 , n18134 );
nand ( n18136 , n18127 , n337995 );
buf ( n337997 , n18136 );
buf ( n337998 , n337997 );
xor ( n18139 , n337970 , n337998 );
xor ( n18140 , n337410 , n17533 );
buf ( n338001 , n18140 );
buf ( n338002 , n14941 );
not ( n18143 , n338002 );
and ( n18144 , n337278 , n334748 );
not ( n18145 , n337278 );
and ( n18146 , n18145 , n578 );
or ( n18147 , n18144 , n18146 );
buf ( n338008 , n18147 );
not ( n18149 , n338008 );
or ( n18150 , n18143 , n18149 );
buf ( n338011 , n578 );
not ( n18152 , n338011 );
buf ( n338013 , n334002 );
not ( n18154 , n338013 );
buf ( n338015 , n18154 );
buf ( n338016 , n338015 );
not ( n18157 , n338016 );
or ( n18158 , n18152 , n18157 );
buf ( n338019 , n17456 );
buf ( n338020 , n334748 );
nand ( n18161 , n338019 , n338020 );
buf ( n338022 , n18161 );
buf ( n338023 , n338022 );
nand ( n18164 , n18158 , n338023 );
buf ( n338025 , n18164 );
buf ( n338026 , n338025 );
buf ( n338027 , n14949 );
nand ( n338028 , n338026 , n338027 );
buf ( n338029 , n338028 );
buf ( n338030 , n338029 );
nand ( n18171 , n18150 , n338030 );
buf ( n338032 , n18171 );
buf ( n338033 , n338032 );
buf ( n338034 , n579 );
buf ( n338035 , n580 );
or ( n18176 , n338034 , n338035 );
buf ( n338037 , n337364 );
nand ( n18178 , n18176 , n338037 );
buf ( n338039 , n18178 );
buf ( n338040 , n338039 );
buf ( n338041 , n579 );
buf ( n338042 , n580 );
and ( n18183 , n338041 , n338042 );
buf ( n338044 , n334748 );
nor ( n18185 , n18183 , n338044 );
buf ( n338046 , n18185 );
buf ( n338047 , n338046 );
nand ( n18188 , n338040 , n338047 );
buf ( n338049 , n18188 );
buf ( n338050 , n338049 );
not ( n18191 , n338050 );
buf ( n338052 , n18191 );
buf ( n338053 , n338052 );
not ( n18194 , n338053 );
buf ( n338055 , n14941 );
not ( n18196 , n338055 );
buf ( n338057 , n338025 );
not ( n18198 , n338057 );
or ( n18199 , n18196 , n18198 );
buf ( n338060 , n334748 );
buf ( n338061 , n337364 );
or ( n18202 , n338060 , n338061 );
buf ( n338063 , n578 );
buf ( n338064 , n337361 );
or ( n18205 , n338063 , n338064 );
nand ( n18206 , n18202 , n18205 );
buf ( n338067 , n18206 );
buf ( n338068 , n338067 );
buf ( n338069 , n14949 );
nand ( n18210 , n338068 , n338069 );
buf ( n338071 , n18210 );
buf ( n338072 , n338071 );
nand ( n18213 , n18199 , n338072 );
buf ( n338074 , n18213 );
buf ( n338075 , n338074 );
not ( n18216 , n338075 );
or ( n18217 , n18194 , n18216 );
buf ( n338078 , n337364 );
buf ( n338079 , n14891 );
nand ( n338080 , n338078 , n338079 );
buf ( n338081 , n338080 );
buf ( n338082 , n338081 );
nand ( n18223 , n18217 , n338082 );
buf ( n338084 , n18223 );
buf ( n338085 , n338084 );
and ( n338086 , n338033 , n338085 );
buf ( n338087 , n338086 );
buf ( n338088 , n338087 );
xor ( n18229 , n338001 , n338088 );
nand ( n338090 , n18131 , n18133 );
buf ( n338091 , n338090 );
buf ( n338092 , n335432 );
not ( n338093 , n338092 );
buf ( n338094 , n338093 );
buf ( n338095 , n338094 );
or ( n338096 , n338091 , n338095 );
buf ( n338097 , n18147 );
buf ( n338098 , n14949 );
nand ( n338099 , n338097 , n338098 );
buf ( n338100 , n338099 );
buf ( n338101 , n338100 );
nand ( n18242 , n338096 , n338101 );
buf ( n338103 , n18242 );
buf ( n338104 , n338103 );
and ( n338105 , n18229 , n338104 );
and ( n18246 , n338001 , n338088 );
or ( n18247 , n338105 , n18246 );
buf ( n338108 , n18247 );
buf ( n338109 , n338108 );
xor ( n18250 , n18139 , n338109 );
buf ( n338111 , n18250 );
buf ( n338112 , n338111 );
xor ( n18253 , n337966 , n338112 );
buf ( n338114 , n334694 );
not ( n338115 , n338114 );
buf ( n338116 , n582 );
not ( n338117 , n338116 );
buf ( n338118 , n336064 );
not ( n338119 , n338118 );
or ( n18260 , n338117 , n338119 );
buf ( n338121 , n336067 );
buf ( n338122 , n334702 );
nand ( n18263 , n338121 , n338122 );
buf ( n338124 , n18263 );
buf ( n338125 , n338124 );
nand ( n18266 , n18260 , n338125 );
buf ( n18267 , n18266 );
buf ( n338128 , n18267 );
not ( n18269 , n338128 );
or ( n338130 , n338115 , n18269 );
and ( n338131 , n336319 , n582 );
not ( n338132 , n336319 );
and ( n338133 , n338132 , n334702 );
or ( n18274 , n338131 , n338133 );
buf ( n18275 , n18274 );
buf ( n338136 , n334727 );
nand ( n338137 , n18275 , n338136 );
buf ( n338138 , n338137 );
buf ( n338139 , n338138 );
nand ( n18280 , n338130 , n338139 );
buf ( n338141 , n18280 );
buf ( n338142 , n338141 );
and ( n338143 , n18253 , n338142 );
and ( n18284 , n337966 , n338112 );
or ( n338145 , n338143 , n18284 );
buf ( n338146 , n338145 );
buf ( n338147 , n338146 );
buf ( n338148 , n334868 );
not ( n338149 , n338148 );
buf ( n338150 , n584 );
not ( n18291 , n338150 );
buf ( n338152 , n335301 );
not ( n18293 , n338152 );
or ( n338154 , n18291 , n18293 );
buf ( n338155 , n335300 );
buf ( n338156 , n334879 );
nand ( n338157 , n338155 , n338156 );
buf ( n338158 , n338157 );
buf ( n338159 , n338158 );
nand ( n338160 , n338154 , n338159 );
buf ( n338161 , n338160 );
buf ( n338162 , n338161 );
not ( n338163 , n338162 );
or ( n338164 , n338149 , n338163 );
buf ( n338165 , n584 );
not ( n338166 , n338165 );
buf ( n338167 , n337680 );
not ( n18308 , n338167 );
buf ( n18309 , n18308 );
buf ( n338170 , n18309 );
not ( n18311 , n338170 );
or ( n18312 , n338166 , n18311 );
buf ( n338173 , n337680 );
buf ( n338174 , n334879 );
nand ( n18315 , n338173 , n338174 );
buf ( n338176 , n18315 );
buf ( n338177 , n338176 );
nand ( n18318 , n18312 , n338177 );
buf ( n18319 , n18318 );
buf ( n338180 , n18319 );
buf ( n338181 , n334917 );
nand ( n338182 , n338180 , n338181 );
buf ( n338183 , n338182 );
buf ( n338184 , n338183 );
nand ( n338185 , n338164 , n338184 );
buf ( n338186 , n338185 );
buf ( n338187 , n338186 );
xor ( n18328 , n338147 , n338187 );
xor ( n338189 , n337970 , n337998 );
and ( n338190 , n338189 , n338109 );
and ( n18331 , n337970 , n337998 );
or ( n338192 , n338190 , n18331 );
buf ( n338193 , n338192 );
buf ( n338194 , n338193 );
and ( n338195 , n337432 , n337320 );
not ( n338196 , n337432 );
and ( n338197 , n338196 , n337323 );
or ( n338198 , n338195 , n338197 );
buf ( n338199 , n338198 );
buf ( n338200 , n337347 );
and ( n338201 , n338199 , n338200 );
not ( n18342 , n338199 );
buf ( n18343 , n337350 );
and ( n18344 , n18342 , n18343 );
nor ( n338205 , n338201 , n18344 );
buf ( n338206 , n338205 );
buf ( n338207 , n338206 );
not ( n338208 , n338207 );
buf ( n338209 , n338208 );
buf ( n338210 , n338209 );
not ( n338211 , n338210 );
not ( n18352 , n14941 );
not ( n18353 , n17771 );
or ( n18354 , n18352 , n18353 );
buf ( n338215 , n337984 );
buf ( n338216 , n14949 );
nand ( n18357 , n338215 , n338216 );
buf ( n338218 , n18357 );
nand ( n18359 , n18354 , n338218 );
buf ( n338220 , n18359 );
not ( n338221 , n338220 );
buf ( n338222 , n338221 );
buf ( n338223 , n338222 );
not ( n18364 , n338223 );
or ( n18365 , n338211 , n18364 );
nand ( n338226 , n18359 , n338206 );
buf ( n338227 , n338226 );
nand ( n338228 , n18365 , n338227 );
buf ( n338229 , n338228 );
buf ( n338230 , n338229 );
xor ( n338231 , n338194 , n338230 );
and ( n338232 , n17798 , n14782 );
and ( n18373 , n18083 , n14822 );
nor ( n338234 , n338232 , n18373 );
buf ( n338235 , n338234 );
buf ( n338236 , n338235 );
xnor ( n18377 , n338231 , n338236 );
buf ( n338238 , n18377 );
buf ( n338239 , n18267 );
not ( n18380 , n338239 );
buf ( n338241 , n18380 );
buf ( n338242 , n338241 );
not ( n338243 , n338242 );
buf ( n338244 , n336910 );
not ( n338245 , n338244 );
and ( n338246 , n338243 , n338245 );
buf ( n338247 , n582 );
not ( n338248 , n338247 );
buf ( n338249 , n335326 );
not ( n18390 , n338249 );
or ( n338251 , n338248 , n18390 );
buf ( n338252 , n15463 );
buf ( n338253 , n334702 );
nand ( n18394 , n338252 , n338253 );
buf ( n338255 , n18394 );
buf ( n338256 , n338255 );
nand ( n338257 , n338251 , n338256 );
buf ( n338258 , n338257 );
buf ( n338259 , n338258 );
buf ( n338260 , n334694 );
and ( n18401 , n338259 , n338260 );
nor ( n338262 , n338246 , n18401 );
buf ( n338263 , n338262 );
xnor ( n18404 , n338238 , n338263 );
buf ( n338265 , n18404 );
xor ( n18406 , n18328 , n338265 );
buf ( n338267 , n18406 );
xor ( n18408 , n338001 , n338088 );
xor ( n338269 , n18408 , n338104 );
buf ( n338270 , n338269 );
buf ( n338271 , n338270 );
buf ( n338272 , n334643 );
not ( n338273 , n338272 );
buf ( n338274 , n337958 );
not ( n338275 , n338274 );
or ( n18416 , n338273 , n338275 );
buf ( n338277 , n580 );
not ( n18418 , n338277 );
buf ( n338279 , n336681 );
not ( n18420 , n338279 );
or ( n338281 , n18418 , n18420 );
buf ( n338282 , n334650 );
buf ( n338283 , n16430 );
nand ( n338284 , n338282 , n338283 );
buf ( n338285 , n338284 );
buf ( n338286 , n338285 );
nand ( n338287 , n338281 , n338286 );
buf ( n338288 , n338287 );
buf ( n338289 , n338288 );
buf ( n338290 , n14822 );
nand ( n338291 , n338289 , n338290 );
buf ( n338292 , n338291 );
buf ( n338293 , n338292 );
nand ( n338294 , n18416 , n338293 );
buf ( n338295 , n338294 );
buf ( n338296 , n338295 );
xor ( n18437 , n338271 , n338296 );
buf ( n338298 , n334694 );
not ( n18439 , n338298 );
buf ( n338300 , n18274 );
not ( n18441 , n338300 );
or ( n338302 , n18439 , n18441 );
buf ( n338303 , n582 );
not ( n18444 , n338303 );
buf ( n338305 , n16843 );
not ( n18446 , n338305 );
or ( n338307 , n18444 , n18446 );
buf ( n338308 , n336463 );
buf ( n338309 , n334702 );
nand ( n338310 , n338308 , n338309 );
buf ( n338311 , n338310 );
buf ( n338312 , n338311 );
nand ( n338313 , n338307 , n338312 );
buf ( n338314 , n338313 );
buf ( n18455 , n338314 );
buf ( n338316 , n334727 );
nand ( n338317 , n18455 , n338316 );
buf ( n338318 , n338317 );
buf ( n338319 , n338318 );
nand ( n18460 , n338302 , n338319 );
buf ( n338321 , n18460 );
buf ( n338322 , n338321 );
and ( n18463 , n18437 , n338322 );
and ( n338324 , n338271 , n338296 );
or ( n338325 , n18463 , n338324 );
buf ( n338326 , n338325 );
buf ( n338327 , n338326 );
buf ( n338328 , n334868 );
not ( n338329 , n338328 );
buf ( n338330 , n18319 );
not ( n18471 , n338330 );
or ( n338332 , n338329 , n18471 );
buf ( n338333 , n584 );
not ( n338334 , n338333 );
buf ( n338335 , n335329 );
not ( n338336 , n338335 );
or ( n338337 , n338334 , n338336 );
buf ( n338338 , n15463 );
buf ( n338339 , n334879 );
nand ( n338340 , n338338 , n338339 );
buf ( n338341 , n338340 );
buf ( n338342 , n338341 );
nand ( n338343 , n338337 , n338342 );
buf ( n338344 , n338343 );
buf ( n338345 , n338344 );
buf ( n338346 , n334914 );
nand ( n338347 , n338345 , n338346 );
buf ( n338348 , n338347 );
buf ( n338349 , n338348 );
nand ( n338350 , n338332 , n338349 );
buf ( n338351 , n338350 );
buf ( n338352 , n338351 );
xor ( n18493 , n338327 , n338352 );
xor ( n338354 , n337966 , n338112 );
xor ( n18495 , n338354 , n338142 );
buf ( n338356 , n18495 );
buf ( n338357 , n338356 );
and ( n338358 , n18493 , n338357 );
and ( n18499 , n338327 , n338352 );
or ( n338360 , n338358 , n18499 );
buf ( n338361 , n338360 );
buf ( n338362 , n338361 );
not ( n18503 , n338362 );
buf ( n338364 , n15163 );
not ( n338365 , n338364 );
buf ( n338366 , n586 );
not ( n18507 , n338366 );
buf ( n338368 , n335361 );
not ( n338369 , n338368 );
buf ( n338370 , n338369 );
buf ( n338371 , n338370 );
not ( n338372 , n338371 );
or ( n18513 , n18507 , n338372 );
buf ( n338374 , n335361 );
buf ( n338375 , n334982 );
nand ( n18516 , n338374 , n338375 );
buf ( n338377 , n18516 );
buf ( n338378 , n338377 );
nand ( n18519 , n18513 , n338378 );
buf ( n338380 , n18519 );
buf ( n338381 , n338380 );
not ( n18522 , n338381 );
or ( n338383 , n338365 , n18522 );
buf ( n338384 , n586 );
not ( n338385 , n338384 );
buf ( n338386 , n15095 );
not ( n18527 , n338386 );
or ( n338388 , n338385 , n18527 );
buf ( n338389 , n15096 );
buf ( n338390 , n334982 );
nand ( n338391 , n338389 , n338390 );
buf ( n338392 , n338391 );
buf ( n338393 , n338392 );
nand ( n338394 , n338388 , n338393 );
buf ( n338395 , n338394 );
buf ( n18536 , n338395 );
buf ( n338397 , n15115 );
nand ( n338398 , n18536 , n338397 );
buf ( n338399 , n338398 );
buf ( n338400 , n338399 );
nand ( n338401 , n338383 , n338400 );
buf ( n338402 , n338401 );
buf ( n338403 , n338402 );
not ( n18544 , n338403 );
buf ( n18545 , n18544 );
buf ( n338406 , n18545 );
nand ( n338407 , n18503 , n338406 );
buf ( n338408 , n338407 );
and ( n338409 , n338267 , n338408 );
and ( n18550 , n338402 , n338361 );
nor ( n338411 , n338409 , n18550 );
buf ( n338412 , n338411 );
buf ( n338413 , n588 );
buf ( n338414 , n17055 );
and ( n338415 , n338413 , n338414 );
not ( n18556 , n338413 );
buf ( n338417 , n15622 );
and ( n338418 , n18556 , n338417 );
nor ( n18559 , n338415 , n338418 );
buf ( n18560 , n18559 );
buf ( n338421 , n18560 );
not ( n18562 , n338421 );
buf ( n338423 , n18562 );
buf ( n18564 , n338423 );
not ( n18565 , n18564 );
buf ( n338426 , n335111 );
not ( n338427 , n338426 );
and ( n18568 , n18565 , n338427 );
buf ( n338429 , n334972 );
not ( n338430 , n338429 );
buf ( n338431 , n14897 );
not ( n18572 , n338431 );
or ( n338433 , n338430 , n18572 );
buf ( n338434 , n14898 );
buf ( n338435 , n588 );
nand ( n338436 , n338434 , n338435 );
buf ( n338437 , n338436 );
buf ( n338438 , n338437 );
nand ( n338439 , n338433 , n338438 );
buf ( n338440 , n338439 );
buf ( n338441 , n338440 );
buf ( n338442 , n15275 );
and ( n338443 , n338441 , n338442 );
nor ( n338444 , n18568 , n338443 );
buf ( n338445 , n338444 );
buf ( n338446 , n338445 );
xor ( n338447 , n338412 , n338446 );
not ( n18588 , n335097 );
not ( n338449 , n16686 );
or ( n18590 , n18588 , n338449 );
or ( n18591 , n16686 , n335097 );
nand ( n338452 , n18590 , n18591 );
buf ( n338453 , n338452 );
not ( n18594 , n338453 );
buf ( n338455 , n335181 );
not ( n18596 , n338455 );
buf ( n338457 , n18596 );
buf ( n338458 , n338457 );
not ( n338459 , n338458 );
and ( n338460 , n18594 , n338459 );
and ( n18601 , n335261 , n590 );
not ( n18602 , n335261 );
and ( n338463 , n18602 , n335097 );
or ( n18604 , n18601 , n338463 );
buf ( n338465 , n18604 );
buf ( n338466 , n591 );
and ( n338467 , n338465 , n338466 );
nor ( n18608 , n338460 , n338467 );
buf ( n18609 , n18608 );
buf ( n338470 , n18609 );
xor ( n18611 , n338447 , n338470 );
buf ( n338472 , n18611 );
buf ( n18613 , n338472 );
not ( n338474 , n18613 );
buf ( n338475 , n338474 );
buf ( n338476 , n338475 );
not ( n338477 , n338476 );
buf ( n338478 , n338361 );
buf ( n338479 , n18545 );
xor ( n338480 , n338478 , n338479 );
buf ( n338481 , n338267 );
xnor ( n18622 , n338480 , n338481 );
buf ( n338483 , n18622 );
buf ( n338484 , n15115 );
not ( n338485 , n338484 );
buf ( n338486 , n338380 );
not ( n18627 , n338486 );
or ( n338488 , n338485 , n18627 );
buf ( n338489 , n586 );
not ( n18630 , n338489 );
buf ( n338491 , n335301 );
not ( n18632 , n338491 );
or ( n338493 , n18630 , n18632 );
buf ( n338494 , n335300 );
buf ( n338495 , n334982 );
nand ( n338496 , n338494 , n338495 );
buf ( n338497 , n338496 );
buf ( n338498 , n338497 );
nand ( n338499 , n338493 , n338498 );
buf ( n338500 , n338499 );
buf ( n338501 , n338500 );
buf ( n338502 , n15163 );
nand ( n338503 , n338501 , n338502 );
buf ( n338504 , n338503 );
buf ( n338505 , n338504 );
nand ( n338506 , n338488 , n338505 );
buf ( n338507 , n338506 );
buf ( n338508 , n338507 );
not ( n338509 , n338508 );
buf ( n338510 , n338509 );
not ( n18651 , n338510 );
xor ( n338512 , n338084 , n338032 );
buf ( n338513 , n338512 );
buf ( n338514 , n334643 );
not ( n338515 , n338514 );
buf ( n338516 , n338288 );
not ( n338517 , n338516 );
or ( n338518 , n338515 , n338517 );
buf ( n338519 , n580 );
not ( n338520 , n338519 );
buf ( n338521 , n336662 );
not ( n338522 , n338521 );
or ( n18663 , n338520 , n338522 );
buf ( n338524 , n16799 );
buf ( n338525 , n334650 );
nand ( n18666 , n338524 , n338525 );
buf ( n18667 , n18666 );
buf ( n338528 , n18667 );
nand ( n338529 , n18663 , n338528 );
buf ( n338530 , n338529 );
buf ( n338531 , n338530 );
buf ( n338532 , n14822 );
nand ( n18673 , n338531 , n338532 );
buf ( n18674 , n18673 );
buf ( n338535 , n18674 );
nand ( n18676 , n338518 , n338535 );
buf ( n338537 , n18676 );
buf ( n338538 , n338537 );
xor ( n18679 , n338513 , n338538 );
buf ( n338540 , n338049 );
not ( n18681 , n338540 );
buf ( n338542 , n338074 );
not ( n338543 , n338542 );
or ( n18684 , n18681 , n338543 );
buf ( n338545 , n338074 );
buf ( n338546 , n338049 );
or ( n338547 , n338545 , n338546 );
nand ( n18688 , n18684 , n338547 );
buf ( n18689 , n18688 );
buf ( n18690 , n18689 );
buf ( n338551 , n334643 );
not ( n18692 , n338551 );
buf ( n338553 , n580 );
not ( n338554 , n338553 );
buf ( n338555 , n337332 );
not ( n338556 , n338555 );
or ( n338557 , n338554 , n338556 );
buf ( n338558 , n334650 );
buf ( n338559 , n337278 );
nand ( n18700 , n338558 , n338559 );
buf ( n338561 , n18700 );
buf ( n338562 , n338561 );
nand ( n18703 , n338557 , n338562 );
buf ( n338564 , n18703 );
buf ( n338565 , n338564 );
not ( n338566 , n338565 );
or ( n338567 , n18692 , n338566 );
and ( n18708 , n337384 , n580 );
not ( n18709 , n337384 );
and ( n18710 , n18709 , n334650 );
or ( n18711 , n18708 , n18710 );
buf ( n338572 , n18711 );
buf ( n338573 , n14822 );
nand ( n338574 , n338572 , n338573 );
buf ( n338575 , n338574 );
buf ( n338576 , n338575 );
nand ( n338577 , n338567 , n338576 );
buf ( n338578 , n338577 );
buf ( n338579 , n338578 );
buf ( n338580 , n581 );
buf ( n338581 , n582 );
or ( n18722 , n338580 , n338581 );
buf ( n338583 , n337364 );
nand ( n18724 , n18722 , n338583 );
buf ( n338585 , n18724 );
buf ( n338586 , n338585 );
buf ( n338587 , n581 );
buf ( n338588 , n582 );
and ( n18729 , n338587 , n338588 );
buf ( n338590 , n334650 );
nor ( n338591 , n18729 , n338590 );
buf ( n338592 , n338591 );
buf ( n338593 , n338592 );
and ( n338594 , n338586 , n338593 );
buf ( n338595 , n338594 );
buf ( n338596 , n338595 );
not ( n338597 , n338596 );
buf ( n338598 , n334643 );
not ( n18739 , n338598 );
buf ( n338600 , n18711 );
not ( n338601 , n338600 );
or ( n18742 , n18739 , n338601 );
buf ( n338603 , n334650 );
buf ( n338604 , n337364 );
or ( n18745 , n338603 , n338604 );
buf ( n338606 , n580 );
buf ( n338607 , n337361 );
or ( n18748 , n338606 , n338607 );
nand ( n338609 , n18745 , n18748 );
buf ( n338610 , n338609 );
buf ( n338611 , n338610 );
buf ( n338612 , n14822 );
nand ( n18753 , n338611 , n338612 );
buf ( n338614 , n18753 );
buf ( n338615 , n338614 );
nand ( n338616 , n18742 , n338615 );
buf ( n338617 , n338616 );
buf ( n338618 , n338617 );
not ( n18759 , n338618 );
or ( n338620 , n338597 , n18759 );
buf ( n338621 , n335432 );
buf ( n338622 , n337364 );
nand ( n338623 , n338621 , n338622 );
buf ( n338624 , n338623 );
buf ( n338625 , n338624 );
nand ( n338626 , n338620 , n338625 );
buf ( n338627 , n338626 );
buf ( n18768 , n338627 );
and ( n18769 , n338579 , n18768 );
buf ( n18770 , n18769 );
buf ( n338631 , n18770 );
xor ( n18772 , n18690 , n338631 );
buf ( n338633 , n334643 );
not ( n338634 , n338633 );
buf ( n338635 , n338530 );
not ( n18776 , n338635 );
or ( n338637 , n338634 , n18776 );
buf ( n338638 , n338564 );
buf ( n338639 , n14822 );
nand ( n338640 , n338638 , n338639 );
buf ( n338641 , n338640 );
buf ( n338642 , n338641 );
nand ( n338643 , n338637 , n338642 );
buf ( n338644 , n338643 );
buf ( n338645 , n338644 );
and ( n338646 , n18772 , n338645 );
and ( n338647 , n18690 , n338631 );
or ( n18788 , n338646 , n338647 );
buf ( n338649 , n18788 );
buf ( n338650 , n338649 );
and ( n18791 , n18679 , n338650 );
and ( n338652 , n338513 , n338538 );
or ( n338653 , n18791 , n338652 );
buf ( n338654 , n338653 );
xor ( n18795 , n338271 , n338296 );
xor ( n338656 , n18795 , n338322 );
buf ( n338657 , n338656 );
xor ( n18798 , n338654 , n338657 );
buf ( n338659 , n334868 );
not ( n338660 , n338659 );
buf ( n338661 , n338344 );
not ( n338662 , n338661 );
or ( n338663 , n338660 , n338662 );
buf ( n338664 , n584 );
not ( n338665 , n338664 );
buf ( n338666 , n336064 );
not ( n18807 , n338666 );
or ( n338668 , n338665 , n18807 );
buf ( n338669 , n336067 );
buf ( n338670 , n334879 );
nand ( n18811 , n338669 , n338670 );
buf ( n338672 , n18811 );
buf ( n338673 , n338672 );
nand ( n338674 , n338668 , n338673 );
buf ( n338675 , n338674 );
buf ( n338676 , n338675 );
buf ( n338677 , n334914 );
nand ( n18818 , n338676 , n338677 );
buf ( n18819 , n18818 );
buf ( n338680 , n18819 );
nand ( n18821 , n338663 , n338680 );
buf ( n338682 , n18821 );
and ( n18823 , n18798 , n338682 );
and ( n338684 , n338654 , n338657 );
or ( n338685 , n18823 , n338684 );
not ( n18826 , n338685 );
not ( n18827 , n18826 );
and ( n18828 , n18651 , n18827 );
nand ( n338689 , n338510 , n18826 );
xor ( n338690 , n338327 , n338352 );
xor ( n18831 , n338690 , n338357 );
buf ( n18832 , n18831 );
and ( n338693 , n338689 , n18832 );
nor ( n18834 , n18828 , n338693 );
buf ( n338695 , n15275 );
not ( n338696 , n338695 );
buf ( n338697 , n18560 );
not ( n338698 , n338697 );
or ( n18839 , n338696 , n338698 );
buf ( n338700 , n335111 );
not ( n338701 , n338700 );
buf ( n338702 , n588 );
not ( n338703 , n338702 );
buf ( n338704 , n14877 );
not ( n18845 , n338704 );
or ( n18846 , n338703 , n18845 );
not ( n18847 , n335434 );
nand ( n18848 , n18847 , n334972 );
buf ( n338709 , n18848 );
nand ( n18850 , n18846 , n338709 );
buf ( n338711 , n18850 );
buf ( n338712 , n338711 );
nand ( n18853 , n338701 , n338712 );
buf ( n338714 , n18853 );
buf ( n338715 , n338714 );
nand ( n338716 , n18839 , n338715 );
buf ( n338717 , n338716 );
buf ( n338718 , n338717 );
not ( n338719 , n338718 );
buf ( n338720 , n338719 );
nand ( n338721 , n18834 , n338720 );
and ( n338722 , n338483 , n338721 );
not ( n338723 , n18834 );
buf ( n338724 , n338723 );
not ( n338725 , n338724 );
buf ( n338726 , n338720 );
nor ( n18867 , n338725 , n338726 );
buf ( n18868 , n18867 );
nor ( n18869 , n338722 , n18868 );
buf ( n338730 , n18869 );
not ( n338731 , n338730 );
xor ( n338732 , n338147 , n338187 );
and ( n18873 , n338732 , n338265 );
and ( n338734 , n338147 , n338187 );
or ( n338735 , n18873 , n338734 );
buf ( n338736 , n338735 );
buf ( n338737 , n338736 );
buf ( n338738 , n15115 );
not ( n338739 , n338738 );
buf ( n338740 , n586 );
not ( n338741 , n338740 );
buf ( n338742 , n14877 );
not ( n18883 , n338742 );
or ( n18884 , n338741 , n18883 );
buf ( n18885 , n334736 );
buf ( n338746 , n334982 );
nand ( n18887 , n18885 , n338746 );
buf ( n338748 , n18887 );
buf ( n338749 , n338748 );
nand ( n18890 , n18884 , n338749 );
buf ( n338751 , n18890 );
buf ( n338752 , n338751 );
not ( n18893 , n338752 );
or ( n338754 , n338739 , n18893 );
buf ( n338755 , n338395 );
buf ( n338756 , n15163 );
nand ( n338757 , n338755 , n338756 );
buf ( n338758 , n338757 );
buf ( n338759 , n338758 );
nand ( n338760 , n338754 , n338759 );
buf ( n338761 , n338760 );
buf ( n338762 , n338761 );
xor ( n338763 , n338737 , n338762 );
buf ( n338764 , n338229 );
not ( n338765 , n338764 );
buf ( n338766 , n338235 );
not ( n338767 , n338766 );
or ( n18908 , n338765 , n338767 );
buf ( n338769 , n338229 );
buf ( n338770 , n338235 );
or ( n18911 , n338769 , n338770 );
nand ( n338772 , n18908 , n18911 );
buf ( n338773 , n338772 );
not ( n338774 , n338773 );
buf ( n338775 , n338263 );
buf ( n338776 , n338193 );
not ( n18917 , n338776 );
buf ( n338778 , n18917 );
buf ( n338779 , n338778 );
nand ( n338780 , n338775 , n338779 );
buf ( n338781 , n338780 );
not ( n338782 , n338781 );
or ( n18923 , n338774 , n338782 );
or ( n18924 , n338263 , n338778 );
nand ( n338785 , n18923 , n18924 );
not ( n338786 , n338785 );
buf ( n338787 , n338786 );
not ( n338788 , n334868 );
buf ( n338789 , n584 );
not ( n18930 , n338789 );
buf ( n338791 , n338370 );
not ( n18932 , n338791 );
or ( n338793 , n18930 , n18932 );
buf ( n338794 , n335355 );
not ( n18935 , n338794 );
buf ( n338796 , n334879 );
nand ( n18937 , n18935 , n338796 );
buf ( n338798 , n18937 );
buf ( n338799 , n338798 );
nand ( n18940 , n338793 , n338799 );
buf ( n338801 , n18940 );
not ( n18942 , n338801 );
or ( n338803 , n338788 , n18942 );
buf ( n338804 , n338161 );
buf ( n338805 , n334917 );
nand ( n18946 , n338804 , n338805 );
buf ( n338807 , n18946 );
nand ( n338808 , n338803 , n338807 );
buf ( n18949 , n338808 );
xor ( n18950 , n338787 , n18949 );
buf ( n338811 , n338222 );
not ( n338812 , n338811 );
buf ( n338813 , n338234 );
not ( n338814 , n338813 );
or ( n338815 , n338812 , n338814 );
buf ( n338816 , n338209 );
nand ( n18957 , n338815 , n338816 );
buf ( n338818 , n18957 );
buf ( n338819 , n338818 );
buf ( n338820 , n338234 );
not ( n338821 , n338820 );
buf ( n338822 , n18359 );
nand ( n18963 , n338821 , n338822 );
buf ( n338824 , n18963 );
buf ( n18965 , n338824 );
and ( n18966 , n338819 , n18965 );
buf ( n18967 , n18966 );
buf ( n338828 , n338258 );
not ( n18969 , n338828 );
buf ( n18970 , n18969 );
buf ( n338831 , n18970 );
not ( n338832 , n338831 );
buf ( n338833 , n336910 );
not ( n338834 , n338833 );
and ( n338835 , n338832 , n338834 );
buf ( n338836 , n17824 );
buf ( n338837 , n334694 );
and ( n338838 , n338836 , n338837 );
nor ( n338839 , n338835 , n338838 );
buf ( n338840 , n338839 );
buf ( n338841 , n338840 );
not ( n338842 , n338841 );
buf ( n338843 , n338842 );
xor ( n18984 , n18967 , n338843 );
xor ( n338845 , n337639 , n337643 );
xor ( n338846 , n338845 , n337666 );
buf ( n338847 , n338846 );
xnor ( n18988 , n18984 , n338847 );
buf ( n338849 , n18988 );
xnor ( n18990 , n18950 , n338849 );
buf ( n338851 , n18990 );
buf ( n338852 , n338851 );
xor ( n338853 , n338763 , n338852 );
buf ( n338854 , n338853 );
buf ( n338855 , n338854 );
not ( n338856 , n338855 );
and ( n18997 , n338731 , n338856 );
buf ( n338858 , n18869 );
buf ( n338859 , n338854 );
and ( n338860 , n338858 , n338859 );
nor ( n338861 , n18997 , n338860 );
buf ( n338862 , n338861 );
buf ( n338863 , n338862 );
not ( n338864 , n338863 );
and ( n19005 , n338477 , n338864 );
buf ( n338866 , n338475 );
buf ( n338867 , n338862 );
and ( n338868 , n338866 , n338867 );
nor ( n19009 , n19005 , n338868 );
buf ( n19010 , n19009 );
buf ( n338871 , n19010 );
buf ( n338872 , n338717 );
buf ( n338873 , n338723 );
xor ( n338874 , n338872 , n338873 );
buf ( n338875 , n338483 );
xnor ( n338876 , n338874 , n338875 );
buf ( n338877 , n338876 );
buf ( n338878 , n338877 );
not ( n19019 , n338878 );
buf ( n338880 , n19019 );
buf ( n338881 , n591 );
not ( n338882 , n338881 );
buf ( n338883 , n338452 );
not ( n19024 , n338883 );
buf ( n338885 , n19024 );
buf ( n338886 , n338885 );
not ( n19027 , n338886 );
or ( n338888 , n338882 , n19027 );
buf ( n338889 , n590 );
not ( n338890 , n338889 );
buf ( n338891 , n14896 );
not ( n19032 , n338891 );
or ( n338893 , n338890 , n19032 );
buf ( n338894 , n14897 );
buf ( n338895 , n335097 );
nand ( n19036 , n338894 , n338895 );
buf ( n338897 , n19036 );
buf ( n338898 , n338897 );
nand ( n338899 , n338893 , n338898 );
buf ( n338900 , n338899 );
buf ( n338901 , n338900 );
buf ( n338902 , n335181 );
nand ( n338903 , n338901 , n338902 );
buf ( n338904 , n338903 );
buf ( n338905 , n338904 );
nand ( n338906 , n338888 , n338905 );
buf ( n338907 , n338906 );
buf ( n338908 , n15275 );
not ( n338909 , n338908 );
buf ( n338910 , n338711 );
not ( n19051 , n338910 );
or ( n338912 , n338909 , n19051 );
and ( n338913 , n15096 , n334972 );
not ( n19054 , n15096 );
and ( n338915 , n19054 , n588 );
or ( n338916 , n338913 , n338915 );
buf ( n338917 , n338916 );
buf ( n338918 , n335114 );
nand ( n19059 , n338917 , n338918 );
buf ( n338920 , n19059 );
buf ( n338921 , n338920 );
nand ( n19062 , n338912 , n338921 );
buf ( n338923 , n19062 );
buf ( n338924 , n338923 );
not ( n338925 , n338924 );
not ( n338926 , n15115 );
not ( n19067 , n338500 );
or ( n338928 , n338926 , n19067 );
buf ( n338929 , n586 );
not ( n19070 , n338929 );
buf ( n338931 , n18309 );
not ( n338932 , n338931 );
or ( n19073 , n19070 , n338932 );
buf ( n338934 , n337680 );
buf ( n338935 , n334982 );
nand ( n19076 , n338934 , n338935 );
buf ( n19077 , n19076 );
buf ( n338938 , n19077 );
nand ( n19079 , n19073 , n338938 );
buf ( n338940 , n19079 );
nand ( n19081 , n338940 , n15163 );
nand ( n338942 , n338928 , n19081 );
not ( n19083 , n338942 );
not ( n19084 , n19083 );
buf ( n338945 , n338314 );
buf ( n338946 , n334694 );
and ( n19087 , n338945 , n338946 );
buf ( n338948 , n582 );
not ( n338949 , n338948 );
buf ( n338950 , n336354 );
not ( n338951 , n338950 );
or ( n338952 , n338949 , n338951 );
buf ( n338953 , n337626 );
buf ( n338954 , n334702 );
nand ( n338955 , n338953 , n338954 );
buf ( n338956 , n338955 );
buf ( n338957 , n338956 );
nand ( n19098 , n338952 , n338957 );
buf ( n338959 , n19098 );
buf ( n338960 , n338959 );
not ( n19101 , n338960 );
buf ( n338962 , n336910 );
nor ( n19103 , n19101 , n338962 );
buf ( n338964 , n19103 );
buf ( n338965 , n338964 );
nor ( n19106 , n19087 , n338965 );
buf ( n338967 , n19106 );
buf ( n338968 , n338967 );
not ( n338969 , n338968 );
buf ( n338970 , n334868 );
not ( n19111 , n338970 );
buf ( n338972 , n338675 );
not ( n19113 , n338972 );
or ( n338974 , n19111 , n19113 );
buf ( n338975 , n584 );
not ( n19116 , n338975 );
buf ( n338977 , n336319 );
not ( n19118 , n338977 );
or ( n19119 , n19116 , n19118 );
buf ( n338980 , n336983 );
buf ( n338981 , n334879 );
nand ( n338982 , n338980 , n338981 );
buf ( n338983 , n338982 );
buf ( n338984 , n338983 );
nand ( n338985 , n19119 , n338984 );
buf ( n338986 , n338985 );
buf ( n338987 , n338986 );
buf ( n338988 , n334914 );
nand ( n338989 , n338987 , n338988 );
buf ( n338990 , n338989 );
buf ( n338991 , n338990 );
nand ( n19132 , n338974 , n338991 );
buf ( n19133 , n19132 );
buf ( n338994 , n19133 );
not ( n19135 , n338994 );
buf ( n19136 , n19135 );
buf ( n338997 , n19136 );
not ( n338998 , n338997 );
or ( n19139 , n338969 , n338998 );
xor ( n19140 , n338513 , n338538 );
xor ( n19141 , n19140 , n338650 );
buf ( n339002 , n19141 );
buf ( n339003 , n339002 );
nand ( n19144 , n19139 , n339003 );
buf ( n339005 , n19144 );
buf ( n339006 , n338967 );
not ( n339007 , n339006 );
buf ( n339008 , n19133 );
nand ( n339009 , n339007 , n339008 );
buf ( n339010 , n339009 );
nand ( n19151 , n339005 , n339010 );
not ( n19152 , n19151 );
not ( n339013 , n19152 );
or ( n19154 , n19084 , n339013 );
xor ( n339015 , n338654 , n338657 );
xor ( n19156 , n339015 , n338682 );
nand ( n339017 , n19154 , n19156 );
buf ( n339018 , n339017 );
nand ( n339019 , n19151 , n338942 );
buf ( n339020 , n339019 );
nand ( n19161 , n339018 , n339020 );
buf ( n339022 , n19161 );
buf ( n339023 , n339022 );
not ( n19164 , n339023 );
buf ( n339025 , n19164 );
buf ( n339026 , n339025 );
nand ( n339027 , n338925 , n339026 );
buf ( n339028 , n339027 );
not ( n19169 , n339028 );
xor ( n339030 , n338685 , n18832 );
xnor ( n339031 , n339030 , n338510 );
not ( n19172 , n339031 );
or ( n339033 , n19169 , n19172 );
buf ( n339034 , n338923 );
buf ( n339035 , n339022 );
nand ( n19176 , n339034 , n339035 );
buf ( n339037 , n19176 );
nand ( n19178 , n339033 , n339037 );
or ( n19179 , n338907 , n19178 );
and ( n19180 , n338880 , n19179 );
buf ( n339041 , n338907 );
buf ( n339042 , n19178 );
and ( n19183 , n339041 , n339042 );
buf ( n339044 , n19183 );
nor ( n19185 , n19180 , n339044 );
buf ( n339046 , n19185 );
nand ( n339047 , n338871 , n339046 );
buf ( n339048 , n339047 );
buf ( n339049 , n339048 );
buf ( n339050 , n15115 );
not ( n19191 , n339050 );
buf ( n339052 , n338940 );
not ( n339053 , n339052 );
or ( n19194 , n19191 , n339053 );
buf ( n339055 , n586 );
not ( n19196 , n339055 );
buf ( n339057 , n335326 );
not ( n339058 , n339057 );
or ( n19199 , n19196 , n339058 );
buf ( n339060 , n15463 );
buf ( n19201 , n334982 );
nand ( n19202 , n339060 , n19201 );
buf ( n339063 , n19202 );
buf ( n339064 , n339063 );
nand ( n19205 , n19199 , n339064 );
buf ( n339066 , n19205 );
buf ( n339067 , n339066 );
buf ( n339068 , n15163 );
nand ( n19209 , n339067 , n339068 );
buf ( n339070 , n19209 );
buf ( n339071 , n339070 );
nand ( n19212 , n19194 , n339071 );
buf ( n339073 , n19212 );
buf ( n339074 , n339073 );
not ( n19215 , n339074 );
xor ( n339076 , n338627 , n338578 );
buf ( n339077 , n339076 );
not ( n339078 , n339077 );
buf ( n339079 , n334694 );
not ( n19220 , n339079 );
and ( n19221 , n16430 , n334702 );
not ( n339082 , n16430 );
and ( n19223 , n339082 , n582 );
or ( n339084 , n19221 , n19223 );
buf ( n339085 , n339084 );
not ( n339086 , n339085 );
or ( n339087 , n19220 , n339086 );
buf ( n339088 , n582 );
not ( n339089 , n339088 );
buf ( n339090 , n18132 );
not ( n339091 , n339090 );
or ( n19232 , n339089 , n339091 );
buf ( n339093 , n336665 );
buf ( n339094 , n334702 );
nand ( n339095 , n339093 , n339094 );
buf ( n339096 , n339095 );
buf ( n339097 , n339096 );
nand ( n339098 , n19232 , n339097 );
buf ( n339099 , n339098 );
buf ( n339100 , n339099 );
buf ( n339101 , n334727 );
nand ( n339102 , n339100 , n339101 );
buf ( n339103 , n339102 );
buf ( n339104 , n339103 );
nand ( n339105 , n339087 , n339104 );
buf ( n339106 , n339105 );
buf ( n339107 , n339106 );
not ( n339108 , n339107 );
or ( n19249 , n339078 , n339108 );
or ( n339110 , n339076 , n339106 );
and ( n339111 , n339099 , n334694 );
buf ( n19252 , n582 );
not ( n19253 , n19252 );
buf ( n339114 , n337332 );
not ( n19255 , n339114 );
or ( n19256 , n19253 , n19255 );
buf ( n339117 , n337278 );
buf ( n339118 , n334702 );
nand ( n339119 , n339117 , n339118 );
buf ( n339120 , n339119 );
buf ( n339121 , n339120 );
nand ( n339122 , n19256 , n339121 );
buf ( n339123 , n339122 );
and ( n19264 , n339123 , n334727 );
nor ( n339125 , n339111 , n19264 );
not ( n339126 , n339125 );
not ( n19267 , n339126 );
xor ( n339128 , n338595 , n338617 );
not ( n339129 , n339128 );
or ( n19270 , n19267 , n339129 );
buf ( n339131 , n339128 );
not ( n19272 , n339131 );
buf ( n339133 , n19272 );
not ( n339134 , n339133 );
not ( n339135 , n339125 );
or ( n19276 , n339134 , n339135 );
buf ( n339137 , n337364 );
buf ( n339138 , n334643 );
and ( n19279 , n339137 , n339138 );
buf ( n339140 , n19279 );
buf ( n339141 , n339140 );
not ( n339142 , n339141 );
buf ( n339143 , n339142 );
buf ( n339144 , n339143 );
not ( n19285 , n339144 );
buf ( n339146 , n334694 );
not ( n339147 , n339146 );
buf ( n339148 , n582 );
not ( n339149 , n339148 );
buf ( n339150 , n337313 );
not ( n19291 , n339150 );
or ( n339152 , n339149 , n19291 );
buf ( n339153 , n17456 );
buf ( n339154 , n334702 );
nand ( n19295 , n339153 , n339154 );
buf ( n339156 , n19295 );
buf ( n339157 , n339156 );
nand ( n339158 , n339152 , n339157 );
buf ( n339159 , n339158 );
buf ( n339160 , n339159 );
not ( n339161 , n339160 );
or ( n339162 , n339147 , n339161 );
buf ( n339163 , n334702 );
buf ( n339164 , n337364 );
or ( n19305 , n339163 , n339164 );
buf ( n339166 , n582 );
buf ( n339167 , n337361 );
or ( n339168 , n339166 , n339167 );
nand ( n339169 , n19305 , n339168 );
buf ( n339170 , n339169 );
buf ( n339171 , n339170 );
buf ( n339172 , n334727 );
nand ( n339173 , n339171 , n339172 );
buf ( n339174 , n339173 );
buf ( n339175 , n339174 );
nand ( n19316 , n339162 , n339175 );
buf ( n339177 , n19316 );
buf ( n339178 , n339177 );
buf ( n339179 , n583 );
buf ( n339180 , n584 );
or ( n339181 , n339179 , n339180 );
buf ( n339182 , n337364 );
nand ( n339183 , n339181 , n339182 );
buf ( n339184 , n339183 );
buf ( n339185 , n339184 );
buf ( n339186 , n583 );
buf ( n339187 , n584 );
and ( n19328 , n339186 , n339187 );
buf ( n339189 , n334702 );
nor ( n19330 , n19328 , n339189 );
buf ( n339191 , n19330 );
buf ( n339192 , n339191 );
and ( n19333 , n339185 , n339192 );
buf ( n339194 , n19333 );
buf ( n339195 , n339194 );
nand ( n19336 , n339178 , n339195 );
buf ( n339197 , n19336 );
buf ( n339198 , n339197 );
not ( n339199 , n339198 );
or ( n339200 , n19285 , n339199 );
buf ( n339201 , n334694 );
not ( n19342 , n339201 );
buf ( n339203 , n339123 );
not ( n339204 , n339203 );
or ( n339205 , n19342 , n339204 );
buf ( n339206 , n339159 );
buf ( n339207 , n334727 );
nand ( n19348 , n339206 , n339207 );
buf ( n339209 , n19348 );
buf ( n339210 , n339209 );
nand ( n339211 , n339205 , n339210 );
buf ( n339212 , n339211 );
buf ( n339213 , n339212 );
nand ( n19354 , n339200 , n339213 );
buf ( n339215 , n19354 );
not ( n19356 , n339215 );
nand ( n19357 , n19276 , n19356 );
nand ( n19358 , n19270 , n19357 );
nand ( n339219 , n339110 , n19358 );
buf ( n339220 , n339219 );
nand ( n19361 , n19249 , n339220 );
buf ( n339222 , n19361 );
buf ( n339223 , n339222 );
not ( n339224 , n339223 );
xor ( n19365 , n18690 , n338631 );
xor ( n19366 , n19365 , n338645 );
buf ( n339227 , n19366 );
buf ( n339228 , n339227 );
not ( n19369 , n339228 );
buf ( n339230 , n334694 );
not ( n339231 , n339230 );
buf ( n339232 , n338959 );
not ( n339233 , n339232 );
or ( n339234 , n339231 , n339233 );
buf ( n339235 , n339084 );
buf ( n339236 , n334727 );
nand ( n339237 , n339235 , n339236 );
buf ( n339238 , n339237 );
buf ( n339239 , n339238 );
nand ( n339240 , n339234 , n339239 );
buf ( n339241 , n339240 );
buf ( n339242 , n339241 );
not ( n19383 , n339242 );
buf ( n339244 , n19383 );
buf ( n339245 , n339244 );
nand ( n19386 , n19369 , n339245 );
buf ( n339247 , n19386 );
buf ( n339248 , n339247 );
not ( n19389 , n339248 );
or ( n19390 , n339224 , n19389 );
buf ( n339251 , n339241 );
buf ( n339252 , n339227 );
nand ( n19393 , n339251 , n339252 );
buf ( n339254 , n19393 );
buf ( n339255 , n339254 );
nand ( n339256 , n19390 , n339255 );
buf ( n339257 , n339256 );
buf ( n339258 , n339257 );
not ( n19399 , n339258 );
buf ( n339260 , n19399 );
buf ( n339261 , n339260 );
nand ( n19402 , n19215 , n339261 );
buf ( n339263 , n19402 );
xor ( n19404 , n338967 , n339002 );
xor ( n19405 , n19404 , n19136 );
and ( n19406 , n339263 , n19405 );
and ( n19407 , n339073 , n339257 );
nor ( n339268 , n19406 , n19407 );
buf ( n339269 , n339268 );
buf ( n339270 , n588 );
not ( n339271 , n339270 );
buf ( n339272 , n338370 );
not ( n19413 , n339272 );
or ( n339274 , n339271 , n19413 );
buf ( n339275 , n335361 );
buf ( n339276 , n334972 );
nand ( n339277 , n339275 , n339276 );
buf ( n339278 , n339277 );
buf ( n339279 , n339278 );
nand ( n19420 , n339274 , n339279 );
buf ( n339281 , n19420 );
buf ( n339282 , n339281 );
not ( n339283 , n339282 );
buf ( n339284 , n339283 );
buf ( n339285 , n339284 );
not ( n339286 , n339285 );
buf ( n339287 , n335111 );
not ( n339288 , n339287 );
and ( n19429 , n339286 , n339288 );
buf ( n339290 , n338916 );
buf ( n339291 , n15275 );
and ( n19432 , n339290 , n339291 );
nor ( n339293 , n19429 , n19432 );
buf ( n339294 , n339293 );
buf ( n339295 , n339294 );
xor ( n19436 , n339269 , n339295 );
buf ( n339297 , n590 );
buf ( n339298 , n335434 );
and ( n339299 , n339297 , n339298 );
not ( n19440 , n339297 );
buf ( n339301 , n334738 );
and ( n19442 , n19440 , n339301 );
nor ( n339303 , n339299 , n19442 );
buf ( n339304 , n339303 );
not ( n19445 , n339304 );
not ( n339306 , n338457 );
and ( n339307 , n19445 , n339306 );
buf ( n339308 , n590 );
not ( n339309 , n339308 );
buf ( n339310 , n15622 );
not ( n19451 , n339310 );
or ( n339312 , n339309 , n19451 );
buf ( n339313 , n17055 );
buf ( n339314 , n335097 );
nand ( n19455 , n339313 , n339314 );
buf ( n339316 , n19455 );
buf ( n339317 , n339316 );
nand ( n19458 , n339312 , n339317 );
buf ( n339319 , n19458 );
and ( n19460 , n339319 , n591 );
nor ( n339321 , n339307 , n19460 );
buf ( n339322 , n339321 );
and ( n19463 , n19436 , n339322 );
and ( n339324 , n339269 , n339295 );
or ( n339325 , n19463 , n339324 );
buf ( n339326 , n339325 );
buf ( n339327 , n339326 );
buf ( n339328 , n339319 );
not ( n19469 , n339328 );
buf ( n19470 , n19469 );
buf ( n339331 , n19470 );
not ( n19472 , n339331 );
buf ( n339333 , n338457 );
not ( n19474 , n339333 );
and ( n19475 , n19472 , n19474 );
buf ( n339336 , n338900 );
buf ( n339337 , n591 );
and ( n339338 , n339336 , n339337 );
nor ( n19479 , n19475 , n339338 );
buf ( n339340 , n19479 );
buf ( n339341 , n339340 );
xor ( n339342 , n339327 , n339341 );
buf ( n339343 , n339031 );
xor ( n339344 , n338923 , n339025 );
buf ( n339345 , n339344 );
xor ( n339346 , n339343 , n339345 );
buf ( n339347 , n339346 );
buf ( n339348 , n339347 );
xor ( n19489 , n339342 , n339348 );
buf ( n339350 , n19489 );
buf ( n19491 , n339350 );
not ( n339352 , n19083 );
not ( n19493 , n19151 );
or ( n339354 , n339352 , n19493 );
nand ( n339355 , n19152 , n338942 );
nand ( n19496 , n339354 , n339355 );
and ( n339357 , n19496 , n19156 );
not ( n339358 , n19496 );
not ( n19499 , n19156 );
and ( n19500 , n339358 , n19499 );
nor ( n339361 , n339357 , n19500 );
not ( n339362 , n339361 );
xor ( n19503 , n339269 , n339295 );
xor ( n339364 , n19503 , n339322 );
buf ( n339365 , n339364 );
buf ( n339366 , n339365 );
buf ( n339367 , n339366 );
buf ( n339368 , n339367 );
nand ( n19509 , n339362 , n339368 );
buf ( n339370 , n334868 );
not ( n19511 , n339370 );
buf ( n339372 , n338986 );
not ( n19513 , n339372 );
or ( n339374 , n19511 , n19513 );
buf ( n339375 , n584 );
not ( n19516 , n339375 );
buf ( n339377 , n16843 );
not ( n339378 , n339377 );
or ( n19519 , n19516 , n339378 );
buf ( n339380 , n336463 );
buf ( n339381 , n334879 );
nand ( n19522 , n339380 , n339381 );
buf ( n19523 , n19522 );
buf ( n339384 , n19523 );
nand ( n339385 , n19519 , n339384 );
buf ( n339386 , n339385 );
buf ( n339387 , n339386 );
buf ( n339388 , n334914 );
nand ( n339389 , n339387 , n339388 );
buf ( n339390 , n339389 );
buf ( n339391 , n339390 );
nand ( n339392 , n339374 , n339391 );
buf ( n339393 , n339392 );
buf ( n339394 , n339393 );
xor ( n339395 , n339227 , n339244 );
xnor ( n339396 , n339395 , n339222 );
buf ( n339397 , n339396 );
xor ( n339398 , n339394 , n339397 );
buf ( n339399 , n15115 );
not ( n339400 , n339399 );
buf ( n339401 , n339066 );
not ( n339402 , n339401 );
or ( n19543 , n339400 , n339402 );
buf ( n339404 , n586 );
not ( n339405 , n339404 );
buf ( n339406 , n336064 );
not ( n339407 , n339406 );
or ( n19548 , n339405 , n339407 );
buf ( n339409 , n336067 );
buf ( n339410 , n334982 );
nand ( n19551 , n339409 , n339410 );
buf ( n339412 , n19551 );
buf ( n339413 , n339412 );
nand ( n19554 , n19548 , n339413 );
buf ( n19555 , n19554 );
buf ( n19556 , n19555 );
buf ( n19557 , n15163 );
nand ( n19558 , n19556 , n19557 );
buf ( n19559 , n19558 );
buf ( n19560 , n19559 );
nand ( n19561 , n19543 , n19560 );
buf ( n19562 , n19561 );
buf ( n339423 , n19562 );
and ( n339424 , n339398 , n339423 );
and ( n19565 , n339394 , n339397 );
or ( n339426 , n339424 , n19565 );
buf ( n339427 , n339426 );
buf ( n339428 , n339427 );
not ( n339429 , n339428 );
buf ( n339430 , n339429 );
buf ( n339431 , n339430 );
not ( n339432 , n339431 );
and ( n19573 , n588 , n335459 );
not ( n339434 , n588 );
and ( n19575 , n339434 , n335301 );
nor ( n19576 , n19573 , n19575 );
not ( n339437 , n19576 );
not ( n19578 , n339437 );
not ( n339439 , n335111 );
and ( n19580 , n19578 , n339439 );
and ( n19581 , n339281 , n15275 );
nor ( n339442 , n19580 , n19581 );
buf ( n339443 , n339442 );
not ( n19584 , n339443 );
or ( n339445 , n339432 , n19584 );
buf ( n339446 , n339260 );
buf ( n339447 , n339073 );
xor ( n339448 , n339446 , n339447 );
buf ( n339449 , n19405 );
xnor ( n339450 , n339448 , n339449 );
buf ( n339451 , n339450 );
buf ( n339452 , n339451 );
nand ( n339453 , n339445 , n339452 );
buf ( n339454 , n339453 );
buf ( n339455 , n339454 );
buf ( n339456 , n339442 );
not ( n19597 , n339456 );
buf ( n339458 , n339427 );
nand ( n19599 , n19597 , n339458 );
buf ( n339460 , n19599 );
buf ( n339461 , n339460 );
nand ( n339462 , n339455 , n339461 );
buf ( n339463 , n339462 );
buf ( n339464 , n339463 );
and ( n19605 , n19509 , n339464 );
not ( n19606 , n339361 );
nor ( n339467 , n339368 , n19606 );
nor ( n19608 , n19605 , n339467 );
buf ( n339469 , n19608 );
nand ( n19610 , n19491 , n339469 );
buf ( n339471 , n19610 );
not ( n339472 , n339471 );
buf ( n339473 , n15275 );
not ( n19614 , n339473 );
and ( n339475 , n588 , n335310 );
not ( n339476 , n588 );
and ( n19617 , n339476 , n337680 );
or ( n339478 , n339475 , n19617 );
buf ( n339479 , n339478 );
not ( n339480 , n339479 );
or ( n19621 , n19614 , n339480 );
and ( n339482 , n588 , n335326 );
not ( n339483 , n588 );
and ( n19624 , n339483 , n15463 );
or ( n339485 , n339482 , n19624 );
buf ( n339486 , n339485 );
buf ( n339487 , n335114 );
nand ( n339488 , n339486 , n339487 );
buf ( n339489 , n339488 );
buf ( n339490 , n339489 );
nand ( n339491 , n19621 , n339490 );
buf ( n339492 , n339491 );
buf ( n339493 , n339492 );
not ( n339494 , n339493 );
xor ( n19635 , n339128 , n339215 );
xnor ( n339496 , n19635 , n339125 );
not ( n339497 , n339496 );
not ( n339498 , n334914 );
buf ( n339499 , n584 );
not ( n339500 , n339499 );
buf ( n339501 , n336296 );
not ( n339502 , n339501 );
or ( n19643 , n339500 , n339502 );
buf ( n339504 , n334879 );
buf ( n339505 , n16430 );
nand ( n19646 , n339504 , n339505 );
buf ( n339507 , n19646 );
buf ( n339508 , n339507 );
nand ( n339509 , n19643 , n339508 );
buf ( n339510 , n339509 );
not ( n339511 , n339510 );
or ( n339512 , n339498 , n339511 );
and ( n19653 , n17762 , n334879 );
not ( n19654 , n17762 );
and ( n339515 , n19654 , n584 );
or ( n339516 , n19653 , n339515 );
nand ( n19657 , n339516 , n334867 );
nand ( n339518 , n339512 , n19657 );
not ( n339519 , n339518 );
buf ( n339520 , n586 );
not ( n339521 , n339520 );
buf ( n339522 , n16411 );
not ( n339523 , n339522 );
or ( n19664 , n339521 , n339523 );
buf ( n339525 , n336275 );
buf ( n339526 , n334982 );
nand ( n19667 , n339525 , n339526 );
buf ( n19668 , n19667 );
buf ( n339529 , n19668 );
nand ( n19670 , n19664 , n339529 );
buf ( n339531 , n19670 );
nand ( n19672 , n339531 , n15163 );
not ( n339533 , n586 );
not ( n19674 , n336319 );
or ( n19675 , n339533 , n19674 );
buf ( n339536 , n16456 );
buf ( n339537 , n334982 );
nand ( n339538 , n339536 , n339537 );
buf ( n339539 , n339538 );
nand ( n19680 , n19675 , n339539 );
nand ( n339541 , n19680 , n15115 );
nand ( n339542 , n339519 , n19672 , n339541 );
nand ( n19683 , n339497 , n339542 );
buf ( n339544 , n19683 );
not ( n339545 , n15163 );
not ( n19686 , n339531 );
or ( n339547 , n339545 , n19686 );
nand ( n339548 , n339547 , n339541 );
buf ( n339549 , n339548 );
buf ( n339550 , n339518 );
nand ( n339551 , n339549 , n339550 );
buf ( n339552 , n339551 );
buf ( n339553 , n339552 );
and ( n339554 , n339544 , n339553 );
buf ( n339555 , n339554 );
buf ( n339556 , n339555 );
buf ( n19697 , n339556 );
buf ( n339558 , n19697 );
buf ( n339559 , n339558 );
nand ( n339560 , n339494 , n339559 );
buf ( n339561 , n339560 );
buf ( n339562 , n339561 );
not ( n339563 , n339106 );
not ( n19704 , n339076 );
and ( n19705 , n339563 , n19704 );
and ( n339566 , n339106 , n339076 );
nor ( n19707 , n19705 , n339566 );
xnor ( n339568 , n19358 , n19707 );
buf ( n339569 , n334868 );
not ( n19710 , n339569 );
buf ( n339571 , n339386 );
not ( n339572 , n339571 );
or ( n19713 , n19710 , n339572 );
buf ( n339574 , n339516 );
buf ( n339575 , n334914 );
nand ( n19716 , n339574 , n339575 );
buf ( n19717 , n19716 );
buf ( n339578 , n19717 );
nand ( n339579 , n19713 , n339578 );
buf ( n339580 , n339579 );
not ( n339581 , n339580 );
and ( n339582 , n339568 , n339581 );
not ( n19723 , n339568 );
and ( n339584 , n19723 , n339580 );
nor ( n339585 , n339582 , n339584 );
buf ( n339586 , n19555 );
buf ( n339587 , n15115 );
and ( n19728 , n339586 , n339587 );
and ( n339589 , n19680 , n15163 );
buf ( n339590 , n339589 );
nor ( n19731 , n19728 , n339590 );
buf ( n339592 , n19731 );
and ( n19733 , n339585 , n339592 );
not ( n339594 , n339585 );
buf ( n339595 , n339592 );
not ( n19736 , n339595 );
buf ( n339597 , n19736 );
and ( n19738 , n339594 , n339597 );
or ( n339599 , n19733 , n19738 );
buf ( n339600 , n339599 );
and ( n19741 , n339562 , n339600 );
buf ( n339602 , n339492 );
not ( n19743 , n339602 );
buf ( n339604 , n339558 );
nor ( n339605 , n19743 , n339604 );
buf ( n339606 , n339605 );
buf ( n339607 , n339606 );
nor ( n19748 , n19741 , n339607 );
buf ( n339609 , n19748 );
buf ( n339610 , n591 );
not ( n19751 , n339610 );
buf ( n339612 , n590 );
buf ( n339613 , n15096 );
and ( n339614 , n339612 , n339613 );
not ( n19755 , n339612 );
buf ( n339616 , n15095 );
and ( n19757 , n19755 , n339616 );
nor ( n339618 , n339614 , n19757 );
buf ( n339619 , n339618 );
buf ( n339620 , n339619 );
not ( n19761 , n339620 );
or ( n19762 , n19751 , n19761 );
buf ( n339623 , n590 );
not ( n19764 , n339623 );
buf ( n339625 , n338370 );
not ( n339626 , n339625 );
or ( n339627 , n19764 , n339626 );
buf ( n339628 , n335361 );
buf ( n339629 , n335097 );
nand ( n339630 , n339628 , n339629 );
buf ( n339631 , n339630 );
buf ( n339632 , n339631 );
nand ( n339633 , n339627 , n339632 );
buf ( n339634 , n339633 );
buf ( n339635 , n339634 );
buf ( n339636 , n335181 );
nand ( n339637 , n339635 , n339636 );
buf ( n339638 , n339637 );
buf ( n339639 , n339638 );
nand ( n19780 , n19762 , n339639 );
buf ( n339641 , n19780 );
xnor ( n19782 , n339609 , n339641 );
buf ( n339643 , n19782 );
buf ( n339644 , n339581 );
not ( n339645 , n339644 );
buf ( n339646 , n339592 );
not ( n19787 , n339646 );
or ( n339648 , n339645 , n19787 );
not ( n339649 , n339568 );
buf ( n339650 , n339649 );
nand ( n339651 , n339648 , n339650 );
buf ( n339652 , n339651 );
buf ( n339653 , n339652 );
buf ( n339654 , n339597 );
buf ( n339655 , n339580 );
nand ( n19796 , n339654 , n339655 );
buf ( n339657 , n19796 );
buf ( n339658 , n339657 );
and ( n339659 , n339653 , n339658 );
buf ( n339660 , n339659 );
buf ( n339661 , n339660 );
not ( n19802 , n15275 );
not ( n19803 , n19576 );
or ( n339664 , n19802 , n19803 );
buf ( n339665 , n339478 );
buf ( n339666 , n335114 );
nand ( n19807 , n339665 , n339666 );
buf ( n339668 , n19807 );
nand ( n339669 , n339664 , n339668 );
buf ( n339670 , n339669 );
xor ( n19811 , n339661 , n339670 );
xor ( n19812 , n339394 , n339397 );
xor ( n19813 , n19812 , n339423 );
buf ( n339674 , n19813 );
buf ( n339675 , n339674 );
xnor ( n19816 , n19811 , n339675 );
buf ( n339677 , n19816 );
buf ( n339678 , n339677 );
not ( n19819 , n339678 );
buf ( n19820 , n19819 );
buf ( n339681 , n19820 );
and ( n19822 , n339643 , n339681 );
not ( n19823 , n339643 );
buf ( n339684 , n339677 );
and ( n19825 , n19823 , n339684 );
nor ( n339686 , n19822 , n19825 );
buf ( n339687 , n339686 );
buf ( n339688 , n339687 );
buf ( n339689 , n591 );
not ( n339690 , n339689 );
buf ( n339691 , n339634 );
not ( n19832 , n339691 );
or ( n339693 , n339690 , n19832 );
buf ( n339694 , n335181 );
buf ( n339695 , n335097 );
buf ( n339696 , n335301 );
and ( n19837 , n339695 , n339696 );
not ( n19838 , n339695 );
buf ( n339699 , n335459 );
and ( n339700 , n19838 , n339699 );
nor ( n339701 , n19837 , n339700 );
buf ( n339702 , n339701 );
buf ( n339703 , n339702 );
nand ( n339704 , n339694 , n339703 );
buf ( n339705 , n339704 );
buf ( n339706 , n339705 );
nand ( n339707 , n339693 , n339706 );
buf ( n339708 , n339707 );
buf ( n339709 , n339708 );
not ( n339710 , n339709 );
buf ( n339711 , n339710 );
not ( n19852 , n339711 );
buf ( n339713 , n339140 );
buf ( n339714 , n339197 );
xor ( n339715 , n339713 , n339714 );
buf ( n339716 , n339212 );
xnor ( n339717 , n339715 , n339716 );
buf ( n339718 , n339717 );
buf ( n339719 , n339718 );
buf ( n339720 , n334868 );
not ( n19861 , n339720 );
buf ( n339722 , n339510 );
not ( n19863 , n339722 );
or ( n339724 , n19861 , n19863 );
buf ( n339725 , n584 );
not ( n19866 , n339725 );
buf ( n339727 , n18132 );
not ( n339728 , n339727 );
or ( n19869 , n19866 , n339728 );
buf ( n339730 , n337990 );
buf ( n339731 , n334879 );
nand ( n19872 , n339730 , n339731 );
buf ( n19873 , n19872 );
buf ( n339734 , n19873 );
nand ( n339735 , n19869 , n339734 );
buf ( n339736 , n339735 );
buf ( n339737 , n339736 );
buf ( n339738 , n334914 );
nand ( n19879 , n339737 , n339738 );
buf ( n19880 , n19879 );
buf ( n339741 , n19880 );
nand ( n19882 , n339724 , n339741 );
buf ( n339743 , n19882 );
buf ( n339744 , n339743 );
xor ( n19885 , n339719 , n339744 );
xor ( n19886 , n339194 , n339177 );
buf ( n339747 , n19886 );
not ( n19888 , n339747 );
buf ( n339749 , n334868 );
not ( n19890 , n339749 );
buf ( n339751 , n339736 );
not ( n339752 , n339751 );
or ( n339753 , n19890 , n339752 );
buf ( n339754 , n584 );
not ( n339755 , n339754 );
buf ( n339756 , n337332 );
not ( n19897 , n339756 );
or ( n339758 , n339755 , n19897 );
buf ( n339759 , n337278 );
buf ( n339760 , n334879 );
nand ( n19901 , n339759 , n339760 );
buf ( n339762 , n19901 );
buf ( n339763 , n339762 );
nand ( n339764 , n339758 , n339763 );
buf ( n339765 , n339764 );
buf ( n339766 , n339765 );
buf ( n339767 , n334914 );
nand ( n339768 , n339766 , n339767 );
buf ( n339769 , n339768 );
buf ( n339770 , n339769 );
nand ( n19911 , n339753 , n339770 );
buf ( n339772 , n19911 );
buf ( n339773 , n339772 );
not ( n19914 , n339773 );
or ( n339775 , n19888 , n19914 );
buf ( n339776 , n19886 );
not ( n339777 , n339776 );
buf ( n339778 , n339777 );
buf ( n339779 , n339778 );
not ( n19920 , n339779 );
buf ( n339781 , n339736 );
buf ( n339782 , n334868 );
and ( n19923 , n339781 , n339782 );
buf ( n19924 , n339769 );
not ( n339785 , n19924 );
buf ( n339786 , n339785 );
buf ( n339787 , n339786 );
nor ( n339788 , n19923 , n339787 );
buf ( n339789 , n339788 );
buf ( n339790 , n339789 );
not ( n339791 , n339790 );
or ( n19932 , n19920 , n339791 );
buf ( n339793 , n337364 );
buf ( n339794 , n334694 );
and ( n339795 , n339793 , n339794 );
buf ( n339796 , n339795 );
buf ( n19937 , n339796 );
not ( n19938 , n19937 );
and ( n339799 , n339765 , n334868 );
and ( n19940 , n334002 , n334879 );
not ( n19941 , n334002 );
and ( n339802 , n19941 , n584 );
or ( n19943 , n19940 , n339802 );
and ( n339804 , n19943 , n334914 );
nor ( n19945 , n339799 , n339804 );
buf ( n339806 , n19945 );
not ( n339807 , n339806 );
buf ( n339808 , n339807 );
buf ( n339809 , n339808 );
not ( n339810 , n339809 );
or ( n339811 , n19938 , n339810 );
buf ( n339812 , n339796 );
not ( n339813 , n339812 );
buf ( n339814 , n339813 );
buf ( n339815 , n339814 );
not ( n339816 , n339815 );
buf ( n339817 , n19945 );
not ( n339818 , n339817 );
or ( n19959 , n339816 , n339818 );
buf ( n339820 , n19943 );
buf ( n339821 , n334868 );
and ( n19962 , n339820 , n339821 );
buf ( n339823 , n334914 );
not ( n339824 , n339823 );
buf ( n339825 , n337361 );
buf ( n339826 , n584 );
and ( n339827 , n339825 , n339826 );
buf ( n339828 , n337364 );
buf ( n339829 , n334879 );
and ( n339830 , n339828 , n339829 );
nor ( n19971 , n339827 , n339830 );
buf ( n19972 , n19971 );
buf ( n339833 , n19972 );
nor ( n19974 , n339824 , n339833 );
buf ( n19975 , n19974 );
buf ( n339836 , n19975 );
nor ( n339837 , n19962 , n339836 );
buf ( n339838 , n339837 );
buf ( n339839 , n339838 );
buf ( n339840 , n585 );
buf ( n339841 , n586 );
or ( n19982 , n339840 , n339841 );
buf ( n339843 , n337364 );
nand ( n19984 , n19982 , n339843 );
buf ( n339845 , n19984 );
buf ( n339846 , n339845 );
buf ( n339847 , n585 );
buf ( n339848 , n586 );
and ( n19989 , n339847 , n339848 );
buf ( n339850 , n334879 );
nor ( n339851 , n19989 , n339850 );
buf ( n339852 , n339851 );
buf ( n339853 , n339852 );
nand ( n339854 , n339846 , n339853 );
buf ( n339855 , n339854 );
buf ( n339856 , n339855 );
nor ( n339857 , n339839 , n339856 );
buf ( n339858 , n339857 );
buf ( n339859 , n339858 );
nand ( n20000 , n19959 , n339859 );
buf ( n20001 , n20000 );
buf ( n20002 , n20001 );
nand ( n20003 , n339811 , n20002 );
buf ( n20004 , n20003 );
buf ( n339865 , n20004 );
nand ( n20006 , n19932 , n339865 );
buf ( n339867 , n20006 );
buf ( n339868 , n339867 );
nand ( n339869 , n339775 , n339868 );
buf ( n339870 , n339869 );
buf ( n339871 , n339870 );
and ( n339872 , n19885 , n339871 );
and ( n20013 , n339719 , n339744 );
or ( n339874 , n339872 , n20013 );
buf ( n339875 , n339874 );
buf ( n339876 , n339875 );
buf ( n339877 , n339518 );
not ( n339878 , n339877 );
buf ( n339879 , n339496 );
not ( n339880 , n339879 );
and ( n339881 , n339878 , n339880 );
buf ( n339882 , n339518 );
buf ( n339883 , n339496 );
and ( n339884 , n339882 , n339883 );
nor ( n339885 , n339881 , n339884 );
buf ( n339886 , n339885 );
xnor ( n339887 , n339548 , n339886 );
buf ( n339888 , n339887 );
xor ( n20029 , n339876 , n339888 );
buf ( n339890 , n15275 );
not ( n339891 , n339890 );
buf ( n339892 , n339485 );
not ( n20033 , n339892 );
or ( n20034 , n339891 , n20033 );
buf ( n339895 , n335114 );
buf ( n339896 , n588 );
not ( n20037 , n339896 );
buf ( n339898 , n336064 );
not ( n339899 , n339898 );
or ( n339900 , n20037 , n339899 );
buf ( n339901 , n336067 );
buf ( n339902 , n334972 );
nand ( n20043 , n339901 , n339902 );
buf ( n339904 , n20043 );
buf ( n339905 , n339904 );
nand ( n20046 , n339900 , n339905 );
buf ( n339907 , n20046 );
buf ( n339908 , n339907 );
nand ( n20049 , n339895 , n339908 );
buf ( n339910 , n20049 );
buf ( n339911 , n339910 );
nand ( n20052 , n20034 , n339911 );
buf ( n20053 , n20052 );
buf ( n339914 , n20053 );
and ( n20055 , n20029 , n339914 );
and ( n339916 , n339876 , n339888 );
or ( n20057 , n20055 , n339916 );
buf ( n339918 , n20057 );
buf ( n339919 , n339918 );
not ( n20060 , n339919 );
buf ( n339921 , n20060 );
not ( n20062 , n339921 );
and ( n339923 , n19852 , n20062 );
buf ( n20064 , n339711 );
buf ( n339925 , n339921 );
nand ( n20066 , n20064 , n339925 );
buf ( n339927 , n20066 );
buf ( n339928 , n339555 );
buf ( n339929 , n339492 );
xor ( n339930 , n339928 , n339929 );
buf ( n339931 , n339599 );
xnor ( n339932 , n339930 , n339931 );
buf ( n339933 , n339932 );
buf ( n339934 , n339933 );
buf ( n339935 , n339934 );
buf ( n339936 , n339935 );
and ( n20077 , n339927 , n339936 );
nor ( n339938 , n339923 , n20077 );
buf ( n339939 , n339938 );
nand ( n20080 , n339688 , n339939 );
buf ( n20081 , n20080 );
buf ( n339942 , n20081 );
not ( n339943 , n339942 );
buf ( n339944 , n591 );
not ( n339945 , n339944 );
buf ( n339946 , n590 );
buf ( n339947 , n337680 );
and ( n339948 , n339946 , n339947 );
not ( n339949 , n339946 );
buf ( n339950 , n18309 );
and ( n20091 , n339949 , n339950 );
nor ( n20092 , n339948 , n20091 );
buf ( n339953 , n20092 );
buf ( n339954 , n339953 );
not ( n20095 , n339954 );
or ( n20096 , n339945 , n20095 );
and ( n20097 , n590 , n335326 );
not ( n339958 , n590 );
and ( n339959 , n339958 , n15463 );
or ( n20100 , n20097 , n339959 );
buf ( n339961 , n20100 );
buf ( n339962 , n335181 );
nand ( n339963 , n339961 , n339962 );
buf ( n339964 , n339963 );
buf ( n339965 , n339964 );
nand ( n20106 , n20096 , n339965 );
buf ( n339967 , n20106 );
buf ( n339968 , n339967 );
buf ( n339969 , n339968 );
buf ( n339970 , n339969 );
not ( n20111 , n339970 );
and ( n20112 , n336259 , n334982 );
not ( n339973 , n336259 );
and ( n339974 , n339973 , n586 );
or ( n20115 , n20112 , n339974 );
and ( n20116 , n20115 , n15115 );
buf ( n339977 , n586 );
not ( n339978 , n339977 );
buf ( n339979 , n16430 );
not ( n20120 , n339979 );
buf ( n339981 , n20120 );
buf ( n339982 , n339981 );
not ( n339983 , n339982 );
or ( n20124 , n339978 , n339983 );
buf ( n339985 , n334982 );
buf ( n339986 , n16430 );
nand ( n339987 , n339985 , n339986 );
buf ( n339988 , n339987 );
buf ( n339989 , n339988 );
nand ( n20130 , n20124 , n339989 );
buf ( n339991 , n20130 );
and ( n339992 , n339991 , n15164 );
nor ( n339993 , n20116 , n339992 );
not ( n20134 , n339993 );
not ( n20135 , n20134 );
buf ( n339996 , n336275 );
not ( n20137 , n339996 );
buf ( n339998 , n334972 );
not ( n20139 , n339998 );
and ( n340000 , n20137 , n20139 );
buf ( n340001 , n336463 );
buf ( n340002 , n334972 );
and ( n340003 , n340001 , n340002 );
nor ( n340004 , n340000 , n340003 );
buf ( n340005 , n340004 );
not ( n340006 , n340005 );
not ( n340007 , n335111 );
and ( n20148 , n340006 , n340007 );
buf ( n340009 , n588 );
not ( n340010 , n340009 );
buf ( n340011 , n14546 );
not ( n20152 , n340011 );
or ( n340013 , n340010 , n20152 );
buf ( n340014 , n16456 );
buf ( n340015 , n334972 );
nand ( n340016 , n340014 , n340015 );
buf ( n340017 , n340016 );
buf ( n340018 , n340017 );
nand ( n20159 , n340013 , n340018 );
buf ( n20160 , n20159 );
and ( n340021 , n20160 , n15275 );
nor ( n20162 , n20148 , n340021 );
not ( n340023 , n20162 );
not ( n20164 , n340023 );
or ( n20165 , n20135 , n20164 );
not ( n20166 , n339993 );
not ( n20167 , n20162 );
or ( n340028 , n20166 , n20167 );
xor ( n20169 , n19886 , n20004 );
and ( n20170 , n20169 , n339772 );
not ( n340031 , n20169 );
and ( n340032 , n340031 , n339789 );
nor ( n20173 , n20170 , n340032 );
nand ( n340034 , n340028 , n20173 );
nand ( n340035 , n20165 , n340034 );
not ( n20176 , n340035 );
or ( n340037 , n20111 , n20176 );
buf ( n20178 , n339970 );
buf ( n340039 , n340035 );
nor ( n20180 , n20178 , n340039 );
buf ( n340041 , n20180 );
buf ( n340042 , n15115 );
not ( n20183 , n340042 );
buf ( n340044 , n339531 );
not ( n20185 , n340044 );
or ( n340046 , n20183 , n20185 );
buf ( n340047 , n20115 );
buf ( n340048 , n15163 );
nand ( n20189 , n340047 , n340048 );
buf ( n340050 , n20189 );
buf ( n340051 , n340050 );
nand ( n20192 , n340046 , n340051 );
buf ( n340053 , n20192 );
buf ( n340054 , n340053 );
xor ( n20195 , n339719 , n339744 );
xor ( n340056 , n20195 , n339871 );
buf ( n340057 , n340056 );
buf ( n340058 , n340057 );
xor ( n340059 , n340054 , n340058 );
buf ( n340060 , n15275 );
not ( n340061 , n340060 );
buf ( n340062 , n339907 );
not ( n340063 , n340062 );
or ( n20204 , n340061 , n340063 );
buf ( n340065 , n335114 );
buf ( n340066 , n20160 );
nand ( n20207 , n340065 , n340066 );
buf ( n340068 , n20207 );
buf ( n340069 , n340068 );
nand ( n20210 , n20204 , n340069 );
buf ( n340071 , n20210 );
buf ( n340072 , n340071 );
xor ( n20213 , n340059 , n340072 );
buf ( n340074 , n20213 );
buf ( n340075 , n340074 );
not ( n20216 , n340075 );
buf ( n20217 , n20216 );
or ( n340078 , n340041 , n20217 );
nand ( n340079 , n340037 , n340078 );
buf ( n340080 , n340079 );
not ( n340081 , n340080 );
xor ( n340082 , n340054 , n340058 );
and ( n20223 , n340082 , n340072 );
and ( n340084 , n340054 , n340058 );
or ( n340085 , n20223 , n340084 );
buf ( n340086 , n340085 );
buf ( n340087 , n340086 );
buf ( n340088 , n591 );
not ( n340089 , n340088 );
buf ( n340090 , n339702 );
not ( n20231 , n340090 );
or ( n340092 , n340089 , n20231 );
buf ( n340093 , n339953 );
buf ( n340094 , n335181 );
nand ( n20235 , n340093 , n340094 );
buf ( n340096 , n20235 );
buf ( n340097 , n340096 );
nand ( n340098 , n340092 , n340097 );
buf ( n340099 , n340098 );
buf ( n340100 , n340099 );
xor ( n340101 , n340087 , n340100 );
buf ( n340102 , n340101 );
buf ( n340103 , n340102 );
xor ( n340104 , n339876 , n339888 );
xor ( n340105 , n340104 , n339914 );
buf ( n340106 , n340105 );
buf ( n340107 , n340106 );
xnor ( n340108 , n340103 , n340107 );
buf ( n340109 , n340108 );
buf ( n340110 , n340109 );
nand ( n340111 , n340081 , n340110 );
buf ( n340112 , n340111 );
not ( n20253 , n340112 );
buf ( n340114 , n340035 );
buf ( n340115 , n339967 );
xor ( n20256 , n340114 , n340115 );
buf ( n340117 , n340074 );
xnor ( n20258 , n20256 , n340117 );
buf ( n340119 , n20258 );
buf ( n340120 , n340119 );
buf ( n340121 , n591 );
not ( n340122 , n340121 );
buf ( n340123 , n20100 );
not ( n20264 , n340123 );
or ( n340125 , n340122 , n20264 );
buf ( n340126 , n590 );
buf ( n340127 , n16201 );
and ( n20268 , n340126 , n340127 );
not ( n340129 , n340126 );
buf ( n340130 , n336064 );
and ( n20271 , n340129 , n340130 );
nor ( n340132 , n20268 , n20271 );
buf ( n340133 , n340132 );
buf ( n340134 , n340133 );
buf ( n340135 , n335181 );
nand ( n20276 , n340134 , n340135 );
buf ( n340137 , n20276 );
buf ( n340138 , n340137 );
nand ( n20279 , n340125 , n340138 );
buf ( n20280 , n20279 );
buf ( n340141 , n20280 );
not ( n20282 , n340141 );
buf ( n20283 , n20282 );
not ( n340144 , n20283 );
buf ( n340145 , n339796 );
buf ( n340146 , n339858 );
xor ( n340147 , n340145 , n340146 );
buf ( n340148 , n339808 );
xor ( n20289 , n340147 , n340148 );
buf ( n20290 , n20289 );
buf ( n340151 , n20290 );
buf ( n340152 , n15115 );
not ( n340153 , n340152 );
buf ( n340154 , n339991 );
not ( n340155 , n340154 );
or ( n20296 , n340153 , n340155 );
buf ( n340157 , n586 );
not ( n340158 , n340157 );
buf ( n340159 , n336662 );
not ( n340160 , n340159 );
or ( n20301 , n340158 , n340160 );
buf ( n340162 , n337990 );
buf ( n340163 , n334982 );
nand ( n340164 , n340162 , n340163 );
buf ( n340165 , n340164 );
buf ( n340166 , n340165 );
nand ( n340167 , n20301 , n340166 );
buf ( n340168 , n340167 );
buf ( n340169 , n340168 );
buf ( n340170 , n15162 );
nand ( n340171 , n340169 , n340170 );
buf ( n340172 , n340171 );
buf ( n340173 , n340172 );
nand ( n340174 , n20296 , n340173 );
buf ( n340175 , n340174 );
buf ( n340176 , n340175 );
xor ( n340177 , n340151 , n340176 );
buf ( n340178 , n339838 );
buf ( n340179 , n339855 );
xor ( n20320 , n340178 , n340179 );
buf ( n340181 , n20320 );
buf ( n340182 , n340181 );
buf ( n340183 , n337364 );
buf ( n340184 , n334868 );
and ( n20325 , n340183 , n340184 );
buf ( n340186 , n20325 );
buf ( n340187 , n340186 );
not ( n20328 , n340187 );
buf ( n340189 , n20328 );
buf ( n340190 , n340189 );
not ( n340191 , n340190 );
and ( n340192 , n337278 , n334982 );
not ( n20333 , n337278 );
and ( n20334 , n20333 , n586 );
or ( n20335 , n340192 , n20334 );
and ( n340196 , n20335 , n15115 );
buf ( n340197 , n586 );
not ( n20338 , n340197 );
buf ( n340199 , n337313 );
not ( n20340 , n340199 );
or ( n340201 , n20338 , n20340 );
buf ( n340202 , n334002 );
buf ( n340203 , n334982 );
nand ( n20344 , n340202 , n340203 );
buf ( n340205 , n20344 );
buf ( n340206 , n340205 );
nand ( n340207 , n340201 , n340206 );
buf ( n340208 , n340207 );
and ( n20349 , n340208 , n15162 );
nor ( n20350 , n340196 , n20349 );
buf ( n340211 , n20350 );
not ( n340212 , n340211 );
or ( n20353 , n340191 , n340212 );
buf ( n340214 , n15115 );
not ( n20355 , n340214 );
buf ( n340216 , n340208 );
not ( n340217 , n340216 );
or ( n20358 , n20355 , n340217 );
buf ( n340219 , n334982 );
buf ( n340220 , n337364 );
or ( n340221 , n340219 , n340220 );
buf ( n340222 , n586 );
buf ( n340223 , n337361 );
or ( n20364 , n340222 , n340223 );
nand ( n20365 , n340221 , n20364 );
buf ( n340226 , n20365 );
buf ( n340227 , n340226 );
buf ( n340228 , n15162 );
nand ( n340229 , n340227 , n340228 );
buf ( n340230 , n340229 );
buf ( n340231 , n340230 );
nand ( n20372 , n20358 , n340231 );
buf ( n340233 , n20372 );
buf ( n340234 , n340233 );
buf ( n340235 , n587 );
buf ( n340236 , n588 );
or ( n20377 , n340235 , n340236 );
buf ( n340238 , n337364 );
nand ( n340239 , n20377 , n340238 );
buf ( n340240 , n340239 );
buf ( n340241 , n340240 );
buf ( n340242 , n587 );
buf ( n340243 , n588 );
and ( n340244 , n340242 , n340243 );
buf ( n340245 , n334982 );
nor ( n340246 , n340244 , n340245 );
buf ( n340247 , n340246 );
buf ( n340248 , n340247 );
and ( n20389 , n340241 , n340248 );
buf ( n340250 , n20389 );
buf ( n340251 , n340250 );
nand ( n20392 , n340234 , n340251 );
buf ( n340253 , n20392 );
buf ( n20394 , n340253 );
not ( n340255 , n20394 );
buf ( n340256 , n340255 );
buf ( n340257 , n340256 );
nand ( n340258 , n20353 , n340257 );
buf ( n340259 , n340258 );
buf ( n340260 , n340259 );
buf ( n340261 , n20350 );
not ( n20402 , n340261 );
buf ( n340263 , n20402 );
buf ( n340264 , n340263 );
buf ( n340265 , n340186 );
nand ( n340266 , n340264 , n340265 );
buf ( n340267 , n340266 );
buf ( n340268 , n340267 );
nand ( n340269 , n340260 , n340268 );
buf ( n340270 , n340269 );
buf ( n340271 , n340270 );
xor ( n20412 , n340182 , n340271 );
buf ( n340273 , n15115 );
not ( n340274 , n340273 );
buf ( n340275 , n340168 );
not ( n340276 , n340275 );
or ( n340277 , n340274 , n340276 );
buf ( n340278 , n20335 );
buf ( n340279 , n15162 );
nand ( n340280 , n340278 , n340279 );
buf ( n340281 , n340280 );
buf ( n340282 , n340281 );
nand ( n20423 , n340277 , n340282 );
buf ( n340284 , n20423 );
buf ( n340285 , n340284 );
and ( n20426 , n20412 , n340285 );
and ( n340287 , n340182 , n340271 );
or ( n20428 , n20426 , n340287 );
buf ( n340289 , n20428 );
buf ( n340290 , n340289 );
and ( n20431 , n340177 , n340290 );
and ( n20432 , n340151 , n340176 );
or ( n340293 , n20431 , n20432 );
buf ( n340294 , n340293 );
buf ( n340295 , n340294 );
not ( n340296 , n340295 );
buf ( n340297 , n340296 );
not ( n20438 , n340297 );
and ( n340299 , n340144 , n20438 );
buf ( n20440 , n20283 );
buf ( n20441 , n340297 );
nand ( n20442 , n20440 , n20441 );
buf ( n20443 , n20442 );
buf ( n340304 , n20162 );
buf ( n340305 , n339993 );
buf ( n340306 , n20173 );
not ( n340307 , n340306 );
buf ( n340308 , n340307 );
buf ( n340309 , n340308 );
and ( n340310 , n340305 , n340309 );
not ( n20451 , n340305 );
buf ( n340312 , n20173 );
and ( n340313 , n20451 , n340312 );
nor ( n20454 , n340310 , n340313 );
buf ( n20455 , n20454 );
buf ( n340316 , n20455 );
not ( n20457 , n340316 );
buf ( n340318 , n20457 );
buf ( n340319 , n340318 );
and ( n340320 , n340304 , n340319 );
not ( n20461 , n340304 );
buf ( n340322 , n20455 );
and ( n20463 , n20461 , n340322 );
nor ( n20464 , n340320 , n20463 );
buf ( n340325 , n20464 );
and ( n340326 , n20443 , n340325 );
nor ( n340327 , n340299 , n340326 );
buf ( n20468 , n340327 );
nand ( n20469 , n340120 , n20468 );
buf ( n20470 , n20469 );
not ( n340331 , n20470 );
not ( n20472 , n15275 );
buf ( n340333 , n340005 );
not ( n340334 , n340333 );
buf ( n340335 , n340334 );
not ( n340336 , n340335 );
or ( n20477 , n20472 , n340336 );
buf ( n340338 , n588 );
not ( n20479 , n340338 );
buf ( n340340 , n17763 );
not ( n340341 , n340340 );
or ( n20482 , n20479 , n340341 );
buf ( n340343 , n336259 );
buf ( n340344 , n334972 );
nand ( n20485 , n340343 , n340344 );
buf ( n340346 , n20485 );
buf ( n340347 , n340346 );
nand ( n340348 , n20482 , n340347 );
buf ( n340349 , n340348 );
nand ( n340350 , n340349 , n335114 );
nand ( n20491 , n20477 , n340350 );
xor ( n340352 , n340151 , n340176 );
xor ( n20493 , n340352 , n340290 );
buf ( n340354 , n20493 );
and ( n20495 , n20491 , n340354 );
not ( n340356 , n20491 );
not ( n20497 , n340354 );
and ( n340358 , n340356 , n20497 );
nor ( n340359 , n20495 , n340358 );
buf ( n340360 , n591 );
not ( n20501 , n340360 );
buf ( n340362 , n340133 );
not ( n340363 , n340362 );
or ( n340364 , n20501 , n340363 );
buf ( n20505 , n590 );
not ( n20506 , n20505 );
buf ( n20507 , n336319 );
not ( n20508 , n20507 );
or ( n20509 , n20506 , n20508 );
buf ( n340370 , n16456 );
buf ( n340371 , n335097 );
nand ( n340372 , n340370 , n340371 );
buf ( n340373 , n340372 );
buf ( n340374 , n340373 );
nand ( n340375 , n20509 , n340374 );
buf ( n340376 , n340375 );
buf ( n340377 , n340376 );
buf ( n340378 , n335181 );
nand ( n340379 , n340377 , n340378 );
buf ( n340380 , n340379 );
buf ( n340381 , n340380 );
nand ( n340382 , n340364 , n340381 );
buf ( n340383 , n340382 );
not ( n20524 , n340383 );
and ( n340385 , n340359 , n20524 );
not ( n340386 , n340359 );
and ( n20527 , n340386 , n340383 );
nor ( n340388 , n340385 , n20527 );
buf ( n340389 , n340388 );
buf ( n340390 , n336275 );
not ( n20531 , n340390 );
buf ( n340392 , n335097 );
not ( n340393 , n340392 );
and ( n340394 , n20531 , n340393 );
buf ( n340395 , n336463 );
buf ( n340396 , n335097 );
and ( n20537 , n340395 , n340396 );
nor ( n340398 , n340394 , n20537 );
buf ( n340399 , n340398 );
buf ( n20540 , n340399 );
not ( n20541 , n20540 );
buf ( n20542 , n338457 );
not ( n20543 , n20542 );
and ( n20544 , n20541 , n20543 );
buf ( n340405 , n340376 );
buf ( n340406 , n591 );
and ( n340407 , n340405 , n340406 );
nor ( n20548 , n20544 , n340407 );
buf ( n340409 , n20548 );
not ( n340410 , n340409 );
and ( n340411 , n588 , n339981 );
not ( n20552 , n588 );
and ( n340413 , n20552 , n16430 );
or ( n340414 , n340411 , n340413 );
buf ( n340415 , n340414 );
not ( n340416 , n340415 );
buf ( n340417 , n340416 );
buf ( n340418 , n340417 );
not ( n20559 , n340418 );
buf ( n340420 , n335111 );
not ( n340421 , n340420 );
and ( n20562 , n20559 , n340421 );
buf ( n340423 , n340349 );
buf ( n340424 , n15275 );
and ( n20565 , n340423 , n340424 );
nor ( n20566 , n20562 , n20565 );
buf ( n340427 , n20566 );
not ( n340428 , n340427 );
and ( n340429 , n340410 , n340428 );
buf ( n340430 , n340427 );
buf ( n340431 , n340409 );
nand ( n20572 , n340430 , n340431 );
buf ( n340433 , n20572 );
xor ( n340434 , n340182 , n340271 );
xor ( n20575 , n340434 , n340285 );
buf ( n340436 , n20575 );
and ( n20577 , n340433 , n340436 );
nor ( n340438 , n340429 , n20577 );
buf ( n340439 , n340438 );
nand ( n20580 , n340389 , n340439 );
buf ( n340441 , n20580 );
buf ( n340442 , n340441 );
buf ( n340443 , n340186 );
buf ( n340444 , n340253 );
xor ( n20585 , n340443 , n340444 );
buf ( n340446 , n340263 );
xnor ( n20587 , n20585 , n340446 );
buf ( n20588 , n20587 );
buf ( n340449 , n20588 );
buf ( n340450 , n15275 );
not ( n20591 , n340450 );
buf ( n340452 , n340414 );
not ( n340453 , n340452 );
or ( n340454 , n20591 , n340453 );
and ( n20595 , n588 , n336662 );
not ( n20596 , n588 );
and ( n20597 , n20596 , n337990 );
or ( n340458 , n20595 , n20597 );
buf ( n340459 , n340458 );
buf ( n340460 , n335114 );
nand ( n20601 , n340459 , n340460 );
buf ( n340462 , n20601 );
buf ( n340463 , n340462 );
nand ( n340464 , n340454 , n340463 );
buf ( n340465 , n340464 );
buf ( n340466 , n340465 );
xor ( n20607 , n340449 , n340466 );
xor ( n340468 , n340250 , n340233 );
buf ( n340469 , n340468 );
buf ( n340470 , n15275 );
not ( n20611 , n340470 );
buf ( n340472 , n340458 );
not ( n340473 , n340472 );
or ( n20614 , n20611 , n340473 );
buf ( n20615 , n588 );
not ( n20616 , n20615 );
buf ( n20617 , n337332 );
not ( n20618 , n20617 );
or ( n20619 , n20616 , n20618 );
buf ( n20620 , n337278 );
buf ( n340481 , n334972 );
nand ( n340482 , n20620 , n340481 );
buf ( n340483 , n340482 );
buf ( n340484 , n340483 );
nand ( n20625 , n20619 , n340484 );
buf ( n340486 , n20625 );
buf ( n20627 , n340486 );
buf ( n340488 , n335114 );
nand ( n340489 , n20627 , n340488 );
buf ( n340490 , n340489 );
buf ( n340491 , n340490 );
nand ( n340492 , n20614 , n340491 );
buf ( n340493 , n340492 );
buf ( n340494 , n340493 );
xor ( n340495 , n340469 , n340494 );
buf ( n340496 , n340486 );
buf ( n340497 , n15275 );
and ( n340498 , n340496 , n340497 );
buf ( n340499 , n588 );
not ( n20640 , n340499 );
buf ( n340501 , n338015 );
not ( n340502 , n340501 );
or ( n20643 , n20640 , n340502 );
buf ( n340504 , n17456 );
buf ( n340505 , n334972 );
nand ( n340506 , n340504 , n340505 );
buf ( n340507 , n340506 );
buf ( n340508 , n340507 );
nand ( n20649 , n20643 , n340508 );
buf ( n340510 , n20649 );
buf ( n340511 , n340510 );
buf ( n340512 , n335114 );
and ( n20653 , n340511 , n340512 );
buf ( n340514 , n20653 );
buf ( n340515 , n340514 );
nor ( n20656 , n340498 , n340515 );
buf ( n340517 , n20656 );
buf ( n340518 , n15115 );
buf ( n340519 , n337364 );
nand ( n340520 , n340518 , n340519 );
buf ( n340521 , n340520 );
xor ( n20662 , n340517 , n340521 );
buf ( n340523 , n588 );
buf ( n340524 , n337361 );
and ( n20665 , n340523 , n340524 );
buf ( n340526 , n337364 );
buf ( n340527 , n334972 );
and ( n20668 , n340526 , n340527 );
nor ( n20669 , n20665 , n20668 );
buf ( n340530 , n20669 );
not ( n20671 , n340530 );
not ( n340532 , n335111 );
and ( n20673 , n20671 , n340532 );
and ( n20674 , n340510 , n15275 );
nor ( n340535 , n20673 , n20674 );
buf ( n340536 , n340535 );
buf ( n340537 , n589 );
buf ( n340538 , n590 );
or ( n340539 , n340537 , n340538 );
buf ( n340540 , n337364 );
nand ( n340541 , n340539 , n340540 );
buf ( n340542 , n340541 );
buf ( n340543 , n340542 );
buf ( n340544 , n589 );
buf ( n340545 , n590 );
and ( n340546 , n340544 , n340545 );
buf ( n340547 , n334972 );
nor ( n20688 , n340546 , n340547 );
buf ( n340549 , n20688 );
buf ( n340550 , n340549 );
nand ( n340551 , n340543 , n340550 );
buf ( n340552 , n340551 );
buf ( n340553 , n340552 );
nor ( n20694 , n340536 , n340553 );
buf ( n340555 , n20694 );
not ( n340556 , n340555 );
and ( n20697 , n20662 , n340556 );
and ( n20698 , n340517 , n340521 );
or ( n20699 , n20697 , n20698 );
not ( n340560 , n20699 );
buf ( n20701 , n340560 );
and ( n20702 , n340495 , n20701 );
and ( n340563 , n340469 , n340494 );
or ( n20704 , n20702 , n340563 );
buf ( n340565 , n20704 );
buf ( n340566 , n340565 );
xnor ( n340567 , n20607 , n340566 );
buf ( n340568 , n340567 );
buf ( n340569 , n340399 );
not ( n340570 , n340569 );
buf ( n340571 , n340570 );
and ( n20712 , n340571 , n591 );
xor ( n340573 , n336259 , n590 );
buf ( n340574 , n340573 );
buf ( n340575 , n335181 );
and ( n20716 , n340574 , n340575 );
buf ( n340577 , n20716 );
nor ( n340578 , n20712 , n340577 );
nand ( n20719 , n340568 , n340578 );
not ( n340580 , n20719 );
buf ( n340581 , n591 );
not ( n20722 , n340581 );
buf ( n340583 , n340573 );
not ( n340584 , n340583 );
or ( n20725 , n20722 , n340584 );
buf ( n340586 , n590 );
not ( n340587 , n340586 );
buf ( n340588 , n336293 );
not ( n340589 , n340588 );
or ( n340590 , n340587 , n340589 );
buf ( n340591 , n16430 );
buf ( n340592 , n335097 );
nand ( n340593 , n340591 , n340592 );
buf ( n340594 , n340593 );
buf ( n340595 , n340594 );
nand ( n340596 , n340590 , n340595 );
buf ( n340597 , n340596 );
buf ( n340598 , n340597 );
buf ( n340599 , n335181 );
nand ( n340600 , n340598 , n340599 );
buf ( n20738 , n340600 );
buf ( n340602 , n20738 );
nand ( n340603 , n20725 , n340602 );
buf ( n340604 , n340603 );
buf ( n340605 , n340604 );
xor ( n20743 , n340469 , n340494 );
xor ( n20744 , n20743 , n20701 );
buf ( n340608 , n20744 );
buf ( n340609 , n340608 );
xor ( n340610 , n340605 , n340609 );
buf ( n340611 , n590 );
not ( n20749 , n340611 );
buf ( n340613 , n336662 );
not ( n340614 , n340613 );
or ( n20752 , n20749 , n340614 );
buf ( n340616 , n16799 );
buf ( n20754 , n335097 );
nand ( n20755 , n340616 , n20754 );
buf ( n340619 , n20755 );
buf ( n340620 , n340619 );
nand ( n340621 , n20752 , n340620 );
buf ( n340622 , n340621 );
buf ( n340623 , n340622 );
not ( n340624 , n340623 );
buf ( n20756 , n340624 );
buf ( n340626 , n20756 );
not ( n340627 , n340626 );
buf ( n340628 , n338457 );
not ( n340629 , n340628 );
and ( n20761 , n340627 , n340629 );
buf ( n340631 , n340597 );
buf ( n340632 , n591 );
and ( n340633 , n340631 , n340632 );
nor ( n340634 , n20761 , n340633 );
buf ( n340635 , n340634 );
buf ( n340636 , n340635 );
not ( n340637 , n340636 );
buf ( n340638 , n340637 );
buf ( n340639 , n340638 );
xor ( n340640 , n340517 , n340521 );
not ( n340641 , n340555 );
xor ( n20766 , n340640 , n340641 );
buf ( n340643 , n20766 );
not ( n20768 , n340643 );
buf ( n340645 , n20768 );
buf ( n340646 , n340645 );
nand ( n340647 , n340639 , n340646 );
buf ( n340648 , n340647 );
buf ( n340649 , n340648 );
buf ( n340650 , n340635 );
buf ( n340651 , n20766 );
nand ( n340652 , n340650 , n340651 );
buf ( n340653 , n340652 );
buf ( n340654 , n340653 );
buf ( n340655 , n590 );
not ( n340656 , n340655 );
buf ( n340657 , n337332 );
not ( n340658 , n340657 );
or ( n340659 , n340656 , n340658 );
buf ( n340660 , n337278 );
buf ( n340661 , n335097 );
nand ( n340662 , n340660 , n340661 );
buf ( n340663 , n340662 );
buf ( n340664 , n340663 );
nand ( n340665 , n340659 , n340664 );
buf ( n340666 , n340665 );
buf ( n340667 , n340666 );
not ( n340668 , n340667 );
buf ( n340669 , n340668 );
buf ( n340670 , n340669 );
not ( n20785 , n340670 );
buf ( n340672 , n338457 );
not ( n340673 , n340672 );
and ( n340674 , n20785 , n340673 );
buf ( n340675 , n340622 );
buf ( n340676 , n591 );
and ( n340677 , n340675 , n340676 );
nor ( n20792 , n340674 , n340677 );
buf ( n20793 , n20792 );
buf ( n340680 , n20793 );
xnor ( n20795 , n340535 , n340552 );
buf ( n340682 , n20795 );
nand ( n340683 , n340680 , n340682 );
buf ( n340684 , n340683 );
not ( n20799 , n340684 );
buf ( n340686 , n15239 );
buf ( n340687 , n337361 );
nor ( n340688 , n340686 , n340687 );
buf ( n340689 , n340688 );
buf ( n340690 , n340689 );
not ( n340691 , n337364 );
not ( n340692 , n338457 );
and ( n20807 , n340691 , n340692 );
buf ( n340694 , n590 );
not ( n20809 , n340694 );
buf ( n340696 , n337313 );
not ( n20811 , n340696 );
or ( n340698 , n20809 , n20811 );
buf ( n340699 , n338015 );
not ( n20814 , n340699 );
buf ( n340701 , n335097 );
nand ( n340702 , n20814 , n340701 );
buf ( n340703 , n340702 );
buf ( n340704 , n340703 );
nand ( n340705 , n340698 , n340704 );
buf ( n340706 , n340705 );
and ( n340707 , n340706 , n591 );
nor ( n20822 , n20807 , n340707 );
buf ( n340709 , n20822 );
nand ( n340710 , n337364 , n591 );
nand ( n340711 , n340710 , n590 );
buf ( n340712 , n340711 );
nor ( n340713 , n340709 , n340712 );
buf ( n340714 , n340713 );
buf ( n340715 , n340714 );
xor ( n340716 , n340690 , n340715 );
buf ( n340717 , n591 );
not ( n20832 , n340717 );
buf ( n340719 , n340666 );
not ( n20833 , n340719 );
or ( n340721 , n20832 , n20833 );
buf ( n340722 , n340706 );
buf ( n340723 , n335181 );
nand ( n340724 , n340722 , n340723 );
buf ( n340725 , n340724 );
buf ( n340726 , n340725 );
nand ( n340727 , n340721 , n340726 );
buf ( n340728 , n340727 );
buf ( n340729 , n340728 );
and ( n340730 , n340716 , n340729 );
and ( n340731 , n340690 , n340715 );
or ( n20844 , n340730 , n340731 );
buf ( n340733 , n20844 );
not ( n20846 , n340733 );
or ( n340735 , n20799 , n20846 );
buf ( n340736 , n20795 );
not ( n20849 , n340736 );
buf ( n340738 , n20849 );
buf ( n340739 , n340738 );
buf ( n340740 , n20793 );
not ( n340741 , n340740 );
buf ( n340742 , n340741 );
buf ( n340743 , n340742 );
nand ( n340744 , n340739 , n340743 );
buf ( n340745 , n340744 );
nand ( n20858 , n340735 , n340745 );
buf ( n340747 , n20858 );
nand ( n20860 , n340654 , n340747 );
buf ( n20861 , n20860 );
buf ( n340750 , n20861 );
nand ( n20863 , n340649 , n340750 );
buf ( n340752 , n20863 );
buf ( n340753 , n340752 );
and ( n340754 , n340610 , n340753 );
and ( n340755 , n340605 , n340609 );
or ( n340756 , n340754 , n340755 );
buf ( n340757 , n340756 );
not ( n340758 , n340757 );
or ( n20871 , n340580 , n340758 );
buf ( n340760 , n340568 );
not ( n340761 , n340760 );
buf ( n340762 , n340761 );
not ( n340763 , n340578 );
nand ( n20876 , n340762 , n340763 );
nand ( n20877 , n20871 , n20876 );
not ( n340766 , n20877 );
buf ( n340767 , n340409 );
buf ( n340768 , n340427 );
buf ( n340769 , n340436 );
not ( n340770 , n340769 );
buf ( n340771 , n340770 );
buf ( n340772 , n340771 );
and ( n340773 , n340768 , n340772 );
not ( n340774 , n340768 );
buf ( n340775 , n340436 );
and ( n340776 , n340774 , n340775 );
nor ( n340777 , n340773 , n340776 );
buf ( n340778 , n340777 );
buf ( n340779 , n340778 );
nand ( n340780 , n340767 , n340779 );
buf ( n340781 , n340780 );
or ( n20894 , n20588 , n340465 );
nand ( n20895 , n20894 , n340565 );
buf ( n340784 , n340465 );
buf ( n340785 , n20588 );
nand ( n20898 , n340784 , n340785 );
buf ( n340787 , n20898 );
nand ( n20900 , n20895 , n340787 );
not ( n340789 , n20900 );
nand ( n340790 , n340781 , n340789 );
buf ( n340791 , n340409 );
not ( n20904 , n340791 );
buf ( n340793 , n20904 );
buf ( n340794 , n340793 );
buf ( n340795 , n340778 );
not ( n20908 , n340795 );
buf ( n340797 , n20908 );
buf ( n340798 , n340797 );
nand ( n340799 , n340794 , n340798 );
buf ( n340800 , n340799 );
buf ( n340801 , n340800 );
not ( n20914 , n340801 );
buf ( n340803 , n20914 );
nor ( n340804 , n340790 , n340803 );
or ( n20917 , n340766 , n340804 );
buf ( n340806 , n340781 );
buf ( n340807 , n340800 );
nand ( n340808 , n340806 , n340807 );
buf ( n340809 , n340808 );
buf ( n340810 , n340809 );
buf ( n340811 , n20900 );
nand ( n20924 , n340810 , n340811 );
buf ( n340813 , n20924 );
nand ( n20926 , n20917 , n340813 );
buf ( n340815 , n20926 );
nand ( n340816 , n340442 , n340815 );
buf ( n340817 , n340816 );
buf ( n340818 , n340817 );
buf ( n340819 , n340388 );
not ( n340820 , n340819 );
buf ( n340821 , n340820 );
buf ( n340822 , n340821 );
buf ( n20935 , n340438 );
not ( n340824 , n20935 );
buf ( n340825 , n340824 );
buf ( n340826 , n340825 );
nand ( n340827 , n340822 , n340826 );
buf ( n340828 , n340827 );
buf ( n340829 , n340828 );
nand ( n340830 , n340818 , n340829 );
buf ( n340831 , n340830 );
not ( n20944 , n340831 );
buf ( n340833 , n340297 );
not ( n340834 , n340833 );
buf ( n340835 , n340325 );
not ( n20948 , n340835 );
or ( n340837 , n340834 , n20948 );
buf ( n340838 , n340297 );
buf ( n340839 , n340325 );
or ( n340840 , n340838 , n340839 );
nand ( n340841 , n340837 , n340840 );
buf ( n340842 , n340841 );
buf ( n340843 , n340842 );
buf ( n20956 , n20283 );
and ( n20957 , n340843 , n20956 );
not ( n340846 , n340843 );
buf ( n340847 , n20280 );
and ( n340848 , n340846 , n340847 );
nor ( n20961 , n20957 , n340848 );
buf ( n340850 , n20961 );
buf ( n340851 , n340850 );
not ( n20964 , n20524 );
not ( n340853 , n20491 );
not ( n20966 , n340853 );
and ( n20967 , n20964 , n20966 );
nand ( n340856 , n20524 , n340853 );
and ( n20969 , n340856 , n340354 );
nor ( n340858 , n20967 , n20969 );
buf ( n340859 , n340858 );
nand ( n340860 , n340851 , n340859 );
buf ( n340861 , n340860 );
not ( n20974 , n340861 );
or ( n340863 , n20944 , n20974 );
buf ( n20976 , n340858 );
not ( n340865 , n20976 );
buf ( n340866 , n340865 );
buf ( n340867 , n340866 );
buf ( n340868 , n340850 );
not ( n20981 , n340868 );
buf ( n20982 , n20981 );
buf ( n340871 , n20982 );
nand ( n340872 , n340867 , n340871 );
buf ( n340873 , n340872 );
nand ( n20986 , n340863 , n340873 );
not ( n340875 , n20986 );
or ( n20988 , n340331 , n340875 );
buf ( n340877 , n340119 );
not ( n340878 , n340877 );
buf ( n340879 , n340878 );
buf ( n340880 , n340327 );
not ( n20993 , n340880 );
buf ( n340882 , n20993 );
nand ( n340883 , n340879 , n340882 );
nand ( n340884 , n20988 , n340883 );
not ( n20997 , n340884 );
or ( n340886 , n20253 , n20997 );
buf ( n340887 , n340109 );
not ( n21000 , n340887 );
buf ( n340889 , n340079 );
nand ( n340890 , n21000 , n340889 );
buf ( n340891 , n340890 );
nand ( n340892 , n340886 , n340891 );
not ( n340893 , n340892 );
buf ( n340894 , n339918 );
buf ( n340895 , n339933 );
xor ( n340896 , n340894 , n340895 );
buf ( n340897 , n339708 );
xnor ( n21010 , n340896 , n340897 );
buf ( n21011 , n21010 );
buf ( n21012 , n21011 );
buf ( n340901 , n340106 );
buf ( n340902 , n340099 );
buf ( n340903 , n340086 );
or ( n340904 , n340902 , n340903 );
buf ( n340905 , n340904 );
buf ( n340906 , n340905 );
and ( n21019 , n340901 , n340906 );
and ( n21020 , n340087 , n340100 );
buf ( n340909 , n21020 );
buf ( n340910 , n340909 );
nor ( n340911 , n21019 , n340910 );
buf ( n340912 , n340911 );
buf ( n340913 , n340912 );
nand ( n340914 , n21012 , n340913 );
buf ( n340915 , n340914 );
not ( n21028 , n340915 );
or ( n340917 , n340893 , n21028 );
buf ( n340918 , n21011 );
not ( n21031 , n340918 );
buf ( n21032 , n21031 );
buf ( n21033 , n21032 );
buf ( n340922 , n340912 );
not ( n21035 , n340922 );
buf ( n21036 , n21035 );
buf ( n340925 , n21036 );
nand ( n340926 , n21033 , n340925 );
buf ( n340927 , n340926 );
nand ( n21040 , n340917 , n340927 );
buf ( n340929 , n21040 );
not ( n340930 , n340929 );
or ( n340931 , n339943 , n340930 );
buf ( n340932 , n339938 );
not ( n21045 , n340932 );
buf ( n340934 , n21045 );
buf ( n340935 , n340934 );
buf ( n340936 , n339687 );
not ( n340937 , n340936 );
buf ( n340938 , n340937 );
buf ( n340939 , n340938 );
nand ( n21052 , n340935 , n340939 );
buf ( n340941 , n21052 );
buf ( n340942 , n340941 );
nand ( n340943 , n340931 , n340942 );
buf ( n340944 , n340943 );
buf ( n340945 , n340944 );
not ( n340946 , n340945 );
buf ( n340947 , n339427 );
buf ( n340948 , n339442 );
xor ( n340949 , n340947 , n340948 );
buf ( n340950 , n339451 );
xnor ( n21063 , n340949 , n340950 );
buf ( n21064 , n21063 );
buf ( n340953 , n21064 );
not ( n21066 , n340953 );
not ( n340955 , n339669 );
not ( n340956 , n340955 );
not ( n21069 , n339660 );
and ( n21070 , n340956 , n21069 );
nand ( n21071 , n339660 , n340955 );
and ( n340960 , n339674 , n21071 );
nor ( n340961 , n21070 , n340960 );
not ( n21074 , n340961 );
not ( n21075 , n21074 );
buf ( n340964 , n591 );
not ( n340965 , n340964 );
buf ( n340966 , n339304 );
not ( n21079 , n340966 );
buf ( n340968 , n21079 );
buf ( n340969 , n340968 );
not ( n340970 , n340969 );
or ( n340971 , n340965 , n340970 );
buf ( n340972 , n339619 );
buf ( n340973 , n335181 );
nand ( n21086 , n340972 , n340973 );
buf ( n340975 , n21086 );
buf ( n340976 , n340975 );
nand ( n21089 , n340971 , n340976 );
buf ( n340978 , n21089 );
not ( n21091 , n340978 );
or ( n340980 , n21075 , n21091 );
or ( n340981 , n340978 , n21074 );
nand ( n21094 , n340980 , n340981 );
buf ( n340983 , n21094 );
not ( n21096 , n340983 );
and ( n340985 , n21066 , n21096 );
buf ( n340986 , n21064 );
buf ( n340987 , n21094 );
and ( n21100 , n340986 , n340987 );
nor ( n21101 , n340985 , n21100 );
buf ( n340990 , n21101 );
buf ( n340991 , n340990 );
buf ( n340992 , n339677 );
buf ( n340993 , n339641 );
not ( n340994 , n340993 );
buf ( n340995 , n339609 );
buf ( n21108 , n340995 );
buf ( n340997 , n21108 );
buf ( n340998 , n340997 );
nand ( n340999 , n340994 , n340998 );
buf ( n341000 , n340999 );
buf ( n341001 , n341000 );
and ( n21114 , n340992 , n341001 );
buf ( n341003 , n339641 );
not ( n21116 , n341003 );
buf ( n341005 , n340997 );
nor ( n341006 , n21116 , n341005 );
buf ( n341007 , n341006 );
buf ( n341008 , n341007 );
nor ( n341009 , n21114 , n341008 );
buf ( n341010 , n341009 );
buf ( n341011 , n341010 );
nand ( n341012 , n340991 , n341011 );
buf ( n341013 , n341012 );
buf ( n341014 , n341013 );
not ( n21127 , n341014 );
or ( n341016 , n340946 , n21127 );
buf ( n341017 , n340990 );
not ( n21130 , n341017 );
buf ( n341019 , n21130 );
buf ( n341020 , n341019 );
buf ( n341021 , n341010 );
not ( n21134 , n341021 );
buf ( n341023 , n21134 );
buf ( n341024 , n341023 );
nand ( n21137 , n341020 , n341024 );
buf ( n341026 , n21137 );
buf ( n341027 , n341026 );
nand ( n341028 , n341016 , n341027 );
buf ( n341029 , n341028 );
buf ( n341030 , n341029 );
not ( n341031 , n339361 );
not ( n341032 , n339463 );
or ( n21145 , n341031 , n341032 );
or ( n341034 , n339361 , n339463 );
nand ( n341035 , n21145 , n341034 );
not ( n341036 , n341035 );
nand ( n21149 , n341036 , n339365 );
not ( n341038 , n339365 );
nand ( n341039 , n341038 , n341035 );
nand ( n21152 , n21149 , n341039 );
buf ( n341041 , n340978 );
not ( n341042 , n341041 );
buf ( n341043 , n340961 );
nand ( n21156 , n341042 , n341043 );
buf ( n341045 , n21156 );
not ( n21158 , n341045 );
not ( n21159 , n21064 );
or ( n341048 , n21158 , n21159 );
buf ( n341049 , n340961 );
not ( n341050 , n341049 );
buf ( n341051 , n340978 );
nand ( n21164 , n341050 , n341051 );
buf ( n341053 , n21164 );
nand ( n341054 , n341048 , n341053 );
or ( n21167 , n21152 , n341054 );
buf ( n341056 , n21167 );
nand ( n341057 , n341030 , n341056 );
buf ( n341058 , n341057 );
buf ( n341059 , n341058 );
not ( n341060 , n21149 );
not ( n341061 , n341039 );
or ( n21174 , n341060 , n341061 );
nand ( n341063 , n21174 , n341054 );
buf ( n341064 , n341063 );
nand ( n21177 , n341059 , n341064 );
buf ( n21178 , n21177 );
not ( n341067 , n21178 );
or ( n341068 , n339472 , n341067 );
buf ( n341069 , n339350 );
not ( n341070 , n341069 );
buf ( n341071 , n341070 );
buf ( n341072 , n341071 );
buf ( n341073 , n19608 );
not ( n21186 , n341073 );
buf ( n341075 , n21186 );
buf ( n341076 , n341075 );
nand ( n21189 , n341072 , n341076 );
buf ( n341078 , n21189 );
nand ( n341079 , n341068 , n341078 );
buf ( n341080 , n341079 );
xor ( n341081 , n339041 , n339042 );
buf ( n341082 , n341081 );
buf ( n341083 , n341082 );
buf ( n341084 , n338877 );
and ( n341085 , n341083 , n341084 );
not ( n341086 , n341083 );
buf ( n341087 , n338880 );
and ( n341088 , n341086 , n341087 );
nor ( n341089 , n341085 , n341088 );
buf ( n341090 , n341089 );
buf ( n341091 , n341090 );
xor ( n341092 , n339327 , n339341 );
and ( n341093 , n341092 , n339348 );
and ( n21206 , n339327 , n339341 );
or ( n341095 , n341093 , n21206 );
buf ( n341096 , n341095 );
buf ( n341097 , n341096 );
nand ( n341098 , n341091 , n341097 );
buf ( n341099 , n341098 );
buf ( n341100 , n341099 );
and ( n21213 , n339049 , n341080 , n341100 );
buf ( n21214 , n21213 );
buf ( n341103 , n21214 );
buf ( n341104 , n339048 );
not ( n21217 , n341104 );
buf ( n341106 , n21217 );
buf ( n341107 , n341106 );
buf ( n341108 , n341090 );
not ( n341109 , n341108 );
buf ( n341110 , n341109 );
buf ( n341111 , n341110 );
buf ( n21224 , n341096 );
not ( n341113 , n21224 );
buf ( n341114 , n341113 );
buf ( n341115 , n341114 );
nand ( n341116 , n341111 , n341115 );
buf ( n341117 , n341116 );
buf ( n341118 , n341117 );
or ( n341119 , n341107 , n341118 );
buf ( n341120 , n19010 );
buf ( n341121 , n19185 );
or ( n341122 , n341120 , n341121 );
buf ( n341123 , n341122 );
buf ( n341124 , n341123 );
nand ( n341125 , n341119 , n341124 );
buf ( n341126 , n341125 );
buf ( n341127 , n341126 );
nor ( n341128 , n341103 , n341127 );
buf ( n341129 , n341128 );
buf ( n341130 , n341129 );
buf ( n341131 , n18967 );
not ( n341132 , n341131 );
buf ( n341133 , n338840 );
not ( n341134 , n341133 );
or ( n21245 , n341132 , n341134 );
buf ( n341136 , n338847 );
nand ( n341137 , n21245 , n341136 );
buf ( n341138 , n341137 );
buf ( n341139 , n341138 );
buf ( n341140 , n18967 );
not ( n21251 , n341140 );
buf ( n341142 , n338843 );
nand ( n341143 , n21251 , n341142 );
buf ( n341144 , n341143 );
buf ( n341145 , n341144 );
nand ( n341146 , n341139 , n341145 );
buf ( n341147 , n341146 );
buf ( n341148 , n341147 );
not ( n341149 , n341148 );
buf ( n341150 , n334868 );
not ( n21261 , n341150 );
buf ( n341152 , n17746 );
not ( n341153 , n341152 );
or ( n21264 , n21261 , n341153 );
buf ( n341155 , n338801 );
buf ( n341156 , n334917 );
nand ( n21267 , n341155 , n341156 );
buf ( n341158 , n21267 );
buf ( n341159 , n341158 );
nand ( n341160 , n21264 , n341159 );
buf ( n341161 , n341160 );
buf ( n341162 , n341161 );
not ( n21272 , n341162 );
buf ( n341164 , n21272 );
buf ( n341165 , n341164 );
nand ( n21275 , n341149 , n341165 );
buf ( n341167 , n21275 );
buf ( n341168 , n341167 );
xor ( n341169 , n337671 , n337691 );
xor ( n21279 , n341169 , n337696 );
buf ( n341171 , n21279 );
buf ( n341172 , n341171 );
and ( n341173 , n341168 , n341172 );
buf ( n341174 , n341161 );
buf ( n341175 , n341147 );
and ( n341176 , n341174 , n341175 );
buf ( n341177 , n341176 );
buf ( n341178 , n341177 );
nor ( n341179 , n341173 , n341178 );
buf ( n341180 , n341179 );
not ( n21290 , n15115 );
not ( n341182 , n337585 );
or ( n341183 , n21290 , n341182 );
buf ( n341184 , n586 );
buf ( n341185 , n15622 );
and ( n341186 , n341184 , n341185 );
not ( n21296 , n341184 );
buf ( n341188 , n17055 );
and ( n21298 , n21296 , n341188 );
nor ( n341190 , n341186 , n21298 );
buf ( n341191 , n341190 );
not ( n21301 , n341191 );
nand ( n21302 , n21301 , n15164 );
nand ( n21303 , n341183 , n21302 );
not ( n341195 , n21303 );
xor ( n341196 , n341180 , n341195 );
and ( n21306 , n337559 , n15275 );
not ( n21307 , n588 );
and ( n21308 , n21307 , n16686 );
not ( n341200 , n21307 );
buf ( n341201 , n335514 );
not ( n21311 , n341201 );
buf ( n341203 , n21311 );
and ( n21313 , n341200 , n341203 );
nor ( n341205 , n21308 , n21313 );
and ( n341206 , n341205 , n335114 );
nor ( n21316 , n21306 , n341206 );
xor ( n21317 , n341196 , n21316 );
buf ( n341209 , n21317 );
not ( n21319 , n341209 );
buf ( n341211 , n21319 );
buf ( n341212 , n341211 );
not ( n341213 , n341212 );
buf ( n341214 , n335114 );
not ( n21324 , n341214 );
buf ( n341216 , n338440 );
not ( n341217 , n341216 );
or ( n21327 , n21324 , n341217 );
buf ( n341219 , n341205 );
buf ( n341220 , n15275 );
nand ( n21330 , n341219 , n341220 );
buf ( n21331 , n21330 );
buf ( n341223 , n21331 );
nand ( n21333 , n21327 , n341223 );
buf ( n341225 , n21333 );
not ( n21335 , n341225 );
buf ( n341227 , n335181 );
not ( n21337 , n341227 );
buf ( n341229 , n18604 );
not ( n341230 , n341229 );
or ( n21340 , n21337 , n341230 );
and ( n21341 , n590 , n336024 );
not ( n21342 , n590 );
and ( n341234 , n21342 , n336030 );
or ( n341235 , n21341 , n341234 );
buf ( n341236 , n341235 );
buf ( n341237 , n591 );
nand ( n21347 , n341236 , n341237 );
buf ( n341239 , n21347 );
buf ( n341240 , n341239 );
nand ( n21350 , n21340 , n341240 );
buf ( n341242 , n21350 );
not ( n21352 , n341242 );
or ( n341244 , n21335 , n21352 );
buf ( n341245 , n341225 );
buf ( n341246 , n341242 );
or ( n21356 , n341245 , n341246 );
xor ( n21357 , n338737 , n338762 );
and ( n341249 , n21357 , n338852 );
and ( n341250 , n338737 , n338762 );
or ( n21360 , n341249 , n341250 );
buf ( n341252 , n21360 );
buf ( n341253 , n341252 );
nand ( n21363 , n21356 , n341253 );
buf ( n21364 , n21363 );
nand ( n21365 , n341244 , n21364 );
not ( n21366 , n21365 );
buf ( n341258 , n21366 );
not ( n341259 , n341258 );
or ( n341260 , n341213 , n341259 );
buf ( n341261 , n21317 );
buf ( n341262 , n21365 );
nand ( n341263 , n341261 , n341262 );
buf ( n341264 , n341263 );
buf ( n341265 , n341264 );
nand ( n21375 , n341260 , n341265 );
buf ( n341267 , n21375 );
buf ( n341268 , n341267 );
buf ( n341269 , n17752 );
buf ( n341270 , n337703 );
and ( n21380 , n341269 , n341270 );
not ( n21381 , n341269 );
buf ( n341273 , n337700 );
and ( n341274 , n21381 , n341273 );
nor ( n341275 , n21380 , n341274 );
buf ( n341276 , n341275 );
and ( n341277 , n341276 , n17740 );
not ( n341278 , n341276 );
not ( n21388 , n17740 );
and ( n341280 , n341278 , n21388 );
nor ( n341281 , n341277 , n341280 );
buf ( n341282 , n341281 );
buf ( n341283 , n341147 );
buf ( n341284 , n341164 );
xor ( n341285 , n341283 , n341284 );
buf ( n341286 , n341171 );
xnor ( n341287 , n341285 , n341286 );
buf ( n341288 , n341287 );
buf ( n341289 , n341288 );
not ( n341290 , n341289 );
not ( n341291 , n338808 );
nand ( n21399 , n341291 , n338786 );
and ( n341293 , n21399 , n18988 );
and ( n21401 , n338808 , n338785 );
nor ( n21402 , n341293 , n21401 );
buf ( n341296 , n21402 );
buf ( n21404 , n341191 );
not ( n21405 , n21404 );
buf ( n21406 , n21405 );
buf ( n341300 , n21406 );
buf ( n341301 , n15115 );
and ( n341302 , n341300 , n341301 );
buf ( n341303 , n338751 );
buf ( n341304 , n15163 );
and ( n341305 , n341303 , n341304 );
buf ( n341306 , n341305 );
buf ( n341307 , n341306 );
nor ( n341308 , n341302 , n341307 );
buf ( n341309 , n341308 );
buf ( n341310 , n341309 );
nand ( n341311 , n341296 , n341310 );
buf ( n341312 , n341311 );
buf ( n341313 , n341312 );
not ( n341314 , n341313 );
or ( n21422 , n341290 , n341314 );
buf ( n341316 , n21402 );
not ( n341317 , n341316 );
buf ( n341318 , n341317 );
buf ( n341319 , n341318 );
buf ( n341320 , n15115 );
not ( n21427 , n341320 );
buf ( n341322 , n21406 );
not ( n21429 , n341322 );
or ( n341324 , n21427 , n21429 );
buf ( n341325 , n341306 );
not ( n21430 , n341325 );
buf ( n341327 , n21430 );
buf ( n341328 , n341327 );
nand ( n341329 , n341324 , n341328 );
buf ( n21431 , n341329 );
buf ( n341331 , n21431 );
nand ( n21433 , n341319 , n341331 );
buf ( n21434 , n21433 );
buf ( n341334 , n21434 );
nand ( n21436 , n21422 , n341334 );
buf ( n341336 , n21436 );
buf ( n341337 , n341336 );
xor ( n341338 , n341282 , n341337 );
buf ( n21440 , n341235 );
not ( n341340 , n21440 );
buf ( n341341 , n341340 );
buf ( n341342 , n341341 );
not ( n21444 , n341342 );
buf ( n341344 , n338457 );
not ( n341345 , n341344 );
and ( n21447 , n21444 , n341345 );
buf ( n341347 , n590 );
buf ( n341348 , n15381 );
and ( n21448 , n341347 , n341348 );
not ( n341350 , n341347 );
buf ( n341351 , n336845 );
and ( n341352 , n341350 , n341351 );
or ( n341353 , n21448 , n341352 );
buf ( n341354 , n341353 );
buf ( n341355 , n341354 );
not ( n341356 , n341355 );
buf ( n341357 , n341356 );
buf ( n341358 , n341357 );
buf ( n341359 , n591 );
and ( n341360 , n341358 , n341359 );
nor ( n341361 , n21447 , n341360 );
buf ( n341362 , n341361 );
buf ( n341363 , n341362 );
not ( n341364 , n341363 );
buf ( n341365 , n341364 );
buf ( n341366 , n341365 );
xor ( n341367 , n341338 , n341366 );
buf ( n341368 , n341367 );
buf ( n341369 , n341368 );
not ( n21466 , n341369 );
buf ( n341371 , n21466 );
buf ( n341372 , n341371 );
and ( n341373 , n341268 , n341372 );
not ( n341374 , n341268 );
buf ( n341375 , n341368 );
and ( n341376 , n341374 , n341375 );
nor ( n341377 , n341373 , n341376 );
buf ( n341378 , n341377 );
buf ( n341379 , n341378 );
buf ( n341380 , n341318 );
buf ( n341381 , n21431 );
and ( n21478 , n341380 , n341381 );
not ( n341383 , n341380 );
buf ( n341384 , n341309 );
and ( n21481 , n341383 , n341384 );
nor ( n21482 , n21478 , n21481 );
buf ( n21483 , n21482 );
buf ( n21484 , n341288 );
buf ( n341389 , n21484 );
buf ( n341390 , n341389 );
xnor ( n341391 , n21483 , n341390 );
buf ( n341392 , n341391 );
xor ( n21489 , n338412 , n338446 );
and ( n341394 , n21489 , n338470 );
and ( n341395 , n338412 , n338446 );
or ( n21492 , n341394 , n341395 );
buf ( n21493 , n21492 );
buf ( n341398 , n21493 );
xor ( n21495 , n341392 , n341398 );
buf ( n341400 , n341225 );
buf ( n341401 , n341242 );
xor ( n341402 , n341400 , n341401 );
buf ( n341403 , n341252 );
xnor ( n341404 , n341402 , n341403 );
buf ( n341405 , n341404 );
buf ( n341406 , n341405 );
and ( n341407 , n21495 , n341406 );
and ( n21503 , n341392 , n341398 );
or ( n341409 , n341407 , n21503 );
buf ( n341410 , n341409 );
buf ( n341411 , n341410 );
nand ( n341412 , n341379 , n341411 );
buf ( n341413 , n341412 );
buf ( n341414 , n341413 );
xor ( n341415 , n341392 , n341398 );
xor ( n341416 , n341415 , n341406 );
buf ( n341417 , n341416 );
buf ( n341418 , n341417 );
buf ( n341419 , n338475 );
buf ( n341420 , n338854 );
not ( n21515 , n341420 );
buf ( n341422 , n18869 );
buf ( n21517 , n341422 );
buf ( n341424 , n21517 );
buf ( n341425 , n341424 );
nand ( n21520 , n21515 , n341425 );
buf ( n341427 , n21520 );
buf ( n341428 , n341427 );
and ( n21523 , n341419 , n341428 );
buf ( n341430 , n338854 );
not ( n341431 , n341430 );
buf ( n341432 , n341424 );
nor ( n341433 , n341431 , n341432 );
buf ( n341434 , n341433 );
buf ( n341435 , n341434 );
nor ( n21530 , n21523 , n341435 );
buf ( n341437 , n21530 );
buf ( n341438 , n341437 );
nand ( n341439 , n341418 , n341438 );
buf ( n341440 , n341439 );
buf ( n341441 , n341440 );
nand ( n341442 , n341414 , n341441 );
buf ( n341443 , n341442 );
buf ( n341444 , n341443 );
or ( n341445 , n341130 , n341444 );
buf ( n341446 , n341413 );
buf ( n341447 , n341417 );
buf ( n341448 , n341437 );
nor ( n21543 , n341447 , n341448 );
buf ( n341450 , n21543 );
buf ( n21545 , n341450 );
nand ( n21546 , n341446 , n21545 );
buf ( n21547 , n21546 );
buf ( n341454 , n21547 );
buf ( n341455 , n341378 );
not ( n341456 , n341455 );
buf ( n341457 , n341456 );
buf ( n341458 , n341457 );
buf ( n341459 , n341410 );
not ( n341460 , n341459 );
buf ( n341461 , n341460 );
buf ( n341462 , n341461 );
nand ( n341463 , n341458 , n341462 );
buf ( n341464 , n341463 );
buf ( n341465 , n341464 );
and ( n21560 , n341454 , n341465 );
buf ( n341467 , n21560 );
buf ( n341468 , n341467 );
nand ( n341469 , n341445 , n341468 );
buf ( n341470 , n341469 );
buf ( n341471 , n341470 );
not ( n21566 , n341471 );
xor ( n341473 , n17677 , n17414 );
xnor ( n341474 , n341473 , n17863 );
buf ( n341475 , n341474 );
and ( n21570 , n336835 , n336854 );
not ( n341477 , n336835 );
and ( n21572 , n341477 , n16998 );
nor ( n21573 , n21570 , n21572 );
xor ( n21574 , n21573 , n17041 );
buf ( n341481 , n21574 );
or ( n21576 , n341475 , n341481 );
buf ( n341483 , n21576 );
buf ( n341484 , n21574 );
not ( n341485 , n341484 );
buf ( n341486 , n341474 );
not ( n341487 , n341486 );
or ( n341488 , n341485 , n341487 );
buf ( n341489 , n341354 );
not ( n341490 , n341489 );
buf ( n341491 , n338457 );
not ( n21586 , n341491 );
and ( n341493 , n341490 , n21586 );
buf ( n341494 , n336878 );
buf ( n341495 , n591 );
and ( n21590 , n341494 , n341495 );
nor ( n21591 , n341493 , n21590 );
buf ( n341498 , n21591 );
buf ( n341499 , n341498 );
not ( n21594 , n341499 );
xor ( n341501 , n341180 , n341195 );
and ( n341502 , n341501 , n21316 );
and ( n21597 , n341180 , n341195 );
or ( n341504 , n341502 , n21597 );
buf ( n341505 , n341504 );
not ( n341506 , n341505 );
or ( n21601 , n21594 , n341506 );
xor ( n341508 , n337277 , n337524 );
xor ( n341509 , n341508 , n337534 );
buf ( n341510 , n341509 );
nand ( n21605 , n21601 , n341510 );
buf ( n341512 , n21605 );
buf ( n341513 , n341504 );
not ( n341514 , n341513 );
buf ( n341515 , n341498 );
not ( n21610 , n341515 );
buf ( n21611 , n21610 );
buf ( n341518 , n21611 );
nand ( n21613 , n341514 , n341518 );
buf ( n341520 , n21613 );
nand ( n21615 , n341512 , n341520 );
buf ( n341522 , n21615 );
nand ( n341523 , n341488 , n341522 );
buf ( n341524 , n341523 );
nand ( n21619 , n341483 , n341524 );
and ( n21620 , n17868 , n17398 );
not ( n341527 , n17868 );
and ( n341528 , n341527 , n17397 );
nor ( n21623 , n21620 , n341528 );
and ( n21624 , n21623 , n17395 );
not ( n21625 , n21623 );
not ( n341532 , n17395 );
and ( n341533 , n21625 , n341532 );
nor ( n21628 , n21624 , n341533 );
nor ( n21629 , n21619 , n21628 );
nand ( n21630 , n341512 , n341520 );
not ( n341537 , n21630 );
not ( n341538 , n21574 );
and ( n21633 , n341537 , n341538 );
and ( n341540 , n21615 , n21574 );
nor ( n341541 , n21633 , n341540 );
and ( n21636 , n341541 , n341474 );
not ( n21637 , n341541 );
not ( n341544 , n341474 );
and ( n21639 , n21637 , n341544 );
nor ( n21640 , n21636 , n21639 );
buf ( n341547 , n21640 );
not ( n341548 , n341547 );
buf ( n341549 , n341548 );
buf ( n341550 , n341549 );
buf ( n341551 , n337714 );
buf ( n341552 , n337592 );
xor ( n341553 , n341551 , n341552 );
buf ( n341554 , n337566 );
xnor ( n21649 , n341553 , n341554 );
buf ( n341556 , n21649 );
buf ( n341557 , n341556 );
buf ( n341558 , n341281 );
not ( n341559 , n341558 );
buf ( n341560 , n341559 );
buf ( n341561 , n341560 );
not ( n341562 , n341561 );
buf ( n341563 , n341362 );
not ( n21658 , n341563 );
or ( n341565 , n341562 , n21658 );
buf ( n341566 , n341336 );
nand ( n21661 , n341565 , n341566 );
buf ( n341568 , n21661 );
buf ( n341569 , n341568 );
buf ( n341570 , n341560 );
not ( n21665 , n341570 );
buf ( n341572 , n341365 );
nand ( n341573 , n21665 , n341572 );
buf ( n341574 , n341573 );
buf ( n341575 , n341574 );
nand ( n21670 , n341569 , n341575 );
buf ( n341577 , n21670 );
buf ( n21672 , n341577 );
not ( n341579 , n21672 );
buf ( n341580 , n341579 );
buf ( n341581 , n341580 );
nand ( n341582 , n341557 , n341581 );
buf ( n341583 , n341582 );
buf ( n341584 , n341583 );
not ( n341585 , n341584 );
xor ( n341586 , n341509 , n21611 );
xnor ( n21681 , n341586 , n341504 );
buf ( n341588 , n21681 );
not ( n341589 , n341588 );
or ( n21684 , n341585 , n341589 );
buf ( n341591 , n341556 );
not ( n341592 , n341591 );
buf ( n341593 , n341577 );
nand ( n21688 , n341592 , n341593 );
buf ( n341595 , n21688 );
buf ( n341596 , n341595 );
nand ( n21691 , n21684 , n341596 );
buf ( n341598 , n21691 );
buf ( n341599 , n341598 );
not ( n341600 , n341599 );
buf ( n341601 , n341600 );
buf ( n341602 , n341601 );
nand ( n341603 , n341550 , n341602 );
buf ( n341604 , n341603 );
buf ( n341605 , n341580 );
not ( n341606 , n341605 );
buf ( n341607 , n341556 );
not ( n21702 , n341607 );
buf ( n21703 , n21702 );
buf ( n341610 , n21703 );
not ( n341611 , n341610 );
or ( n21706 , n341606 , n341611 );
not ( n341613 , n341362 );
nand ( n341614 , n341613 , n341281 );
not ( n21709 , n341614 );
not ( n341616 , n341568 );
or ( n341617 , n21709 , n341616 );
nand ( n21712 , n341617 , n341556 );
buf ( n341619 , n21712 );
nand ( n341620 , n21706 , n341619 );
buf ( n341621 , n341620 );
and ( n21716 , n341621 , n21681 );
not ( n341623 , n341621 );
not ( n21718 , n21681 );
and ( n341625 , n341623 , n21718 );
nor ( n21720 , n21716 , n341625 );
not ( n21721 , n21720 );
buf ( n21722 , n341211 );
not ( n21723 , n21722 );
buf ( n341630 , n21365 );
not ( n21725 , n341630 );
or ( n341632 , n21723 , n21725 );
buf ( n341633 , n341368 );
buf ( n341634 , n21366 );
buf ( n341635 , n21317 );
nand ( n21730 , n341634 , n341635 );
buf ( n341637 , n21730 );
buf ( n341638 , n341637 );
nand ( n341639 , n341633 , n341638 );
buf ( n341640 , n341639 );
buf ( n341641 , n341640 );
nand ( n21736 , n341632 , n341641 );
buf ( n21737 , n21736 );
not ( n341644 , n21737 );
nand ( n21739 , n21721 , n341644 );
nand ( n341646 , n341604 , n21739 );
nor ( n341647 , n21629 , n341646 );
buf ( n341648 , n341647 );
not ( n21743 , n341648 );
or ( n21744 , n21566 , n21743 );
buf ( n341651 , n21720 );
buf ( n341652 , n21737 );
nand ( n341653 , n341651 , n341652 );
buf ( n341654 , n341653 );
buf ( n341655 , n341654 );
buf ( n341656 , n21640 );
buf ( n341657 , n341598 );
nand ( n21752 , n341656 , n341657 );
buf ( n341659 , n21752 );
buf ( n341660 , n341659 );
nand ( n21755 , n341655 , n341660 );
buf ( n341662 , n21755 );
buf ( n341663 , n341662 );
buf ( n341664 , n341604 );
nand ( n341665 , n341663 , n341664 );
buf ( n341666 , n341665 );
nor ( n21761 , n21629 , n341666 );
buf ( n341668 , n21761 );
not ( n341669 , n21619 );
not ( n21764 , n21628 );
nor ( n21765 , n341669 , n21764 );
buf ( n341672 , n21765 );
nor ( n341673 , n341668 , n341672 );
buf ( n341674 , n341673 );
buf ( n341675 , n341674 );
nand ( n21770 , n21744 , n341675 );
buf ( n341677 , n21770 );
not ( n341678 , n341677 );
or ( n341679 , n18077 , n341678 );
nor ( n21774 , n17393 , n337738 );
not ( n21775 , n21774 );
not ( n21776 , n18075 );
or ( n341683 , n21775 , n21776 );
not ( n341684 , n18070 );
buf ( n341685 , n18074 );
not ( n21780 , n341685 );
buf ( n341687 , n21780 );
nand ( n341688 , n341684 , n341687 );
nand ( n341689 , n341683 , n341688 );
buf ( n341690 , n341689 );
not ( n21785 , n341690 );
buf ( n341692 , n21785 );
nand ( n341693 , n341679 , n341692 );
buf ( n341694 , n341693 );
buf ( n21789 , n341694 );
buf ( n341696 , n21789 );
buf ( n341697 , n341696 );
not ( n341698 , n341697 );
xor ( n341699 , n335932 , n336204 );
buf ( n341700 , n341699 );
buf ( n341701 , n341700 );
buf ( n341702 , n335924 );
and ( n341703 , n341701 , n341702 );
not ( n21798 , n341701 );
buf ( n341705 , n335921 );
and ( n21800 , n21798 , n341705 );
nor ( n341707 , n341703 , n21800 );
buf ( n341708 , n341707 );
buf ( n341709 , n341708 );
buf ( n341710 , n335556 );
buf ( n341711 , n335457 );
xor ( n341712 , n341710 , n341711 );
buf ( n341713 , n335653 );
xnor ( n341714 , n341712 , n341713 );
buf ( n341715 , n341714 );
buf ( n341716 , n341715 );
xor ( n341717 , n15515 , n335408 );
xor ( n21812 , n341717 , n335445 );
buf ( n341719 , n21812 );
not ( n341720 , n341719 );
buf ( n341721 , n341720 );
buf ( n341722 , n341721 );
not ( n341723 , n341722 );
not ( n21818 , n15164 );
not ( n341725 , n337781 );
or ( n341726 , n21818 , n341725 );
not ( n341727 , n335936 );
not ( n21822 , n335941 );
or ( n341729 , n341727 , n21822 );
nand ( n341730 , n341729 , n15115 );
nand ( n21825 , n341726 , n341730 );
not ( n341732 , n21825 );
buf ( n21827 , n341732 );
nand ( n21828 , n341723 , n21827 );
buf ( n21829 , n21828 );
buf ( n341736 , n21829 );
xor ( n21831 , n337860 , n337873 );
and ( n21832 , n21831 , n337887 );
and ( n21833 , n337860 , n337873 );
or ( n21834 , n21832 , n21833 );
buf ( n341741 , n21834 );
buf ( n341742 , n341741 );
and ( n21837 , n341736 , n341742 );
and ( n341744 , n341721 , n21825 );
buf ( n341745 , n341744 );
nor ( n21840 , n21837 , n341745 );
buf ( n21841 , n21840 );
not ( n341748 , n16086 );
not ( n341749 , n335964 );
or ( n21844 , n341748 , n341749 );
xor ( n341751 , n15764 , n15784 );
xnor ( n21846 , n341751 , n15772 );
nand ( n21847 , n21846 , n335945 );
nand ( n341754 , n21844 , n21847 );
not ( n21849 , n16099 );
and ( n341756 , n341754 , n21849 );
not ( n21851 , n341754 );
not ( n21852 , n21849 );
and ( n341759 , n21851 , n21852 );
nor ( n341760 , n341756 , n341759 );
xor ( n21855 , n21841 , n341760 );
not ( n341762 , n591 );
not ( n341763 , n336177 );
or ( n21858 , n341762 , n341763 );
or ( n341765 , n337907 , n338457 );
nand ( n341766 , n21858 , n341765 );
buf ( n341767 , n341766 );
buf ( n341768 , n15275 );
not ( n341769 , n341768 );
buf ( n341770 , n16094 );
not ( n21865 , n341770 );
or ( n341772 , n341769 , n21865 );
buf ( n21867 , n337799 );
buf ( n341774 , n335114 );
nand ( n21869 , n21867 , n341774 );
buf ( n341776 , n21869 );
buf ( n341777 , n341776 );
nand ( n21872 , n341772 , n341777 );
buf ( n341779 , n21872 );
buf ( n341780 , n341779 );
or ( n341781 , n341767 , n341780 );
buf ( n341782 , n341781 );
buf ( n341783 , n341782 );
buf ( n21878 , n336152 );
buf ( n21879 , n336014 );
xor ( n21880 , n21878 , n21879 );
buf ( n341787 , n336042 );
xor ( n341788 , n21880 , n341787 );
buf ( n341789 , n341788 );
buf ( n341790 , n341789 );
and ( n341791 , n341783 , n341790 );
buf ( n341792 , n341766 );
buf ( n341793 , n341779 );
and ( n341794 , n341792 , n341793 );
buf ( n341795 , n341794 );
buf ( n341796 , n341795 );
nor ( n341797 , n341791 , n341796 );
buf ( n341798 , n341797 );
and ( n21893 , n21855 , n341798 );
and ( n21894 , n21841 , n341760 );
or ( n341801 , n21893 , n21894 );
buf ( n21896 , n341801 );
xor ( n21897 , n341716 , n21896 );
buf ( n341804 , n335971 );
buf ( n341805 , n336198 );
xor ( n341806 , n341804 , n341805 );
buf ( n341807 , n16118 );
xor ( n21902 , n341806 , n341807 );
buf ( n341809 , n21902 );
buf ( n341810 , n341809 );
and ( n341811 , n21897 , n341810 );
and ( n21906 , n341716 , n21896 );
or ( n341813 , n341811 , n21906 );
buf ( n341814 , n341813 );
buf ( n341815 , n341814 );
nand ( n21910 , n341709 , n341815 );
buf ( n341817 , n21910 );
buf ( n341818 , n341817 );
xor ( n21913 , n336157 , n336185 );
xor ( n341820 , n21913 , n336194 );
buf ( n341821 , n341820 );
buf ( n341822 , n341821 );
not ( n341823 , n341822 );
buf ( n341824 , n341823 );
buf ( n341825 , n341824 );
not ( n21920 , n341825 );
xor ( n341827 , n21841 , n341760 );
xor ( n341828 , n341827 , n341798 );
buf ( n341829 , n341828 );
not ( n341830 , n341829 );
or ( n341831 , n21920 , n341830 );
xor ( n21926 , n337767 , n17931 );
and ( n21927 , n21926 , n337806 );
and ( n21928 , n337767 , n17931 );
or ( n341835 , n21927 , n21928 );
not ( n341836 , n341835 );
not ( n21931 , n341741 );
not ( n21932 , n21931 );
buf ( n341839 , n341721 );
not ( n21934 , n341839 );
buf ( n341841 , n341732 );
not ( n341842 , n341841 );
or ( n341843 , n21934 , n341842 );
nand ( n21938 , n21825 , n21812 );
buf ( n341845 , n21938 );
nand ( n21940 , n341843 , n341845 );
buf ( n341847 , n21940 );
not ( n21942 , n341847 );
not ( n21943 , n21942 );
or ( n21944 , n21932 , n21943 );
nand ( n341851 , n341741 , n341847 );
nand ( n341852 , n21944 , n341851 );
not ( n21947 , n341852 );
not ( n21948 , n21947 );
or ( n21949 , n341836 , n21948 );
not ( n341856 , n341835 );
not ( n341857 , n341856 );
not ( n21952 , n341852 );
or ( n21953 , n341857 , n21952 );
buf ( n341860 , n337917 );
not ( n341861 , n341860 );
buf ( n341862 , n341861 );
not ( n21957 , n341862 );
not ( n21958 , n17993 );
or ( n21959 , n21957 , n21958 );
buf ( n341866 , n341862 );
buf ( n341867 , n17993 );
or ( n21962 , n341866 , n341867 );
buf ( n341869 , n337889 );
nand ( n21964 , n21962 , n341869 );
buf ( n341871 , n21964 );
nand ( n21966 , n21959 , n341871 );
nand ( n21967 , n21953 , n21966 );
nand ( n21968 , n21949 , n21967 );
buf ( n341875 , n21968 );
nand ( n21970 , n341831 , n341875 );
buf ( n341877 , n21970 );
buf ( n21972 , n341877 );
not ( n341879 , n341828 );
buf ( n341880 , n341879 );
buf ( n341881 , n341821 );
nand ( n341882 , n341880 , n341881 );
buf ( n341883 , n341882 );
buf ( n341884 , n341883 );
nand ( n341885 , n21972 , n341884 );
buf ( n341886 , n341885 );
buf ( n341887 , n341886 );
not ( n21982 , n341887 );
xor ( n341889 , n341716 , n21896 );
xor ( n341890 , n341889 , n341810 );
buf ( n341891 , n341890 );
buf ( n341892 , n341891 );
nand ( n341893 , n21982 , n341892 );
buf ( n341894 , n341893 );
buf ( n341895 , n341894 );
and ( n21990 , n341818 , n341895 );
buf ( n341897 , n21990 );
buf ( n341898 , n341897 );
not ( n341899 , n341898 );
buf ( n341900 , n341899 );
buf ( n341901 , n341900 );
not ( n21996 , n337920 );
not ( n341903 , n17971 );
or ( n341904 , n21996 , n341903 );
buf ( n21999 , n17988 );
nand ( n341906 , n341904 , n21999 );
buf ( n341907 , n341906 );
or ( n22002 , n17971 , n337920 );
buf ( n341909 , n22002 );
nand ( n22004 , n341907 , n341909 );
buf ( n341911 , n22004 );
not ( n341912 , n341911 );
buf ( n341913 , n337761 );
not ( n341914 , n341913 );
buf ( n341915 , n17947 );
buf ( n341916 , n341915 );
not ( n341917 , n341916 );
or ( n341918 , n341914 , n341917 );
xor ( n22011 , n337767 , n17931 );
xnor ( n341920 , n22011 , n337806 );
not ( n22013 , n341920 );
not ( n22014 , n337761 );
not ( n22015 , n22014 );
or ( n22016 , n22013 , n22015 );
nand ( n22017 , n22016 , n337830 );
buf ( n341926 , n22017 );
nand ( n341927 , n341918 , n341926 );
buf ( n341928 , n341927 );
buf ( n341929 , n341928 );
buf ( n341930 , n341779 );
buf ( n341931 , n341789 );
xor ( n22024 , n341930 , n341931 );
buf ( n341933 , n341766 );
xor ( n341934 , n22024 , n341933 );
buf ( n341935 , n341934 );
buf ( n341936 , n341935 );
xor ( n341937 , n341929 , n341936 );
buf ( n341938 , n341937 );
not ( n341939 , n21931 );
not ( n22031 , n21942 );
or ( n341941 , n341939 , n22031 );
nand ( n22033 , n341941 , n341851 );
xor ( n22034 , n341835 , n22033 );
xnor ( n341944 , n22034 , n21966 );
xor ( n22036 , n341938 , n341944 );
not ( n341946 , n22036 );
nand ( n341947 , n341912 , n341946 );
not ( n22037 , n341879 );
and ( n341949 , n341821 , n21968 );
not ( n341950 , n341821 );
not ( n341951 , n21968 );
and ( n341952 , n341950 , n341951 );
nor ( n341953 , n341949 , n341952 );
not ( n22040 , n341953 );
or ( n341955 , n22037 , n22040 );
not ( n341956 , n341953 );
not ( n341957 , n341879 );
nand ( n22044 , n341956 , n341957 );
nand ( n341959 , n341955 , n22044 );
buf ( n341960 , n341959 );
buf ( n341961 , n341935 );
buf ( n341962 , n341928 );
or ( n341963 , n341961 , n341962 );
buf ( n341964 , n341963 );
and ( n341965 , n341964 , n341944 );
and ( n341966 , n341929 , n341936 );
buf ( n341967 , n341966 );
nor ( n22054 , n341965 , n341967 );
buf ( n341969 , n22054 );
nand ( n22056 , n341960 , n341969 );
buf ( n341971 , n22056 );
nand ( n341972 , n341947 , n341971 );
buf ( n341973 , n341972 );
nor ( n341974 , n341901 , n341973 );
buf ( n341975 , n341974 );
buf ( n341976 , n341975 );
not ( n341977 , n341976 );
or ( n341978 , n341698 , n341977 );
not ( n341979 , n341971 );
nand ( n341980 , n22036 , n341911 );
not ( n341981 , n341980 );
not ( n22063 , n341981 );
or ( n341983 , n341979 , n22063 );
or ( n341984 , n341959 , n22054 );
nand ( n341985 , n341983 , n341984 );
buf ( n341986 , n341985 );
not ( n341987 , n341986 );
buf ( n341988 , n341897 );
not ( n22070 , n341988 );
or ( n341990 , n341987 , n22070 );
not ( n341991 , n341817 );
not ( n22073 , n341886 );
nor ( n341993 , n22073 , n341891 );
not ( n22075 , n341993 );
or ( n341995 , n341991 , n22075 );
or ( n22077 , n341708 , n341814 );
nand ( n22078 , n341995 , n22077 );
not ( n341998 , n22078 );
buf ( n341999 , n341998 );
nand ( n22081 , n341990 , n341999 );
buf ( n342001 , n22081 );
buf ( n342002 , n342001 );
not ( n342003 , n342002 );
buf ( n342004 , n342003 );
buf ( n342005 , n342004 );
nand ( n342006 , n341978 , n342005 );
buf ( n342007 , n342006 );
buf ( n342008 , n342007 );
buf ( n342009 , n342008 );
buf ( n342010 , n342009 );
buf ( n342011 , n342010 );
buf ( n342012 , n342011 );
buf ( n342013 , n342012 );
not ( n342014 , n342013 );
not ( n342015 , n342014 );
or ( n22097 , n336229 , n342015 );
nand ( n342017 , n342013 , n336227 );
nand ( n342018 , n22097 , n342017 );
buf ( n342019 , n342018 );
buf ( n342020 , n342019 );
xor ( n342021 , n334637 , n334638 );
xor ( n342022 , n342021 , n342020 );
buf ( n342023 , n342022 );
xor ( n342024 , n334637 , n334638 );
and ( n342025 , n342024 , n342020 );
and ( n22107 , n334637 , n334638 );
or ( n22108 , n342025 , n22107 );
buf ( n22109 , n22108 );
buf ( n342029 , n332653 );
buf ( n342030 , n332625 );
xor ( n342031 , n335801 , n335829 );
and ( n22112 , n342031 , n335870 );
and ( n342033 , n335801 , n335829 );
or ( n342034 , n22112 , n342033 );
buf ( n342035 , n342034 );
buf ( n342036 , n342035 );
buf ( n342037 , n334862 );
not ( n342038 , n342037 );
buf ( n342039 , n335033 );
not ( n22119 , n342039 );
or ( n22120 , n342038 , n22119 );
buf ( n342042 , n335033 );
buf ( n342043 , n334862 );
or ( n22123 , n342042 , n342043 );
buf ( n342045 , n335086 );
nand ( n22125 , n22123 , n342045 );
buf ( n342047 , n22125 );
buf ( n342048 , n342047 );
nand ( n22128 , n22120 , n342048 );
buf ( n342050 , n22128 );
buf ( n342051 , n342050 );
and ( n342052 , n342036 , n342051 );
not ( n22132 , n342036 );
buf ( n342054 , n342050 );
not ( n342055 , n342054 );
buf ( n342056 , n342055 );
buf ( n342057 , n342056 );
and ( n342058 , n22132 , n342057 );
nor ( n342059 , n342052 , n342058 );
buf ( n342060 , n342059 );
not ( n342061 , n342060 );
xor ( n342062 , n334689 , n334734 );
and ( n342063 , n342062 , n334860 );
and ( n22143 , n334689 , n334734 );
or ( n342065 , n342063 , n22143 );
buf ( n342066 , n342065 );
buf ( n342067 , n342066 );
not ( n342068 , n15275 );
buf ( n342069 , n588 );
not ( n22149 , n342069 );
not ( n22150 , n14199 );
buf ( n342072 , n22150 );
not ( n342073 , n342072 );
or ( n342074 , n22149 , n342073 );
buf ( n342075 , n14199 );
buf ( n342076 , n334972 );
nand ( n342077 , n342075 , n342076 );
buf ( n342078 , n342077 );
buf ( n342079 , n342078 );
nand ( n342080 , n342074 , n342079 );
buf ( n342081 , n342080 );
not ( n342082 , n342081 );
or ( n22162 , n342068 , n342082 );
buf ( n342084 , n335818 );
buf ( n342085 , n335114 );
nand ( n342086 , n342084 , n342085 );
buf ( n342087 , n342086 );
nand ( n22167 , n22162 , n342087 );
buf ( n342089 , n22167 );
xor ( n22169 , n342067 , n342089 );
buf ( n342091 , n335181 );
not ( n342092 , n342091 );
buf ( n342093 , n16002 );
not ( n342094 , n342093 );
or ( n22174 , n342092 , n342094 );
nand ( n342096 , n334043 , n334037 );
buf ( n342097 , n342096 );
and ( n22177 , n342097 , n335097 );
not ( n342099 , n342097 );
and ( n342100 , n342099 , n590 );
or ( n22180 , n22177 , n342100 );
buf ( n342102 , n22180 );
buf ( n342103 , n591 );
nand ( n342104 , n342102 , n342103 );
buf ( n342105 , n342104 );
buf ( n342106 , n342105 );
nand ( n22186 , n22174 , n342106 );
buf ( n342108 , n22186 );
buf ( n342109 , n342108 );
xor ( n22189 , n22169 , n342109 );
buf ( n342111 , n22189 );
not ( n342112 , n342111 );
or ( n342113 , n342061 , n342112 );
not ( n22193 , n342060 );
not ( n342115 , n342111 );
nand ( n342116 , n22193 , n342115 );
nand ( n22196 , n342113 , n342116 );
not ( n342118 , n335872 );
buf ( n342119 , n15925 );
buf ( n22199 , n342119 );
buf ( n342121 , n22199 );
not ( n22201 , n342121 );
or ( n22202 , n342118 , n22201 );
buf ( n342124 , n342121 );
buf ( n342125 , n335872 );
or ( n22205 , n342124 , n342125 );
buf ( n342127 , n16048 );
nand ( n22207 , n22205 , n342127 );
buf ( n342129 , n22207 );
nand ( n342130 , n22202 , n342129 );
xor ( n342131 , n335047 , n335072 );
and ( n22211 , n342131 , n335084 );
and ( n342133 , n335047 , n335072 );
or ( n342134 , n22211 , n342133 );
buf ( n342135 , n342134 );
not ( n342136 , n342135 );
not ( n342137 , n342136 );
buf ( n342138 , n334643 );
not ( n22218 , n342138 );
buf ( n342140 , n580 );
not ( n342141 , n342140 );
buf ( n342142 , n334715 );
not ( n22222 , n342142 );
or ( n22223 , n342141 , n22222 );
buf ( n342145 , n334709 );
buf ( n342146 , n334650 );
nand ( n342147 , n342145 , n342146 );
buf ( n342148 , n342147 );
buf ( n342149 , n342148 );
nand ( n22229 , n22223 , n342149 );
buf ( n342151 , n22229 );
buf ( n342152 , n342151 );
not ( n342153 , n342152 );
or ( n342154 , n22218 , n342153 );
buf ( n342155 , n334654 );
buf ( n342156 , n14822 );
nand ( n342157 , n342155 , n342156 );
buf ( n342158 , n342157 );
buf ( n342159 , n342158 );
nand ( n22239 , n342154 , n342159 );
buf ( n342161 , n22239 );
buf ( n342162 , n334727 );
not ( n22242 , n342162 );
buf ( n342164 , n14844 );
not ( n342165 , n342164 );
or ( n22245 , n22242 , n342165 );
buf ( n342167 , n582 );
not ( n342168 , n342167 );
buf ( n342169 , n334873 );
not ( n342170 , n342169 );
or ( n342171 , n342168 , n342170 );
nand ( n342172 , n15012 , n334702 );
buf ( n342173 , n342172 );
nand ( n342174 , n342171 , n342173 );
buf ( n342175 , n342174 );
buf ( n342176 , n342175 );
buf ( n342177 , n334694 );
nand ( n22257 , n342176 , n342177 );
buf ( n342179 , n22257 );
buf ( n342180 , n342179 );
nand ( n342181 , n22245 , n342180 );
buf ( n342182 , n342181 );
xor ( n22262 , n342161 , n342182 );
xor ( n22263 , n334743 , n334793 );
and ( n342185 , n22263 , n334857 );
and ( n342186 , n334743 , n334793 );
or ( n22266 , n342185 , n342186 );
buf ( n342188 , n22266 );
xor ( n342189 , n22262 , n342188 );
not ( n22269 , n342189 );
or ( n342191 , n342137 , n22269 );
not ( n342192 , n342189 );
nand ( n342193 , n342192 , n342135 );
nand ( n22273 , n342191 , n342193 );
and ( n342195 , n334772 , n334774 );
buf ( n342196 , n342195 );
buf ( n342197 , n342196 );
buf ( n342198 , n14891 );
not ( n342199 , n342198 );
buf ( n342200 , n576 );
not ( n22280 , n342200 );
buf ( n342202 , n335514 );
not ( n342203 , n342202 );
or ( n22283 , n22280 , n342203 );
buf ( n342205 , n332672 );
buf ( n342206 , n14958 );
nand ( n342207 , n342205 , n342206 );
buf ( n342208 , n342207 );
buf ( n342209 , n342208 );
nand ( n342210 , n22283 , n342209 );
buf ( n342211 , n342210 );
buf ( n22291 , n342211 );
not ( n22292 , n22291 );
or ( n22293 , n342199 , n22292 );
buf ( n22294 , n334768 );
buf ( n22295 , n334786 );
nand ( n22296 , n22294 , n22295 );
buf ( n22297 , n22296 );
buf ( n22298 , n22297 );
nand ( n22299 , n22293 , n22298 );
buf ( n22300 , n22299 );
buf ( n342222 , n22300 );
xor ( n342223 , n342197 , n342222 );
buf ( n342224 , n14949 );
not ( n342225 , n342224 );
buf ( n342226 , n334847 );
not ( n22306 , n342226 );
or ( n342228 , n342225 , n22306 );
buf ( n342229 , n578 );
not ( n22309 , n342229 );
buf ( n342231 , n334564 );
not ( n22311 , n342231 );
or ( n342233 , n22309 , n22311 );
buf ( n22313 , n334561 );
buf ( n342235 , n334748 );
nand ( n22315 , n22313 , n342235 );
buf ( n342237 , n22315 );
buf ( n342238 , n342237 );
nand ( n22318 , n342233 , n342238 );
buf ( n342240 , n22318 );
buf ( n342241 , n342240 );
buf ( n342242 , n335432 );
nand ( n22322 , n342241 , n342242 );
buf ( n342244 , n22322 );
buf ( n342245 , n342244 );
nand ( n22325 , n342228 , n342245 );
buf ( n22326 , n22325 );
buf ( n342248 , n22326 );
xor ( n22328 , n342223 , n342248 );
buf ( n342250 , n22328 );
not ( n342251 , n334978 );
buf ( n342252 , n586 );
not ( n22332 , n342252 );
buf ( n342254 , n335163 );
not ( n342255 , n342254 );
or ( n342256 , n22332 , n342255 );
buf ( n342257 , n15300 );
buf ( n342258 , n334982 );
nand ( n22338 , n342257 , n342258 );
buf ( n342260 , n22338 );
buf ( n342261 , n342260 );
nand ( n22341 , n342256 , n342261 );
buf ( n342263 , n22341 );
not ( n22343 , n342263 );
or ( n342265 , n342251 , n22343 );
nand ( n342266 , n15221 , n15164 );
nand ( n22346 , n342265 , n342266 );
xor ( n22347 , n342250 , n22346 );
not ( n22348 , n334868 );
not ( n342270 , n334879 );
not ( n342271 , n335121 );
or ( n22351 , n342270 , n342271 );
buf ( n342273 , n15264 );
buf ( n342274 , n584 );
nand ( n342275 , n342273 , n342274 );
buf ( n342276 , n342275 );
nand ( n22356 , n22351 , n342276 );
not ( n22357 , n22356 );
or ( n22358 , n22348 , n22357 );
nand ( n342280 , n334917 , n335061 );
nand ( n22360 , n22358 , n342280 );
xor ( n22361 , n22347 , n22360 );
not ( n22362 , n22361 );
and ( n22363 , n22273 , n22362 );
not ( n342285 , n22273 );
and ( n342286 , n342285 , n22361 );
nor ( n22366 , n22363 , n342286 );
not ( n22367 , n22366 );
and ( n22368 , n342130 , n22367 );
not ( n22369 , n342130 );
and ( n342291 , n22369 , n22366 );
nor ( n342292 , n22368 , n342291 );
xor ( n22372 , n22196 , n342292 );
buf ( n342294 , n22372 );
buf ( n342295 , n15908 );
buf ( n342296 , n335092 );
or ( n22376 , n342295 , n342296 );
buf ( n342298 , n22376 );
and ( n342299 , n335914 , n342298 );
and ( n22379 , n335092 , n15908 );
nor ( n342301 , n342299 , n22379 );
buf ( n342302 , n342301 );
nand ( n342303 , n342294 , n342302 );
buf ( n342304 , n342303 );
buf ( n22384 , n342304 );
buf ( n342306 , n22372 );
not ( n22386 , n342306 );
buf ( n342308 , n22386 );
buf ( n342309 , n342308 );
buf ( n22389 , n342301 );
not ( n342311 , n22389 );
buf ( n342312 , n342311 );
buf ( n342313 , n342312 );
nand ( n342314 , n342309 , n342313 );
buf ( n342315 , n342314 );
nand ( n342316 , n22384 , n342315 );
and ( n342317 , n336219 , n342316 );
not ( n342318 , n342317 );
not ( n22398 , n342010 );
not ( n342320 , n22398 );
not ( n22400 , n342320 );
or ( n22401 , n342318 , n22400 );
not ( n22402 , n336224 );
nor ( n22403 , n22402 , n342316 );
and ( n22404 , n22398 , n22403 );
not ( n22405 , n336219 );
not ( n342327 , n22405 );
not ( n342328 , n22403 );
or ( n22408 , n342327 , n342328 );
nand ( n342330 , n22402 , n342316 );
nand ( n342331 , n22408 , n342330 );
nor ( n22411 , n22404 , n342331 );
nand ( n342333 , n22401 , n22411 );
not ( n342334 , n342333 );
buf ( n342335 , n342334 );
buf ( n342336 , n342335 );
not ( n342337 , n342336 );
buf ( n342338 , n342337 );
buf ( n342339 , n342338 );
xor ( n342340 , n342029 , n342030 );
xor ( n22420 , n342340 , n342339 );
buf ( n342342 , n22420 );
xor ( n22422 , n342029 , n342030 );
and ( n22423 , n22422 , n342339 );
and ( n342345 , n342029 , n342030 );
or ( n342346 , n22423 , n342345 );
buf ( n342347 , n342346 );
buf ( n342348 , n320925 );
buf ( n342349 , n321236 );
xor ( n22429 , n340605 , n340609 );
xor ( n342351 , n22429 , n340753 );
buf ( n342352 , n342351 );
buf ( n342353 , n342352 );
xor ( n22433 , n342348 , n342349 );
xor ( n342355 , n22433 , n342353 );
buf ( n342356 , n342355 );
xor ( n22436 , n342348 , n342349 );
and ( n342358 , n22436 , n342353 );
and ( n342359 , n342348 , n342349 );
or ( n22439 , n342358 , n342359 );
buf ( n342361 , n22439 );
buf ( n342362 , n320889 );
buf ( n22442 , n320596 );
nand ( n22443 , n20876 , n20719 );
not ( n342365 , n340757 );
xor ( n342366 , n22443 , n342365 );
buf ( n342367 , n342366 );
xor ( n342368 , n342362 , n22442 );
xor ( n342369 , n342368 , n342367 );
buf ( n342370 , n342369 );
xor ( n342371 , n342362 , n22442 );
and ( n22449 , n342371 , n342367 );
and ( n22450 , n342362 , n22442 );
or ( n22451 , n22449 , n22450 );
buf ( n342375 , n22451 );
buf ( n342376 , n321119 );
buf ( n342377 , n334017 );
buf ( n22455 , n340828 );
buf ( n22456 , n340441 );
nand ( n22457 , n22455 , n22456 );
buf ( n22458 , n22457 );
buf ( n342382 , n22458 );
buf ( n342383 , n20926 );
xnor ( n342384 , n342382 , n342383 );
buf ( n342385 , n342384 );
buf ( n342386 , n342385 );
xor ( n342387 , n342376 , n342377 );
xor ( n342388 , n342387 , n342386 );
buf ( n342389 , n342388 );
xor ( n342390 , n342376 , n342377 );
and ( n342391 , n342390 , n342386 );
and ( n342392 , n342376 , n342377 );
or ( n342393 , n342391 , n342392 );
buf ( n342394 , n342393 );
buf ( n342395 , n334012 );
buf ( n342396 , n321945 );
buf ( n22465 , n340892 );
not ( n342398 , n22465 );
buf ( n342399 , n342398 );
buf ( n342400 , n342399 );
not ( n22469 , n342400 );
buf ( n342402 , n340927 );
buf ( n342403 , n340915 );
buf ( n22472 , n342403 );
buf ( n342405 , n22472 );
buf ( n342406 , n342405 );
nand ( n22473 , n342402 , n342406 );
buf ( n342408 , n22473 );
buf ( n342409 , n342408 );
not ( n342410 , n342409 );
buf ( n22474 , n342410 );
buf ( n342412 , n22474 );
not ( n22476 , n342412 );
or ( n342414 , n22469 , n22476 );
buf ( n22478 , n342408 );
buf ( n22479 , n340892 );
nand ( n22480 , n22478 , n22479 );
buf ( n22481 , n22480 );
buf ( n22482 , n22481 );
nand ( n22483 , n342414 , n22482 );
buf ( n22484 , n22483 );
buf ( n342422 , n22484 );
xor ( n22486 , n342395 , n342396 );
xor ( n342424 , n22486 , n342422 );
buf ( n342425 , n342424 );
xor ( n342426 , n342395 , n342396 );
and ( n22490 , n342426 , n342422 );
and ( n342428 , n342395 , n342396 );
or ( n22492 , n22490 , n342428 );
buf ( n342430 , n22492 );
buf ( n342431 , n324325 );
buf ( n342432 , n342431 );
buf ( n342433 , n324372 );
nand ( n342434 , n341026 , n341013 );
buf ( n342435 , n340944 );
buf ( n342436 , n342435 );
buf ( n342437 , n342436 );
buf ( n342438 , n342437 );
not ( n342439 , n342438 );
buf ( n342440 , n342439 );
and ( n342441 , n342434 , n342440 );
not ( n342442 , n342434 );
and ( n342443 , n342442 , n342437 );
nor ( n22499 , n342441 , n342443 );
buf ( n342445 , n22499 );
buf ( n342446 , n342445 );
xor ( n342447 , n342432 , n342433 );
xor ( n22503 , n342447 , n342446 );
buf ( n342449 , n22503 );
xor ( n342450 , n342432 , n342433 );
and ( n22506 , n342450 , n342446 );
and ( n342452 , n342432 , n342433 );
or ( n342453 , n22506 , n342452 );
buf ( n342454 , n342453 );
buf ( n342455 , n7688 );
buf ( n342456 , n7672 );
buf ( n342457 , n341099 );
not ( n22513 , n342457 );
buf ( n22514 , n341079 );
buf ( n342460 , n22514 );
not ( n342461 , n342460 );
or ( n22517 , n22513 , n342461 );
buf ( n342463 , n341117 );
nand ( n342464 , n22517 , n342463 );
buf ( n342465 , n342464 );
buf ( n342466 , n341123 );
buf ( n342467 , n339048 );
nand ( n342468 , n342466 , n342467 );
buf ( n342469 , n342468 );
or ( n22525 , n342465 , n342469 );
buf ( n342471 , n342465 );
buf ( n342472 , n342469 );
nand ( n22528 , n342471 , n342472 );
buf ( n22529 , n22528 );
nand ( n342475 , n22525 , n22529 );
buf ( n342476 , n342475 );
xor ( n342477 , n342455 , n342456 );
xor ( n22533 , n342477 , n342476 );
buf ( n342479 , n22533 );
xor ( n22535 , n342455 , n342456 );
and ( n342481 , n22535 , n342476 );
and ( n342482 , n342455 , n342456 );
or ( n22538 , n342481 , n342482 );
buf ( n342484 , n22538 );
buf ( n22540 , n326366 );
buf ( n342486 , n326487 );
nand ( n342487 , n21721 , n341644 );
buf ( n342488 , n341654 );
buf ( n22544 , n342488 );
buf ( n22545 , n22544 );
nand ( n342491 , n342487 , n22545 );
not ( n22547 , n342491 );
not ( n22548 , n22547 );
buf ( n342494 , n341470 );
buf ( n342495 , n342494 );
buf ( n342496 , n342495 );
buf ( n342497 , n342496 );
not ( n22552 , n342497 );
buf ( n342499 , n22552 );
not ( n342500 , n342499 );
or ( n22555 , n22548 , n342500 );
nand ( n342502 , n342496 , n342491 );
nand ( n22556 , n22555 , n342502 );
buf ( n342504 , n22556 );
xor ( n342505 , n22540 , n342486 );
xor ( n22559 , n342505 , n342504 );
buf ( n342507 , n22559 );
xor ( n22560 , n22540 , n342486 );
and ( n342509 , n22560 , n342504 );
and ( n342510 , n22540 , n342486 );
or ( n342511 , n342509 , n342510 );
buf ( n342512 , n342511 );
buf ( n342513 , n5166 );
buf ( n342514 , n325355 );
nand ( n22567 , n342487 , n341470 );
buf ( n342516 , n22567 );
buf ( n342517 , n22545 );
nand ( n342518 , n342516 , n342517 );
buf ( n342519 , n342518 );
buf ( n342520 , n342519 );
buf ( n22573 , n341549 );
buf ( n22574 , n341601 );
nand ( n22575 , n22573 , n22574 );
buf ( n22576 , n22575 );
nand ( n342525 , n341659 , n22576 );
buf ( n342526 , n342525 );
xnor ( n342527 , n342520 , n342526 );
buf ( n342528 , n342527 );
buf ( n342529 , n342528 );
xor ( n22582 , n342513 , n342514 );
xor ( n342531 , n22582 , n342529 );
buf ( n342532 , n342531 );
xor ( n22585 , n342513 , n342514 );
and ( n342534 , n22585 , n342529 );
and ( n342535 , n342513 , n342514 );
or ( n22588 , n342534 , n342535 );
buf ( n342537 , n22588 );
buf ( n342538 , n7106 );
buf ( n342539 , n327272 );
buf ( n342540 , n22576 );
not ( n22593 , n342540 );
buf ( n342542 , n22593 );
or ( n22595 , n22567 , n342542 );
buf ( n342544 , n341666 );
not ( n342545 , n342544 );
buf ( n342546 , n342545 );
not ( n22599 , n342546 );
nand ( n22600 , n22595 , n22599 );
not ( n342549 , n22600 );
buf ( n342550 , n21619 );
not ( n22603 , n342550 );
not ( n22604 , n21764 );
not ( n22605 , n22604 );
and ( n342554 , n22603 , n22605 );
and ( n342555 , n22604 , n342550 );
nor ( n22608 , n342554 , n342555 );
buf ( n342557 , n22608 );
not ( n22610 , n342557 );
buf ( n342559 , n22610 );
and ( n342560 , n342549 , n342559 );
not ( n22613 , n342549 );
and ( n22614 , n22613 , n22608 );
nor ( n22615 , n342560 , n22614 );
buf ( n342564 , n22615 );
buf ( n22617 , n342564 );
buf ( n22618 , n22617 );
buf ( n22619 , n22618 );
buf ( n342568 , n22619 );
xor ( n22621 , n342538 , n342539 );
xor ( n342570 , n22621 , n342568 );
buf ( n342571 , n342570 );
xor ( n22624 , n342538 , n342539 );
and ( n342573 , n22624 , n342568 );
and ( n22626 , n342538 , n342539 );
or ( n22627 , n342573 , n22626 );
buf ( n342576 , n22627 );
buf ( n342577 , n326948 );
buf ( n342578 , n327265 );
buf ( n342579 , n337739 );
not ( n22632 , n21774 );
nand ( n22633 , n342579 , n22632 );
buf ( n342582 , n341677 );
not ( n22635 , n342582 );
buf ( n342584 , n22635 );
buf ( n22637 , n342584 );
and ( n342586 , n22633 , n22637 );
not ( n342587 , n22633 );
not ( n22640 , n22637 );
and ( n342589 , n342587 , n22640 );
nor ( n342590 , n342586 , n342589 );
buf ( n342591 , n342590 );
xor ( n342592 , n342577 , n342578 );
xor ( n342593 , n342592 , n342591 );
buf ( n342594 , n342593 );
xor ( n22647 , n342577 , n342578 );
and ( n22648 , n22647 , n342591 );
and ( n22649 , n342577 , n342578 );
or ( n22650 , n22648 , n22649 );
buf ( n342599 , n22650 );
buf ( n342600 , n327799 );
buf ( n342601 , n14148 );
and ( n22654 , n341688 , n18075 );
not ( n342603 , n22654 );
not ( n22656 , n342579 );
or ( n342605 , n342584 , n22656 );
nand ( n22658 , n342605 , n22632 );
buf ( n342607 , n22658 );
not ( n342608 , n342607 );
buf ( n342609 , n342608 );
not ( n22662 , n342609 );
or ( n342611 , n342603 , n22662 );
not ( n342612 , n22654 );
nand ( n22665 , n342612 , n22658 );
nand ( n342614 , n342611 , n22665 );
buf ( n22667 , n342614 );
buf ( n342616 , n22667 );
buf ( n342617 , n342616 );
buf ( n342618 , n342617 );
xor ( n342619 , n342600 , n342601 );
xor ( n22672 , n342619 , n342618 );
buf ( n342621 , n22672 );
xor ( n342622 , n342600 , n342601 );
and ( n22675 , n342622 , n342618 );
and ( n22676 , n342600 , n342601 );
or ( n342625 , n22675 , n22676 );
buf ( n342626 , n342625 );
buf ( n342627 , n331818 );
buf ( n342628 , n331731 );
buf ( n342629 , n341971 );
buf ( n342630 , n341984 );
nand ( n22683 , n342629 , n342630 );
buf ( n342632 , n22683 );
buf ( n342633 , n342632 );
not ( n22686 , n342633 );
buf ( n342635 , n22686 );
not ( n342636 , n342635 );
not ( n22689 , n341911 );
nand ( n342638 , n22689 , n341946 );
not ( n342639 , n342638 );
not ( n22692 , n341693 );
or ( n342641 , n342639 , n22692 );
buf ( n342642 , n341980 );
buf ( n22695 , n342642 );
buf ( n342644 , n22695 );
nand ( n342645 , n342641 , n342644 );
not ( n22698 , n342645 );
not ( n342647 , n22698 );
or ( n22700 , n342636 , n342647 );
buf ( n342649 , n342645 );
buf ( n342650 , n342632 );
nand ( n22703 , n342649 , n342650 );
buf ( n22704 , n22703 );
nand ( n342653 , n22700 , n22704 );
buf ( n342654 , n342653 );
not ( n22707 , n342654 );
not ( n342656 , n22707 );
not ( n342657 , n342656 );
not ( n22710 , n342657 );
buf ( n342659 , n22710 );
xor ( n342660 , n342627 , n342628 );
xor ( n342661 , n342660 , n342659 );
buf ( n342662 , n342661 );
xor ( n342663 , n342627 , n342628 );
and ( n342664 , n342663 , n342659 );
and ( n22717 , n342627 , n342628 );
or ( n342666 , n342664 , n22717 );
buf ( n342667 , n342666 );
buf ( n342668 , n332041 );
buf ( n342669 , n331971 );
not ( n22722 , n341972 );
not ( n342671 , n22722 );
not ( n342672 , n341693 );
or ( n342673 , n342671 , n342672 );
not ( n22726 , n341985 );
nand ( n342675 , n342673 , n22726 );
not ( n22728 , n342675 );
buf ( n342677 , n341993 );
not ( n22730 , n342677 );
buf ( n342679 , n22730 );
buf ( n342680 , n342679 );
buf ( n342681 , n341894 );
buf ( n342682 , n342681 );
buf ( n342683 , n342682 );
buf ( n342684 , n342683 );
nand ( n342685 , n342680 , n342684 );
buf ( n342686 , n342685 );
xor ( n342687 , n22728 , n342686 );
buf ( n342688 , n342687 );
buf ( n342689 , n342688 );
xor ( n22742 , n342668 , n342669 );
xor ( n22743 , n22742 , n342689 );
buf ( n342692 , n22743 );
xor ( n22745 , n342668 , n342669 );
and ( n22746 , n22745 , n342689 );
and ( n22747 , n342668 , n342669 );
or ( n22748 , n22746 , n22747 );
buf ( n342697 , n22748 );
buf ( n342698 , n332472 );
buf ( n342699 , n332348 );
not ( n342700 , n342683 );
not ( n342701 , n342675 );
or ( n22754 , n342700 , n342701 );
buf ( n342703 , n342679 );
nand ( n22756 , n22754 , n342703 );
buf ( n342705 , n341817 );
buf ( n342706 , n22077 );
nand ( n22759 , n342705 , n342706 );
buf ( n342708 , n22759 );
not ( n342709 , n342708 );
or ( n22762 , n22756 , n342709 );
buf ( n342711 , n342708 );
not ( n342712 , n342711 );
nand ( n22765 , n342712 , n22756 );
nand ( n342714 , n22762 , n22765 );
not ( n342715 , n342714 );
not ( n22768 , n342715 );
not ( n22769 , n22768 );
not ( n342718 , n22769 );
not ( n342719 , n342718 );
buf ( n22772 , n342719 );
buf ( n342721 , n22772 );
xor ( n22774 , n342698 , n342699 );
xor ( n342723 , n22774 , n342721 );
buf ( n342724 , n342723 );
xor ( n22777 , n342698 , n342699 );
and ( n342726 , n22777 , n342721 );
and ( n342727 , n342698 , n342699 );
or ( n22780 , n342726 , n342727 );
buf ( n342729 , n22780 );
buf ( n342730 , n332816 );
buf ( n342731 , n332781 );
xor ( n342732 , n342730 , n342731 );
buf ( n342733 , n342732 );
buf ( n342734 , n22109 );
buf ( n342735 , n342342 );
buf ( n342736 , n342023 );
buf ( n342737 , n342729 );
xor ( n22790 , n342736 , n342737 );
buf ( n342739 , n342697 );
buf ( n342740 , n342724 );
xor ( n342741 , n342739 , n342740 );
buf ( n342742 , n342692 );
buf ( n342743 , n342667 );
xor ( n22796 , n342742 , n342743 );
buf ( n342745 , n331348 );
buf ( n342746 , n331575 );
xor ( n342747 , n342745 , n342746 );
buf ( n22800 , n342644 );
buf ( n342749 , n342638 );
nand ( n22802 , n22800 , n342749 );
buf ( n342751 , n22802 );
not ( n342752 , n342751 );
not ( n22805 , n342752 );
not ( n342754 , n341696 );
not ( n22807 , n342754 );
or ( n342756 , n22805 , n22807 );
nand ( n22809 , n342751 , n341696 );
nand ( n22810 , n342756 , n22809 );
buf ( n342759 , n22810 );
buf ( n342760 , n342759 );
buf ( n342761 , n342760 );
and ( n342762 , n342747 , n342761 );
and ( n342763 , n342745 , n342746 );
or ( n22816 , n342762 , n342763 );
buf ( n342765 , n22816 );
buf ( n342766 , n342765 );
buf ( n342767 , n342662 );
xor ( n342768 , n342766 , n342767 );
xor ( n342769 , n342745 , n342746 );
xor ( n22822 , n342769 , n342761 );
buf ( n342771 , n22822 );
buf ( n342772 , n342771 );
not ( n342773 , n342772 );
buf ( n342774 , n342621 );
buf ( n342775 , n342599 );
nand ( n22828 , n342774 , n342775 );
buf ( n342777 , n22828 );
buf ( n342778 , n342777 );
buf ( n342779 , n342626 );
not ( n342780 , n342779 );
buf ( n342781 , n342780 );
buf ( n342782 , n342781 );
and ( n342783 , n342778 , n342782 );
buf ( n342784 , n342783 );
buf ( n342785 , n342784 );
buf ( n342786 , n342599 );
not ( n342787 , n342786 );
buf ( n342788 , n342621 );
not ( n342789 , n342788 );
buf ( n342790 , n342789 );
buf ( n342791 , n342790 );
nand ( n342792 , n342787 , n342791 );
buf ( n342793 , n342792 );
buf ( n342794 , n342793 );
buf ( n342795 , n342594 );
buf ( n342796 , n342576 );
nor ( n342797 , n342795 , n342796 );
buf ( n342798 , n342797 );
buf ( n342799 , n342798 );
buf ( n342800 , n342571 );
buf ( n342801 , n342537 );
nand ( n22854 , n342800 , n342801 );
buf ( n342803 , n22854 );
buf ( n342804 , n342803 );
or ( n342805 , n342799 , n342804 );
buf ( n22858 , n342594 );
buf ( n342807 , n342576 );
nand ( n22860 , n22858 , n342807 );
buf ( n342809 , n22860 );
buf ( n342810 , n342809 );
nand ( n22863 , n342805 , n342810 );
buf ( n342812 , n22863 );
buf ( n342813 , n342812 );
nand ( n342814 , n342794 , n342813 );
buf ( n342815 , n342814 );
buf ( n342816 , n342815 );
buf ( n22869 , n342532 );
buf ( n342818 , n342512 );
xor ( n22871 , n22869 , n342818 );
not ( n342820 , n6646 );
not ( n342821 , n6709 );
or ( n22874 , n342820 , n342821 );
nand ( n342823 , n22874 , n326566 );
buf ( n342824 , n342823 );
buf ( n342825 , n327287 );
xor ( n342826 , n342824 , n342825 );
buf ( n22879 , n341129 );
buf ( n342828 , n22879 );
buf ( n342829 , n342828 );
buf ( n342830 , n341413 );
buf ( n342831 , n341464 );
and ( n22884 , n342830 , n342831 );
buf ( n22885 , n22884 );
buf ( n22886 , n341450 );
not ( n342835 , n22886 );
buf ( n342836 , n342835 );
nand ( n342837 , n342829 , n22885 , n342836 );
not ( n22890 , n342829 );
buf ( n22891 , n341440 );
not ( n342840 , n22885 );
nand ( n22893 , n22890 , n22891 , n342840 );
not ( n342842 , n342836 );
nor ( n22895 , n342842 , n22891 );
nand ( n22896 , n22885 , n22895 );
or ( n342845 , n22885 , n342836 );
nand ( n342846 , n342837 , n22893 , n22896 , n342845 );
not ( n22899 , n342846 );
not ( n342848 , n22899 );
buf ( n342849 , n342848 );
and ( n22902 , n342826 , n342849 );
and ( n342851 , n342824 , n342825 );
or ( n342852 , n22902 , n342851 );
buf ( n342853 , n342852 );
buf ( n342854 , n342853 );
buf ( n342855 , n342507 );
xor ( n342856 , n342854 , n342855 );
xor ( n22909 , n342824 , n342825 );
xor ( n342858 , n22909 , n342849 );
buf ( n342859 , n342858 );
buf ( n342860 , n342859 );
buf ( n342861 , n327338 );
xor ( n342862 , n342861 , n327584 );
buf ( n342863 , n342829 );
buf ( n342864 , n22891 );
buf ( n342865 , n342836 );
nand ( n22916 , n342864 , n342865 );
buf ( n342867 , n22916 );
buf ( n342868 , n342867 );
and ( n22919 , n342863 , n342868 );
not ( n342870 , n342863 );
buf ( n342871 , n342867 );
not ( n342872 , n342871 );
buf ( n342873 , n342872 );
buf ( n342874 , n342873 );
and ( n342875 , n342870 , n342874 );
nor ( n342876 , n22919 , n342875 );
buf ( n342877 , n342876 );
not ( n342878 , n342877 );
not ( n342879 , n342878 );
buf ( n22930 , n342879 );
buf ( n342881 , n22930 );
and ( n342882 , n342862 , n342881 );
and ( n342883 , n342861 , n327584 );
or ( n22934 , n342882 , n342883 );
buf ( n342885 , n22934 );
xor ( n342886 , n342860 , n342885 );
buf ( n342887 , n342484 );
buf ( n342888 , n7603 );
nand ( n342889 , n327482 , n342888 );
buf ( n342890 , n341117 );
buf ( n342891 , n341099 );
nand ( n22941 , n342890 , n342891 );
buf ( n342893 , n22941 );
buf ( n22943 , n342893 );
not ( n22944 , n22943 );
buf ( n342896 , n22944 );
not ( n22946 , n342896 );
not ( n22947 , n22514 );
not ( n22948 , n22947 );
or ( n22949 , n22946 , n22948 );
buf ( n342901 , n22514 );
buf ( n342902 , n342893 );
nand ( n22952 , n342901 , n342902 );
buf ( n342904 , n22952 );
nand ( n22954 , n22949 , n342904 );
buf ( n22955 , n22954 );
not ( n22956 , n22955 );
buf ( n342908 , n22956 );
buf ( n342909 , n342908 );
not ( n22959 , n342909 );
nand ( n22960 , n327482 , n22959 );
not ( n22961 , n342909 );
nand ( n342913 , n342888 , n22961 );
nand ( n342914 , n342889 , n22960 , n342913 );
buf ( n342915 , n342914 );
buf ( n342916 , n342479 );
xor ( n22966 , n342915 , n342916 );
buf ( n342918 , n324050 );
buf ( n342919 , n323395 );
xor ( n22969 , n342918 , n342919 );
buf ( n342921 , n341078 );
buf ( n342922 , n339471 );
nand ( n342923 , n342921 , n342922 );
buf ( n342924 , n342923 );
buf ( n342925 , n342924 );
buf ( n342926 , n21178 );
buf ( n22976 , n342926 );
buf ( n342928 , n22976 );
buf ( n342929 , n342928 );
xnor ( n342930 , n342925 , n342929 );
buf ( n342931 , n342930 );
buf ( n342932 , n342931 );
buf ( n342933 , n342932 );
buf ( n342934 , n342933 );
buf ( n342935 , n342934 );
and ( n342936 , n22969 , n342935 );
and ( n342937 , n342918 , n342919 );
or ( n22985 , n342936 , n342937 );
buf ( n342939 , n22985 );
buf ( n342940 , n342939 );
buf ( n342941 , n323484 );
buf ( n342942 , n21152 );
buf ( n342943 , n341054 );
nor ( n342944 , n342942 , n342943 );
buf ( n342945 , n342944 );
buf ( n342946 , n342945 );
not ( n342947 , n342946 );
buf ( n22995 , n341063 );
nand ( n22996 , n342947 , n22995 );
buf ( n22997 , n22996 );
buf ( n342951 , n22997 );
not ( n22999 , n342951 );
buf ( n23000 , n22999 );
not ( n342954 , n23000 );
buf ( n342955 , n341029 );
not ( n23003 , n342955 );
buf ( n23004 , n23003 );
not ( n342958 , n23004 );
or ( n23006 , n342954 , n342958 );
buf ( n342960 , n22997 );
buf ( n23008 , n341029 );
nand ( n23009 , n342960 , n23008 );
buf ( n342963 , n23009 );
nand ( n342964 , n23006 , n342963 );
buf ( n342965 , n342964 );
buf ( n342966 , n342965 );
xor ( n342967 , n342941 , n342966 );
buf ( n342968 , n4436 );
and ( n342969 , n342967 , n342968 );
and ( n342970 , n342941 , n342966 );
or ( n342971 , n342969 , n342970 );
buf ( n342972 , n342971 );
buf ( n23013 , n342972 );
xor ( n342974 , n342918 , n342919 );
xor ( n23015 , n342974 , n342935 );
buf ( n342976 , n23015 );
buf ( n342977 , n342976 );
xor ( n23016 , n23013 , n342977 );
buf ( n342979 , n342454 );
xor ( n342980 , n342941 , n342966 );
xor ( n342981 , n342980 , n342968 );
buf ( n342982 , n342981 );
buf ( n342983 , n342982 );
xor ( n23019 , n342979 , n342983 );
buf ( n342985 , n324383 );
buf ( n342986 , n14153 );
xor ( n23022 , n342985 , n342986 );
buf ( n342988 , n340941 );
buf ( n342989 , n20081 );
nand ( n342990 , n342988 , n342989 );
buf ( n342991 , n342990 );
buf ( n342992 , n21040 );
and ( n342993 , n342991 , n342992 );
not ( n342994 , n342991 );
not ( n23027 , n340915 );
not ( n342996 , n340892 );
or ( n342997 , n23027 , n342996 );
nand ( n23030 , n342997 , n340927 );
not ( n342999 , n23030 );
and ( n23032 , n342994 , n342999 );
nor ( n343001 , n342993 , n23032 );
not ( n23034 , n343001 );
buf ( n343003 , n23034 );
buf ( n23036 , n343003 );
buf ( n23037 , n23036 );
buf ( n343006 , n23037 );
and ( n343007 , n23022 , n343006 );
and ( n343008 , n342985 , n342986 );
or ( n23041 , n343007 , n343008 );
buf ( n343010 , n23041 );
buf ( n343011 , n343010 );
buf ( n343012 , n342449 );
xor ( n343013 , n343011 , n343012 );
buf ( n343014 , n342430 );
not ( n343015 , n343014 );
xor ( n343016 , n342985 , n342986 );
xor ( n343017 , n343016 , n343006 );
buf ( n343018 , n343017 );
buf ( n343019 , n343018 );
not ( n343020 , n343019 );
or ( n343021 , n343015 , n343020 );
buf ( n343022 , n343018 );
buf ( n343023 , n342430 );
or ( n343024 , n343022 , n343023 );
buf ( n23057 , n322691 );
buf ( n23058 , n322744 );
xor ( n23059 , n23057 , n23058 );
buf ( n343028 , n340873 );
buf ( n343029 , n340861 );
nand ( n23062 , n343028 , n343029 );
buf ( n343031 , n23062 );
buf ( n343032 , n340831 );
not ( n343033 , n343032 );
buf ( n343034 , n343033 );
and ( n343035 , n343031 , n343034 );
not ( n343036 , n343031 );
buf ( n23069 , n340831 );
and ( n343038 , n343036 , n23069 );
nor ( n343039 , n343035 , n343038 );
buf ( n343040 , n343039 );
and ( n23073 , n23059 , n343040 );
and ( n343042 , n23057 , n23058 );
or ( n343043 , n23073 , n343042 );
buf ( n343044 , n343043 );
buf ( n343045 , n343044 );
xor ( n23078 , n322679 , n2787 );
nand ( n343047 , n340883 , n20470 );
buf ( n23080 , n20986 );
not ( n23081 , n23080 );
and ( n343050 , n343047 , n23081 );
not ( n343051 , n343047 );
and ( n23084 , n343051 , n23080 );
nor ( n343053 , n343050 , n23084 );
xor ( n343054 , n23078 , n343053 );
buf ( n343055 , n343054 );
xor ( n343056 , n343045 , n343055 );
buf ( n343057 , n342394 );
not ( n23090 , n343057 );
xor ( n343059 , n23057 , n23058 );
xor ( n23091 , n343059 , n343040 );
buf ( n343061 , n23091 );
buf ( n343062 , n343061 );
not ( n23094 , n343062 );
or ( n343064 , n23090 , n23094 );
buf ( n343065 , n342389 );
buf ( n343066 , n320797 );
buf ( n343067 , n14158 );
xor ( n23098 , n343066 , n343067 );
not ( n23099 , n340790 );
not ( n343070 , n23099 );
not ( n343071 , n340800 );
or ( n23102 , n343070 , n343071 );
nand ( n343073 , n23102 , n340813 );
xor ( n23104 , n340766 , n343073 );
buf ( n343075 , n23104 );
and ( n23106 , n23098 , n343075 );
and ( n23107 , n343066 , n343067 );
or ( n23108 , n23106 , n23107 );
buf ( n343079 , n23108 );
buf ( n343080 , n343079 );
nor ( n23111 , n343065 , n343080 );
buf ( n343082 , n23111 );
buf ( n343083 , n343082 );
buf ( n343084 , n342361 );
buf ( n343085 , n1531 );
buf ( n343086 , n343085 );
buf ( n343087 , n321317 );
buf ( n343088 , n321351 );
xor ( n343089 , n343087 , n343088 );
buf ( n343090 , n321432 );
buf ( n343091 , n321340 );
xor ( n23122 , n343090 , n343091 );
buf ( n343093 , n321467 );
buf ( n343094 , n1771 );
and ( n23125 , n343093 , n343094 );
buf ( n343096 , n23125 );
buf ( n343097 , n343096 );
and ( n343098 , n23122 , n343097 );
and ( n23129 , n343090 , n343091 );
or ( n343100 , n343098 , n23129 );
buf ( n343101 , n343100 );
buf ( n343102 , n343101 );
and ( n23133 , n343089 , n343102 );
and ( n23134 , n343087 , n343088 );
or ( n343105 , n23133 , n23134 );
buf ( n343106 , n343105 );
buf ( n343107 , n343106 );
xor ( n23138 , n343086 , n343107 );
buf ( n343109 , n342356 );
and ( n343110 , n23138 , n343109 );
and ( n23141 , n343086 , n343107 );
or ( n343112 , n343110 , n23141 );
buf ( n343113 , n343112 );
buf ( n343114 , n343113 );
xor ( n343115 , n343084 , n343114 );
buf ( n343116 , n342370 );
and ( n343117 , n343115 , n343116 );
and ( n343118 , n343084 , n343114 );
or ( n343119 , n343117 , n343118 );
buf ( n343120 , n343119 );
buf ( n343121 , n343120 );
not ( n343122 , n343121 );
buf ( n343123 , n343122 );
buf ( n343124 , n343123 );
xor ( n343125 , n343066 , n343067 );
xor ( n23156 , n343125 , n343075 );
buf ( n343127 , n23156 );
buf ( n343128 , n343127 );
buf ( n343129 , n342375 );
nor ( n343130 , n343128 , n343129 );
buf ( n343131 , n343130 );
buf ( n343132 , n343131 );
or ( n343133 , n343124 , n343132 );
buf ( n343134 , n343127 );
buf ( n343135 , n342375 );
nand ( n23166 , n343134 , n343135 );
buf ( n343137 , n23166 );
buf ( n343138 , n343137 );
nand ( n343139 , n343133 , n343138 );
buf ( n343140 , n343139 );
buf ( n343141 , n343140 );
not ( n23170 , n343141 );
buf ( n343143 , n23170 );
buf ( n343144 , n343143 );
or ( n343145 , n343083 , n343144 );
buf ( n343146 , n342389 );
buf ( n343147 , n343079 );
nand ( n343148 , n343146 , n343147 );
buf ( n343149 , n343148 );
buf ( n343150 , n343149 );
nand ( n343151 , n343145 , n343150 );
buf ( n343152 , n343151 );
buf ( n343153 , n343152 );
buf ( n343154 , n343061 );
buf ( n343155 , n342394 );
or ( n23184 , n343154 , n343155 );
buf ( n343157 , n23184 );
buf ( n343158 , n343157 );
nand ( n23187 , n343153 , n343158 );
buf ( n343160 , n23187 );
buf ( n343161 , n343160 );
nand ( n23190 , n343064 , n343161 );
buf ( n343163 , n23190 );
buf ( n343164 , n343163 );
and ( n23193 , n343056 , n343164 );
and ( n343166 , n343045 , n343055 );
or ( n343167 , n23193 , n343166 );
buf ( n343168 , n343167 );
buf ( n343169 , n343168 );
not ( n343170 , n343169 );
buf ( n343171 , n343170 );
buf ( n343172 , n343171 );
buf ( n343173 , n334009 );
buf ( n343174 , n322587 );
xor ( n23203 , n343173 , n343174 );
buf ( n343176 , n340891 );
buf ( n23205 , n340112 );
nand ( n23206 , n343176 , n23205 );
buf ( n343179 , n23206 );
buf ( n343180 , n343179 );
buf ( n23208 , n340884 );
buf ( n343182 , n23208 );
buf ( n343183 , n343182 );
buf ( n343184 , n343183 );
not ( n343185 , n343184 );
buf ( n343186 , n343185 );
buf ( n343187 , n343186 );
and ( n23213 , n343180 , n343187 );
not ( n343189 , n343180 );
buf ( n343190 , n343183 );
and ( n23215 , n343189 , n343190 );
nor ( n343192 , n23213 , n23215 );
buf ( n343193 , n343192 );
buf ( n343194 , n343193 );
xor ( n343195 , n23203 , n343194 );
buf ( n343196 , n343195 );
buf ( n343197 , n343196 );
xor ( n343198 , n322679 , n2787 );
and ( n343199 , n343198 , n343053 );
and ( n23219 , n322679 , n2787 );
or ( n343201 , n343199 , n23219 );
buf ( n343202 , n343201 );
nor ( n23222 , n343197 , n343202 );
buf ( n343204 , n23222 );
buf ( n343205 , n343204 );
or ( n343206 , n343172 , n343205 );
buf ( n23226 , n343201 );
buf ( n343208 , n343196 );
nand ( n343209 , n23226 , n343208 );
buf ( n343210 , n343209 );
buf ( n23230 , n343210 );
nand ( n23231 , n343206 , n23230 );
buf ( n23232 , n23231 );
buf ( n343214 , n23232 );
not ( n23234 , n343214 );
buf ( n23235 , n23234 );
buf ( n343217 , n23235 );
buf ( n343218 , n342425 );
xor ( n343219 , n343173 , n343174 );
and ( n343220 , n343219 , n343194 );
and ( n23240 , n343173 , n343174 );
or ( n343222 , n343220 , n23240 );
buf ( n343223 , n343222 );
buf ( n343224 , n343223 );
nor ( n23244 , n343218 , n343224 );
buf ( n23245 , n23244 );
buf ( n343227 , n23245 );
or ( n343228 , n343217 , n343227 );
buf ( n343229 , n342425 );
buf ( n343230 , n343223 );
nand ( n343231 , n343229 , n343230 );
buf ( n343232 , n343231 );
buf ( n343233 , n343232 );
nand ( n343234 , n343228 , n343233 );
buf ( n343235 , n343234 );
buf ( n343236 , n343235 );
nand ( n343237 , n343024 , n343236 );
buf ( n343238 , n343237 );
buf ( n343239 , n343238 );
nand ( n343240 , n343021 , n343239 );
buf ( n343241 , n343240 );
buf ( n343242 , n343241 );
and ( n343243 , n343013 , n343242 );
and ( n343244 , n343011 , n343012 );
or ( n23264 , n343243 , n343244 );
buf ( n343246 , n23264 );
buf ( n343247 , n343246 );
and ( n343248 , n23019 , n343247 );
and ( n23268 , n342979 , n342983 );
or ( n23269 , n343248 , n23268 );
buf ( n343251 , n23269 );
buf ( n343252 , n343251 );
and ( n343253 , n23016 , n343252 );
and ( n23271 , n23013 , n342977 );
or ( n23272 , n343253 , n23271 );
buf ( n343256 , n23272 );
buf ( n343257 , n343256 );
xor ( n343258 , n342940 , n343257 );
xor ( n343259 , n327482 , n342888 );
xnor ( n23277 , n343259 , n342909 );
buf ( n343261 , n23277 );
and ( n23278 , n343258 , n343261 );
and ( n343263 , n342940 , n343257 );
or ( n343264 , n23278 , n343263 );
buf ( n343265 , n343264 );
buf ( n343266 , n343265 );
and ( n23282 , n22966 , n343266 );
and ( n343268 , n342915 , n342916 );
or ( n343269 , n23282 , n343268 );
buf ( n343270 , n343269 );
buf ( n343271 , n343270 );
xor ( n343272 , n342887 , n343271 );
xor ( n23288 , n342861 , n327584 );
xor ( n343274 , n23288 , n342881 );
buf ( n343275 , n343274 );
and ( n23291 , n343272 , n343275 );
and ( n343277 , n342887 , n343271 );
or ( n343278 , n23291 , n343277 );
buf ( n343279 , n343278 );
buf ( n343280 , n343279 );
and ( n343281 , n342886 , n343280 );
and ( n23297 , n342860 , n342885 );
or ( n343283 , n343281 , n23297 );
buf ( n343284 , n343283 );
buf ( n343285 , n343284 );
and ( n23301 , n342856 , n343285 );
and ( n343287 , n342854 , n342855 );
or ( n343288 , n23301 , n343287 );
buf ( n343289 , n343288 );
buf ( n343290 , n343289 );
and ( n343291 , n22871 , n343290 );
and ( n23307 , n22869 , n342818 );
or ( n343293 , n343291 , n23307 );
buf ( n343294 , n343293 );
buf ( n343295 , n343294 );
buf ( n343296 , n342793 );
buf ( n343297 , n342798 );
buf ( n343298 , n342571 );
buf ( n343299 , n342537 );
nor ( n343300 , n343298 , n343299 );
buf ( n343301 , n343300 );
buf ( n343302 , n343301 );
nor ( n343303 , n343297 , n343302 );
buf ( n343304 , n343303 );
buf ( n343305 , n343304 );
nand ( n343306 , n343295 , n343296 , n343305 );
buf ( n343307 , n343306 );
buf ( n343308 , n343307 );
nand ( n23322 , n342785 , n342816 , n343308 );
buf ( n343310 , n23322 );
buf ( n343311 , n343310 );
not ( n23325 , n343311 );
or ( n343313 , n342773 , n23325 );
buf ( n343314 , n343307 );
buf ( n343315 , n342815 );
buf ( n343316 , n342777 );
nand ( n23330 , n343314 , n343315 , n343316 );
buf ( n23331 , n23330 );
buf ( n23332 , n23331 );
buf ( n23333 , n342626 );
nand ( n23334 , n23332 , n23333 );
buf ( n23335 , n23334 );
buf ( n23336 , n23335 );
nand ( n23337 , n343313 , n23336 );
buf ( n23338 , n23337 );
buf ( n23339 , n23338 );
and ( n23340 , n342768 , n23339 );
and ( n343328 , n342766 , n342767 );
or ( n343329 , n23340 , n343328 );
buf ( n343330 , n343329 );
buf ( n343331 , n343330 );
and ( n23345 , n22796 , n343331 );
and ( n23346 , n342742 , n342743 );
or ( n23347 , n23345 , n23346 );
buf ( n343335 , n23347 );
buf ( n343336 , n343335 );
and ( n343337 , n342741 , n343336 );
and ( n23351 , n342739 , n342740 );
or ( n23352 , n343337 , n23351 );
buf ( n343340 , n23352 );
buf ( n343341 , n343340 );
and ( n343342 , n22790 , n343341 );
and ( n23356 , n342736 , n342737 );
or ( n23357 , n343342 , n23356 );
buf ( n343345 , n23357 );
buf ( n343346 , n343345 );
xor ( n343347 , n342734 , n342735 );
xor ( n23361 , n343347 , n343346 );
buf ( n343349 , n23361 );
xor ( n343350 , n342734 , n342735 );
and ( n23364 , n343350 , n343346 );
and ( n343352 , n342734 , n342735 );
or ( n343353 , n23364 , n343352 );
buf ( n343354 , n343353 );
xor ( n23368 , n342736 , n342737 );
xor ( n343356 , n23368 , n343341 );
buf ( n343357 , n343356 );
xor ( n23371 , n342739 , n342740 );
xor ( n343359 , n23371 , n343336 );
buf ( n343360 , n343359 );
xor ( n23374 , n342742 , n342743 );
xor ( n343362 , n23374 , n343331 );
buf ( n343363 , n343362 );
xor ( n343364 , n342766 , n342767 );
xor ( n23378 , n343364 , n23339 );
buf ( n343366 , n23378 );
buf ( n343367 , n342793 );
buf ( n343368 , n342798 );
not ( n23382 , n343368 );
buf ( n343370 , n23382 );
buf ( n343371 , n343370 );
not ( n23385 , n343371 );
buf ( n23386 , n343301 );
not ( n343374 , n23386 );
buf ( n343375 , n343374 );
buf ( n343376 , n343375 );
not ( n343377 , n343376 );
buf ( n343378 , n343294 );
not ( n343379 , n343378 );
or ( n343380 , n343377 , n343379 );
buf ( n343381 , n342803 );
nand ( n23395 , n343380 , n343381 );
buf ( n343383 , n23395 );
buf ( n343384 , n343383 );
not ( n23398 , n343384 );
or ( n343386 , n23385 , n23398 );
buf ( n343387 , n342809 );
nand ( n343388 , n343386 , n343387 );
buf ( n343389 , n343388 );
buf ( n343390 , n343389 );
buf ( n343391 , n342777 );
not ( n23405 , n343367 );
not ( n23406 , n343390 );
or ( n23407 , n23405 , n23406 );
nand ( n343395 , n23407 , n343391 );
buf ( n343396 , n343395 );
xor ( n23410 , n22869 , n342818 );
xor ( n343398 , n23410 , n343290 );
buf ( n343399 , n343398 );
xor ( n23413 , n342854 , n342855 );
xor ( n343401 , n23413 , n343285 );
buf ( n343402 , n343401 );
xor ( n23416 , n23013 , n342977 );
xor ( n23417 , n23416 , n343252 );
buf ( n343405 , n23417 );
xor ( n343406 , n342979 , n342983 );
xor ( n23420 , n343406 , n343247 );
buf ( n343408 , n23420 );
xor ( n343409 , n343011 , n343012 );
xor ( n23423 , n343409 , n343242 );
buf ( n343411 , n23423 );
buf ( n23424 , n23235 );
buf ( n343413 , n23232 );
buf ( n343414 , n342425 );
buf ( n343415 , n343223 );
xor ( n343416 , n343414 , n343415 );
buf ( n343417 , n343416 );
buf ( n343418 , n343417 );
and ( n343419 , n343418 , n343413 );
not ( n23430 , n343418 );
and ( n23431 , n23430 , n23424 );
nor ( n343422 , n343419 , n23431 );
buf ( n343423 , n343422 );
buf ( n343424 , n343171 );
buf ( n343425 , n343168 );
buf ( n343426 , n343196 );
buf ( n343427 , n343201 );
xor ( n343428 , n343426 , n343427 );
buf ( n343429 , n343428 );
buf ( n343430 , n343429 );
and ( n343431 , n343430 , n343425 );
not ( n23440 , n343430 );
and ( n343433 , n23440 , n343424 );
nor ( n343434 , n343431 , n343433 );
buf ( n343435 , n343434 );
xor ( n343436 , n343045 , n343055 );
xor ( n343437 , n343436 , n343164 );
buf ( n343438 , n343437 );
buf ( n343439 , n343061 );
buf ( n343440 , n342394 );
xor ( n23448 , n343439 , n343440 );
buf ( n343442 , n23448 );
buf ( n343443 , n343442 );
buf ( n343444 , n343152 );
xor ( n23452 , n343443 , n343444 );
buf ( n343446 , n23452 );
buf ( n343447 , n343143 );
buf ( n343448 , n343140 );
buf ( n343449 , n342389 );
buf ( n343450 , n343079 );
xor ( n343451 , n343449 , n343450 );
buf ( n343452 , n343451 );
buf ( n343453 , n343452 );
and ( n23459 , n343453 , n343448 );
not ( n23460 , n343453 );
and ( n343456 , n23460 , n343447 );
nor ( n23462 , n23459 , n343456 );
buf ( n23463 , n23462 );
buf ( n23464 , n343123 );
buf ( n343460 , n343120 );
buf ( n343461 , n343127 );
buf ( n343462 , n342375 );
xor ( n343463 , n343461 , n343462 );
buf ( n343464 , n343463 );
buf ( n343465 , n343464 );
and ( n23471 , n343465 , n343460 );
not ( n343467 , n343465 );
and ( n343468 , n343467 , n23464 );
nor ( n23474 , n23471 , n343468 );
buf ( n23475 , n23474 );
xor ( n343471 , n343084 , n343114 );
xor ( n23477 , n343471 , n343116 );
buf ( n343473 , n23477 );
xor ( n23479 , n343087 , n343088 );
xor ( n343475 , n23479 , n343102 );
buf ( n343476 , n343475 );
buf ( n343477 , n342781 );
buf ( n343478 , n342626 );
buf ( n343479 , n342771 );
and ( n23485 , n343479 , n343478 );
not ( n343481 , n343479 );
and ( n343482 , n343481 , n343477 );
nor ( n23488 , n23485 , n343482 );
buf ( n23489 , n23488 );
buf ( n343485 , n342790 );
buf ( n343486 , n342621 );
buf ( n343487 , n342599 );
and ( n343488 , n343487 , n343486 );
not ( n343489 , n343487 );
and ( n343490 , n343489 , n343485 );
nor ( n343491 , n343488 , n343490 );
buf ( n343492 , n343491 );
buf ( n343493 , n343294 );
buf ( n343494 , n342571 );
buf ( n343495 , n342537 );
xor ( n23499 , n343494 , n343495 );
buf ( n343497 , n23499 );
buf ( n343498 , n343497 );
xor ( n23502 , n343493 , n343498 );
buf ( n343500 , n23502 );
buf ( n343501 , n343383 );
buf ( n343502 , n342576 );
buf ( n343503 , n342594 );
xor ( n343504 , n343502 , n343503 );
buf ( n343505 , n343504 );
buf ( n343506 , n343505 );
xor ( n343507 , n343501 , n343506 );
buf ( n343508 , n343507 );
buf ( n343509 , n343389 );
buf ( n343510 , n343492 );
xor ( n343511 , n343509 , n343510 );
buf ( n343512 , n343511 );
buf ( n343513 , n343396 );
buf ( n343514 , n23489 );
xor ( n23518 , n343513 , n343514 );
buf ( n23519 , n23518 );
buf ( n343517 , n342347 );
buf ( n343518 , n342733 );
xor ( n23522 , n343517 , n343518 );
buf ( n343520 , n23522 );
buf ( n343521 , n332409 );
buf ( n23525 , n332479 );
and ( n23526 , n603 , n604 );
not ( n343524 , n603 );
buf ( n343525 , n604 );
not ( n23529 , n343525 );
buf ( n23530 , n23529 );
and ( n343528 , n343524 , n23530 );
nor ( n23532 , n23526 , n343528 );
buf ( n343530 , n23532 );
buf ( n343531 , n343530 );
buf ( n343532 , n343531 );
not ( n343533 , n343532 );
buf ( n343534 , n602 );
not ( n343535 , n343534 );
not ( n343536 , n14255 );
nand ( n343537 , n343536 , n14327 );
not ( n343538 , n343537 );
nor ( n23540 , n14665 , n14837 );
nand ( n343540 , n343538 , n23540 , n14680 );
and ( n23542 , n343540 , n17937 );
not ( n343542 , n343540 );
and ( n343543 , n343542 , n15012 );
nor ( n23545 , n23542 , n343543 );
buf ( n343545 , n23545 );
buf ( n343546 , n343545 );
not ( n343547 , n343546 );
buf ( n343548 , n343547 );
buf ( n23550 , n343548 );
not ( n23551 , n23550 );
or ( n23552 , n343535 , n23551 );
buf ( n343552 , n343545 );
not ( n343553 , n602 );
buf ( n343554 , n343553 );
nand ( n23553 , n343552 , n343554 );
buf ( n23554 , n23553 );
buf ( n343557 , n23554 );
nand ( n23556 , n23552 , n343557 );
buf ( n23557 , n23556 );
buf ( n343560 , n23557 );
not ( n23559 , n343560 );
or ( n343562 , n343533 , n23559 );
buf ( n343563 , n602 );
not ( n343564 , n343563 );
buf ( n343565 , n14695 );
buf ( n343566 , n343565 );
buf ( n343567 , n343566 );
buf ( n343568 , n343567 );
not ( n343569 , n343568 );
buf ( n343570 , n343569 );
buf ( n343571 , n343570 );
not ( n343572 , n343571 );
or ( n343573 , n343564 , n343572 );
buf ( n343574 , n343567 );
buf ( n343575 , n343553 );
nand ( n343576 , n343574 , n343575 );
buf ( n343577 , n343576 );
buf ( n343578 , n343577 );
nand ( n343579 , n343573 , n343578 );
buf ( n343580 , n343579 );
buf ( n343581 , n343580 );
buf ( n343582 , n602 );
buf ( n343583 , n603 );
and ( n343584 , n343582 , n343583 );
buf ( n343585 , n23532 );
buf ( n343586 , n602 );
buf ( n343587 , n603 );
nor ( n23575 , n343586 , n343587 );
buf ( n343589 , n23575 );
buf ( n343590 , n343589 );
nor ( n343591 , n343584 , n343585 , n343590 );
buf ( n343592 , n343591 );
buf ( n343593 , n343592 );
buf ( n343594 , n343593 );
buf ( n343595 , n343594 );
buf ( n343596 , n343595 );
nand ( n343597 , n343581 , n343596 );
buf ( n343598 , n343597 );
buf ( n343599 , n343598 );
nand ( n343600 , n343562 , n343599 );
buf ( n343601 , n343600 );
buf ( n343602 , n343601 );
not ( n23590 , n334505 );
not ( n343604 , n334495 );
or ( n343605 , n23590 , n343604 );
nand ( n23593 , n343605 , n334369 );
not ( n343607 , n23593 );
not ( n343608 , n343607 );
not ( n23596 , n323949 );
not ( n343610 , n15462 );
not ( n23598 , n343610 );
or ( n343612 , n23596 , n23598 );
nand ( n343613 , n343612 , n14511 );
not ( n23601 , n343613 );
not ( n23602 , n23601 );
or ( n23603 , n343608 , n23602 );
nand ( n23604 , n343613 , n23593 );
nand ( n23605 , n23603 , n23604 );
buf ( n23606 , n23605 );
buf ( n343620 , n23606 );
not ( n23608 , n343620 );
buf ( n343622 , n592 );
not ( n343623 , n343622 );
buf ( n343624 , n343623 );
buf ( n343625 , n343624 );
nor ( n343626 , n23608 , n343625 );
buf ( n343627 , n343626 );
buf ( n343628 , n343627 );
not ( n343629 , n343628 );
buf ( n343630 , n594 );
not ( n343631 , n343630 );
buf ( n343632 , n343631 );
and ( n343633 , n593 , n343632 );
not ( n343634 , n593 );
and ( n343635 , n343634 , n594 );
or ( n23612 , n343633 , n343635 );
buf ( n23613 , n23612 );
not ( n23614 , n23613 );
nand ( n343639 , n14729 , n334614 , n14774 );
buf ( n23615 , n334334 );
not ( n23616 , n23615 );
not ( n343642 , n5821 );
and ( n23618 , n23616 , n343642 );
and ( n343644 , n23615 , n14475 );
nor ( n23620 , n23618 , n343644 );
and ( n23621 , n343639 , n23620 );
not ( n23622 , n343639 );
not ( n343648 , n23620 );
and ( n343649 , n23622 , n343648 );
nor ( n343650 , n23621 , n343649 );
not ( n343651 , n343650 );
and ( n343652 , n343651 , n592 );
not ( n23626 , n343651 );
and ( n343654 , n23626 , n343624 );
or ( n343655 , n343652 , n343654 );
not ( n23629 , n343655 );
or ( n23630 , n23614 , n23629 );
buf ( n343658 , n592 );
not ( n23632 , n343658 );
not ( n23633 , n334497 );
not ( n343661 , n14647 );
or ( n343662 , n23633 , n343661 );
nand ( n23636 , n343662 , n334373 );
not ( n23637 , n14455 );
not ( n343665 , n334317 );
or ( n343666 , n23637 , n343665 );
nand ( n23640 , n343666 , n334375 );
and ( n343668 , n23636 , n23640 );
not ( n343669 , n23636 );
not ( n23643 , n23640 );
and ( n343671 , n343669 , n23643 );
nor ( n343672 , n343668 , n343671 );
buf ( n343673 , n343672 );
not ( n23647 , n343673 );
buf ( n343675 , n23647 );
buf ( n343676 , n343675 );
not ( n23649 , n343676 );
buf ( n343678 , n23649 );
buf ( n343679 , n343678 );
not ( n23652 , n343679 );
or ( n343681 , n23632 , n23652 );
buf ( n343682 , n343675 );
buf ( n343683 , n343624 );
nand ( n23656 , n343682 , n343683 );
buf ( n343685 , n23656 );
buf ( n343686 , n343685 );
nand ( n23659 , n343681 , n343686 );
buf ( n343688 , n23659 );
buf ( n343689 , n592 );
buf ( n343690 , n593 );
and ( n343691 , n343689 , n343690 );
buf ( n23664 , n23613 );
buf ( n343693 , n592 );
buf ( n343694 , n593 );
nor ( n23667 , n343693 , n343694 );
buf ( n343696 , n23667 );
buf ( n343697 , n343696 );
nor ( n23670 , n343691 , n23664 , n343697 );
buf ( n343699 , n23670 );
nand ( n23672 , n343688 , n343699 );
nand ( n343701 , n23630 , n23672 );
not ( n23674 , n343701 );
buf ( n343703 , n23674 );
nand ( n343704 , n343629 , n343703 );
buf ( n343705 , n343704 );
buf ( n343706 , n343705 );
not ( n343707 , n343706 );
xnor ( n23680 , n596 , n595 );
not ( n23681 , n23680 );
not ( n343710 , n23681 );
not ( n343711 , n594 );
not ( n23684 , n14766 );
nand ( n343713 , n14751 , n14721 );
and ( n343714 , n334508 , n334497 );
not ( n23687 , n334337 );
nand ( n343716 , n343714 , n23687 , n14721 );
nand ( n343717 , n343713 , n343716 , n14722 );
not ( n343718 , n343717 );
not ( n343719 , n343718 );
or ( n343720 , n23684 , n343719 );
nand ( n343721 , n343717 , n334625 );
nand ( n23692 , n343720 , n343721 );
buf ( n343723 , n23692 );
not ( n23694 , n343723 );
not ( n343725 , n23694 );
or ( n23696 , n343711 , n343725 );
buf ( n343727 , n343723 );
buf ( n343728 , n343632 );
nand ( n343729 , n343727 , n343728 );
buf ( n343730 , n343729 );
nand ( n343731 , n23696 , n343730 );
not ( n343732 , n343731 );
or ( n23703 , n343710 , n343732 );
buf ( n343734 , n594 );
not ( n343735 , n343734 );
buf ( n343736 , n334588 );
not ( n343737 , n343736 );
buf ( n343738 , n343737 );
buf ( n343739 , n343738 );
not ( n343740 , n343739 );
or ( n343741 , n343735 , n343740 );
buf ( n343742 , n343738 );
not ( n23713 , n343742 );
buf ( n343744 , n23713 );
buf ( n343745 , n343744 );
buf ( n343746 , n343632 );
nand ( n343747 , n343745 , n343746 );
buf ( n343748 , n343747 );
buf ( n343749 , n343748 );
nand ( n343750 , n343741 , n343749 );
buf ( n343751 , n343750 );
buf ( n343752 , n594 );
buf ( n343753 , n595 );
and ( n23723 , n343752 , n343753 );
buf ( n343755 , n23681 );
buf ( n343756 , n594 );
buf ( n343757 , n595 );
nor ( n343758 , n343756 , n343757 );
buf ( n343759 , n343758 );
buf ( n343760 , n343759 );
nor ( n23730 , n23723 , n343755 , n343760 );
buf ( n343762 , n23730 );
buf ( n343763 , n343762 );
buf ( n23733 , n343763 );
buf ( n343765 , n23733 );
nand ( n23735 , n343751 , n343765 );
nand ( n343767 , n23703 , n23735 );
buf ( n343768 , n343767 );
not ( n343769 , n343768 );
or ( n343770 , n343707 , n343769 );
buf ( n343771 , n23674 );
not ( n343772 , n343771 );
buf ( n343773 , n343627 );
nand ( n343774 , n343772 , n343773 );
buf ( n343775 , n343774 );
buf ( n343776 , n343775 );
nand ( n343777 , n343770 , n343776 );
buf ( n343778 , n343777 );
buf ( n343779 , n343778 );
buf ( n343780 , n343675 );
buf ( n343781 , n592 );
and ( n23750 , n343780 , n343781 );
buf ( n23751 , n23750 );
buf ( n343784 , n23751 );
buf ( n343785 , n23613 );
not ( n23754 , n343785 );
buf ( n23755 , n592 );
buf ( n343788 , n334588 );
buf ( n23757 , n343788 );
buf ( n23758 , n23757 );
buf ( n343791 , n23758 );
xor ( n23760 , n23755 , n343791 );
buf ( n343793 , n23760 );
buf ( n343794 , n343793 );
not ( n23763 , n343794 );
or ( n23764 , n23754 , n23763 );
buf ( n343797 , n343655 );
buf ( n343798 , n343699 );
nand ( n23766 , n343797 , n343798 );
buf ( n343800 , n23766 );
buf ( n343801 , n343800 );
nand ( n343802 , n23764 , n343801 );
buf ( n343803 , n343802 );
buf ( n343804 , n343803 );
xor ( n23772 , n343784 , n343804 );
buf ( n343806 , n23681 );
not ( n23774 , n343806 );
buf ( n343808 , n594 );
not ( n23776 , n343808 );
and ( n23777 , n334302 , n334313 );
not ( n343811 , n23777 );
not ( n343812 , n334612 );
or ( n23780 , n343811 , n343812 );
not ( n343814 , n334509 );
and ( n343815 , n23777 , n343814 );
not ( n23783 , n334302 );
not ( n343817 , n334304 );
or ( n343818 , n23783 , n343817 );
nand ( n23786 , n343818 , n334309 );
nor ( n343820 , n343815 , n23786 );
nand ( n23788 , n23780 , n343820 );
and ( n343822 , n23788 , n14768 );
not ( n23790 , n23788 );
and ( n23791 , n23790 , n334629 );
nor ( n343825 , n343822 , n23791 );
buf ( n343826 , n343825 );
buf ( n23794 , n343826 );
buf ( n23795 , n23794 );
buf ( n343829 , n23795 );
not ( n23797 , n343829 );
buf ( n23798 , n23797 );
buf ( n343832 , n23798 );
not ( n23800 , n343832 );
or ( n23801 , n23776 , n23800 );
buf ( n343835 , n23795 );
buf ( n343836 , n343835 );
buf ( n343837 , n343836 );
buf ( n343838 , n343837 );
buf ( n343839 , n343632 );
nand ( n343840 , n343838 , n343839 );
buf ( n343841 , n343840 );
buf ( n343842 , n343841 );
nand ( n343843 , n23801 , n343842 );
buf ( n343844 , n343843 );
buf ( n343845 , n343844 );
not ( n343846 , n343845 );
or ( n343847 , n23774 , n343846 );
buf ( n343848 , n343731 );
buf ( n343849 , n343765 );
nand ( n343850 , n343848 , n343849 );
buf ( n343851 , n343850 );
buf ( n343852 , n343851 );
nand ( n343853 , n343847 , n343852 );
buf ( n343854 , n343853 );
buf ( n343855 , n343854 );
xor ( n23823 , n23772 , n343855 );
buf ( n343857 , n23823 );
buf ( n343858 , n343857 );
xor ( n23826 , n343779 , n343858 );
buf ( n343860 , n597 );
buf ( n343861 , n598 );
xor ( n343862 , n343860 , n343861 );
buf ( n343863 , n343862 );
buf ( n343864 , n343863 );
not ( n343865 , n343864 );
buf ( n343866 , n596 );
not ( n23834 , n343866 );
not ( n343868 , n14254 );
xor ( n343869 , n343868 , n14665 );
buf ( n343870 , n343869 );
not ( n343871 , n343870 );
buf ( n343872 , n343871 );
buf ( n343873 , n343872 );
not ( n23841 , n343873 );
or ( n343875 , n23834 , n23841 );
buf ( n343876 , n343872 );
not ( n23844 , n343876 );
buf ( n343878 , n23844 );
buf ( n343879 , n343878 );
buf ( n343880 , n596 );
not ( n343881 , n343880 );
buf ( n343882 , n343881 );
buf ( n343883 , n343882 );
nand ( n343884 , n343879 , n343883 );
buf ( n343885 , n343884 );
buf ( n343886 , n343885 );
nand ( n23854 , n343875 , n343886 );
buf ( n343888 , n23854 );
buf ( n343889 , n343888 );
not ( n343890 , n343889 );
or ( n343891 , n343865 , n343890 );
not ( n23859 , n14661 );
nand ( n23860 , n23859 , n14656 );
not ( n23861 , n23860 );
or ( n343895 , n334612 , n343814 );
nand ( n343896 , n343895 , n14767 );
not ( n23864 , n334314 );
or ( n343898 , n343896 , n23864 );
and ( n343899 , n14767 , n23786 );
nor ( n23867 , n343899 , n334519 );
nand ( n23868 , n343898 , n23867 );
not ( n23869 , n23868 );
or ( n23870 , n23861 , n23869 );
or ( n343904 , n23860 , n23868 );
nand ( n343905 , n23870 , n343904 );
buf ( n343906 , n343905 );
buf ( n343907 , n343906 );
buf ( n343908 , n343907 );
buf ( n343909 , n343908 );
not ( n343910 , n343909 );
buf ( n343911 , n343910 );
not ( n23879 , n343911 );
not ( n343913 , n596 );
or ( n23881 , n23879 , n343913 );
nand ( n343915 , n343908 , n343882 );
nand ( n23883 , n23881 , n343915 );
buf ( n343917 , n23883 );
and ( n23885 , n596 , n597 );
nor ( n343919 , n23885 , n343863 );
or ( n23887 , n596 , n597 );
and ( n343921 , n343919 , n23887 );
buf ( n23889 , n343921 );
buf ( n343923 , n23889 );
nand ( n23891 , n343917 , n343923 );
buf ( n343925 , n23891 );
buf ( n343926 , n343925 );
nand ( n343927 , n343891 , n343926 );
buf ( n343928 , n343927 );
buf ( n343929 , n343928 );
and ( n343930 , n23826 , n343929 );
and ( n23898 , n343779 , n343858 );
or ( n343932 , n343930 , n23898 );
buf ( n343933 , n343932 );
buf ( n343934 , n343933 );
xor ( n23902 , n343602 , n343934 );
xnor ( n343936 , n598 , n599 );
buf ( n343937 , n600 );
not ( n23905 , n343937 );
buf ( n23906 , n23905 );
and ( n343940 , n599 , n23906 );
not ( n23908 , n599 );
and ( n343942 , n23908 , n600 );
or ( n23910 , n343940 , n343942 );
buf ( n23911 , n23910 );
nor ( n343945 , n343936 , n23911 );
buf ( n343946 , n343945 );
buf ( n343947 , n343946 );
buf ( n343948 , n343947 );
buf ( n343949 , n343948 );
not ( n23917 , n343949 );
buf ( n343951 , n598 );
not ( n23919 , n343951 );
buf ( n343953 , n23919 );
not ( n23921 , n343953 );
nand ( n343955 , n334556 , n14897 );
buf ( n23923 , n14958 );
and ( n343957 , n343955 , n23923 );
not ( n23925 , n343955 );
not ( n343959 , n23923 );
and ( n343960 , n23925 , n343959 );
nor ( n23928 , n343957 , n343960 );
buf ( n343962 , n23928 );
not ( n23930 , n343962 );
not ( n343964 , n23930 );
or ( n23932 , n23921 , n343964 );
not ( n343966 , n23928 );
buf ( n23934 , n343966 );
not ( n343968 , n23934 );
buf ( n343969 , n343968 );
nand ( n343970 , n343969 , n598 );
nand ( n343971 , n23932 , n343970 );
buf ( n343972 , n343971 );
not ( n343973 , n343972 );
or ( n23941 , n23917 , n343973 );
buf ( n343975 , n598 );
not ( n343976 , n343975 );
nand ( n343977 , n334556 , n14697 );
and ( n23945 , n343977 , n335261 );
not ( n343979 , n343977 );
and ( n23947 , n343979 , n337552 );
nor ( n23948 , n23945 , n23947 );
buf ( n343982 , n23948 );
buf ( n343983 , n343982 );
not ( n23951 , n343983 );
buf ( n343985 , n23951 );
buf ( n343986 , n343985 );
not ( n23954 , n343986 );
or ( n23955 , n343976 , n23954 );
buf ( n343989 , n343982 );
buf ( n23957 , n343989 );
buf ( n343991 , n23957 );
buf ( n343992 , n343991 );
buf ( n343993 , n343953 );
nand ( n343994 , n343992 , n343993 );
buf ( n343995 , n343994 );
buf ( n343996 , n343995 );
nand ( n343997 , n23955 , n343996 );
buf ( n343998 , n343997 );
buf ( n343999 , n343998 );
buf ( n344000 , n23911 );
nand ( n344001 , n343999 , n344000 );
buf ( n344002 , n344001 );
buf ( n344003 , n344002 );
nand ( n23971 , n23941 , n344003 );
buf ( n23972 , n23971 );
buf ( n344006 , n23972 );
not ( n23974 , n344006 );
or ( n344008 , n600 , n601 );
and ( n344009 , n600 , n601 );
not ( n23977 , n602 );
and ( n344011 , n601 , n23977 );
not ( n344012 , n601 );
and ( n23980 , n344012 , n602 );
nor ( n344014 , n344011 , n23980 );
not ( n344015 , n344014 );
nor ( n23983 , n344009 , n344015 );
nand ( n344017 , n344008 , n23983 );
not ( n344018 , n344017 );
buf ( n344019 , n344018 );
not ( n344020 , n344019 );
buf ( n344021 , n600 );
not ( n23989 , n344021 );
not ( n344023 , n334561 );
not ( n23991 , n14699 );
or ( n344025 , n344023 , n23991 );
nand ( n23993 , n344025 , n14705 );
buf ( n344027 , n23993 );
not ( n23995 , n344027 );
buf ( n23996 , n23995 );
buf ( n344030 , n23996 );
not ( n344031 , n344030 );
or ( n344032 , n23989 , n344031 );
buf ( n344033 , n23993 );
buf ( n344034 , n344033 );
buf ( n344035 , n344034 );
buf ( n24003 , n344035 );
buf ( n24004 , n23906 );
nand ( n24005 , n24003 , n24004 );
buf ( n24006 , n24005 );
buf ( n344040 , n24006 );
nand ( n24008 , n344032 , n344040 );
buf ( n24009 , n24008 );
buf ( n344043 , n24009 );
not ( n344044 , n344043 );
or ( n24012 , n344020 , n344044 );
buf ( n344046 , n600 );
not ( n24014 , n344046 );
not ( n24015 , n343537 );
nand ( n24016 , n24015 , n334579 );
not ( n24017 , n337183 );
and ( n344051 , n24016 , n24017 );
not ( n24019 , n24016 );
and ( n344053 , n24019 , n15381 );
nor ( n344054 , n344051 , n344053 );
not ( n344055 , n344054 );
buf ( n344056 , n344055 );
not ( n344057 , n344056 );
or ( n344058 , n24014 , n344057 );
not ( n24026 , n344054 );
not ( n344060 , n24026 );
buf ( n344061 , n344060 );
buf ( n344062 , n23906 );
nand ( n24030 , n344061 , n344062 );
buf ( n344064 , n24030 );
buf ( n344065 , n344064 );
nand ( n344066 , n344058 , n344065 );
buf ( n344067 , n344066 );
buf ( n344068 , n344067 );
buf ( n344069 , n344015 );
nand ( n344070 , n344068 , n344069 );
buf ( n344071 , n344070 );
buf ( n344072 , n344071 );
nand ( n344073 , n24012 , n344072 );
buf ( n344074 , n344073 );
buf ( n344075 , n344074 );
not ( n344076 , n344075 );
or ( n24044 , n23974 , n344076 );
buf ( n344078 , n344074 );
buf ( n344079 , n23972 );
or ( n24047 , n344078 , n344079 );
buf ( n344081 , n23613 );
not ( n344082 , n344081 );
buf ( n344083 , n343688 );
not ( n24051 , n344083 );
or ( n344085 , n344082 , n24051 );
buf ( n344086 , n592 );
not ( n24054 , n344086 );
not ( n24055 , n343613 );
not ( n24056 , n23593 );
and ( n24057 , n24055 , n24056 );
and ( n24058 , n343613 , n23593 );
nor ( n24059 , n24057 , n24058 );
buf ( n344093 , n24059 );
not ( n24061 , n344093 );
or ( n24062 , n24054 , n24061 );
buf ( n344096 , n343624 );
buf ( n344097 , n23605 );
nand ( n24065 , n344096 , n344097 );
buf ( n344099 , n24065 );
buf ( n344100 , n344099 );
nand ( n24068 , n24062 , n344100 );
buf ( n344102 , n24068 );
buf ( n344103 , n344102 );
buf ( n344104 , n343699 );
nand ( n24072 , n344103 , n344104 );
buf ( n344106 , n24072 );
buf ( n344107 , n344106 );
nand ( n24075 , n344085 , n344107 );
buf ( n344109 , n24075 );
buf ( n344110 , n344109 );
not ( n24078 , n344110 );
buf ( n344112 , n24078 );
buf ( n344113 , n344112 );
not ( n344114 , n323556 );
not ( n24082 , n14644 );
or ( n344116 , n344114 , n24082 );
nand ( n344117 , n344116 , n334369 );
not ( n24085 , n344117 );
not ( n344119 , n334497 );
or ( n24087 , n24085 , n344119 );
not ( n24088 , n344117 );
nand ( n24089 , n24088 , n14636 );
nand ( n24090 , n24087 , n24089 );
not ( n24091 , n24090 );
not ( n24092 , n24091 );
buf ( n344126 , n24092 );
buf ( n344127 , n592 );
nand ( n24095 , n344126 , n344127 );
buf ( n344129 , n24095 );
buf ( n344130 , n344129 );
nand ( n24098 , n344113 , n344130 );
buf ( n344132 , n24098 );
buf ( n344133 , n344132 );
not ( n344134 , n344133 );
nand ( n344135 , n14634 , n14547 );
not ( n344136 , n14535 );
not ( n344137 , n14613 );
or ( n24105 , n344136 , n344137 );
nand ( n24106 , n24105 , n14753 );
xor ( n344140 , n344135 , n24106 );
not ( n24108 , n344140 );
not ( n24109 , n24108 );
not ( n24110 , n24109 );
buf ( n344144 , n24110 );
not ( n24112 , n344144 );
buf ( n344146 , n343624 );
nor ( n24114 , n24112 , n344146 );
buf ( n344148 , n24114 );
not ( n344149 , n23613 );
not ( n24117 , n344102 );
or ( n344151 , n344149 , n24117 );
not ( n344152 , n344117 );
not ( n24120 , n334497 );
or ( n344154 , n344152 , n24120 );
nand ( n344155 , n344154 , n24089 );
and ( n344156 , n344155 , n343624 );
not ( n24124 , n344155 );
and ( n344158 , n24124 , n592 );
or ( n24126 , n344156 , n344158 );
buf ( n344160 , n24126 );
buf ( n344161 , n343699 );
nand ( n344162 , n344160 , n344161 );
buf ( n344163 , n344162 );
nand ( n344164 , n344151 , n344163 );
or ( n344165 , n344148 , n344164 );
buf ( n344166 , n344165 );
not ( n344167 , n344166 );
buf ( n344168 , n23681 );
not ( n344169 , n344168 );
and ( n24137 , n343650 , n343632 );
not ( n344171 , n343650 );
and ( n24139 , n344171 , n594 );
or ( n344173 , n24137 , n24139 );
buf ( n344174 , n344173 );
not ( n344175 , n344174 );
or ( n344176 , n344169 , n344175 );
buf ( n344177 , n594 );
not ( n344178 , n344177 );
buf ( n344179 , n343672 );
not ( n24147 , n344179 );
or ( n344181 , n344178 , n24147 );
and ( n24149 , n23636 , n23643 );
not ( n24150 , n23636 );
and ( n344184 , n24150 , n23640 );
nor ( n344185 , n24149 , n344184 );
nand ( n24153 , n344185 , n343632 );
buf ( n344187 , n24153 );
nand ( n344188 , n344181 , n344187 );
buf ( n344189 , n344188 );
buf ( n344190 , n344189 );
buf ( n344191 , n343762 );
nand ( n344192 , n344190 , n344191 );
buf ( n344193 , n344192 );
buf ( n344194 , n344193 );
nand ( n24162 , n344176 , n344194 );
buf ( n344196 , n24162 );
buf ( n344197 , n344196 );
not ( n24165 , n344197 );
or ( n344199 , n344167 , n24165 );
buf ( n24167 , n344164 );
buf ( n344201 , n344148 );
nand ( n24169 , n24167 , n344201 );
buf ( n344203 , n24169 );
buf ( n344204 , n344203 );
nand ( n24172 , n344199 , n344204 );
buf ( n344206 , n24172 );
buf ( n344207 , n344206 );
not ( n24175 , n344207 );
or ( n24176 , n344134 , n24175 );
buf ( n24177 , n344109 );
buf ( n344211 , n344129 );
not ( n24179 , n344211 );
buf ( n24180 , n24179 );
buf ( n344214 , n24180 );
nand ( n24182 , n24177 , n344214 );
buf ( n24183 , n24182 );
buf ( n344217 , n24183 );
nand ( n24185 , n24176 , n344217 );
buf ( n344219 , n24185 );
buf ( n344220 , n344219 );
buf ( n344221 , n343863 );
not ( n344222 , n344221 );
buf ( n344223 , n23883 );
not ( n344224 , n344223 );
or ( n344225 , n344222 , n344224 );
buf ( n344226 , n596 );
not ( n24194 , n344226 );
buf ( n24195 , n23795 );
not ( n344229 , n24195 );
buf ( n344230 , n344229 );
buf ( n344231 , n344230 );
not ( n344232 , n344231 );
or ( n24200 , n24194 , n344232 );
buf ( n344234 , n23795 );
buf ( n344235 , n343882 );
nand ( n24203 , n344234 , n344235 );
buf ( n344237 , n24203 );
buf ( n344238 , n344237 );
nand ( n344239 , n24200 , n344238 );
buf ( n344240 , n344239 );
buf ( n344241 , n344240 );
buf ( n344242 , n23889 );
nand ( n344243 , n344241 , n344242 );
buf ( n344244 , n344243 );
buf ( n344245 , n344244 );
nand ( n344246 , n344225 , n344245 );
buf ( n344247 , n344246 );
buf ( n344248 , n344247 );
xor ( n24216 , n344220 , n344248 );
not ( n344250 , n343627 );
and ( n24218 , n343701 , n344250 );
not ( n344252 , n343701 );
and ( n24220 , n344252 , n343627 );
or ( n24221 , n24218 , n24220 );
xor ( n344255 , n24221 , n343767 );
buf ( n344256 , n344255 );
and ( n24224 , n24216 , n344256 );
and ( n344258 , n344220 , n344248 );
or ( n344259 , n24224 , n344258 );
buf ( n344260 , n344259 );
buf ( n344261 , n344260 );
nand ( n344262 , n24047 , n344261 );
buf ( n344263 , n344262 );
buf ( n344264 , n344263 );
nand ( n344265 , n24044 , n344264 );
buf ( n344266 , n344265 );
buf ( n344267 , n344266 );
and ( n344268 , n23902 , n344267 );
and ( n344269 , n343602 , n343934 );
or ( n24237 , n344268 , n344269 );
buf ( n344271 , n24237 );
buf ( n344272 , n23911 );
not ( n344273 , n344272 );
and ( n344274 , n598 , n23996 );
not ( n24242 , n598 );
and ( n24243 , n24242 , n344035 );
or ( n344277 , n344274 , n24243 );
buf ( n344278 , n344277 );
not ( n24246 , n344278 );
or ( n344280 , n344273 , n24246 );
buf ( n344281 , n343948 );
buf ( n344282 , n343998 );
nand ( n24250 , n344281 , n344282 );
buf ( n344284 , n24250 );
buf ( n344285 , n344284 );
nand ( n24253 , n344280 , n344285 );
buf ( n24254 , n24253 );
not ( n344288 , n24254 );
buf ( n344289 , n344015 );
not ( n344290 , n344289 );
buf ( n344291 , n600 );
not ( n24259 , n344291 );
nand ( n24260 , n334632 , n334556 , n334647 );
not ( n24261 , n334709 );
and ( n344295 , n24260 , n24261 );
not ( n344296 , n24260 );
and ( n24264 , n344296 , n334709 );
nor ( n24265 , n344295 , n24264 );
buf ( n344299 , n24265 );
not ( n344300 , n344299 );
buf ( n344301 , n344300 );
buf ( n344302 , n344301 );
not ( n344303 , n344302 );
or ( n24271 , n24259 , n344303 );
buf ( n344305 , n23906 );
buf ( n344306 , n24265 );
not ( n24274 , n344306 );
buf ( n344308 , n24274 );
buf ( n344309 , n344308 );
not ( n24277 , n344309 );
buf ( n24278 , n24277 );
buf ( n344312 , n24278 );
nand ( n24280 , n344305 , n344312 );
buf ( n344314 , n24280 );
buf ( n24282 , n344314 );
nand ( n24283 , n24271 , n24282 );
buf ( n24284 , n24283 );
buf ( n344318 , n24284 );
not ( n24286 , n344318 );
or ( n24287 , n344290 , n24286 );
buf ( n344321 , n344067 );
buf ( n344322 , n344018 );
nand ( n24290 , n344321 , n344322 );
buf ( n344324 , n24290 );
buf ( n344325 , n344324 );
nand ( n24293 , n24287 , n344325 );
buf ( n24294 , n24293 );
not ( n24295 , n24294 );
not ( n24296 , n24295 );
or ( n24297 , n344288 , n24296 );
not ( n344331 , n24254 );
nand ( n344332 , n24294 , n344331 );
nand ( n24300 , n24297 , n344332 );
buf ( n344334 , n605 );
buf ( n344335 , n606 );
xor ( n344336 , n344334 , n344335 );
buf ( n344337 , n344336 );
buf ( n344338 , n344337 );
buf ( n344339 , n344338 );
not ( n344340 , n344339 );
buf ( n344341 , n604 );
not ( n344342 , n344341 );
not ( n344343 , n15128 );
not ( n24311 , n344343 );
not ( n344345 , n24311 );
not ( n344346 , n14709 );
not ( n24314 , n344346 );
or ( n344348 , n344345 , n24314 );
nand ( n344349 , n14709 , n344343 );
nand ( n344350 , n344348 , n344349 );
buf ( n344351 , n344350 );
not ( n344352 , n344351 );
buf ( n344353 , n344352 );
buf ( n344354 , n344353 );
not ( n344355 , n344354 );
or ( n24323 , n344342 , n344355 );
buf ( n344357 , n23530 );
not ( n344358 , n344346 );
not ( n24326 , n15129 );
or ( n344360 , n344358 , n24326 );
nand ( n344361 , n344360 , n344349 );
buf ( n344362 , n344361 );
nand ( n24330 , n344357 , n344362 );
buf ( n344364 , n24330 );
buf ( n344365 , n344364 );
nand ( n344366 , n24323 , n344365 );
buf ( n344367 , n344366 );
buf ( n344368 , n344367 );
not ( n24336 , n344368 );
or ( n344370 , n344340 , n24336 );
not ( n344371 , n14711 );
not ( n24339 , n334615 );
or ( n24340 , n344371 , n24339 );
not ( n24341 , n14711 );
not ( n24342 , n334623 );
or ( n24343 , n24341 , n24342 );
nand ( n344377 , n24343 , n14706 );
nand ( n24345 , n24340 , n344377 );
buf ( n24346 , n24345 );
not ( n344380 , n24346 );
not ( n24348 , n23530 );
or ( n24349 , n344380 , n24348 );
not ( n344383 , n24345 );
nand ( n344384 , n604 , n344383 );
nand ( n24352 , n24349 , n344384 );
buf ( n344386 , n24352 );
buf ( n344387 , n604 );
buf ( n344388 , n605 );
and ( n344389 , n344387 , n344388 );
buf ( n344390 , n344338 );
buf ( n344391 , n604 );
buf ( n344392 , n605 );
nor ( n24360 , n344391 , n344392 );
buf ( n344394 , n24360 );
buf ( n344395 , n344394 );
nor ( n24363 , n344389 , n344390 , n344395 );
buf ( n344397 , n24363 );
buf ( n24365 , n344397 );
buf ( n24366 , n24365 );
buf ( n344400 , n24366 );
buf ( n344401 , n344400 );
nand ( n24369 , n344386 , n344401 );
buf ( n344403 , n24369 );
buf ( n344404 , n344403 );
nand ( n24372 , n344370 , n344404 );
buf ( n344406 , n24372 );
and ( n24374 , n24300 , n344406 );
not ( n24375 , n24300 );
not ( n24376 , n344406 );
and ( n24377 , n24375 , n24376 );
nor ( n24378 , n24374 , n24377 );
buf ( n344412 , n24378 );
not ( n344413 , n344412 );
buf ( n344414 , n607 );
not ( n24382 , n344414 );
not ( n24383 , n334578 );
and ( n24384 , n14214 , n14329 );
not ( n344418 , n24384 );
or ( n344419 , n24383 , n344418 );
not ( n24387 , n15300 );
not ( n24388 , n24387 );
nand ( n24389 , n344419 , n24388 );
nand ( n24390 , n24384 , n24387 , n334578 );
nand ( n24391 , n24389 , n24390 );
not ( n24392 , n24391 );
or ( n24393 , n606 , n24392 );
nand ( n24394 , n606 , n24392 );
nand ( n24395 , n24393 , n24394 );
buf ( n344429 , n24395 );
not ( n344430 , n344429 );
or ( n24398 , n24382 , n344430 );
not ( n344432 , n606 );
not ( n24400 , n334576 );
nand ( n24401 , n24384 , n14720 );
xor ( n344435 , n24400 , n24401 );
buf ( n344436 , n344435 );
not ( n24404 , n344436 );
or ( n344438 , n344432 , n24404 );
buf ( n344439 , n344435 );
not ( n24407 , n344439 );
buf ( n24408 , n24407 );
buf ( n344442 , n24408 );
buf ( n344443 , n606 );
not ( n24411 , n344443 );
buf ( n344445 , n24411 );
buf ( n344446 , n344445 );
nand ( n24414 , n344442 , n344446 );
buf ( n344448 , n24414 );
nand ( n344449 , n344438 , n344448 );
buf ( n344450 , n607 );
not ( n344451 , n344450 );
buf ( n344452 , n344451 );
nand ( n24420 , n344452 , n606 );
not ( n344454 , n24420 );
nand ( n344455 , n344449 , n344454 );
buf ( n344456 , n344455 );
nand ( n24424 , n24398 , n344456 );
buf ( n344458 , n24424 );
buf ( n344459 , n344458 );
not ( n24427 , n344459 );
or ( n344461 , n344413 , n24427 );
buf ( n344462 , n24378 );
buf ( n344463 , n344458 );
or ( n24431 , n344462 , n344463 );
xor ( n24432 , n343784 , n343804 );
and ( n344466 , n24432 , n343855 );
and ( n344467 , n343784 , n343804 );
or ( n24435 , n344466 , n344467 );
buf ( n344469 , n24435 );
buf ( n344470 , n344469 );
not ( n24438 , n23613 );
not ( n24439 , n592 );
not ( n344473 , n23694 );
or ( n344474 , n24439 , n344473 );
nand ( n344475 , n343723 , n343624 );
nand ( n24443 , n344474 , n344475 );
not ( n344477 , n24443 );
or ( n344478 , n24438 , n344477 );
buf ( n344479 , n343793 );
buf ( n344480 , n343699 );
nand ( n344481 , n344479 , n344480 );
buf ( n344482 , n344481 );
nand ( n344483 , n344478 , n344482 );
buf ( n344484 , n343651 );
not ( n24452 , n344484 );
buf ( n344486 , n24452 );
buf ( n344487 , n592 );
and ( n344488 , n344486 , n344487 );
buf ( n344489 , n344488 );
not ( n24457 , n344489 );
xor ( n344491 , n344483 , n24457 );
buf ( n344492 , n23681 );
not ( n344493 , n344492 );
buf ( n344494 , n594 );
not ( n344495 , n344494 );
buf ( n24463 , n343911 );
not ( n24464 , n24463 );
or ( n24465 , n344495 , n24464 );
buf ( n344499 , n343908 );
buf ( n344500 , n343632 );
nand ( n344501 , n344499 , n344500 );
buf ( n344502 , n344501 );
buf ( n344503 , n344502 );
nand ( n344504 , n24465 , n344503 );
buf ( n344505 , n344504 );
buf ( n344506 , n344505 );
not ( n344507 , n344506 );
or ( n344508 , n344493 , n344507 );
buf ( n344509 , n343844 );
buf ( n344510 , n343765 );
nand ( n344511 , n344509 , n344510 );
buf ( n344512 , n344511 );
buf ( n344513 , n344512 );
nand ( n344514 , n344508 , n344513 );
buf ( n344515 , n344514 );
not ( n24483 , n344515 );
and ( n24484 , n344491 , n24483 );
not ( n24485 , n344491 );
and ( n344519 , n24485 , n344515 );
nor ( n344520 , n24484 , n344519 );
buf ( n344521 , n344520 );
xor ( n344522 , n344470 , n344521 );
buf ( n24490 , n343863 );
not ( n24491 , n24490 );
not ( n24492 , n343882 );
not ( n24493 , n23930 );
or ( n24494 , n24492 , n24493 );
nand ( n24495 , n343969 , n596 );
nand ( n24496 , n24494 , n24495 );
not ( n24497 , n24496 );
or ( n24498 , n24491 , n24497 );
buf ( n344532 , n343888 );
buf ( n344533 , n23889 );
nand ( n24501 , n344532 , n344533 );
buf ( n344535 , n24501 );
nand ( n24503 , n24498 , n344535 );
buf ( n344537 , n24503 );
xor ( n24505 , n344522 , n344537 );
buf ( n344539 , n24505 );
buf ( n344540 , n344539 );
nand ( n24508 , n24431 , n344540 );
buf ( n344542 , n24508 );
buf ( n344543 , n344542 );
nand ( n24511 , n344461 , n344543 );
buf ( n24512 , n24511 );
xor ( n24513 , n344271 , n24512 );
xor ( n24514 , n344470 , n344521 );
and ( n24515 , n24514 , n344537 );
and ( n24516 , n344470 , n344521 );
or ( n344550 , n24515 , n24516 );
buf ( n344551 , n344550 );
buf ( n344552 , n344515 );
not ( n344553 , n344552 );
buf ( n344554 , n344489 );
not ( n344555 , n344554 );
not ( n24523 , n344483 );
buf ( n344557 , n24523 );
nand ( n344558 , n344555 , n344557 );
buf ( n344559 , n344558 );
buf ( n344560 , n344559 );
not ( n24528 , n344560 );
or ( n344562 , n344553 , n24528 );
buf ( n344563 , n24523 );
not ( n24531 , n344563 );
buf ( n344565 , n344489 );
nand ( n344566 , n24531 , n344565 );
buf ( n344567 , n344566 );
buf ( n344568 , n344567 );
nand ( n344569 , n344562 , n344568 );
buf ( n344570 , n344569 );
not ( n344571 , n23889 );
not ( n344572 , n24496 );
or ( n24540 , n344571 , n344572 );
and ( n24541 , n343982 , n343882 );
not ( n24542 , n343982 );
and ( n24543 , n24542 , n596 );
or ( n344577 , n24541 , n24543 );
nand ( n344578 , n24490 , n344577 );
nand ( n24546 , n24540 , n344578 );
xor ( n24547 , n344570 , n24546 );
buf ( n344581 , n23911 );
not ( n344582 , n344581 );
buf ( n344583 , n598 );
not ( n24551 , n344583 );
buf ( n344585 , n24026 );
not ( n24553 , n344585 );
or ( n344587 , n24551 , n24553 );
buf ( n344588 , n344054 );
buf ( n344589 , n344588 );
buf ( n344590 , n343953 );
nand ( n344591 , n344589 , n344590 );
buf ( n344592 , n344591 );
buf ( n344593 , n344592 );
nand ( n344594 , n344587 , n344593 );
buf ( n344595 , n344594 );
buf ( n344596 , n344595 );
not ( n344597 , n344596 );
or ( n344598 , n344582 , n344597 );
buf ( n344599 , n344277 );
buf ( n344600 , n343948 );
nand ( n24568 , n344599 , n344600 );
buf ( n344602 , n24568 );
buf ( n344603 , n344602 );
nand ( n344604 , n344598 , n344603 );
buf ( n344605 , n344604 );
xor ( n24573 , n24547 , n344605 );
buf ( n24574 , n24573 );
xor ( n344608 , n344551 , n24574 );
not ( n344609 , n607 );
not ( n24577 , n606 );
not ( n24578 , n14710 );
nand ( n24579 , n24578 , n14762 , n344343 , n334618 );
not ( n344613 , n15289 );
and ( n344614 , n24579 , n344613 );
not ( n24582 , n24579 );
and ( n344616 , n24582 , n15290 );
nor ( n344617 , n344614 , n344616 );
buf ( n344618 , n344617 );
not ( n24586 , n344618 );
not ( n344620 , n24586 );
or ( n24588 , n24577 , n344620 );
buf ( n344622 , n344618 );
buf ( n344623 , n344445 );
nand ( n24591 , n344622 , n344623 );
buf ( n344625 , n24591 );
nand ( n344626 , n24588 , n344625 );
not ( n24594 , n344626 );
or ( n24595 , n344609 , n24594 );
buf ( n344629 , n344454 );
not ( n24597 , n344629 );
buf ( n344631 , n24597 );
not ( n344632 , n344631 );
nand ( n24600 , n344632 , n24395 );
nand ( n24601 , n24595 , n24600 );
not ( n344635 , n24601 );
xnor ( n344636 , n344608 , n344635 );
xnor ( n24604 , n24513 , n344636 );
not ( n344638 , n24604 );
not ( n24606 , n344638 );
buf ( n344640 , n344015 );
not ( n344641 , n344640 );
and ( n24609 , n14695 , n23906 );
not ( n24610 , n14695 );
and ( n24611 , n24610 , n600 );
or ( n24612 , n24609 , n24611 );
buf ( n344646 , n24612 );
not ( n344647 , n344646 );
or ( n344648 , n344641 , n344647 );
buf ( n344649 , n24284 );
buf ( n344650 , n344018 );
nand ( n344651 , n344649 , n344650 );
buf ( n344652 , n344651 );
buf ( n344653 , n344652 );
nand ( n344654 , n344648 , n344653 );
buf ( n344655 , n344654 );
buf ( n24623 , n344655 );
buf ( n344657 , n344505 );
not ( n24625 , n344657 );
buf ( n24626 , n24625 );
buf ( n344660 , n24626 );
not ( n24628 , n344660 );
buf ( n24629 , n343765 );
not ( n24630 , n24629 );
buf ( n24631 , n24630 );
buf ( n344665 , n24631 );
not ( n24633 , n344665 );
and ( n344667 , n24628 , n24633 );
buf ( n344668 , n594 );
not ( n24636 , n344668 );
buf ( n344670 , n343872 );
not ( n24638 , n344670 );
or ( n344672 , n24636 , n24638 );
buf ( n344673 , n343869 );
buf ( n344674 , n343632 );
nand ( n344675 , n344673 , n344674 );
buf ( n344676 , n344675 );
buf ( n344677 , n344676 );
nand ( n24645 , n344672 , n344677 );
buf ( n344679 , n24645 );
buf ( n344680 , n344679 );
buf ( n344681 , n23681 );
and ( n344682 , n344680 , n344681 );
nor ( n24650 , n344667 , n344682 );
buf ( n344684 , n24650 );
and ( n344685 , n23755 , n343791 );
buf ( n344686 , n344685 );
buf ( n344687 , n344686 );
buf ( n344688 , n23613 );
not ( n344689 , n344688 );
buf ( n344690 , n592 );
buf ( n344691 , n344230 );
and ( n24659 , n344690 , n344691 );
not ( n24660 , n344690 );
buf ( n344694 , n343837 );
and ( n344695 , n24660 , n344694 );
nor ( n24663 , n24659 , n344695 );
buf ( n344697 , n24663 );
not ( n344698 , n344697 );
buf ( n344699 , n344698 );
not ( n24667 , n344699 );
or ( n24668 , n344689 , n24667 );
buf ( n344702 , n24443 );
buf ( n344703 , n343699 );
buf ( n344704 , n344703 );
buf ( n344705 , n344704 );
buf ( n344706 , n344705 );
nand ( n24674 , n344702 , n344706 );
buf ( n344708 , n24674 );
buf ( n344709 , n344708 );
nand ( n344710 , n24668 , n344709 );
buf ( n344711 , n344710 );
buf ( n344712 , n344711 );
and ( n344713 , n344687 , n344712 );
not ( n24681 , n344687 );
buf ( n344715 , n344711 );
not ( n344716 , n344715 );
buf ( n344717 , n344716 );
buf ( n344718 , n344717 );
and ( n344719 , n24681 , n344718 );
nor ( n24687 , n344713 , n344719 );
buf ( n344721 , n24687 );
xor ( n344722 , n344684 , n344721 );
buf ( n344723 , n344722 );
xor ( n24691 , n24623 , n344723 );
buf ( n344725 , n343531 );
not ( n344726 , n344725 );
buf ( n344727 , n602 );
not ( n24695 , n344727 );
buf ( n344729 , n344383 );
not ( n24697 , n344729 );
or ( n344731 , n24695 , n24697 );
buf ( n24699 , n24346 );
buf ( n24700 , n343553 );
nand ( n24701 , n24699 , n24700 );
buf ( n344735 , n24701 );
buf ( n344736 , n344735 );
nand ( n344737 , n344731 , n344736 );
buf ( n344738 , n344737 );
buf ( n344739 , n344738 );
not ( n24707 , n344739 );
or ( n24708 , n344726 , n24707 );
buf ( n344742 , n23557 );
buf ( n344743 , n343595 );
nand ( n24711 , n344742 , n344743 );
buf ( n344745 , n24711 );
buf ( n344746 , n344745 );
nand ( n24714 , n24708 , n344746 );
buf ( n344748 , n24714 );
buf ( n344749 , n344748 );
not ( n24717 , n344749 );
buf ( n344751 , n24717 );
buf ( n344752 , n344751 );
xor ( n24720 , n24691 , n344752 );
buf ( n344754 , n24720 );
buf ( n344755 , n344754 );
buf ( n344756 , n344338 );
not ( n344757 , n344756 );
not ( n344758 , n23530 );
not ( n344759 , n24408 );
or ( n24727 , n344758 , n344759 );
nand ( n344761 , n344436 , n604 );
nand ( n24729 , n24727 , n344761 );
buf ( n344763 , n24729 );
not ( n24731 , n344763 );
or ( n344765 , n344757 , n24731 );
buf ( n24733 , n344367 );
buf ( n24734 , n344400 );
nand ( n24735 , n24733 , n24734 );
buf ( n24736 , n24735 );
buf ( n344770 , n24736 );
nand ( n24738 , n344765 , n344770 );
buf ( n344772 , n24738 );
buf ( n344773 , n344772 );
and ( n24741 , n344755 , n344773 );
not ( n344775 , n344755 );
not ( n24743 , n344772 );
buf ( n344777 , n24743 );
and ( n344778 , n344775 , n344777 );
nor ( n24746 , n24741 , n344778 );
buf ( n24747 , n24746 );
buf ( n344781 , n24747 );
not ( n24749 , n344406 );
nand ( n344783 , n24295 , n344331 );
not ( n344784 , n344783 );
or ( n24752 , n24749 , n344784 );
nand ( n24753 , n24254 , n24294 );
nand ( n344787 , n24752 , n24753 );
buf ( n344788 , n344787 );
not ( n24756 , n344788 );
buf ( n344790 , n24756 );
buf ( n344791 , n344790 );
and ( n344792 , n344781 , n344791 );
not ( n24760 , n344781 );
buf ( n24761 , n344787 );
and ( n344795 , n24760 , n24761 );
nor ( n344796 , n344792 , n344795 );
buf ( n344797 , n344796 );
not ( n344798 , n344797 );
not ( n344799 , n344798 );
buf ( n344800 , n343531 );
not ( n344801 , n344800 );
buf ( n24769 , n343580 );
not ( n24770 , n24769 );
or ( n24771 , n344801 , n24770 );
buf ( n344805 , n602 );
not ( n24773 , n344805 );
buf ( n344807 , n344308 );
not ( n344808 , n344807 );
or ( n344809 , n24773 , n344808 );
buf ( n344810 , n24278 );
buf ( n344811 , n343553 );
nand ( n344812 , n344810 , n344811 );
buf ( n344813 , n344812 );
buf ( n344814 , n344813 );
nand ( n344815 , n344809 , n344814 );
buf ( n344816 , n344815 );
buf ( n344817 , n344816 );
buf ( n344818 , n343595 );
nand ( n24786 , n344817 , n344818 );
buf ( n344820 , n24786 );
buf ( n344821 , n344820 );
nand ( n24789 , n24771 , n344821 );
buf ( n344823 , n24789 );
buf ( n344824 , n344823 );
not ( n24792 , n344824 );
not ( n344826 , n344338 );
not ( n344827 , n24352 );
or ( n344828 , n344826 , n344827 );
buf ( n344829 , n604 );
not ( n344830 , n344829 );
buf ( n344831 , n343545 );
not ( n24799 , n344831 );
buf ( n24800 , n24799 );
buf ( n344834 , n24800 );
not ( n24802 , n344834 );
or ( n344836 , n344830 , n24802 );
buf ( n344837 , n604 );
not ( n344838 , n344837 );
buf ( n344839 , n343545 );
nand ( n344840 , n344838 , n344839 );
buf ( n344841 , n344840 );
buf ( n344842 , n344841 );
nand ( n344843 , n344836 , n344842 );
buf ( n344844 , n344843 );
buf ( n344845 , n344844 );
buf ( n344846 , n344400 );
nand ( n24814 , n344845 , n344846 );
buf ( n344848 , n24814 );
nand ( n24816 , n344828 , n344848 );
not ( n24817 , n24816 );
not ( n24818 , n24817 );
buf ( n344852 , n24818 );
not ( n344853 , n344852 );
or ( n344854 , n24792 , n344853 );
buf ( n344855 , n344823 );
not ( n344856 , n344855 );
buf ( n344857 , n344856 );
buf ( n344858 , n344857 );
not ( n344859 , n344858 );
buf ( n344860 , n24817 );
not ( n24828 , n344860 );
or ( n24829 , n344859 , n24828 );
xor ( n24830 , n343779 , n343858 );
xor ( n24831 , n24830 , n343929 );
buf ( n344865 , n24831 );
buf ( n344866 , n344865 );
nand ( n24834 , n24829 , n344866 );
buf ( n344868 , n24834 );
buf ( n344869 , n344868 );
nand ( n24837 , n344854 , n344869 );
buf ( n344871 , n24837 );
not ( n344872 , n344871 );
not ( n24840 , n344872 );
xor ( n24841 , n343602 , n343934 );
xor ( n24842 , n24841 , n344267 );
buf ( n344876 , n24842 );
not ( n344877 , n344876 );
not ( n344878 , n344877 );
or ( n344879 , n24840 , n344878 );
not ( n344880 , n344338 );
not ( n24848 , n344844 );
or ( n344882 , n344880 , n24848 );
xor ( n344883 , n604 , n14695 );
buf ( n24851 , n344883 );
buf ( n24852 , n344400 );
nand ( n24853 , n24851 , n24852 );
buf ( n24854 , n24853 );
nand ( n24855 , n344882 , n24854 );
not ( n344889 , n24855 );
not ( n24857 , n343531 );
not ( n24858 , n344816 );
or ( n344892 , n24857 , n24858 );
buf ( n344893 , n602 );
not ( n24861 , n344893 );
not ( n344895 , n344055 );
not ( n344896 , n344895 );
buf ( n344897 , n344896 );
not ( n24865 , n344897 );
or ( n344899 , n24861 , n24865 );
buf ( n344900 , n344895 );
buf ( n344901 , n343553 );
nand ( n24869 , n344900 , n344901 );
buf ( n344903 , n24869 );
buf ( n344904 , n344903 );
nand ( n344905 , n344899 , n344904 );
buf ( n344906 , n344905 );
buf ( n24874 , n344906 );
buf ( n24875 , n343595 );
nand ( n24876 , n24874 , n24875 );
buf ( n24877 , n24876 );
nand ( n344911 , n344892 , n24877 );
not ( n344912 , n344911 );
or ( n24880 , n344889 , n344912 );
buf ( n344914 , n24855 );
not ( n24882 , n344914 );
buf ( n344916 , n24882 );
not ( n24884 , n344916 );
buf ( n344918 , n344911 );
not ( n344919 , n344918 );
buf ( n344920 , n344919 );
not ( n24888 , n344920 );
or ( n344922 , n24884 , n24888 );
xor ( n24890 , n344220 , n344248 );
xor ( n24891 , n24890 , n344256 );
buf ( n344925 , n24891 );
nand ( n24893 , n344922 , n344925 );
nand ( n344927 , n24880 , n24893 );
not ( n344928 , n344927 );
buf ( n344929 , n344015 );
not ( n24897 , n344929 );
buf ( n344931 , n24009 );
not ( n24899 , n344931 );
or ( n344933 , n24897 , n24899 );
nand ( n24901 , n343985 , n600 );
not ( n344935 , n24901 );
buf ( n344936 , n343991 );
buf ( n344937 , n23906 );
nand ( n344938 , n344936 , n344937 );
buf ( n344939 , n344938 );
not ( n344940 , n344939 );
or ( n24908 , n344935 , n344940 );
nand ( n344942 , n24908 , n344018 );
buf ( n344943 , n344942 );
nand ( n24911 , n344933 , n344943 );
buf ( n24912 , n24911 );
not ( n344946 , n24912 );
not ( n24914 , n23911 );
not ( n344948 , n343971 );
or ( n24916 , n24914 , n344948 );
buf ( n344950 , n598 );
not ( n344951 , n344950 );
buf ( n344952 , n343872 );
not ( n24920 , n344952 );
or ( n344954 , n344951 , n24920 );
buf ( n344955 , n343869 );
buf ( n24923 , n344955 );
buf ( n344957 , n24923 );
buf ( n344958 , n344957 );
buf ( n344959 , n343953 );
nand ( n344960 , n344958 , n344959 );
buf ( n344961 , n344960 );
buf ( n344962 , n344961 );
nand ( n344963 , n344954 , n344962 );
buf ( n344964 , n344963 );
nand ( n24932 , n344964 , n343948 );
nand ( n24933 , n24916 , n24932 );
not ( n24934 , n24933 );
or ( n344968 , n344946 , n24934 );
buf ( n344969 , n23911 );
not ( n344970 , n344969 );
buf ( n344971 , n343971 );
not ( n24939 , n344971 );
or ( n24940 , n344970 , n24939 );
buf ( n344974 , n24932 );
nand ( n24942 , n24940 , n344974 );
buf ( n344976 , n24942 );
buf ( n344977 , n344976 );
buf ( n344978 , n24912 );
or ( n24946 , n344977 , n344978 );
buf ( n344980 , n23681 );
not ( n24948 , n344980 );
buf ( n344982 , n343751 );
not ( n24950 , n344982 );
or ( n24951 , n24948 , n24950 );
buf ( n344985 , n344173 );
buf ( n344986 , n343765 );
nand ( n24954 , n344985 , n344986 );
buf ( n344988 , n24954 );
buf ( n344989 , n344988 );
nand ( n24957 , n24951 , n344989 );
buf ( n344991 , n24957 );
buf ( n344992 , n344991 );
buf ( n344993 , n343863 );
not ( n344994 , n344993 );
buf ( n344995 , n344240 );
not ( n344996 , n344995 );
or ( n24964 , n344994 , n344996 );
buf ( n344998 , n596 );
not ( n344999 , n344998 );
buf ( n345000 , n23694 );
not ( n24968 , n345000 );
or ( n345002 , n344999 , n24968 );
buf ( n24970 , n343723 );
buf ( n345004 , n343882 );
nand ( n345005 , n24970 , n345004 );
buf ( n345006 , n345005 );
buf ( n345007 , n345006 );
nand ( n345008 , n345002 , n345007 );
buf ( n345009 , n345008 );
buf ( n345010 , n345009 );
buf ( n345011 , n23889 );
nand ( n345012 , n345010 , n345011 );
buf ( n345013 , n345012 );
buf ( n345014 , n345013 );
nand ( n345015 , n24964 , n345014 );
buf ( n345016 , n345015 );
buf ( n345017 , n345016 );
xor ( n24985 , n344992 , n345017 );
buf ( n345019 , n344112 );
buf ( n345020 , n344129 );
and ( n345021 , n345019 , n345020 );
not ( n345022 , n345019 );
buf ( n24990 , n24180 );
and ( n345024 , n345022 , n24990 );
nor ( n24992 , n345021 , n345024 );
buf ( n24993 , n24992 );
xor ( n24994 , n344206 , n24993 );
buf ( n345028 , n24994 );
and ( n24996 , n24985 , n345028 );
and ( n24997 , n344992 , n345017 );
or ( n24998 , n24996 , n24997 );
buf ( n345032 , n24998 );
buf ( n345033 , n345032 );
nand ( n25001 , n24946 , n345033 );
buf ( n345035 , n25001 );
nand ( n25003 , n344968 , n345035 );
not ( n345037 , n25003 );
or ( n25005 , n344928 , n345037 );
buf ( n345039 , n344927 );
buf ( n345040 , n25003 );
or ( n25008 , n345039 , n345040 );
buf ( n345042 , n344260 );
buf ( n345043 , n23972 );
xor ( n345044 , n345042 , n345043 );
buf ( n345045 , n344074 );
xor ( n25013 , n345044 , n345045 );
buf ( n25014 , n25013 );
buf ( n345048 , n25014 );
nand ( n25016 , n25008 , n345048 );
buf ( n345050 , n25016 );
nand ( n25018 , n25005 , n345050 );
nand ( n345052 , n344879 , n25018 );
buf ( n25020 , n344876 );
buf ( n25021 , n344871 );
nand ( n25022 , n25020 , n25021 );
buf ( n345056 , n25022 );
nand ( n25024 , n345052 , n345056 );
not ( n25025 , n25024 );
not ( n345059 , n25025 );
or ( n25027 , n344799 , n345059 );
not ( n345061 , n344797 );
or ( n345062 , n25025 , n345061 );
nand ( n25030 , n25027 , n345062 );
not ( n25031 , n25030 );
or ( n345065 , n24606 , n25031 );
or ( n25033 , n25030 , n344638 );
nand ( n25034 , n345065 , n25033 );
not ( n25035 , n344539 );
not ( n25036 , n344458 );
not ( n345070 , n25036 );
or ( n345071 , n25035 , n345070 );
not ( n345072 , n344539 );
nand ( n345073 , n345072 , n344458 );
nand ( n25041 , n345071 , n345073 );
buf ( n345075 , n24378 );
and ( n345076 , n25041 , n345075 );
not ( n25044 , n25041 );
not ( n345078 , n345075 );
and ( n345079 , n25044 , n345078 );
nor ( n25047 , n345076 , n345079 );
buf ( n345081 , n25047 );
buf ( n345082 , n607 );
not ( n25050 , n345082 );
buf ( n345084 , n344449 );
not ( n345085 , n345084 );
or ( n25053 , n25050 , n345085 );
buf ( n345087 , n606 );
not ( n25055 , n345087 );
buf ( n345089 , n344350 );
not ( n25057 , n345089 );
buf ( n345091 , n25057 );
buf ( n345092 , n345091 );
not ( n345093 , n345092 );
or ( n25061 , n25055 , n345093 );
buf ( n345095 , n345091 );
not ( n345096 , n345095 );
buf ( n345097 , n345096 );
buf ( n345098 , n345097 );
buf ( n345099 , n344445 );
nand ( n25067 , n345098 , n345099 );
buf ( n345101 , n25067 );
buf ( n345102 , n345101 );
nand ( n25070 , n25061 , n345102 );
buf ( n345104 , n25070 );
buf ( n345105 , n345104 );
buf ( n345106 , n344454 );
nand ( n345107 , n345105 , n345106 );
buf ( n345108 , n345107 );
buf ( n345109 , n345108 );
nand ( n25077 , n25053 , n345109 );
buf ( n345111 , n25077 );
buf ( n345112 , n345111 );
not ( n345113 , n345112 );
xor ( n345114 , n344823 , n24817 );
xor ( n25082 , n345114 , n344865 );
buf ( n345116 , n25082 );
not ( n25084 , n345116 );
buf ( n345118 , n25084 );
buf ( n345119 , n345118 );
not ( n25087 , n345119 );
or ( n345121 , n345113 , n25087 );
buf ( n345122 , n345118 );
buf ( n345123 , n345111 );
or ( n25091 , n345122 , n345123 );
buf ( n345125 , n607 );
not ( n25093 , n345125 );
buf ( n345127 , n345104 );
not ( n25095 , n345127 );
or ( n25096 , n25093 , n25095 );
buf ( n345130 , n344454 );
buf ( n345131 , n606 );
not ( n345132 , n345131 );
buf ( n345133 , n344383 );
not ( n25101 , n345133 );
or ( n345135 , n345132 , n25101 );
buf ( n345136 , n24346 );
buf ( n345137 , n344445 );
nand ( n25105 , n345136 , n345137 );
buf ( n345139 , n25105 );
buf ( n345140 , n345139 );
nand ( n345141 , n345135 , n345140 );
buf ( n345142 , n345141 );
buf ( n345143 , n345142 );
nand ( n345144 , n345130 , n345143 );
buf ( n345145 , n345144 );
buf ( n345146 , n345145 );
nand ( n345147 , n25096 , n345146 );
buf ( n345148 , n345147 );
buf ( n345149 , n345148 );
not ( n25117 , n345149 );
not ( n25118 , n23613 );
not ( n345152 , n24126 );
or ( n345153 , n25118 , n345152 );
and ( n345154 , n24108 , n592 );
not ( n25122 , n24108 );
and ( n345156 , n25122 , n343624 );
nor ( n25124 , n345154 , n345156 );
buf ( n345158 , n25124 );
buf ( n345159 , n343699 );
nand ( n345160 , n345158 , n345159 );
buf ( n345161 , n345160 );
nand ( n345162 , n345153 , n345161 );
buf ( n345163 , n345162 );
not ( n25131 , n345163 );
nand ( n25132 , n334490 , n14535 );
not ( n25133 , n25132 );
not ( n25134 , n334482 );
not ( n25135 , n14613 );
nand ( n25136 , n25134 , n25135 );
not ( n25137 , n25136 );
or ( n25138 , n25133 , n25137 );
nand ( n25139 , n14535 , n25134 , n25135 , n334490 );
nand ( n25140 , n25138 , n25139 );
not ( n25141 , n25140 );
buf ( n345175 , n25141 );
not ( n345176 , n345175 );
nand ( n25144 , n345176 , n592 );
buf ( n345178 , n25144 );
nand ( n345179 , n25131 , n345178 );
buf ( n345180 , n345179 );
buf ( n345181 , n345180 );
not ( n25149 , n345181 );
buf ( n345183 , n23681 );
not ( n25151 , n345183 );
buf ( n345185 , n344189 );
not ( n25153 , n345185 );
or ( n25154 , n25151 , n25153 );
buf ( n345188 , n594 );
not ( n25156 , n345188 );
buf ( n345190 , n24059 );
not ( n25158 , n345190 );
or ( n25159 , n25156 , n25158 );
nand ( n25160 , n23605 , n343632 );
buf ( n345194 , n25160 );
nand ( n25162 , n25159 , n345194 );
buf ( n345196 , n25162 );
buf ( n345197 , n345196 );
buf ( n345198 , n343762 );
nand ( n345199 , n345197 , n345198 );
buf ( n345200 , n345199 );
buf ( n345201 , n345200 );
nand ( n345202 , n25154 , n345201 );
buf ( n345203 , n345202 );
buf ( n345204 , n345203 );
not ( n345205 , n345204 );
or ( n25173 , n25149 , n345205 );
buf ( n345207 , n25144 );
not ( n25175 , n345207 );
buf ( n345209 , n345162 );
nand ( n25177 , n25175 , n345209 );
buf ( n345211 , n25177 );
buf ( n345212 , n345211 );
nand ( n25180 , n25173 , n345212 );
buf ( n345214 , n25180 );
buf ( n345215 , n345214 );
not ( n25183 , n344196 );
not ( n25184 , n344148 );
not ( n345218 , n344164 );
or ( n25186 , n25184 , n345218 );
or ( n25187 , n344164 , n344148 );
nand ( n25188 , n25186 , n25187 );
not ( n345222 , n25188 );
or ( n345223 , n25183 , n345222 );
or ( n345224 , n344196 , n25188 );
nand ( n25192 , n345223 , n345224 );
buf ( n345226 , n25192 );
xor ( n25194 , n345215 , n345226 );
buf ( n345228 , n343863 );
not ( n345229 , n345228 );
buf ( n345230 , n345009 );
not ( n25198 , n345230 );
or ( n345232 , n345229 , n25198 );
and ( n345233 , n334588 , n343882 );
not ( n25201 , n334588 );
and ( n345235 , n25201 , n596 );
or ( n345236 , n345233 , n345235 );
buf ( n345237 , n345236 );
buf ( n345238 , n23889 );
nand ( n345239 , n345237 , n345238 );
buf ( n345240 , n345239 );
buf ( n345241 , n345240 );
nand ( n345242 , n345232 , n345241 );
buf ( n345243 , n345242 );
buf ( n345244 , n345243 );
and ( n345245 , n25194 , n345244 );
and ( n25213 , n345215 , n345226 );
or ( n345247 , n345245 , n25213 );
buf ( n345248 , n345247 );
buf ( n345249 , n345248 );
buf ( n345250 , n23911 );
not ( n345251 , n345250 );
buf ( n345252 , n344964 );
not ( n345253 , n345252 );
or ( n25221 , n345251 , n345253 );
buf ( n345255 , n598 );
not ( n345256 , n345255 );
buf ( n345257 , n343911 );
not ( n345258 , n345257 );
or ( n25226 , n345256 , n345258 );
buf ( n345260 , n343908 );
buf ( n345261 , n343953 );
nand ( n345262 , n345260 , n345261 );
buf ( n345263 , n345262 );
buf ( n345264 , n345263 );
nand ( n25232 , n25226 , n345264 );
buf ( n345266 , n25232 );
buf ( n25234 , n345266 );
buf ( n25235 , n343948 );
nand ( n25236 , n25234 , n25235 );
buf ( n345270 , n25236 );
buf ( n345271 , n345270 );
nand ( n25239 , n25221 , n345271 );
buf ( n345273 , n25239 );
buf ( n345274 , n345273 );
xor ( n345275 , n345249 , n345274 );
not ( n345276 , n344018 );
not ( n345277 , n600 );
not ( n345278 , n343962 );
or ( n25246 , n345277 , n345278 );
nand ( n345280 , n23906 , n343966 );
nand ( n345281 , n25246 , n345280 );
not ( n25249 , n345281 );
or ( n345283 , n345276 , n25249 );
not ( n345284 , n24901 );
not ( n25252 , n344939 );
or ( n25253 , n345284 , n25252 );
nand ( n345287 , n25253 , n344015 );
nand ( n25255 , n345283 , n345287 );
buf ( n345289 , n25255 );
and ( n345290 , n345275 , n345289 );
and ( n345291 , n345249 , n345274 );
or ( n25259 , n345290 , n345291 );
buf ( n345293 , n25259 );
buf ( n345294 , n345293 );
not ( n345295 , n345294 );
or ( n345296 , n25117 , n345295 );
buf ( n345297 , n345148 );
not ( n25265 , n345297 );
buf ( n345299 , n25265 );
buf ( n345300 , n345299 );
not ( n25268 , n345300 );
buf ( n345302 , n345293 );
not ( n25270 , n345302 );
buf ( n345304 , n25270 );
buf ( n345305 , n345304 );
not ( n25273 , n345305 );
or ( n25274 , n25268 , n25273 );
xor ( n345308 , n344992 , n345017 );
xor ( n25276 , n345308 , n345028 );
buf ( n345310 , n25276 );
buf ( n25278 , n345310 );
not ( n345312 , n25278 );
buf ( n345313 , n344400 );
not ( n345314 , n345313 );
buf ( n345315 , n604 );
not ( n25283 , n345315 );
buf ( n345317 , n344308 );
not ( n345318 , n345317 );
or ( n25286 , n25283 , n345318 );
buf ( n345320 , n24265 );
buf ( n345321 , n345320 );
buf ( n345322 , n345321 );
buf ( n345323 , n345322 );
buf ( n345324 , n23530 );
nand ( n25292 , n345323 , n345324 );
buf ( n25293 , n25292 );
buf ( n345327 , n25293 );
nand ( n25295 , n25286 , n345327 );
buf ( n345329 , n25295 );
buf ( n345330 , n345329 );
not ( n345331 , n345330 );
or ( n25299 , n345314 , n345331 );
buf ( n345333 , n344883 );
buf ( n345334 , n344338 );
nand ( n25302 , n345333 , n345334 );
buf ( n25303 , n25302 );
buf ( n345337 , n25303 );
nand ( n25305 , n25299 , n345337 );
buf ( n25306 , n25305 );
not ( n25307 , n25306 );
or ( n25308 , n345312 , n25307 );
or ( n25309 , n25306 , n25278 );
buf ( n345343 , n343531 );
not ( n345344 , n345343 );
buf ( n345345 , n344906 );
not ( n345346 , n345345 );
or ( n25314 , n345344 , n345346 );
buf ( n345348 , n602 );
not ( n345349 , n345348 );
buf ( n345350 , n23996 );
not ( n345351 , n345350 );
or ( n345352 , n345349 , n345351 );
buf ( n345353 , n344035 );
buf ( n345354 , n343553 );
nand ( n25322 , n345353 , n345354 );
buf ( n345356 , n25322 );
buf ( n345357 , n345356 );
nand ( n25325 , n345352 , n345357 );
buf ( n345359 , n25325 );
buf ( n345360 , n345359 );
buf ( n345361 , n343595 );
nand ( n25329 , n345360 , n345361 );
buf ( n345363 , n25329 );
buf ( n345364 , n345363 );
nand ( n25332 , n25314 , n345364 );
buf ( n345366 , n25332 );
nand ( n25334 , n25309 , n345366 );
nand ( n25335 , n25308 , n25334 );
buf ( n345369 , n25335 );
nand ( n25337 , n25274 , n345369 );
buf ( n345371 , n25337 );
buf ( n345372 , n345371 );
nand ( n345373 , n345296 , n345372 );
buf ( n345374 , n345373 );
buf ( n345375 , n345374 );
nand ( n345376 , n25091 , n345375 );
buf ( n345377 , n345376 );
buf ( n345378 , n345377 );
nand ( n345379 , n345121 , n345378 );
buf ( n345380 , n345379 );
buf ( n345381 , n345380 );
xor ( n25349 , n345081 , n345381 );
buf ( n25350 , n344871 );
buf ( n25351 , n344876 );
xor ( n25352 , n25350 , n25351 );
buf ( n345386 , n25018 );
xor ( n345387 , n25352 , n345386 );
buf ( n345388 , n345387 );
buf ( n345389 , n345388 );
and ( n345390 , n25349 , n345389 );
and ( n345391 , n345081 , n345381 );
or ( n25359 , n345390 , n345391 );
buf ( n345393 , n25359 );
buf ( n345394 , n345393 );
not ( n345395 , n345394 );
buf ( n345396 , n345395 );
nand ( n345397 , n25034 , n345396 );
not ( n25365 , n345397 );
xor ( n345399 , n25003 , n25014 );
xnor ( n25367 , n345399 , n344927 );
buf ( n345401 , n25367 );
not ( n25369 , n345401 );
buf ( n345403 , n25369 );
not ( n25371 , n345403 );
buf ( n345405 , n23911 );
not ( n345406 , n345405 );
buf ( n345407 , n345266 );
not ( n345408 , n345407 );
or ( n25376 , n345406 , n345408 );
buf ( n345410 , n598 );
not ( n25378 , n345410 );
buf ( n345412 , n344230 );
not ( n345413 , n345412 );
or ( n25381 , n25378 , n345413 );
buf ( n345415 , n23795 );
buf ( n345416 , n343953 );
nand ( n25384 , n345415 , n345416 );
buf ( n25385 , n25384 );
buf ( n345419 , n25385 );
nand ( n25387 , n25381 , n345419 );
buf ( n345421 , n25387 );
buf ( n345422 , n345421 );
buf ( n345423 , n343945 );
nand ( n345424 , n345422 , n345423 );
buf ( n345425 , n345424 );
buf ( n345426 , n345425 );
nand ( n345427 , n25376 , n345426 );
buf ( n345428 , n345427 );
buf ( n345429 , n345428 );
nand ( n25397 , n25124 , n23613 );
buf ( n345431 , n592 );
not ( n25399 , n345431 );
buf ( n345433 , n25141 );
not ( n25401 , n345433 );
or ( n25402 , n25399 , n25401 );
not ( n25403 , n25141 );
buf ( n345437 , n25403 );
buf ( n345438 , n343624 );
nand ( n25406 , n345437 , n345438 );
buf ( n345440 , n25406 );
buf ( n345441 , n345440 );
nand ( n345442 , n25402 , n345441 );
buf ( n345443 , n345442 );
nand ( n345444 , n345443 , n343699 );
buf ( n345445 , n592 );
not ( n345446 , n14734 );
not ( n345447 , n345446 );
not ( n345448 , n334590 );
not ( n25416 , n345448 );
or ( n345450 , n345447 , n25416 );
nand ( n345451 , n345450 , n14735 );
buf ( n345452 , n345451 );
not ( n345453 , n345452 );
buf ( n345454 , n345453 );
buf ( n25422 , n345454 );
not ( n25423 , n25422 );
buf ( n25424 , n25423 );
buf ( n25425 , n25424 );
and ( n25426 , n345445 , n25425 );
buf ( n345460 , n25426 );
not ( n345461 , n345460 );
nand ( n25429 , n25397 , n345444 , n345461 );
buf ( n345463 , n25429 );
not ( n345464 , n345463 );
buf ( n345465 , n23681 );
not ( n25433 , n345465 );
buf ( n345467 , n345196 );
not ( n25435 , n345467 );
or ( n345469 , n25433 , n25435 );
buf ( n345470 , n594 );
not ( n25438 , n345470 );
buf ( n345472 , n24091 );
not ( n25440 , n345472 );
or ( n345474 , n25438 , n25440 );
buf ( n345475 , n343632 );
buf ( n345476 , n344155 );
nand ( n345477 , n345475 , n345476 );
buf ( n345478 , n345477 );
buf ( n345479 , n345478 );
nand ( n25447 , n345474 , n345479 );
buf ( n345481 , n25447 );
buf ( n25449 , n345481 );
buf ( n345483 , n343762 );
nand ( n345484 , n25449 , n345483 );
buf ( n345485 , n345484 );
buf ( n345486 , n345485 );
nand ( n25454 , n345469 , n345486 );
buf ( n25455 , n25454 );
buf ( n345489 , n25455 );
not ( n25457 , n345489 );
or ( n345491 , n345464 , n25457 );
not ( n25459 , n23613 );
not ( n345493 , n25124 );
or ( n345494 , n25459 , n345493 );
nand ( n25462 , n345494 , n345444 );
nand ( n345496 , n25462 , n345460 );
buf ( n345497 , n345496 );
nand ( n345498 , n345491 , n345497 );
buf ( n345499 , n345498 );
buf ( n345500 , n345499 );
not ( n345501 , n345500 );
buf ( n345502 , n345501 );
buf ( n345503 , n345502 );
not ( n345504 , n345503 );
buf ( n345505 , n343863 );
not ( n345506 , n345505 );
buf ( n345507 , n345236 );
not ( n25475 , n345507 );
or ( n345509 , n345506 , n25475 );
buf ( n345510 , n23889 );
and ( n345511 , n343650 , n343882 );
not ( n25479 , n343650 );
and ( n25480 , n25479 , n596 );
or ( n345514 , n345511 , n25480 );
buf ( n345515 , n345514 );
nand ( n345516 , n345510 , n345515 );
buf ( n345517 , n345516 );
buf ( n345518 , n345517 );
nand ( n345519 , n345509 , n345518 );
buf ( n345520 , n345519 );
buf ( n345521 , n345520 );
not ( n25489 , n345521 );
buf ( n345523 , n25489 );
buf ( n345524 , n345523 );
not ( n25492 , n345524 );
or ( n25493 , n345504 , n25492 );
buf ( n345527 , n345203 );
not ( n345528 , n345527 );
not ( n345529 , n25144 );
not ( n345530 , n345529 );
not ( n25498 , n345162 );
or ( n345532 , n345530 , n25498 );
or ( n345533 , n345529 , n345162 );
nand ( n25501 , n345532 , n345533 );
buf ( n345535 , n25501 );
not ( n345536 , n345535 );
or ( n25504 , n345528 , n345536 );
buf ( n345538 , n345203 );
buf ( n345539 , n25501 );
or ( n25507 , n345538 , n345539 );
nand ( n345541 , n25504 , n25507 );
buf ( n345542 , n345541 );
buf ( n345543 , n345542 );
nand ( n25511 , n25493 , n345543 );
buf ( n345545 , n25511 );
buf ( n345546 , n345545 );
buf ( n345547 , n345520 );
buf ( n345548 , n345499 );
nand ( n25516 , n345547 , n345548 );
buf ( n345550 , n25516 );
buf ( n345551 , n345550 );
nand ( n345552 , n345546 , n345551 );
buf ( n345553 , n345552 );
buf ( n345554 , n345553 );
xor ( n345555 , n345429 , n345554 );
xor ( n25523 , n345215 , n345226 );
xor ( n345557 , n25523 , n345244 );
buf ( n345558 , n345557 );
buf ( n345559 , n345558 );
and ( n345560 , n345555 , n345559 );
and ( n25528 , n345429 , n345554 );
or ( n25529 , n345560 , n25528 );
buf ( n345563 , n25529 );
buf ( n345564 , n345563 );
buf ( n345565 , n607 );
not ( n25533 , n345565 );
buf ( n345567 , n345142 );
not ( n345568 , n345567 );
or ( n25536 , n25533 , n345568 );
buf ( n345570 , n606 );
not ( n345571 , n345570 );
buf ( n345572 , n343548 );
not ( n25540 , n345572 );
or ( n345574 , n345571 , n25540 );
buf ( n345575 , n343545 );
buf ( n345576 , n344445 );
nand ( n345577 , n345575 , n345576 );
buf ( n345578 , n345577 );
buf ( n345579 , n345578 );
nand ( n25547 , n345574 , n345579 );
buf ( n345581 , n25547 );
buf ( n345582 , n345581 );
buf ( n345583 , n344454 );
nand ( n345584 , n345582 , n345583 );
buf ( n345585 , n345584 );
buf ( n345586 , n345585 );
nand ( n345587 , n25536 , n345586 );
buf ( n345588 , n345587 );
buf ( n345589 , n345588 );
xor ( n25557 , n345564 , n345589 );
xor ( n345591 , n345249 , n345274 );
xor ( n345592 , n345591 , n345289 );
buf ( n345593 , n345592 );
buf ( n345594 , n345593 );
and ( n345595 , n25557 , n345594 );
and ( n25563 , n345564 , n345589 );
or ( n345597 , n345595 , n25563 );
buf ( n345598 , n345597 );
not ( n25566 , n345598 );
buf ( n345600 , n345032 );
buf ( n345601 , n24933 );
xor ( n345602 , n345600 , n345601 );
buf ( n345603 , n24912 );
xnor ( n345604 , n345602 , n345603 );
buf ( n345605 , n345604 );
nor ( n25573 , n25566 , n345605 );
not ( n345607 , n25573 );
buf ( n345608 , n345605 );
not ( n25576 , n345608 );
buf ( n345610 , n345598 );
not ( n345611 , n345610 );
buf ( n345612 , n345611 );
buf ( n345613 , n345612 );
not ( n345614 , n345613 );
or ( n345615 , n25576 , n345614 );
buf ( n345616 , n344925 );
buf ( n345617 , n24855 );
xor ( n345618 , n345616 , n345617 );
buf ( n345619 , n344920 );
xnor ( n25587 , n345618 , n345619 );
buf ( n345621 , n25587 );
buf ( n345622 , n345621 );
nand ( n345623 , n345615 , n345622 );
buf ( n345624 , n345623 );
nand ( n25592 , n345607 , n345624 );
not ( n25593 , n25592 );
not ( n345627 , n25593 );
or ( n345628 , n25371 , n345627 );
nand ( n25596 , n25592 , n25367 );
nand ( n25597 , n345628 , n25596 );
buf ( n345631 , n345111 );
buf ( n345632 , n25082 );
xor ( n345633 , n345631 , n345632 );
buf ( n345634 , n345374 );
xor ( n25602 , n345633 , n345634 );
buf ( n345636 , n25602 );
buf ( n345637 , n345636 );
not ( n345638 , n345637 );
buf ( n345639 , n345638 );
and ( n25607 , n25597 , n345639 );
not ( n25608 , n25597 );
and ( n345642 , n25608 , n345636 );
nor ( n345643 , n25607 , n345642 );
buf ( n345644 , n345643 );
not ( n25612 , n25335 );
and ( n25613 , n345293 , n345148 );
not ( n345647 , n345293 );
and ( n345648 , n345647 , n345299 );
nor ( n25616 , n25613 , n345648 );
not ( n25617 , n25616 );
not ( n25618 , n25617 );
or ( n345652 , n25612 , n25618 );
not ( n345653 , n25335 );
nand ( n25621 , n345653 , n25616 );
nand ( n25622 , n345652 , n25621 );
buf ( n345656 , n25622 );
not ( n345657 , n345656 );
buf ( n345658 , n345514 );
buf ( n345659 , n343863 );
and ( n25627 , n345658 , n345659 );
buf ( n345661 , n23889 );
not ( n345662 , n345661 );
buf ( n345663 , n344185 );
not ( n25631 , n345663 );
buf ( n345665 , n343882 );
not ( n25633 , n345665 );
and ( n345667 , n25631 , n25633 );
buf ( n345668 , n343675 );
buf ( n345669 , n343882 );
and ( n25637 , n345668 , n345669 );
nor ( n25638 , n345667 , n25637 );
buf ( n345672 , n25638 );
buf ( n345673 , n345672 );
nor ( n25641 , n345662 , n345673 );
buf ( n345675 , n25641 );
buf ( n345676 , n345675 );
nor ( n345677 , n25627 , n345676 );
buf ( n345678 , n345677 );
buf ( n25646 , n345678 );
buf ( n345680 , n23613 );
not ( n345681 , n345680 );
buf ( n345682 , n345443 );
not ( n25650 , n345682 );
or ( n25651 , n345681 , n25650 );
xor ( n25652 , n345445 , n25425 );
buf ( n345686 , n25652 );
buf ( n25654 , n345686 );
buf ( n345688 , n343699 );
nand ( n345689 , n25654 , n345688 );
buf ( n345690 , n345689 );
buf ( n345691 , n345690 );
nand ( n345692 , n25651 , n345691 );
buf ( n345693 , n345692 );
buf ( n345694 , n345693 );
not ( n345695 , n345694 );
buf ( n345696 , n14776 );
not ( n25664 , n345696 );
buf ( n25665 , n25664 );
buf ( n345699 , n25665 );
not ( n25667 , n345699 );
buf ( n25668 , n25667 );
buf ( n25669 , n25668 );
buf ( n345703 , n592 );
nand ( n25671 , n25669 , n345703 );
buf ( n345705 , n25671 );
buf ( n345706 , n345705 );
nand ( n25674 , n345695 , n345706 );
buf ( n345708 , n25674 );
buf ( n345709 , n345708 );
not ( n345710 , n345709 );
buf ( n345711 , n23681 );
not ( n25679 , n345711 );
buf ( n345713 , n345481 );
not ( n345714 , n345713 );
or ( n345715 , n25679 , n345714 );
buf ( n345716 , n594 );
not ( n25684 , n345716 );
buf ( n345718 , n24109 );
not ( n345719 , n345718 );
or ( n25687 , n25684 , n345719 );
buf ( n345721 , n24108 );
buf ( n345722 , n343632 );
nand ( n25690 , n345721 , n345722 );
buf ( n25691 , n25690 );
buf ( n345725 , n25691 );
nand ( n345726 , n25687 , n345725 );
buf ( n345727 , n345726 );
buf ( n345728 , n345727 );
buf ( n345729 , n343762 );
nand ( n25697 , n345728 , n345729 );
buf ( n345731 , n25697 );
buf ( n345732 , n345731 );
nand ( n345733 , n345715 , n345732 );
buf ( n345734 , n345733 );
buf ( n345735 , n345734 );
not ( n345736 , n345735 );
or ( n25704 , n345710 , n345736 );
buf ( n345738 , n345705 );
not ( n25706 , n345738 );
buf ( n345740 , n345693 );
nand ( n25708 , n25706 , n345740 );
buf ( n25709 , n25708 );
buf ( n345743 , n25709 );
nand ( n25711 , n25704 , n345743 );
buf ( n345745 , n25711 );
buf ( n345746 , n345745 );
not ( n25714 , n345746 );
buf ( n345748 , n25714 );
buf ( n345749 , n345748 );
nand ( n25717 , n25646 , n345749 );
buf ( n345751 , n25717 );
buf ( n345752 , n345751 );
not ( n25720 , n345752 );
xor ( n345754 , n345461 , n25462 );
buf ( n25722 , n25455 );
xnor ( n25723 , n345754 , n25722 );
buf ( n345757 , n25723 );
not ( n25725 , n345757 );
or ( n25726 , n25720 , n25725 );
buf ( n345760 , n345678 );
not ( n25728 , n345760 );
buf ( n345762 , n345745 );
nand ( n345763 , n25728 , n345762 );
buf ( n345764 , n345763 );
buf ( n345765 , n345764 );
nand ( n345766 , n25726 , n345765 );
buf ( n345767 , n345766 );
buf ( n345768 , n345767 );
buf ( n345769 , n23911 );
not ( n25737 , n345769 );
buf ( n345771 , n345421 );
not ( n345772 , n345771 );
or ( n25740 , n25737 , n345772 );
buf ( n345774 , n598 );
not ( n345775 , n345774 );
buf ( n345776 , n23694 );
not ( n25744 , n345776 );
or ( n345778 , n345775 , n25744 );
buf ( n345779 , n343953 );
buf ( n345780 , n343723 );
nand ( n345781 , n345779 , n345780 );
buf ( n345782 , n345781 );
buf ( n345783 , n345782 );
nand ( n345784 , n345778 , n345783 );
buf ( n345785 , n345784 );
buf ( n345786 , n345785 );
buf ( n345787 , n343945 );
nand ( n25755 , n345786 , n345787 );
buf ( n345789 , n25755 );
buf ( n345790 , n345789 );
nand ( n25758 , n25740 , n345790 );
buf ( n25759 , n25758 );
buf ( n345793 , n25759 );
xor ( n25761 , n345768 , n345793 );
xor ( n25762 , n345502 , n345542 );
xnor ( n25763 , n25762 , n345520 );
buf ( n345797 , n25763 );
and ( n345798 , n25761 , n345797 );
and ( n345799 , n345768 , n345793 );
or ( n345800 , n345798 , n345799 );
buf ( n345801 , n345800 );
buf ( n345802 , n345801 );
buf ( n345803 , n344015 );
not ( n25771 , n345803 );
buf ( n345805 , n345281 );
not ( n345806 , n345805 );
or ( n345807 , n25771 , n345806 );
buf ( n345808 , n600 );
not ( n345809 , n345808 );
buf ( n345810 , n343872 );
not ( n345811 , n345810 );
or ( n345812 , n345809 , n345811 );
buf ( n345813 , n343869 );
buf ( n345814 , n23906 );
nand ( n25782 , n345813 , n345814 );
buf ( n345816 , n25782 );
buf ( n345817 , n345816 );
nand ( n25785 , n345812 , n345817 );
buf ( n345819 , n25785 );
buf ( n345820 , n345819 );
buf ( n345821 , n344018 );
nand ( n345822 , n345820 , n345821 );
buf ( n345823 , n345822 );
buf ( n345824 , n345823 );
nand ( n345825 , n345807 , n345824 );
buf ( n345826 , n345825 );
buf ( n345827 , n345826 );
xor ( n345828 , n345802 , n345827 );
buf ( n345829 , n343531 );
not ( n345830 , n345829 );
buf ( n345831 , n345359 );
not ( n25799 , n345831 );
or ( n345833 , n345830 , n25799 );
and ( n345834 , n343982 , n343553 );
not ( n25802 , n343982 );
and ( n345836 , n25802 , n602 );
or ( n345837 , n345834 , n345836 );
buf ( n345838 , n345837 );
buf ( n345839 , n343595 );
nand ( n345840 , n345838 , n345839 );
buf ( n345841 , n345840 );
buf ( n345842 , n345841 );
nand ( n345843 , n345833 , n345842 );
buf ( n345844 , n345843 );
buf ( n345845 , n345844 );
and ( n25813 , n345828 , n345845 );
and ( n25814 , n345802 , n345827 );
or ( n345848 , n25813 , n25814 );
buf ( n345849 , n345848 );
not ( n345850 , n345849 );
buf ( n345851 , n345850 );
not ( n25819 , n345851 );
buf ( n345853 , n345310 );
buf ( n25821 , n25306 );
xor ( n25822 , n345853 , n25821 );
buf ( n345856 , n345366 );
xnor ( n25824 , n25822 , n345856 );
buf ( n345858 , n25824 );
buf ( n345859 , n345858 );
not ( n345860 , n345859 );
or ( n345861 , n25819 , n345860 );
buf ( n345862 , n344338 );
not ( n345863 , n345862 );
buf ( n345864 , n345329 );
not ( n345865 , n345864 );
or ( n25833 , n345863 , n345865 );
buf ( n345867 , n604 );
not ( n25835 , n345867 );
buf ( n345869 , n344055 );
not ( n345870 , n345869 );
or ( n345871 , n25835 , n345870 );
buf ( n345872 , n344588 );
buf ( n345873 , n23530 );
nand ( n25841 , n345872 , n345873 );
buf ( n345875 , n25841 );
buf ( n345876 , n345875 );
nand ( n25844 , n345871 , n345876 );
buf ( n345878 , n25844 );
buf ( n345879 , n345878 );
buf ( n345880 , n344400 );
nand ( n345881 , n345879 , n345880 );
buf ( n345882 , n345881 );
buf ( n345883 , n345882 );
nand ( n25851 , n25833 , n345883 );
buf ( n345885 , n25851 );
buf ( n345886 , n345885 );
not ( n25854 , n345886 );
buf ( n345888 , n25854 );
buf ( n345889 , n345888 );
not ( n25857 , n345889 );
and ( n345891 , n14695 , n344445 );
not ( n345892 , n14695 );
and ( n345893 , n345892 , n606 );
or ( n25861 , n345891 , n345893 );
buf ( n345895 , n25861 );
not ( n345896 , n345895 );
buf ( n345897 , n345896 );
buf ( n345898 , n345897 );
not ( n345899 , n345898 );
buf ( n345900 , n344631 );
not ( n345901 , n345900 );
and ( n25869 , n345899 , n345901 );
buf ( n345903 , n345581 );
buf ( n345904 , n607 );
and ( n345905 , n345903 , n345904 );
nor ( n25873 , n25869 , n345905 );
buf ( n25874 , n25873 );
buf ( n345908 , n25874 );
not ( n345909 , n345908 );
or ( n25877 , n25857 , n345909 );
xor ( n25878 , n345429 , n345554 );
xor ( n345912 , n25878 , n345559 );
buf ( n345913 , n345912 );
buf ( n25881 , n345913 );
buf ( n345915 , n25881 );
nand ( n345916 , n25877 , n345915 );
buf ( n345917 , n345916 );
buf ( n345918 , n345917 );
buf ( n345919 , n25874 );
not ( n25887 , n345919 );
buf ( n345921 , n345885 );
nand ( n345922 , n25887 , n345921 );
buf ( n345923 , n345922 );
buf ( n345924 , n345923 );
nand ( n25892 , n345918 , n345924 );
buf ( n345926 , n25892 );
buf ( n345927 , n345926 );
nand ( n25895 , n345861 , n345927 );
buf ( n345929 , n25895 );
buf ( n345930 , n345858 );
not ( n25898 , n345930 );
buf ( n345932 , n25898 );
buf ( n345933 , n345932 );
not ( n345934 , n345850 );
buf ( n345935 , n345934 );
nand ( n25903 , n345933 , n345935 );
buf ( n345937 , n25903 );
nand ( n25905 , n345929 , n345937 );
not ( n25906 , n25905 );
buf ( n345940 , n25906 );
nand ( n25908 , n345657 , n345940 );
buf ( n345942 , n25908 );
buf ( n345943 , n345942 );
not ( n345944 , n345943 );
buf ( n345945 , n345605 );
buf ( n345946 , n345621 );
xor ( n345947 , n345945 , n345946 );
buf ( n345948 , n345598 );
xnor ( n345949 , n345947 , n345948 );
buf ( n345950 , n345949 );
buf ( n345951 , n345950 );
not ( n25919 , n345951 );
buf ( n345953 , n25919 );
buf ( n345954 , n345953 );
not ( n345955 , n345954 );
buf ( n345956 , n345955 );
buf ( n345957 , n345956 );
not ( n345958 , n345957 );
or ( n345959 , n345944 , n345958 );
buf ( n345960 , n25906 );
not ( n25928 , n345960 );
buf ( n345962 , n25622 );
nand ( n25930 , n25928 , n345962 );
buf ( n345964 , n25930 );
buf ( n345965 , n345964 );
nand ( n25933 , n345959 , n345965 );
buf ( n345967 , n25933 );
buf ( n345968 , n345967 );
nor ( n345969 , n345644 , n345968 );
buf ( n345970 , n345969 );
buf ( n345971 , n345970 );
and ( n345972 , n25622 , n25905 );
not ( n25940 , n25622 );
and ( n25941 , n25940 , n25906 );
nor ( n345975 , n345972 , n25941 );
or ( n25943 , n345953 , n345975 );
buf ( n345977 , n345950 );
not ( n25945 , n345977 );
buf ( n345979 , n25945 );
nand ( n345980 , n345975 , n345979 );
nand ( n345981 , n25943 , n345980 );
buf ( n345982 , n345981 );
buf ( n25950 , n345982 );
buf ( n345984 , n25950 );
buf ( n345985 , n345984 );
buf ( n345986 , n345849 );
buf ( n345987 , n345858 );
xor ( n345988 , n345986 , n345987 );
buf ( n345989 , n345926 );
xnor ( n25957 , n345988 , n345989 );
buf ( n345991 , n25957 );
buf ( n345992 , n345991 );
not ( n345993 , n345992 );
buf ( n345994 , n345993 );
buf ( n345995 , n345994 );
not ( n345996 , n345995 );
xor ( n345997 , n345564 , n345589 );
xor ( n25965 , n345997 , n345594 );
buf ( n345999 , n25965 );
not ( n346000 , n345999 );
not ( n25968 , n346000 );
buf ( n346002 , n25968 );
nand ( n25970 , n345996 , n346002 );
buf ( n346004 , n25970 );
buf ( n346005 , n346004 );
buf ( n346006 , n346000 );
not ( n25974 , n346006 );
buf ( n346008 , n345994 );
not ( n25976 , n346008 );
or ( n346010 , n25974 , n25976 );
xor ( n346011 , n345802 , n345827 );
xor ( n25979 , n346011 , n345845 );
buf ( n346013 , n25979 );
buf ( n346014 , n346013 );
not ( n25982 , n346014 );
not ( n25983 , n607 );
not ( n25984 , n25861 );
or ( n25985 , n25983 , n25984 );
not ( n346019 , n606 );
not ( n346020 , n344301 );
or ( n346021 , n346019 , n346020 );
buf ( n346022 , n345322 );
buf ( n346023 , n344445 );
nand ( n25991 , n346022 , n346023 );
buf ( n346025 , n25991 );
nand ( n25993 , n346021 , n346025 );
nand ( n25994 , n25993 , n344454 );
nand ( n25995 , n25985 , n25994 );
not ( n25996 , n25995 );
not ( n25997 , n344338 );
not ( n346031 , n345878 );
or ( n25999 , n25997 , n346031 );
and ( n26000 , n23993 , n23530 );
not ( n346034 , n23993 );
and ( n26002 , n346034 , n604 );
or ( n26003 , n26000 , n26002 );
buf ( n346037 , n26003 );
buf ( n346038 , n344400 );
nand ( n346039 , n346037 , n346038 );
buf ( n346040 , n346039 );
nand ( n346041 , n25999 , n346040 );
not ( n346042 , n346041 );
xor ( n26010 , n345768 , n345793 );
xor ( n346044 , n26010 , n345797 );
buf ( n346045 , n346044 );
not ( n26013 , n346045 );
nand ( n346047 , n346042 , n26013 );
not ( n346048 , n346047 );
or ( n26016 , n25996 , n346048 );
not ( n346050 , n346042 );
nand ( n26018 , n346050 , n346045 );
nand ( n346052 , n26016 , n26018 );
buf ( n26020 , n346052 );
not ( n26021 , n26020 );
or ( n26022 , n25982 , n26021 );
buf ( n346056 , n346013 );
buf ( n346057 , n346052 );
or ( n346058 , n346056 , n346057 );
buf ( n346059 , n600 );
buf ( n346060 , n343908 );
and ( n346061 , n346059 , n346060 );
not ( n26029 , n346059 );
buf ( n346063 , n343911 );
and ( n346064 , n26029 , n346063 );
or ( n26032 , n346061 , n346064 );
buf ( n26033 , n26032 );
buf ( n346067 , n26033 );
not ( n26035 , n346067 );
buf ( n346069 , n344017 );
not ( n346070 , n346069 );
and ( n26038 , n26035 , n346070 );
buf ( n346072 , n345819 );
buf ( n346073 , n344015 );
and ( n26041 , n346072 , n346073 );
nor ( n346075 , n26038 , n26041 );
buf ( n346076 , n346075 );
buf ( n346077 , n346076 );
not ( n346078 , n346077 );
and ( n26046 , n345837 , n343531 );
buf ( n346080 , n602 );
buf ( n346081 , n343962 );
and ( n26049 , n346080 , n346081 );
not ( n26050 , n346080 );
buf ( n346084 , n343966 );
and ( n26052 , n26050 , n346084 );
nor ( n26053 , n26049 , n26052 );
buf ( n346087 , n26053 );
buf ( n346088 , n343595 );
not ( n346089 , n346088 );
buf ( n346090 , n346089 );
nor ( n26058 , n346087 , n346090 );
nor ( n26059 , n26046 , n26058 );
buf ( n346093 , n26059 );
not ( n26061 , n346093 );
or ( n346095 , n346078 , n26061 );
buf ( n346096 , n345678 );
buf ( n346097 , n345748 );
and ( n346098 , n346096 , n346097 );
not ( n346099 , n346096 );
buf ( n346100 , n345745 );
and ( n26068 , n346099 , n346100 );
nor ( n346102 , n346098 , n26068 );
buf ( n346103 , n346102 );
buf ( n346104 , n346103 );
buf ( n346105 , n25723 );
not ( n346106 , n346105 );
buf ( n346107 , n346106 );
buf ( n346108 , n346107 );
and ( n346109 , n346104 , n346108 );
not ( n26077 , n346104 );
buf ( n346111 , n25723 );
and ( n26079 , n26077 , n346111 );
nor ( n26080 , n346109 , n26079 );
buf ( n346114 , n26080 );
buf ( n346115 , n346114 );
not ( n26083 , n346115 );
buf ( n346117 , n345785 );
buf ( n346118 , n23911 );
and ( n346119 , n346117 , n346118 );
buf ( n346120 , n343945 );
not ( n346121 , n346120 );
buf ( n346122 , n598 );
buf ( n346123 , n343738 );
and ( n26091 , n346122 , n346123 );
not ( n346125 , n346122 );
buf ( n346126 , n343744 );
and ( n346127 , n346125 , n346126 );
nor ( n346128 , n26091 , n346127 );
buf ( n346129 , n346128 );
buf ( n346130 , n346129 );
nor ( n346131 , n346121 , n346130 );
buf ( n346132 , n346131 );
buf ( n346133 , n346132 );
nor ( n346134 , n346119 , n346133 );
buf ( n346135 , n346134 );
buf ( n346136 , n346135 );
not ( n26104 , n346136 );
or ( n346138 , n26083 , n26104 );
not ( n346139 , n14740 );
not ( n26107 , n334630 );
or ( n346141 , n346139 , n26107 );
nand ( n346142 , n346141 , n14739 );
buf ( n26110 , n346142 );
buf ( n26111 , n592 );
and ( n26112 , n26110 , n26111 );
buf ( n26113 , n26112 );
buf ( n26114 , n26113 );
buf ( n26115 , n23613 );
not ( n26116 , n26115 );
buf ( n346150 , n345686 );
not ( n26118 , n346150 );
or ( n346152 , n26116 , n26118 );
buf ( n346153 , n592 );
not ( n26121 , n346153 );
buf ( n26122 , n25668 );
not ( n346156 , n26122 );
buf ( n346157 , n346156 );
buf ( n346158 , n346157 );
not ( n346159 , n346158 );
or ( n26127 , n26121 , n346159 );
buf ( n346161 , n25668 );
buf ( n346162 , n343624 );
nand ( n26130 , n346161 , n346162 );
buf ( n346164 , n26130 );
buf ( n346165 , n346164 );
nand ( n26133 , n26127 , n346165 );
buf ( n346167 , n26133 );
buf ( n346168 , n346167 );
buf ( n346169 , n343699 );
nand ( n346170 , n346168 , n346169 );
buf ( n346171 , n346170 );
buf ( n346172 , n346171 );
nand ( n346173 , n346152 , n346172 );
buf ( n346174 , n346173 );
buf ( n346175 , n346174 );
xor ( n346176 , n26114 , n346175 );
buf ( n26144 , n14746 );
buf ( n346178 , n26144 );
buf ( n346179 , n346178 );
buf ( n346180 , n346179 );
buf ( n346181 , n592 );
and ( n26149 , n346180 , n346181 );
buf ( n26150 , n26149 );
buf ( n346184 , n26150 );
buf ( n346185 , n23613 );
not ( n346186 , n346185 );
buf ( n346187 , n346167 );
not ( n346188 , n346187 );
or ( n26156 , n346186 , n346188 );
buf ( n346190 , n592 );
not ( n26158 , n346190 );
not ( n26159 , n346142 );
buf ( n346193 , n26159 );
not ( n346194 , n346193 );
or ( n26162 , n26158 , n346194 );
not ( n346196 , n14740 );
not ( n346197 , n334630 );
or ( n26165 , n346196 , n346197 );
nand ( n346199 , n26165 , n14739 );
buf ( n346200 , n346199 );
not ( n26168 , n346200 );
buf ( n346202 , n26168 );
buf ( n346203 , n346202 );
not ( n26171 , n346203 );
buf ( n346205 , n26171 );
buf ( n346206 , n346205 );
buf ( n346207 , n343624 );
nand ( n26175 , n346206 , n346207 );
buf ( n346209 , n26175 );
buf ( n346210 , n346209 );
nand ( n26178 , n26162 , n346210 );
buf ( n26179 , n26178 );
buf ( n346213 , n26179 );
buf ( n346214 , n343699 );
nand ( n346215 , n346213 , n346214 );
buf ( n346216 , n346215 );
buf ( n346217 , n346216 );
nand ( n26185 , n26156 , n346217 );
buf ( n26186 , n26185 );
buf ( n346220 , n26186 );
xor ( n26188 , n346184 , n346220 );
buf ( n346222 , n23613 );
not ( n346223 , n346222 );
buf ( n346224 , n26179 );
not ( n26192 , n346224 );
or ( n26193 , n346223 , n26192 );
buf ( n346227 , n592 );
not ( n346228 , n346227 );
buf ( n346229 , n346179 );
not ( n26197 , n346229 );
buf ( n346231 , n26197 );
buf ( n346232 , n346231 );
not ( n346233 , n346232 );
or ( n346234 , n346228 , n346233 );
buf ( n346235 , n346179 );
buf ( n346236 , n343624 );
nand ( n346237 , n346235 , n346236 );
buf ( n346238 , n346237 );
buf ( n346239 , n346238 );
nand ( n26207 , n346234 , n346239 );
buf ( n346241 , n26207 );
buf ( n26209 , n346241 );
buf ( n26210 , n343699 );
nand ( n26211 , n26209 , n26210 );
buf ( n26212 , n26211 );
buf ( n26213 , n26212 );
nand ( n26214 , n26193 , n26213 );
buf ( n26215 , n26214 );
not ( n346249 , n26215 );
buf ( n346250 , n592 );
not ( n26218 , n346250 );
buf ( n26219 , n14749 );
not ( n346253 , n26219 );
buf ( n346254 , n346253 );
buf ( n346255 , n346254 );
nor ( n346256 , n26218 , n346255 );
buf ( n346257 , n346256 );
not ( n346258 , n346257 );
or ( n346259 , n346249 , n346258 );
buf ( n346260 , n26215 );
buf ( n346261 , n346257 );
nor ( n26229 , n346260 , n346261 );
buf ( n346263 , n26229 );
buf ( n346264 , n592 );
xnor ( n26232 , n14599 , n591 );
not ( n26233 , n26232 );
buf ( n346267 , n26233 );
and ( n26235 , n346264 , n346267 );
buf ( n346269 , n26235 );
buf ( n26237 , n346269 );
buf ( n346271 , n23613 );
not ( n26239 , n346271 );
buf ( n346273 , n592 );
not ( n346274 , n346273 );
buf ( n346275 , n346254 );
not ( n346276 , n346275 );
or ( n346277 , n346274 , n346276 );
buf ( n346278 , n14749 );
buf ( n346279 , n343624 );
nand ( n346280 , n346278 , n346279 );
buf ( n346281 , n346280 );
buf ( n346282 , n346281 );
nand ( n26250 , n346277 , n346282 );
buf ( n346284 , n26250 );
buf ( n346285 , n346284 );
not ( n346286 , n346285 );
or ( n26254 , n26239 , n346286 );
xor ( n26255 , n346264 , n346267 );
buf ( n346289 , n26255 );
buf ( n346290 , n346289 );
buf ( n346291 , n343699 );
nand ( n346292 , n346290 , n346291 );
buf ( n346293 , n346292 );
buf ( n346294 , n346293 );
nand ( n26262 , n26254 , n346294 );
buf ( n346296 , n26262 );
buf ( n346297 , n346296 );
buf ( n346298 , n593 );
buf ( n346299 , n594 );
or ( n26267 , n346298 , n346299 );
buf ( n346301 , n26233 );
nand ( n346302 , n26267 , n346301 );
buf ( n346303 , n346302 );
buf ( n346304 , n346303 );
buf ( n346305 , n593 );
buf ( n346306 , n594 );
and ( n346307 , n346305 , n346306 );
buf ( n346308 , n343624 );
nor ( n346309 , n346307 , n346308 );
buf ( n346310 , n346309 );
buf ( n346311 , n346310 );
and ( n346312 , n346304 , n346311 );
buf ( n346313 , n346312 );
buf ( n346314 , n346313 );
and ( n346315 , n346297 , n346314 );
buf ( n346316 , n346315 );
buf ( n346317 , n346316 );
xor ( n346318 , n26237 , n346317 );
buf ( n346319 , n23613 );
not ( n26287 , n346319 );
buf ( n346321 , n346241 );
not ( n346322 , n346321 );
or ( n346323 , n26287 , n346322 );
buf ( n346324 , n346284 );
buf ( n346325 , n343699 );
nand ( n26293 , n346324 , n346325 );
buf ( n346327 , n26293 );
buf ( n346328 , n346327 );
nand ( n26296 , n346323 , n346328 );
buf ( n346330 , n26296 );
buf ( n346331 , n346330 );
and ( n346332 , n346318 , n346331 );
and ( n26300 , n26237 , n346317 );
or ( n26301 , n346332 , n26300 );
buf ( n346335 , n26301 );
buf ( n346336 , n346335 );
not ( n26304 , n346336 );
buf ( n346338 , n26304 );
or ( n346339 , n346263 , n346338 );
nand ( n26307 , n346259 , n346339 );
buf ( n346341 , n26307 );
and ( n346342 , n26188 , n346341 );
and ( n26310 , n346184 , n346220 );
or ( n346344 , n346342 , n26310 );
buf ( n346345 , n346344 );
buf ( n346346 , n346345 );
and ( n26314 , n346176 , n346346 );
and ( n346348 , n26114 , n346175 );
or ( n26316 , n26314 , n346348 );
buf ( n346350 , n26316 );
buf ( n346351 , n346350 );
buf ( n346352 , n343863 );
not ( n26320 , n346352 );
buf ( n346354 , n345672 );
not ( n26322 , n346354 );
buf ( n346356 , n26322 );
buf ( n346357 , n346356 );
not ( n26325 , n346357 );
or ( n26326 , n26320 , n26325 );
buf ( n346360 , n596 );
not ( n346361 , n346360 );
buf ( n346362 , n23605 );
not ( n26330 , n346362 );
buf ( n26331 , n26330 );
buf ( n346365 , n26331 );
not ( n26333 , n346365 );
or ( n346367 , n346361 , n26333 );
buf ( n346368 , n23605 );
buf ( n346369 , n343882 );
nand ( n346370 , n346368 , n346369 );
buf ( n346371 , n346370 );
buf ( n346372 , n346371 );
nand ( n26340 , n346367 , n346372 );
buf ( n346374 , n26340 );
buf ( n346375 , n346374 );
buf ( n346376 , n23889 );
nand ( n346377 , n346375 , n346376 );
buf ( n346378 , n346377 );
buf ( n346379 , n346378 );
nand ( n346380 , n26326 , n346379 );
buf ( n346381 , n346380 );
buf ( n346382 , n346381 );
xor ( n346383 , n346351 , n346382 );
xor ( n26351 , n345693 , n345705 );
xnor ( n346385 , n26351 , n345734 );
buf ( n346386 , n346385 );
and ( n26354 , n346383 , n346386 );
and ( n346388 , n346351 , n346382 );
or ( n346389 , n26354 , n346388 );
buf ( n346390 , n346389 );
buf ( n346391 , n346390 );
nand ( n346392 , n346138 , n346391 );
buf ( n346393 , n346392 );
buf ( n346394 , n346135 );
not ( n346395 , n346394 );
not ( n26363 , n346114 );
buf ( n346397 , n26363 );
nand ( n346398 , n346395 , n346397 );
buf ( n346399 , n346398 );
nand ( n26367 , n346393 , n346399 );
buf ( n346401 , n26367 );
nand ( n346402 , n346095 , n346401 );
buf ( n346403 , n346402 );
buf ( n346404 , n346403 );
buf ( n346405 , n346076 );
not ( n26373 , n346405 );
buf ( n26374 , n26059 );
not ( n346408 , n26374 );
buf ( n346409 , n346408 );
buf ( n346410 , n346409 );
nand ( n26378 , n26373 , n346410 );
buf ( n346412 , n26378 );
buf ( n26380 , n346412 );
nand ( n26381 , n346404 , n26380 );
buf ( n26382 , n26381 );
buf ( n346416 , n26382 );
nand ( n346417 , n346058 , n346416 );
buf ( n346418 , n346417 );
buf ( n346419 , n346418 );
nand ( n26387 , n26022 , n346419 );
buf ( n346421 , n26387 );
buf ( n346422 , n346421 );
nand ( n26390 , n346010 , n346422 );
buf ( n346424 , n26390 );
buf ( n346425 , n346424 );
nand ( n26393 , n346005 , n346425 );
buf ( n346427 , n26393 );
buf ( n346428 , n346427 );
nor ( n26396 , n345985 , n346428 );
buf ( n346430 , n26396 );
buf ( n346431 , n346430 );
nor ( n346432 , n345971 , n346431 );
buf ( n346433 , n346432 );
not ( n26401 , n346433 );
xor ( n26402 , n345999 , n346421 );
xnor ( n26403 , n26402 , n345991 );
not ( n26404 , n26382 );
not ( n26405 , n346052 );
xor ( n346439 , n26404 , n26405 );
xnor ( n346440 , n346439 , n346013 );
not ( n26408 , n346440 );
not ( n26409 , n345885 );
not ( n26410 , n345913 );
not ( n26411 , n26410 );
or ( n346445 , n26409 , n26411 );
nand ( n26413 , n345888 , n345913 );
nand ( n346447 , n346445 , n26413 );
and ( n26415 , n346447 , n25874 );
not ( n26416 , n346447 );
not ( n26417 , n25874 );
and ( n26418 , n26416 , n26417 );
nor ( n26419 , n26415 , n26418 );
buf ( n26420 , n26419 );
not ( n26421 , n26420 );
and ( n26422 , n26408 , n26421 );
xor ( n26423 , n26404 , n346013 );
xnor ( n346457 , n26423 , n26405 );
nand ( n26425 , n346457 , n26419 );
buf ( n346459 , n344015 );
not ( n26427 , n346459 );
buf ( n346461 , n26033 );
not ( n26429 , n346461 );
buf ( n346463 , n26429 );
buf ( n346464 , n346463 );
not ( n346465 , n346464 );
or ( n26433 , n26427 , n346465 );
buf ( n346467 , n600 );
not ( n346468 , n346467 );
buf ( n346469 , n23798 );
not ( n26437 , n346469 );
or ( n346471 , n346468 , n26437 );
buf ( n346472 , n343837 );
buf ( n346473 , n23906 );
nand ( n346474 , n346472 , n346473 );
buf ( n346475 , n346474 );
buf ( n346476 , n346475 );
nand ( n26444 , n346471 , n346476 );
buf ( n26445 , n26444 );
buf ( n346479 , n26445 );
buf ( n346480 , n344018 );
nand ( n26448 , n346479 , n346480 );
buf ( n346482 , n26448 );
buf ( n346483 , n346482 );
nand ( n26451 , n26433 , n346483 );
buf ( n346485 , n26451 );
buf ( n346486 , n346485 );
not ( n26454 , n346486 );
buf ( n346488 , n598 );
not ( n346489 , n346488 );
buf ( n346490 , n343651 );
not ( n346491 , n346490 );
or ( n346492 , n346489 , n346491 );
not ( n346493 , n343651 );
buf ( n346494 , n346493 );
buf ( n346495 , n343953 );
nand ( n26463 , n346494 , n346495 );
buf ( n346497 , n26463 );
buf ( n346498 , n346497 );
nand ( n26466 , n346492 , n346498 );
buf ( n346500 , n26466 );
not ( n346501 , n346500 );
not ( n26469 , n343945 );
or ( n346503 , n346501 , n26469 );
not ( n346504 , n346129 );
nand ( n26472 , n346504 , n23911 );
nand ( n346506 , n346503 , n26472 );
not ( n346507 , n346506 );
not ( n26475 , n594 );
not ( n346509 , n345175 );
or ( n26477 , n26475 , n346509 );
buf ( n346511 , n25403 );
buf ( n346512 , n343632 );
nand ( n346513 , n346511 , n346512 );
buf ( n346514 , n346513 );
nand ( n26482 , n26477 , n346514 );
buf ( n346516 , n26482 );
buf ( n346517 , n343762 );
and ( n26485 , n346516 , n346517 );
buf ( n346519 , n345727 );
buf ( n346520 , n23681 );
and ( n26488 , n346519 , n346520 );
nor ( n346522 , n26485 , n26488 );
buf ( n346523 , n346522 );
buf ( n346524 , n346523 );
not ( n26492 , n346524 );
buf ( n346526 , n26492 );
buf ( n346527 , n346526 );
not ( n26495 , n346527 );
buf ( n346529 , n343863 );
not ( n346530 , n346529 );
buf ( n346531 , n346374 );
not ( n26499 , n346531 );
or ( n346533 , n346530 , n26499 );
and ( n346534 , n24091 , n596 );
not ( n26502 , n24091 );
and ( n346536 , n26502 , n343882 );
or ( n346537 , n346534 , n346536 );
buf ( n346538 , n346537 );
buf ( n346539 , n23889 );
nand ( n346540 , n346538 , n346539 );
buf ( n346541 , n346540 );
buf ( n346542 , n346541 );
nand ( n346543 , n346533 , n346542 );
buf ( n346544 , n346543 );
buf ( n346545 , n346544 );
not ( n346546 , n346545 );
or ( n26514 , n26495 , n346546 );
buf ( n346548 , n346544 );
buf ( n346549 , n346526 );
or ( n346550 , n346548 , n346549 );
xor ( n346551 , n26114 , n346175 );
xor ( n346552 , n346551 , n346346 );
buf ( n346553 , n346552 );
buf ( n346554 , n346553 );
nand ( n26522 , n346550 , n346554 );
buf ( n346556 , n26522 );
buf ( n346557 , n346556 );
nand ( n346558 , n26514 , n346557 );
buf ( n346559 , n346558 );
buf ( n346560 , n346559 );
buf ( n346561 , n346560 );
buf ( n346562 , n346561 );
not ( n26530 , n346562 );
or ( n346564 , n346507 , n26530 );
buf ( n346565 , n346506 );
buf ( n346566 , n346562 );
nor ( n346567 , n346565 , n346566 );
buf ( n346568 , n346567 );
xor ( n26536 , n346351 , n346382 );
xor ( n346570 , n26536 , n346386 );
buf ( n346571 , n346570 );
buf ( n346572 , n346571 );
not ( n346573 , n346572 );
buf ( n346574 , n346573 );
or ( n346575 , n346568 , n346574 );
nand ( n26543 , n346564 , n346575 );
buf ( n346577 , n26543 );
not ( n346578 , n346577 );
or ( n26546 , n26454 , n346578 );
buf ( n346580 , n346463 );
buf ( n346581 , n344015 );
and ( n26549 , n346580 , n346581 );
buf ( n346583 , n26445 );
not ( n346584 , n346583 );
buf ( n346585 , n344017 );
nor ( n26553 , n346584 , n346585 );
buf ( n346587 , n26553 );
buf ( n346588 , n346587 );
nor ( n26556 , n26549 , n346588 );
buf ( n346590 , n26556 );
buf ( n346591 , n346590 );
not ( n346592 , n346591 );
buf ( n346593 , n26543 );
not ( n26561 , n346593 );
buf ( n346595 , n26561 );
buf ( n346596 , n346595 );
not ( n26564 , n346596 );
or ( n346598 , n346592 , n26564 );
not ( n346599 , n346135 );
xor ( n26567 , n346390 , n346599 );
not ( n346601 , n26363 );
xnor ( n346602 , n26567 , n346601 );
buf ( n346603 , n346602 );
nand ( n26571 , n346598 , n346603 );
buf ( n26572 , n26571 );
buf ( n26573 , n26572 );
nand ( n26574 , n26546 , n26573 );
buf ( n26575 , n26574 );
buf ( n346609 , n26575 );
not ( n26577 , n346609 );
not ( n346611 , n346409 );
not ( n26579 , n346076 );
nand ( n346613 , n346393 , n346399 );
not ( n26581 , n346613 );
or ( n26582 , n26579 , n26581 );
or ( n346616 , n346076 , n26367 );
nand ( n26584 , n26582 , n346616 );
not ( n346618 , n26584 );
or ( n26586 , n346611 , n346618 );
or ( n26587 , n346409 , n26584 );
nand ( n346621 , n26586 , n26587 );
buf ( n346622 , n346621 );
not ( n26590 , n346622 );
buf ( n26591 , n26590 );
not ( n346625 , n26591 );
or ( n26593 , n26577 , n346625 );
buf ( n346627 , n26575 );
not ( n346628 , n346627 );
buf ( n346629 , n346628 );
not ( n26597 , n346629 );
not ( n346631 , n346621 );
or ( n346632 , n26597 , n346631 );
not ( n26600 , n344454 );
buf ( n346634 , n606 );
not ( n346635 , n346634 );
buf ( n346636 , n24026 );
not ( n26604 , n346636 );
or ( n26605 , n346635 , n26604 );
buf ( n346639 , n344060 );
buf ( n346640 , n344445 );
nand ( n26608 , n346639 , n346640 );
buf ( n346642 , n26608 );
buf ( n346643 , n346642 );
nand ( n346644 , n26605 , n346643 );
buf ( n346645 , n346644 );
not ( n346646 , n346645 );
or ( n26614 , n26600 , n346646 );
nand ( n346648 , n25993 , n607 );
nand ( n26616 , n26614 , n346648 );
not ( n26617 , n26616 );
not ( n26618 , n343595 );
buf ( n346652 , n602 );
not ( n26620 , n346652 );
buf ( n346654 , n343872 );
not ( n346655 , n346654 );
or ( n346656 , n26620 , n346655 );
buf ( n346657 , n343878 );
buf ( n346658 , n343553 );
nand ( n346659 , n346657 , n346658 );
buf ( n346660 , n346659 );
buf ( n346661 , n346660 );
nand ( n346662 , n346656 , n346661 );
buf ( n346663 , n346662 );
not ( n26631 , n346663 );
or ( n26632 , n26618 , n26631 );
buf ( n346666 , n346087 );
not ( n346667 , n346666 );
buf ( n346668 , n343531 );
nand ( n26636 , n346667 , n346668 );
buf ( n346670 , n26636 );
nand ( n26638 , n26632 , n346670 );
not ( n26639 , n26638 );
or ( n346673 , n26617 , n26639 );
nor ( n26641 , n26616 , n26638 );
buf ( n346675 , n346559 );
buf ( n346676 , n346571 );
xor ( n26644 , n346675 , n346676 );
buf ( n346678 , n346506 );
xnor ( n346679 , n26644 , n346678 );
buf ( n346680 , n346679 );
buf ( n346681 , n346680 );
not ( n346682 , n346681 );
buf ( n346683 , n346682 );
buf ( n346684 , n346683 );
not ( n346685 , n346684 );
buf ( n346686 , n23681 );
not ( n26654 , n346686 );
buf ( n346688 , n26482 );
not ( n346689 , n346688 );
or ( n26657 , n26654 , n346689 );
buf ( n346691 , n594 );
not ( n346692 , n346691 );
buf ( n346693 , n25424 );
not ( n26661 , n346693 );
buf ( n346695 , n26661 );
buf ( n346696 , n346695 );
not ( n346697 , n346696 );
or ( n26665 , n346692 , n346697 );
buf ( n346699 , n25424 );
buf ( n346700 , n343632 );
nand ( n346701 , n346699 , n346700 );
buf ( n346702 , n346701 );
buf ( n346703 , n346702 );
nand ( n26671 , n26665 , n346703 );
buf ( n346705 , n26671 );
buf ( n346706 , n346705 );
buf ( n346707 , n343762 );
nand ( n26675 , n346706 , n346707 );
buf ( n346709 , n26675 );
buf ( n346710 , n346709 );
nand ( n26678 , n26657 , n346710 );
buf ( n346712 , n26678 );
buf ( n346713 , n346712 );
xor ( n26681 , n346184 , n346220 );
xor ( n346715 , n26681 , n346341 );
buf ( n346716 , n346715 );
buf ( n346717 , n346716 );
xor ( n346718 , n346713 , n346717 );
buf ( n346719 , n343863 );
not ( n26687 , n346719 );
buf ( n346721 , n346537 );
not ( n346722 , n346721 );
or ( n346723 , n26687 , n346722 );
buf ( n346724 , n596 );
not ( n26692 , n346724 );
buf ( n346726 , n24109 );
not ( n346727 , n346726 );
or ( n26695 , n26692 , n346727 );
buf ( n346729 , n343882 );
buf ( n346730 , n24108 );
nand ( n346731 , n346729 , n346730 );
buf ( n346732 , n346731 );
buf ( n346733 , n346732 );
nand ( n346734 , n26695 , n346733 );
buf ( n346735 , n346734 );
buf ( n346736 , n346735 );
buf ( n346737 , n23889 );
nand ( n346738 , n346736 , n346737 );
buf ( n346739 , n346738 );
buf ( n346740 , n346739 );
nand ( n346741 , n346723 , n346740 );
buf ( n346742 , n346741 );
buf ( n346743 , n346742 );
and ( n346744 , n346718 , n346743 );
and ( n346745 , n346713 , n346717 );
or ( n26713 , n346744 , n346745 );
buf ( n346747 , n26713 );
buf ( n346748 , n346747 );
not ( n26716 , n346748 );
buf ( n26717 , n26716 );
buf ( n346751 , n26717 );
not ( n26719 , n346751 );
buf ( n346753 , n23911 );
not ( n26721 , n346753 );
buf ( n346755 , n346500 );
not ( n346756 , n346755 );
or ( n346757 , n26721 , n346756 );
buf ( n346758 , n598 );
not ( n346759 , n346758 );
buf ( n346760 , n343678 );
not ( n346761 , n346760 );
or ( n346762 , n346759 , n346761 );
buf ( n346763 , n343675 );
buf ( n346764 , n343953 );
nand ( n346765 , n346763 , n346764 );
buf ( n346766 , n346765 );
buf ( n346767 , n346766 );
nand ( n26735 , n346762 , n346767 );
buf ( n346769 , n26735 );
buf ( n346770 , n346769 );
buf ( n346771 , n343945 );
nand ( n26739 , n346770 , n346771 );
buf ( n26740 , n26739 );
buf ( n346774 , n26740 );
nand ( n346775 , n346757 , n346774 );
buf ( n346776 , n346775 );
buf ( n346777 , n346776 );
not ( n346778 , n346777 );
buf ( n346779 , n346778 );
buf ( n346780 , n346779 );
not ( n346781 , n346780 );
or ( n26749 , n26719 , n346781 );
buf ( n346783 , n346553 );
not ( n26751 , n346783 );
buf ( n346785 , n346523 );
not ( n26753 , n346785 );
and ( n346787 , n26751 , n26753 );
buf ( n346788 , n346523 );
buf ( n346789 , n346553 );
and ( n346790 , n346788 , n346789 );
nor ( n26758 , n346787 , n346790 );
buf ( n346792 , n26758 );
xor ( n346793 , n346544 , n346792 );
buf ( n346794 , n346793 );
not ( n26762 , n346794 );
buf ( n26763 , n26762 );
buf ( n346797 , n26763 );
nand ( n26765 , n26749 , n346797 );
buf ( n346799 , n26765 );
buf ( n346800 , n346799 );
buf ( n346801 , n346776 );
buf ( n346802 , n346747 );
nand ( n26770 , n346801 , n346802 );
buf ( n346804 , n26770 );
buf ( n346805 , n346804 );
nand ( n26773 , n346800 , n346805 );
buf ( n346807 , n26773 );
buf ( n346808 , n346807 );
not ( n26776 , n346808 );
buf ( n346810 , n344015 );
not ( n26778 , n346810 );
buf ( n346812 , n26445 );
not ( n26780 , n346812 );
or ( n26781 , n26778 , n26780 );
buf ( n346815 , n600 );
not ( n346816 , n346815 );
buf ( n346817 , n23694 );
not ( n26785 , n346817 );
or ( n26786 , n346816 , n26785 );
buf ( n26787 , n343723 );
buf ( n346821 , n23906 );
nand ( n346822 , n26787 , n346821 );
buf ( n346823 , n346822 );
buf ( n346824 , n346823 );
nand ( n346825 , n26786 , n346824 );
buf ( n346826 , n346825 );
buf ( n346827 , n346826 );
buf ( n346828 , n344018 );
nand ( n26796 , n346827 , n346828 );
buf ( n26797 , n26796 );
buf ( n346831 , n26797 );
nand ( n26799 , n26781 , n346831 );
buf ( n346833 , n26799 );
buf ( n346834 , n346833 );
not ( n26802 , n346834 );
buf ( n346836 , n26802 );
buf ( n346837 , n346836 );
nand ( n26805 , n26776 , n346837 );
buf ( n346839 , n26805 );
buf ( n346840 , n346839 );
not ( n26808 , n346840 );
or ( n26809 , n346685 , n26808 );
buf ( n346843 , n346836 );
not ( n26811 , n346843 );
buf ( n346845 , n346807 );
nand ( n26813 , n26811 , n346845 );
buf ( n346847 , n26813 );
buf ( n346848 , n346847 );
nand ( n26816 , n26809 , n346848 );
buf ( n346850 , n26816 );
buf ( n346851 , n346850 );
not ( n346852 , n346851 );
buf ( n346853 , n346852 );
or ( n346854 , n26641 , n346853 );
nand ( n346855 , n346673 , n346854 );
nand ( n26823 , n346632 , n346855 );
nand ( n346857 , n26593 , n26823 );
buf ( n26825 , n346857 );
and ( n346859 , n26425 , n26825 );
nor ( n26827 , n26422 , n346859 );
nand ( n346861 , n26403 , n26827 );
buf ( n346862 , n346861 );
not ( n26830 , n346862 );
not ( n26831 , n346857 );
and ( n26832 , n26419 , n26831 );
not ( n346866 , n26419 );
and ( n26834 , n346866 , n346857 );
nor ( n26835 , n26832 , n26834 );
not ( n346869 , n346440 );
and ( n346870 , n26835 , n346869 );
not ( n26838 , n26835 );
and ( n346872 , n26838 , n346440 );
nor ( n346873 , n346870 , n346872 );
not ( n26841 , n346045 );
buf ( n346875 , n25995 );
not ( n346876 , n346875 );
nand ( n346877 , n26841 , n346876 , n346050 );
nor ( n26845 , n346050 , n26013 );
nand ( n346879 , n346876 , n26845 );
not ( n26847 , n26018 );
nand ( n26848 , n26847 , n346875 );
not ( n346882 , n346047 );
nand ( n26850 , n346882 , n346875 );
nand ( n26851 , n346877 , n346879 , n26848 , n26850 );
buf ( n346885 , n344338 );
not ( n26853 , n346885 );
buf ( n346887 , n26003 );
not ( n346888 , n346887 );
or ( n346889 , n26853 , n346888 );
buf ( n346890 , n604 );
not ( n346891 , n346890 );
buf ( n346892 , n343985 );
not ( n26860 , n346892 );
or ( n346894 , n346891 , n26860 );
buf ( n26862 , n343982 );
buf ( n26863 , n23530 );
nand ( n26864 , n26862 , n26863 );
buf ( n26865 , n26864 );
buf ( n26866 , n26865 );
nand ( n26867 , n346894 , n26866 );
buf ( n26868 , n26867 );
buf ( n346902 , n26868 );
buf ( n346903 , n344400 );
nand ( n26871 , n346902 , n346903 );
buf ( n346905 , n26871 );
buf ( n346906 , n346905 );
nand ( n346907 , n346889 , n346906 );
buf ( n346908 , n346907 );
not ( n26876 , n346908 );
buf ( n346910 , n344015 );
not ( n346911 , n346910 );
buf ( n346912 , n346826 );
not ( n26880 , n346912 );
or ( n26881 , n346911 , n26880 );
not ( n26882 , n600 );
buf ( n346916 , n23758 );
not ( n346917 , n346916 );
buf ( n346918 , n346917 );
not ( n26886 , n346918 );
or ( n26887 , n26882 , n26886 );
buf ( n346921 , n343744 );
buf ( n346922 , n23906 );
nand ( n346923 , n346921 , n346922 );
buf ( n346924 , n346923 );
nand ( n26892 , n26887 , n346924 );
buf ( n346926 , n26892 );
buf ( n346927 , n344018 );
nand ( n26895 , n346926 , n346927 );
buf ( n346929 , n26895 );
buf ( n346930 , n346929 );
nand ( n346931 , n26881 , n346930 );
buf ( n346932 , n346931 );
buf ( n346933 , n346932 );
not ( n26901 , n346933 );
buf ( n346935 , n23681 );
not ( n26903 , n346935 );
buf ( n346937 , n346705 );
not ( n26905 , n346937 );
or ( n346939 , n26903 , n26905 );
buf ( n346940 , n594 );
not ( n26908 , n346940 );
buf ( n346942 , n346157 );
not ( n346943 , n346942 );
or ( n26911 , n26908 , n346943 );
buf ( n346945 , n25668 );
buf ( n346946 , n343632 );
nand ( n26914 , n346945 , n346946 );
buf ( n346948 , n26914 );
buf ( n346949 , n346948 );
nand ( n346950 , n26911 , n346949 );
buf ( n346951 , n346950 );
buf ( n346952 , n346951 );
buf ( n346953 , n343762 );
nand ( n26921 , n346952 , n346953 );
buf ( n346955 , n26921 );
buf ( n346956 , n346955 );
nand ( n26924 , n346939 , n346956 );
buf ( n346958 , n26924 );
buf ( n346959 , n346958 );
buf ( n346960 , n346257 );
buf ( n346961 , n346335 );
xor ( n346962 , n346960 , n346961 );
buf ( n346963 , n26215 );
xor ( n346964 , n346962 , n346963 );
buf ( n346965 , n346964 );
buf ( n346966 , n346965 );
xor ( n26934 , n346959 , n346966 );
buf ( n26935 , n23681 );
not ( n26936 , n26935 );
buf ( n26937 , n346951 );
not ( n26938 , n26937 );
or ( n26939 , n26936 , n26938 );
buf ( n346973 , n594 );
not ( n346974 , n346973 );
buf ( n346975 , n346202 );
not ( n26943 , n346975 );
or ( n346977 , n346974 , n26943 );
buf ( n346978 , n346205 );
buf ( n346979 , n343632 );
nand ( n346980 , n346978 , n346979 );
buf ( n346981 , n346980 );
buf ( n346982 , n346981 );
nand ( n346983 , n346977 , n346982 );
buf ( n346984 , n346983 );
buf ( n346985 , n346984 );
buf ( n346986 , n343762 );
nand ( n346987 , n346985 , n346986 );
buf ( n346988 , n346987 );
buf ( n346989 , n346988 );
nand ( n26957 , n26939 , n346989 );
buf ( n346991 , n26957 );
not ( n346992 , n346991 );
xor ( n346993 , n26237 , n346317 );
xor ( n26961 , n346993 , n346331 );
buf ( n346995 , n26961 );
not ( n346996 , n346995 );
nand ( n26964 , n346992 , n346996 );
not ( n346998 , n26964 );
xnor ( n346999 , n346296 , n346313 );
buf ( n347000 , n346999 );
not ( n26968 , n347000 );
buf ( n347002 , n23681 );
not ( n26970 , n347002 );
buf ( n347004 , n346984 );
not ( n26972 , n347004 );
or ( n26973 , n26970 , n26972 );
buf ( n347007 , n594 );
not ( n26975 , n347007 );
buf ( n347009 , n346231 );
not ( n26977 , n347009 );
or ( n26978 , n26975 , n26977 );
buf ( n347012 , n14746 );
buf ( n347013 , n343632 );
nand ( n347014 , n347012 , n347013 );
buf ( n347015 , n347014 );
buf ( n347016 , n347015 );
nand ( n26984 , n26978 , n347016 );
buf ( n347018 , n26984 );
buf ( n347019 , n347018 );
buf ( n347020 , n343762 );
nand ( n26988 , n347019 , n347020 );
buf ( n347022 , n26988 );
buf ( n347023 , n347022 );
nand ( n26991 , n26973 , n347023 );
buf ( n347025 , n26991 );
buf ( n347026 , n347025 );
not ( n26994 , n347026 );
buf ( n347028 , n26994 );
buf ( n347029 , n347028 );
not ( n26997 , n347029 );
or ( n347031 , n26968 , n26997 );
buf ( n347032 , n23681 );
not ( n347033 , n347032 );
buf ( n27001 , n347018 );
not ( n27002 , n27001 );
or ( n27003 , n347033 , n27002 );
buf ( n347037 , n594 );
not ( n347038 , n347037 );
buf ( n347039 , n346254 );
not ( n347040 , n347039 );
or ( n347041 , n347038 , n347040 );
buf ( n347042 , n14749 );
buf ( n347043 , n343632 );
nand ( n27011 , n347042 , n347043 );
buf ( n347045 , n27011 );
buf ( n347046 , n347045 );
nand ( n27014 , n347041 , n347046 );
buf ( n347048 , n27014 );
buf ( n347049 , n347048 );
buf ( n347050 , n343762 );
nand ( n347051 , n347049 , n347050 );
buf ( n347052 , n347051 );
buf ( n347053 , n347052 );
nand ( n27021 , n27003 , n347053 );
buf ( n347055 , n27021 );
buf ( n347056 , n347055 );
buf ( n347057 , n26233 );
buf ( n347058 , n23613 );
nand ( n347059 , n347057 , n347058 );
buf ( n347060 , n347059 );
buf ( n347061 , n347060 );
not ( n347062 , n347061 );
buf ( n347063 , n347062 );
buf ( n347064 , n347063 );
or ( n27032 , n347056 , n347064 );
buf ( n27033 , n23681 );
not ( n27034 , n27033 );
buf ( n27035 , n347048 );
not ( n27036 , n27035 );
or ( n27037 , n27034 , n27036 );
buf ( n347071 , n26233 );
buf ( n347072 , n343632 );
or ( n27040 , n347071 , n347072 );
not ( n347074 , n26233 );
buf ( n27042 , n347074 );
buf ( n347076 , n594 );
or ( n347077 , n27042 , n347076 );
nand ( n347078 , n27040 , n347077 );
buf ( n347079 , n347078 );
buf ( n347080 , n347079 );
buf ( n347081 , n343762 );
nand ( n347082 , n347080 , n347081 );
buf ( n347083 , n347082 );
buf ( n347084 , n347083 );
nand ( n347085 , n27037 , n347084 );
buf ( n347086 , n347085 );
buf ( n347087 , n347086 );
buf ( n347088 , n595 );
buf ( n347089 , n596 );
or ( n347090 , n347088 , n347089 );
buf ( n347091 , n26233 );
nand ( n27059 , n347090 , n347091 );
buf ( n347093 , n27059 );
buf ( n347094 , n347093 );
buf ( n347095 , n595 );
buf ( n347096 , n596 );
and ( n27064 , n347095 , n347096 );
buf ( n347098 , n343632 );
nor ( n347099 , n27064 , n347098 );
buf ( n347100 , n347099 );
buf ( n347101 , n347100 );
and ( n347102 , n347094 , n347101 );
buf ( n347103 , n347102 );
buf ( n347104 , n347103 );
and ( n347105 , n347087 , n347104 );
buf ( n347106 , n347105 );
buf ( n347107 , n347106 );
nand ( n347108 , n27032 , n347107 );
buf ( n347109 , n347108 );
buf ( n347110 , n347109 );
buf ( n347111 , n347063 );
buf ( n347112 , n347055 );
nand ( n27080 , n347111 , n347112 );
buf ( n347114 , n27080 );
buf ( n347115 , n347114 );
and ( n347116 , n347110 , n347115 );
buf ( n347117 , n347116 );
buf ( n347118 , n347117 );
not ( n27086 , n347118 );
buf ( n347120 , n27086 );
buf ( n347121 , n347120 );
nand ( n27089 , n347031 , n347121 );
buf ( n347123 , n27089 );
buf ( n347124 , n346999 );
not ( n27092 , n347124 );
buf ( n347126 , n347025 );
nand ( n347127 , n27092 , n347126 );
buf ( n347128 , n347127 );
nand ( n347129 , n347123 , n347128 );
not ( n347130 , n347129 );
or ( n27098 , n346998 , n347130 );
nand ( n27099 , n346991 , n346995 );
nand ( n27100 , n27098 , n27099 );
buf ( n347134 , n27100 );
and ( n347135 , n26934 , n347134 );
and ( n347136 , n346959 , n346966 );
or ( n27104 , n347135 , n347136 );
buf ( n347138 , n27104 );
buf ( n347139 , n347138 );
buf ( n347140 , n23911 );
not ( n27108 , n347140 );
buf ( n347142 , n346769 );
not ( n347143 , n347142 );
or ( n27111 , n27108 , n347143 );
buf ( n347145 , n598 );
not ( n347146 , n347145 );
buf ( n347147 , n26331 );
not ( n347148 , n347147 );
or ( n347149 , n347146 , n347148 );
buf ( n347150 , n23606 );
buf ( n347151 , n343953 );
nand ( n347152 , n347150 , n347151 );
buf ( n347153 , n347152 );
buf ( n347154 , n347153 );
nand ( n347155 , n347149 , n347154 );
buf ( n347156 , n347155 );
buf ( n347157 , n347156 );
buf ( n347158 , n343945 );
nand ( n27126 , n347157 , n347158 );
buf ( n347160 , n27126 );
buf ( n347161 , n347160 );
nand ( n347162 , n27111 , n347161 );
buf ( n347163 , n347162 );
buf ( n347164 , n347163 );
xor ( n347165 , n347139 , n347164 );
xor ( n27133 , n346713 , n346717 );
xor ( n347167 , n27133 , n346743 );
buf ( n347168 , n347167 );
buf ( n347169 , n347168 );
and ( n347170 , n347165 , n347169 );
and ( n347171 , n347139 , n347164 );
or ( n27139 , n347170 , n347171 );
buf ( n347173 , n27139 );
buf ( n347174 , n347173 );
not ( n27142 , n347174 );
buf ( n27143 , n27142 );
buf ( n347177 , n27143 );
nand ( n347178 , n26901 , n347177 );
buf ( n347179 , n347178 );
buf ( n347180 , n347179 );
buf ( n347181 , n346747 );
buf ( n347182 , n346776 );
xor ( n347183 , n347181 , n347182 );
buf ( n347184 , n346793 );
xor ( n347185 , n347183 , n347184 );
buf ( n347186 , n347185 );
buf ( n347187 , n347186 );
not ( n27155 , n347187 );
buf ( n27156 , n27155 );
buf ( n347190 , n27156 );
and ( n347191 , n347180 , n347190 );
buf ( n347192 , n346932 );
not ( n347193 , n347192 );
buf ( n347194 , n27143 );
nor ( n27162 , n347193 , n347194 );
buf ( n347196 , n27162 );
buf ( n347197 , n347196 );
nor ( n27165 , n347191 , n347197 );
buf ( n27166 , n27165 );
buf ( n347200 , n27166 );
buf ( n347201 , n346663 );
buf ( n347202 , n343531 );
and ( n347203 , n347201 , n347202 );
not ( n27171 , n343908 );
not ( n27172 , n343553 );
or ( n27173 , n27171 , n27172 );
buf ( n347207 , n343908 );
buf ( n27175 , n347207 );
buf ( n347209 , n27175 );
not ( n27177 , n347209 );
nand ( n347211 , n27177 , n602 );
nand ( n27179 , n27173 , n347211 );
buf ( n347213 , n27179 );
not ( n27181 , n347213 );
buf ( n347215 , n346090 );
nor ( n347216 , n27181 , n347215 );
buf ( n347217 , n347216 );
buf ( n347218 , n347217 );
nor ( n27186 , n347203 , n347218 );
buf ( n347220 , n27186 );
buf ( n347221 , n347220 );
xor ( n27189 , n347200 , n347221 );
buf ( n347223 , n604 );
not ( n27191 , n347223 );
buf ( n347225 , n343962 );
not ( n347226 , n347225 );
or ( n347227 , n27191 , n347226 );
buf ( n347228 , n343966 );
buf ( n347229 , n23530 );
nand ( n27197 , n347228 , n347229 );
buf ( n347231 , n27197 );
buf ( n347232 , n347231 );
nand ( n27200 , n347227 , n347232 );
buf ( n347234 , n27200 );
buf ( n347235 , n347234 );
buf ( n347236 , n344400 );
and ( n347237 , n347235 , n347236 );
buf ( n347238 , n26868 );
buf ( n347239 , n344338 );
and ( n347240 , n347238 , n347239 );
nor ( n27208 , n347237 , n347240 );
buf ( n27209 , n27208 );
buf ( n347243 , n27209 );
and ( n27211 , n27189 , n347243 );
and ( n27212 , n347200 , n347221 );
or ( n27213 , n27211 , n27212 );
buf ( n347247 , n27213 );
buf ( n347248 , n347247 );
not ( n27216 , n347248 );
buf ( n347250 , n27216 );
not ( n27218 , n347250 );
or ( n347252 , n26876 , n27218 );
buf ( n27220 , n346908 );
not ( n347254 , n27220 );
buf ( n347255 , n347254 );
buf ( n347256 , n347255 );
not ( n27224 , n347256 );
buf ( n347258 , n347247 );
not ( n27226 , n347258 );
or ( n27227 , n27224 , n27226 );
buf ( n347261 , n346595 );
buf ( n347262 , n346590 );
and ( n27230 , n347261 , n347262 );
not ( n27231 , n347261 );
buf ( n27232 , n346485 );
and ( n347266 , n27231 , n27232 );
nor ( n27234 , n27230 , n347266 );
buf ( n27235 , n27234 );
and ( n347269 , n27235 , n346602 );
not ( n27237 , n27235 );
not ( n347271 , n346602 );
and ( n347272 , n27237 , n347271 );
nor ( n27240 , n347269 , n347272 );
buf ( n347274 , n27240 );
nand ( n27242 , n27227 , n347274 );
buf ( n347276 , n27242 );
nand ( n347277 , n347252 , n347276 );
xor ( n27245 , n26851 , n347277 );
xor ( n27246 , n26575 , n26591 );
xor ( n27247 , n27246 , n346855 );
and ( n347281 , n27245 , n27247 );
and ( n347282 , n26851 , n347277 );
or ( n27250 , n347281 , n347282 );
nor ( n27251 , n346873 , n27250 );
not ( n347285 , n27251 );
not ( n347286 , n26616 );
and ( n27254 , n26638 , n346853 );
not ( n347288 , n26638 );
and ( n27256 , n347288 , n346850 );
nor ( n347290 , n27254 , n27256 );
not ( n27258 , n347290 );
not ( n347292 , n27258 );
or ( n27260 , n347286 , n347292 );
not ( n27261 , n26616 );
nand ( n347295 , n27261 , n347290 );
nand ( n347296 , n27260 , n347295 );
not ( n27264 , n347296 );
and ( n347298 , n27240 , n346908 );
not ( n347299 , n27240 );
and ( n27267 , n347299 , n347255 );
nor ( n347301 , n347298 , n27267 );
and ( n347302 , n347301 , n347247 );
not ( n27270 , n347301 );
and ( n27271 , n27270 , n347250 );
nor ( n347305 , n347302 , n27271 );
not ( n347306 , n347305 );
or ( n27274 , n27264 , n347306 );
buf ( n347308 , n346807 );
buf ( n347309 , n346833 );
xor ( n27277 , n347308 , n347309 );
buf ( n347311 , n346680 );
xnor ( n347312 , n27277 , n347311 );
buf ( n347313 , n347312 );
buf ( n347314 , n347313 );
buf ( n347315 , n347314 );
buf ( n347316 , n347315 );
buf ( n347317 , n347316 );
not ( n27285 , n347317 );
buf ( n347319 , n607 );
not ( n347320 , n347319 );
buf ( n347321 , n346645 );
not ( n27289 , n347321 );
or ( n347323 , n347320 , n27289 );
buf ( n347324 , n606 );
not ( n27292 , n347324 );
buf ( n347326 , n23996 );
not ( n347327 , n347326 );
or ( n27295 , n27292 , n347327 );
buf ( n347329 , n344035 );
buf ( n347330 , n344445 );
nand ( n347331 , n347329 , n347330 );
buf ( n347332 , n347331 );
buf ( n347333 , n347332 );
nand ( n347334 , n27295 , n347333 );
buf ( n347335 , n347334 );
buf ( n347336 , n347335 );
buf ( n27304 , n344454 );
nand ( n27305 , n347336 , n27304 );
buf ( n347339 , n27305 );
buf ( n347340 , n347339 );
nand ( n27308 , n347323 , n347340 );
buf ( n347342 , n27308 );
buf ( n347343 , n347342 );
not ( n27311 , n347343 );
or ( n347345 , n27285 , n27311 );
buf ( n347346 , n347316 );
buf ( n347347 , n347342 );
or ( n347348 , n347346 , n347347 );
buf ( n347349 , n343531 );
not ( n27317 , n347349 );
buf ( n347351 , n27179 );
not ( n347352 , n347351 );
or ( n27320 , n27317 , n347352 );
buf ( n347354 , n602 );
not ( n347355 , n347354 );
buf ( n347356 , n343837 );
not ( n347357 , n347356 );
buf ( n347358 , n347357 );
buf ( n347359 , n347358 );
not ( n27327 , n347359 );
or ( n27328 , n347355 , n27327 );
buf ( n347362 , n23798 );
not ( n347363 , n347362 );
buf ( n347364 , n343553 );
nand ( n27332 , n347363 , n347364 );
buf ( n347366 , n27332 );
buf ( n347367 , n347366 );
nand ( n347368 , n27328 , n347367 );
buf ( n347369 , n347368 );
buf ( n347370 , n347369 );
buf ( n347371 , n343595 );
nand ( n347372 , n347370 , n347371 );
buf ( n347373 , n347372 );
buf ( n347374 , n347373 );
nand ( n27342 , n27320 , n347374 );
buf ( n347376 , n27342 );
buf ( n347377 , n347376 );
not ( n27345 , n347377 );
buf ( n347379 , n347173 );
buf ( n347380 , n346932 );
xor ( n347381 , n347379 , n347380 );
buf ( n347382 , n347186 );
xnor ( n27350 , n347381 , n347382 );
buf ( n27351 , n27350 );
buf ( n347385 , n27351 );
not ( n27353 , n347385 );
or ( n347387 , n27345 , n27353 );
buf ( n347388 , n27351 );
buf ( n347389 , n347376 );
or ( n347390 , n347388 , n347389 );
buf ( n347391 , n343863 );
not ( n27359 , n347391 );
buf ( n347393 , n346735 );
not ( n347394 , n347393 );
or ( n347395 , n27359 , n347394 );
buf ( n347396 , n596 );
not ( n27364 , n347396 );
buf ( n347398 , n345175 );
not ( n27366 , n347398 );
or ( n347400 , n27364 , n27366 );
buf ( n27368 , n25403 );
buf ( n347402 , n343882 );
nand ( n27370 , n27368 , n347402 );
buf ( n347404 , n27370 );
buf ( n347405 , n347404 );
nand ( n27373 , n347400 , n347405 );
buf ( n347407 , n27373 );
buf ( n347408 , n347407 );
buf ( n347409 , n23889 );
nand ( n347410 , n347408 , n347409 );
buf ( n347411 , n347410 );
buf ( n347412 , n347411 );
nand ( n347413 , n347395 , n347412 );
buf ( n347414 , n347413 );
buf ( n347415 , n347414 );
xor ( n27383 , n346959 , n346966 );
xor ( n27384 , n27383 , n347134 );
buf ( n27385 , n27384 );
buf ( n347419 , n27385 );
xor ( n27387 , n347415 , n347419 );
buf ( n347421 , n23911 );
not ( n27389 , n347421 );
buf ( n347423 , n347156 );
not ( n347424 , n347423 );
or ( n347425 , n27389 , n347424 );
buf ( n347426 , n598 );
not ( n347427 , n347426 );
buf ( n347428 , n24091 );
not ( n27396 , n347428 );
or ( n347430 , n347427 , n27396 );
buf ( n347431 , n24092 );
buf ( n347432 , n343953 );
nand ( n27400 , n347431 , n347432 );
buf ( n347434 , n27400 );
buf ( n347435 , n347434 );
nand ( n347436 , n347430 , n347435 );
buf ( n347437 , n347436 );
buf ( n347438 , n347437 );
buf ( n347439 , n343945 );
nand ( n27407 , n347438 , n347439 );
buf ( n27408 , n27407 );
buf ( n347442 , n27408 );
nand ( n347443 , n347425 , n347442 );
buf ( n347444 , n347443 );
buf ( n347445 , n347444 );
and ( n347446 , n27387 , n347445 );
and ( n27414 , n347415 , n347419 );
or ( n347448 , n347446 , n27414 );
buf ( n347449 , n347448 );
not ( n27417 , n347449 );
not ( n27418 , n600 );
not ( n27419 , n344484 );
or ( n347453 , n27418 , n27419 );
buf ( n347454 , n346493 );
buf ( n347455 , n23906 );
nand ( n27423 , n347454 , n347455 );
buf ( n347457 , n27423 );
nand ( n347458 , n347453 , n347457 );
not ( n347459 , n347458 );
not ( n27427 , n347459 );
not ( n27428 , n344017 );
and ( n27429 , n27427 , n27428 );
and ( n347463 , n26892 , n344015 );
nor ( n27431 , n27429 , n347463 );
nand ( n347465 , n27417 , n27431 );
not ( n27433 , n347465 );
xor ( n27434 , n347139 , n347164 );
xor ( n347468 , n27434 , n347169 );
buf ( n347469 , n347468 );
not ( n27437 , n347469 );
or ( n347471 , n27433 , n27437 );
buf ( n347472 , n27431 );
not ( n27440 , n347472 );
buf ( n347474 , n347449 );
nand ( n27442 , n27440 , n347474 );
buf ( n347476 , n27442 );
nand ( n347477 , n347471 , n347476 );
buf ( n347478 , n347477 );
nand ( n27446 , n347390 , n347478 );
buf ( n347480 , n27446 );
buf ( n347481 , n347480 );
nand ( n347482 , n347387 , n347481 );
buf ( n347483 , n347482 );
buf ( n347484 , n347483 );
nand ( n27452 , n347348 , n347484 );
buf ( n347486 , n27452 );
buf ( n347487 , n347486 );
nand ( n27455 , n347345 , n347487 );
buf ( n347489 , n27455 );
nand ( n347490 , n27274 , n347489 );
buf ( n347491 , n347490 );
not ( n27459 , n347296 );
buf ( n347493 , n347305 );
not ( n27461 , n347493 );
buf ( n347495 , n27461 );
nand ( n27463 , n27459 , n347495 );
buf ( n347497 , n27463 );
nand ( n27465 , n347491 , n347497 );
buf ( n347499 , n27465 );
buf ( n27467 , n347499 );
not ( n347501 , n27467 );
buf ( n347502 , n347501 );
xor ( n347503 , n26851 , n347277 );
xor ( n347504 , n347503 , n27247 );
not ( n27472 , n347504 );
nand ( n347506 , n347502 , n27472 );
nand ( n347507 , n347285 , n347506 );
buf ( n347508 , n347507 );
nor ( n27476 , n26830 , n347508 );
buf ( n347510 , n27476 );
not ( n347511 , n347510 );
xor ( n27479 , n347376 , n347477 );
buf ( n347513 , n27479 );
buf ( n347514 , n27351 );
buf ( n27482 , n347514 );
buf ( n27483 , n27482 );
buf ( n347517 , n27483 );
xnor ( n347518 , n347513 , n347517 );
buf ( n347519 , n347518 );
buf ( n347520 , n347519 );
buf ( n347521 , n344338 );
not ( n27489 , n347521 );
buf ( n347523 , n344957 );
not ( n347524 , n347523 );
buf ( n347525 , n347524 );
and ( n27493 , n604 , n347525 );
not ( n347527 , n604 );
and ( n27495 , n347527 , n343878 );
or ( n27496 , n27493 , n27495 );
buf ( n347530 , n27496 );
not ( n347531 , n347530 );
or ( n347532 , n27489 , n347531 );
buf ( n347533 , n344400 );
buf ( n347534 , n604 );
not ( n347535 , n347534 );
buf ( n347536 , n343911 );
not ( n347537 , n347536 );
or ( n347538 , n347535 , n347537 );
buf ( n347539 , n347209 );
buf ( n347540 , n23530 );
nand ( n27508 , n347539 , n347540 );
buf ( n347542 , n27508 );
buf ( n347543 , n347542 );
nand ( n347544 , n347538 , n347543 );
buf ( n347545 , n347544 );
buf ( n347546 , n347545 );
nand ( n347547 , n347533 , n347546 );
buf ( n347548 , n347547 );
buf ( n347549 , n347548 );
nand ( n347550 , n347532 , n347549 );
buf ( n347551 , n347550 );
not ( n27519 , n347551 );
buf ( n347553 , n27519 );
not ( n347554 , n347553 );
buf ( n347555 , n607 );
not ( n347556 , n347555 );
and ( n347557 , n343985 , n606 );
not ( n27525 , n343985 );
and ( n27526 , n27525 , n344445 );
or ( n27527 , n347557 , n27526 );
buf ( n347561 , n27527 );
not ( n347562 , n347561 );
or ( n27530 , n347556 , n347562 );
buf ( n347564 , n606 );
not ( n27532 , n347564 );
buf ( n347566 , n343969 );
not ( n347567 , n347566 );
or ( n27535 , n27532 , n347567 );
buf ( n347569 , n343966 );
buf ( n347570 , n344445 );
nand ( n347571 , n347569 , n347570 );
buf ( n347572 , n347571 );
buf ( n347573 , n347572 );
nand ( n27541 , n27535 , n347573 );
buf ( n347575 , n27541 );
buf ( n347576 , n347575 );
buf ( n27544 , n344454 );
nand ( n27545 , n347576 , n27544 );
buf ( n347579 , n27545 );
buf ( n347580 , n347579 );
nand ( n347581 , n27530 , n347580 );
buf ( n347582 , n347581 );
buf ( n347583 , n347582 );
not ( n347584 , n347583 );
buf ( n347585 , n347584 );
buf ( n347586 , n347585 );
not ( n27554 , n347586 );
or ( n27555 , n347554 , n27554 );
not ( n27556 , n23911 );
not ( n27557 , n347437 );
or ( n27558 , n27556 , n27557 );
not ( n347592 , n343953 );
not ( n347593 , n24110 );
or ( n27561 , n347592 , n347593 );
not ( n347595 , n24109 );
buf ( n347596 , n347595 );
not ( n347597 , n347596 );
buf ( n347598 , n598 );
nand ( n27566 , n347597 , n347598 );
buf ( n347600 , n27566 );
nand ( n347601 , n27561 , n347600 );
nand ( n347602 , n347601 , n343945 );
nand ( n27570 , n27558 , n347602 );
buf ( n347604 , n344015 );
not ( n27572 , n347604 );
buf ( n347606 , n600 );
not ( n347607 , n347606 );
buf ( n347608 , n343678 );
not ( n27576 , n347608 );
or ( n27577 , n347607 , n27576 );
buf ( n347611 , n343675 );
buf ( n347612 , n23906 );
nand ( n27580 , n347611 , n347612 );
buf ( n347614 , n27580 );
buf ( n347615 , n347614 );
nand ( n347616 , n27577 , n347615 );
buf ( n347617 , n347616 );
buf ( n347618 , n347617 );
not ( n27586 , n347618 );
or ( n27587 , n27572 , n27586 );
buf ( n347621 , n600 );
not ( n27589 , n347621 );
buf ( n347623 , n26331 );
not ( n27591 , n347623 );
or ( n27592 , n27589 , n27591 );
buf ( n347626 , n23606 );
buf ( n347627 , n23906 );
nand ( n347628 , n347626 , n347627 );
buf ( n347629 , n347628 );
buf ( n347630 , n347629 );
nand ( n27598 , n27592 , n347630 );
buf ( n347632 , n27598 );
buf ( n347633 , n347632 );
buf ( n347634 , n344018 );
nand ( n347635 , n347633 , n347634 );
buf ( n347636 , n347635 );
buf ( n347637 , n347636 );
nand ( n347638 , n27587 , n347637 );
buf ( n347639 , n347638 );
nor ( n27607 , n27570 , n347639 );
buf ( n347641 , n347407 );
buf ( n347642 , n343863 );
and ( n27610 , n347641 , n347642 );
buf ( n347644 , n343882 );
not ( n347645 , n347644 );
buf ( n347646 , n25424 );
not ( n27614 , n347646 );
or ( n347648 , n347645 , n27614 );
buf ( n347649 , n345451 );
not ( n27617 , n347649 );
buf ( n347651 , n596 );
nand ( n347652 , n27617 , n347651 );
buf ( n347653 , n347652 );
buf ( n347654 , n347653 );
nand ( n27622 , n347648 , n347654 );
buf ( n347656 , n27622 );
buf ( n347657 , n347656 );
not ( n347658 , n347657 );
buf ( n27626 , n23889 );
not ( n347660 , n27626 );
buf ( n347661 , n347660 );
buf ( n347662 , n347661 );
nor ( n27630 , n347658 , n347662 );
buf ( n347664 , n27630 );
buf ( n347665 , n347664 );
nor ( n347666 , n27610 , n347665 );
buf ( n347667 , n347666 );
buf ( n347668 , n347667 );
not ( n347669 , n346996 );
not ( n27637 , n346992 );
or ( n347671 , n347669 , n27637 );
nand ( n347672 , n347671 , n27099 );
xor ( n27640 , n347672 , n347129 );
buf ( n347674 , n27640 );
xor ( n27642 , n347668 , n347674 );
buf ( n347676 , n596 );
not ( n347677 , n347676 );
buf ( n347678 , n346157 );
not ( n347679 , n347678 );
or ( n347680 , n347677 , n347679 );
buf ( n347681 , n25668 );
buf ( n347682 , n343882 );
nand ( n347683 , n347681 , n347682 );
buf ( n347684 , n347683 );
buf ( n347685 , n347684 );
nand ( n27653 , n347680 , n347685 );
buf ( n347687 , n27653 );
buf ( n347688 , n347687 );
not ( n347689 , n347688 );
buf ( n347690 , n347689 );
not ( n347691 , n347690 );
not ( n27659 , n347661 );
and ( n347693 , n347691 , n27659 );
and ( n27661 , n347656 , n343863 );
nor ( n347695 , n347693 , n27661 );
not ( n27663 , n347695 );
buf ( n347697 , n346999 );
buf ( n347698 , n347117 );
xor ( n27666 , n347697 , n347698 );
buf ( n347700 , n347025 );
xnor ( n27668 , n27666 , n347700 );
buf ( n27669 , n27668 );
not ( n347703 , n27669 );
and ( n27671 , n27663 , n347703 );
buf ( n347705 , n343863 );
not ( n347706 , n347705 );
buf ( n347707 , n347687 );
not ( n27675 , n347707 );
or ( n347709 , n347706 , n27675 );
buf ( n347710 , n596 );
not ( n27678 , n347710 );
buf ( n347712 , n26159 );
not ( n347713 , n347712 );
or ( n27681 , n27678 , n347713 );
buf ( n347715 , n346142 );
buf ( n347716 , n343882 );
nand ( n27684 , n347715 , n347716 );
buf ( n347718 , n27684 );
buf ( n347719 , n347718 );
nand ( n27687 , n27681 , n347719 );
buf ( n347721 , n27687 );
buf ( n347722 , n347721 );
buf ( n347723 , n23889 );
nand ( n347724 , n347722 , n347723 );
buf ( n347725 , n347724 );
buf ( n347726 , n347725 );
nand ( n27694 , n347709 , n347726 );
buf ( n347728 , n27694 );
buf ( n347729 , n347728 );
buf ( n347730 , n347055 );
buf ( n347731 , n347060 );
not ( n347732 , n347731 );
buf ( n347733 , n347106 );
not ( n347734 , n347733 );
or ( n347735 , n347732 , n347734 );
buf ( n347736 , n347106 );
buf ( n347737 , n347060 );
or ( n347738 , n347736 , n347737 );
nand ( n27706 , n347735 , n347738 );
buf ( n347740 , n27706 );
buf ( n347741 , n347740 );
xor ( n347742 , n347730 , n347741 );
buf ( n347743 , n347742 );
buf ( n347744 , n347743 );
nor ( n347745 , n347729 , n347744 );
buf ( n347746 , n347745 );
buf ( n347747 , n347746 );
buf ( n347748 , n347086 );
buf ( n347749 , n347103 );
xor ( n347750 , n347748 , n347749 );
buf ( n347751 , n347750 );
buf ( n347752 , n347751 );
buf ( n347753 , n343863 );
not ( n347754 , n347753 );
buf ( n347755 , n596 );
not ( n27723 , n347755 );
buf ( n347757 , n346231 );
not ( n27725 , n347757 );
or ( n347759 , n27723 , n27725 );
buf ( n347760 , n346179 );
buf ( n347761 , n343882 );
nand ( n347762 , n347760 , n347761 );
buf ( n347763 , n347762 );
buf ( n347764 , n347763 );
nand ( n347765 , n347759 , n347764 );
buf ( n347766 , n347765 );
buf ( n347767 , n347766 );
not ( n347768 , n347767 );
or ( n27736 , n347754 , n347768 );
buf ( n347770 , n596 );
not ( n347771 , n347770 );
buf ( n347772 , n14749 );
not ( n347773 , n347772 );
buf ( n347774 , n347773 );
buf ( n347775 , n347774 );
not ( n27743 , n347775 );
or ( n347777 , n347771 , n27743 );
buf ( n347778 , n14749 );
buf ( n347779 , n343882 );
nand ( n347780 , n347778 , n347779 );
buf ( n347781 , n347780 );
buf ( n347782 , n347781 );
nand ( n347783 , n347777 , n347782 );
buf ( n347784 , n347783 );
buf ( n347785 , n347784 );
buf ( n347786 , n23889 );
nand ( n27754 , n347785 , n347786 );
buf ( n347788 , n27754 );
buf ( n347789 , n347788 );
nand ( n347790 , n27736 , n347789 );
buf ( n347791 , n347790 );
not ( n27759 , n347791 );
buf ( n347793 , n26233 );
buf ( n347794 , n23681 );
nand ( n27762 , n347793 , n347794 );
buf ( n27763 , n27762 );
buf ( n347797 , n597 );
buf ( n347798 , n598 );
or ( n347799 , n347797 , n347798 );
buf ( n347800 , n26233 );
nand ( n27768 , n347799 , n347800 );
buf ( n347802 , n27768 );
buf ( n347803 , n347802 );
buf ( n347804 , n597 );
buf ( n347805 , n598 );
and ( n27773 , n347804 , n347805 );
buf ( n347807 , n343882 );
nor ( n347808 , n27773 , n347807 );
buf ( n347809 , n347808 );
buf ( n347810 , n347809 );
nand ( n347811 , n347803 , n347810 );
buf ( n347812 , n347811 );
buf ( n347813 , n347812 );
not ( n27781 , n347813 );
buf ( n347815 , n343863 );
not ( n27783 , n347815 );
buf ( n347817 , n347784 );
not ( n347818 , n347817 );
or ( n27786 , n27783 , n347818 );
buf ( n347820 , n26233 );
buf ( n347821 , n343882 );
or ( n27789 , n347820 , n347821 );
buf ( n347823 , n347074 );
buf ( n347824 , n596 );
or ( n347825 , n347823 , n347824 );
nand ( n347826 , n27789 , n347825 );
buf ( n347827 , n347826 );
buf ( n347828 , n347827 );
buf ( n347829 , n23889 );
nand ( n27797 , n347828 , n347829 );
buf ( n27798 , n27797 );
buf ( n347832 , n27798 );
nand ( n27800 , n27786 , n347832 );
buf ( n347834 , n27800 );
buf ( n347835 , n347834 );
nand ( n347836 , n27781 , n347835 );
buf ( n347837 , n347836 );
and ( n27805 , n27763 , n347837 );
nor ( n27806 , n27759 , n27805 );
buf ( n347840 , n27806 );
xor ( n27808 , n347752 , n347840 );
buf ( n347842 , n343863 );
not ( n347843 , n347842 );
buf ( n347844 , n347721 );
not ( n27812 , n347844 );
or ( n347846 , n347843 , n27812 );
buf ( n347847 , n347766 );
buf ( n347848 , n23889 );
nand ( n347849 , n347847 , n347848 );
buf ( n347850 , n347849 );
buf ( n347851 , n347850 );
nand ( n347852 , n347846 , n347851 );
buf ( n347853 , n347852 );
buf ( n347854 , n347853 );
and ( n347855 , n27808 , n347854 );
and ( n347856 , n347752 , n347840 );
or ( n27824 , n347855 , n347856 );
buf ( n347858 , n27824 );
buf ( n347859 , n347858 );
not ( n347860 , n347859 );
buf ( n347861 , n347860 );
buf ( n347862 , n347861 );
or ( n347863 , n347747 , n347862 );
buf ( n347864 , n347728 );
buf ( n347865 , n347743 );
nand ( n347866 , n347864 , n347865 );
buf ( n347867 , n347866 );
buf ( n347868 , n347867 );
nand ( n347869 , n347863 , n347868 );
buf ( n347870 , n347869 );
nand ( n27838 , n347695 , n27669 );
and ( n27839 , n347870 , n27838 );
nor ( n27840 , n27671 , n27839 );
buf ( n347874 , n27840 );
xor ( n347875 , n27642 , n347874 );
buf ( n347876 , n347875 );
or ( n27844 , n27607 , n347876 );
buf ( n347878 , n347639 );
buf ( n347879 , n27570 );
nand ( n347880 , n347878 , n347879 );
buf ( n347881 , n347880 );
nand ( n27849 , n27844 , n347881 );
buf ( n347883 , n27849 );
buf ( n347884 , n343592 );
not ( n347885 , n347884 );
buf ( n347886 , n602 );
not ( n27854 , n347886 );
buf ( n347888 , n346918 );
not ( n347889 , n347888 );
or ( n347890 , n27854 , n347889 );
buf ( n347891 , n23758 );
buf ( n347892 , n343553 );
nand ( n347893 , n347891 , n347892 );
buf ( n347894 , n347893 );
buf ( n347895 , n347894 );
nand ( n347896 , n347890 , n347895 );
buf ( n347897 , n347896 );
buf ( n347898 , n347897 );
not ( n347899 , n347898 );
or ( n347900 , n347885 , n347899 );
not ( n27868 , n602 );
not ( n27869 , n23694 );
or ( n27870 , n27868 , n27869 );
not ( n347904 , n343723 );
or ( n347905 , n347904 , n602 );
nand ( n27873 , n27870 , n347905 );
nand ( n27874 , n27873 , n343531 );
buf ( n347908 , n27874 );
nand ( n347909 , n347900 , n347908 );
buf ( n347910 , n347909 );
buf ( n347911 , n347910 );
xor ( n347912 , n347883 , n347911 );
xor ( n27880 , n347668 , n347674 );
and ( n27881 , n27880 , n347874 );
and ( n347915 , n347668 , n347674 );
or ( n347916 , n27881 , n347915 );
buf ( n347917 , n347916 );
buf ( n347918 , n347917 );
buf ( n347919 , n344015 );
not ( n27887 , n347919 );
buf ( n347921 , n347458 );
not ( n347922 , n347921 );
or ( n347923 , n27887 , n347922 );
buf ( n347924 , n347617 );
buf ( n347925 , n344018 );
nand ( n347926 , n347924 , n347925 );
buf ( n347927 , n347926 );
buf ( n347928 , n347927 );
nand ( n347929 , n347923 , n347928 );
buf ( n347930 , n347929 );
buf ( n347931 , n347930 );
xor ( n27899 , n347918 , n347931 );
xor ( n27900 , n347415 , n347419 );
xor ( n27901 , n27900 , n347445 );
buf ( n347935 , n27901 );
buf ( n347936 , n347935 );
xnor ( n347937 , n27899 , n347936 );
buf ( n347938 , n347937 );
buf ( n347939 , n347938 );
and ( n27907 , n347912 , n347939 );
and ( n347941 , n347883 , n347911 );
or ( n347942 , n27907 , n347941 );
buf ( n347943 , n347942 );
buf ( n347944 , n347943 );
nand ( n27912 , n27555 , n347944 );
buf ( n347946 , n27912 );
buf ( n347947 , n347946 );
buf ( n347948 , n347582 );
buf ( n347949 , n347551 );
nand ( n27917 , n347948 , n347949 );
buf ( n347951 , n27917 );
buf ( n347952 , n347951 );
and ( n27920 , n347947 , n347952 );
buf ( n27921 , n27920 );
buf ( n27922 , n27921 );
xor ( n27923 , n347520 , n27922 );
buf ( n347957 , n343531 );
not ( n347958 , n347957 );
buf ( n347959 , n347369 );
not ( n347960 , n347959 );
or ( n347961 , n347958 , n347960 );
buf ( n347962 , n27873 );
buf ( n347963 , n343592 );
nand ( n347964 , n347962 , n347963 );
buf ( n347965 , n347964 );
buf ( n347966 , n347965 );
nand ( n27934 , n347961 , n347966 );
buf ( n347968 , n27934 );
buf ( n347969 , n347968 );
not ( n347970 , n347969 );
buf ( n347971 , n347930 );
not ( n27939 , n347971 );
buf ( n347973 , n27939 );
not ( n347974 , n347973 );
not ( n27942 , n347917 );
and ( n27943 , n347974 , n27942 );
buf ( n347977 , n347973 );
buf ( n347978 , n347917 );
nand ( n347979 , n347977 , n347978 );
buf ( n347980 , n347979 );
and ( n27948 , n347980 , n347935 );
nor ( n27949 , n27943 , n27948 );
buf ( n347983 , n27949 );
nand ( n27951 , n347970 , n347983 );
buf ( n347985 , n27951 );
buf ( n347986 , n347985 );
not ( n347987 , n347986 );
buf ( n347988 , n347449 );
buf ( n347989 , n347469 );
xor ( n27957 , n347988 , n347989 );
buf ( n347991 , n27431 );
xnor ( n27959 , n27957 , n347991 );
buf ( n347993 , n27959 );
buf ( n347994 , n347993 );
not ( n347995 , n347994 );
or ( n27963 , n347987 , n347995 );
buf ( n347997 , n27949 );
not ( n347998 , n347997 );
buf ( n347999 , n347968 );
nand ( n348000 , n347998 , n347999 );
buf ( n348001 , n348000 );
buf ( n348002 , n348001 );
nand ( n27970 , n27963 , n348002 );
buf ( n27971 , n27970 );
buf ( n348005 , n344338 );
not ( n27973 , n348005 );
buf ( n348007 , n347234 );
not ( n27975 , n348007 );
or ( n348009 , n27973 , n27975 );
buf ( n348010 , n27496 );
buf ( n348011 , n344400 );
nand ( n348012 , n348010 , n348011 );
buf ( n348013 , n348012 );
buf ( n348014 , n348013 );
nand ( n348015 , n348009 , n348014 );
buf ( n348016 , n348015 );
xor ( n348017 , n27971 , n348016 );
buf ( n348018 , n607 );
not ( n348019 , n348018 );
buf ( n348020 , n347335 );
not ( n27988 , n348020 );
or ( n348022 , n348019 , n27988 );
buf ( n348023 , n27527 );
buf ( n348024 , n344454 );
nand ( n348025 , n348023 , n348024 );
buf ( n348026 , n348025 );
buf ( n348027 , n348026 );
nand ( n348028 , n348022 , n348027 );
buf ( n348029 , n348028 );
not ( n27997 , n348029 );
xor ( n348031 , n348017 , n27997 );
buf ( n348032 , n348031 );
and ( n348033 , n27923 , n348032 );
and ( n348034 , n347520 , n27922 );
or ( n348035 , n348033 , n348034 );
buf ( n348036 , n348035 );
not ( n348037 , n348036 );
xor ( n348038 , n347200 , n347221 );
xor ( n28006 , n348038 , n347243 );
buf ( n348040 , n28006 );
buf ( n348041 , n348040 );
buf ( n348042 , n348029 );
not ( n348043 , n348042 );
buf ( n28011 , n348016 );
not ( n28012 , n28011 );
or ( n28013 , n348043 , n28012 );
buf ( n348047 , n348029 );
buf ( n348048 , n348016 );
or ( n348049 , n348047 , n348048 );
buf ( n348050 , n27971 );
nand ( n348051 , n348049 , n348050 );
buf ( n348052 , n348051 );
buf ( n348053 , n348052 );
nand ( n348054 , n28013 , n348053 );
buf ( n348055 , n348054 );
buf ( n348056 , n348055 );
not ( n28024 , n348056 );
buf ( n348058 , n28024 );
buf ( n348059 , n348058 );
xor ( n28027 , n348041 , n348059 );
buf ( n28028 , n347313 );
buf ( n348062 , n347376 );
not ( n28030 , n348062 );
buf ( n348064 , n27351 );
not ( n28032 , n348064 );
or ( n348066 , n28030 , n28032 );
buf ( n348067 , n347480 );
nand ( n28035 , n348066 , n348067 );
buf ( n28036 , n28035 );
buf ( n348070 , n28036 );
xor ( n28038 , n28028 , n348070 );
buf ( n348072 , n347342 );
xnor ( n28040 , n28038 , n348072 );
buf ( n348074 , n28040 );
buf ( n348075 , n348074 );
xor ( n28043 , n28027 , n348075 );
buf ( n348077 , n28043 );
not ( n348078 , n348077 );
or ( n348079 , n348037 , n348078 );
xor ( n28047 , n347520 , n27922 );
xor ( n348081 , n28047 , n348032 );
buf ( n348082 , n348081 );
buf ( n348083 , n348082 );
buf ( n28051 , n347943 );
not ( n28052 , n28051 );
buf ( n28053 , n27519 );
not ( n28054 , n28053 );
or ( n28055 , n28052 , n28054 );
buf ( n348089 , n347943 );
not ( n348090 , n348089 );
buf ( n348091 , n347551 );
nand ( n348092 , n348090 , n348091 );
buf ( n348093 , n348092 );
buf ( n348094 , n348093 );
nand ( n348095 , n28055 , n348094 );
buf ( n348096 , n348095 );
buf ( n348097 , n348096 );
buf ( n348098 , n347582 );
and ( n348099 , n348097 , n348098 );
not ( n348100 , n348097 );
buf ( n348101 , n347585 );
and ( n348102 , n348100 , n348101 );
nor ( n348103 , n348099 , n348102 );
buf ( n348104 , n348103 );
buf ( n348105 , n348104 );
buf ( n348106 , n348105 );
buf ( n348107 , n347993 );
not ( n348108 , n348107 );
buf ( n348109 , n347968 );
not ( n28077 , n348109 );
buf ( n28078 , n27949 );
not ( n28079 , n28078 );
and ( n28080 , n28077 , n28079 );
buf ( n348114 , n347968 );
buf ( n348115 , n27949 );
and ( n28083 , n348114 , n348115 );
nor ( n348117 , n28080 , n28083 );
buf ( n348118 , n348117 );
buf ( n348119 , n348118 );
not ( n348120 , n348119 );
or ( n348121 , n348108 , n348120 );
buf ( n348122 , n348118 );
buf ( n348123 , n347993 );
or ( n348124 , n348122 , n348123 );
nand ( n28092 , n348121 , n348124 );
buf ( n348126 , n28092 );
buf ( n348127 , n348126 );
not ( n348128 , n348127 );
xor ( n28096 , n347883 , n347911 );
xor ( n28097 , n28096 , n347939 );
buf ( n348131 , n28097 );
not ( n28099 , n348131 );
buf ( n348133 , n344338 );
not ( n28101 , n348133 );
buf ( n348135 , n347545 );
not ( n348136 , n348135 );
or ( n348137 , n28101 , n348136 );
buf ( n348138 , n604 );
not ( n348139 , n348138 );
buf ( n348140 , n347358 );
not ( n28108 , n348140 );
or ( n348142 , n348139 , n28108 );
buf ( n28110 , n343837 );
buf ( n28111 , n23530 );
nand ( n28112 , n28110 , n28111 );
buf ( n28113 , n28112 );
buf ( n28114 , n28113 );
nand ( n28115 , n348142 , n28114 );
buf ( n28116 , n28115 );
buf ( n348150 , n28116 );
buf ( n348151 , n344400 );
nand ( n348152 , n348150 , n348151 );
buf ( n348153 , n348152 );
buf ( n348154 , n348153 );
nand ( n28122 , n348137 , n348154 );
buf ( n348156 , n28122 );
or ( n28124 , n27669 , n347695 );
nand ( n348158 , n28124 , n27838 );
xnor ( n348159 , n348158 , n347870 );
buf ( n348160 , n348159 );
not ( n28128 , n23911 );
not ( n28129 , n347601 );
or ( n28130 , n28128 , n28129 );
and ( n28131 , n345176 , n343953 );
not ( n348165 , n345176 );
and ( n348166 , n348165 , n598 );
or ( n28134 , n28131 , n348166 );
buf ( n348168 , n28134 );
buf ( n348169 , n343945 );
nand ( n348170 , n348168 , n348169 );
buf ( n348171 , n348170 );
nand ( n348172 , n28130 , n348171 );
buf ( n348173 , n348172 );
xor ( n28141 , n348160 , n348173 );
buf ( n28142 , n344015 );
not ( n28143 , n28142 );
buf ( n28144 , n347632 );
not ( n28145 , n28144 );
or ( n28146 , n28143 , n28145 );
buf ( n348180 , n600 );
not ( n348181 , n348180 );
buf ( n348182 , n24091 );
not ( n28150 , n348182 );
or ( n348184 , n348181 , n28150 );
buf ( n348185 , n24092 );
buf ( n348186 , n23906 );
nand ( n348187 , n348185 , n348186 );
buf ( n348188 , n348187 );
buf ( n348189 , n348188 );
nand ( n28157 , n348184 , n348189 );
buf ( n348191 , n28157 );
buf ( n348192 , n348191 );
buf ( n348193 , n344018 );
nand ( n28161 , n348192 , n348193 );
buf ( n28162 , n28161 );
buf ( n348196 , n28162 );
nand ( n28164 , n28146 , n348196 );
buf ( n348198 , n28164 );
buf ( n348199 , n348198 );
and ( n348200 , n28141 , n348199 );
and ( n28168 , n348160 , n348173 );
or ( n348202 , n348200 , n28168 );
buf ( n348203 , n348202 );
buf ( n348204 , n348203 );
buf ( n348205 , n347639 );
not ( n348206 , n348205 );
xor ( n28174 , n347876 , n27570 );
buf ( n348208 , n28174 );
not ( n28176 , n348208 );
or ( n348210 , n348206 , n28176 );
buf ( n348211 , n347639 );
buf ( n348212 , n28174 );
or ( n348213 , n348211 , n348212 );
nand ( n348214 , n348210 , n348213 );
buf ( n348215 , n348214 );
buf ( n348216 , n348215 );
xor ( n348217 , n348204 , n348216 );
buf ( n348218 , n343531 );
not ( n28186 , n348218 );
buf ( n348220 , n347897 );
not ( n348221 , n348220 );
or ( n28189 , n28186 , n348221 );
and ( n28190 , n344484 , n602 );
not ( n348224 , n344484 );
and ( n348225 , n348224 , n343553 );
or ( n28193 , n28190 , n348225 );
buf ( n348227 , n28193 );
buf ( n348228 , n343592 );
nand ( n28196 , n348227 , n348228 );
buf ( n28197 , n28196 );
buf ( n348231 , n28197 );
nand ( n28199 , n28189 , n348231 );
buf ( n348233 , n28199 );
buf ( n348234 , n348233 );
and ( n348235 , n348217 , n348234 );
and ( n28203 , n348204 , n348216 );
or ( n348237 , n348235 , n28203 );
buf ( n348238 , n348237 );
or ( n28206 , n348156 , n348238 );
not ( n28207 , n28206 );
or ( n28208 , n28099 , n28207 );
nand ( n348242 , n348238 , n348156 );
nand ( n28210 , n28208 , n348242 );
not ( n348244 , n28210 );
buf ( n348245 , n348244 );
nand ( n28213 , n348128 , n348245 );
buf ( n348247 , n28213 );
buf ( n348248 , n348247 );
and ( n28216 , n348106 , n348248 );
buf ( n348250 , n348126 );
not ( n348251 , n348250 );
buf ( n348252 , n348244 );
nor ( n348253 , n348251 , n348252 );
buf ( n348254 , n348253 );
buf ( n348255 , n348254 );
nor ( n28223 , n28216 , n348255 );
buf ( n348257 , n28223 );
buf ( n348258 , n348257 );
nand ( n348259 , n348083 , n348258 );
buf ( n348260 , n348259 );
nand ( n28228 , n348079 , n348260 );
not ( n348262 , n28228 );
buf ( n348263 , n343530 );
not ( n348264 , n348263 );
and ( n28232 , n602 , n345454 );
not ( n28233 , n602 );
and ( n28234 , n28233 , n345451 );
or ( n28235 , n28232 , n28234 );
buf ( n348269 , n28235 );
not ( n28237 , n348269 );
or ( n28238 , n348264 , n28237 );
and ( n28239 , n602 , n25665 );
not ( n28240 , n602 );
buf ( n348274 , n25665 );
not ( n28242 , n348274 );
buf ( n348276 , n28242 );
and ( n28244 , n28240 , n348276 );
or ( n28245 , n28239 , n28244 );
buf ( n348279 , n28245 );
buf ( n348280 , n343592 );
nand ( n28248 , n348279 , n348280 );
buf ( n348282 , n28248 );
buf ( n348283 , n348282 );
nand ( n348284 , n28238 , n348283 );
buf ( n348285 , n348284 );
buf ( n348286 , n348285 );
buf ( n348287 , n599 );
buf ( n348288 , n600 );
or ( n348289 , n348287 , n348288 );
buf ( n348290 , n26233 );
nand ( n28258 , n348289 , n348290 );
buf ( n348292 , n28258 );
buf ( n348293 , n348292 );
buf ( n348294 , n599 );
buf ( n348295 , n600 );
and ( n28263 , n348294 , n348295 );
buf ( n348297 , n343953 );
nor ( n28265 , n28263 , n348297 );
buf ( n348299 , n28265 );
buf ( n348300 , n348299 );
nand ( n28268 , n348293 , n348300 );
buf ( n348302 , n28268 );
buf ( n348303 , n348302 );
not ( n28271 , n348303 );
buf ( n348305 , n23911 );
not ( n28273 , n348305 );
and ( n28274 , n14749 , n343953 );
not ( n28275 , n14749 );
and ( n348309 , n28275 , n598 );
or ( n348310 , n28274 , n348309 );
buf ( n348311 , n348310 );
not ( n348312 , n348311 );
or ( n348313 , n28273 , n348312 );
buf ( n348314 , n26233 );
buf ( n348315 , n343953 );
or ( n348316 , n348314 , n348315 );
buf ( n348317 , n347074 );
buf ( n348318 , n598 );
or ( n28286 , n348317 , n348318 );
nand ( n28287 , n348316 , n28286 );
buf ( n348321 , n28287 );
buf ( n28289 , n348321 );
buf ( n348323 , n343945 );
nand ( n348324 , n28289 , n348323 );
buf ( n348325 , n348324 );
buf ( n348326 , n348325 );
nand ( n348327 , n348313 , n348326 );
buf ( n348328 , n348327 );
buf ( n348329 , n348328 );
not ( n28297 , n348329 );
or ( n348331 , n28271 , n28297 );
buf ( n348332 , n348328 );
buf ( n348333 , n348302 );
or ( n348334 , n348332 , n348333 );
nand ( n28302 , n348331 , n348334 );
buf ( n28303 , n28302 );
buf ( n348337 , n28303 );
buf ( n348338 , n344015 );
not ( n28306 , n348338 );
buf ( n348340 , n600 );
not ( n28308 , n348340 );
buf ( n348342 , n346231 );
not ( n348343 , n348342 );
or ( n28311 , n28308 , n348343 );
buf ( n348345 , n14746 );
not ( n28313 , n348345 );
buf ( n348347 , n28313 );
buf ( n348348 , n348347 );
not ( n348349 , n348348 );
buf ( n28317 , n23906 );
nand ( n348351 , n348349 , n28317 );
buf ( n348352 , n348351 );
buf ( n348353 , n348352 );
nand ( n348354 , n28311 , n348353 );
buf ( n348355 , n348354 );
buf ( n348356 , n348355 );
not ( n28324 , n348356 );
or ( n28325 , n28306 , n28324 );
and ( n348359 , n14749 , n23906 );
not ( n348360 , n14749 );
and ( n348361 , n348360 , n600 );
or ( n28329 , n348359 , n348361 );
buf ( n348363 , n28329 );
buf ( n348364 , n344018 );
nand ( n28332 , n348363 , n348364 );
buf ( n348366 , n28332 );
buf ( n348367 , n348366 );
nand ( n348368 , n28325 , n348367 );
buf ( n348369 , n348368 );
not ( n348370 , n348369 );
buf ( n348371 , n26233 );
buf ( n348372 , n23911 );
nand ( n348373 , n348371 , n348372 );
buf ( n348374 , n348373 );
not ( n28342 , n348374 );
buf ( n348376 , n347074 );
buf ( n348377 , n600 );
and ( n348378 , n348376 , n348377 );
buf ( n348379 , n26233 );
buf ( n348380 , n23906 );
and ( n348381 , n348379 , n348380 );
nor ( n28349 , n348378 , n348381 );
buf ( n348383 , n28349 );
not ( n28351 , n348383 );
not ( n28352 , n344017 );
and ( n348386 , n28351 , n28352 );
and ( n348387 , n28329 , n344015 );
nor ( n348388 , n348386 , n348387 );
buf ( n348389 , n348388 );
buf ( n348390 , n601 );
buf ( n348391 , n602 );
or ( n28359 , n348390 , n348391 );
buf ( n348393 , n26233 );
nand ( n28361 , n28359 , n348393 );
buf ( n348395 , n28361 );
buf ( n28363 , n348395 );
buf ( n348397 , n601 );
buf ( n348398 , n602 );
and ( n28366 , n348397 , n348398 );
buf ( n348400 , n23906 );
nor ( n28368 , n28366 , n348400 );
buf ( n348402 , n28368 );
buf ( n348403 , n348402 );
nand ( n28371 , n28363 , n348403 );
buf ( n348405 , n28371 );
buf ( n348406 , n348405 );
nor ( n28374 , n348389 , n348406 );
buf ( n348408 , n28374 );
nor ( n28376 , n28342 , n348408 );
nor ( n348410 , n348370 , n28376 );
buf ( n348411 , n348410 );
xor ( n348412 , n348337 , n348411 );
buf ( n348413 , n344015 );
not ( n348414 , n348413 );
not ( n28382 , n600 );
not ( n348416 , n26159 );
or ( n28384 , n28382 , n348416 );
buf ( n348418 , n346205 );
buf ( n348419 , n23906 );
nand ( n28387 , n348418 , n348419 );
buf ( n28388 , n28387 );
nand ( n28389 , n28384 , n28388 );
buf ( n348423 , n28389 );
not ( n348424 , n348423 );
or ( n348425 , n348414 , n348424 );
buf ( n348426 , n348355 );
buf ( n348427 , n344018 );
nand ( n348428 , n348426 , n348427 );
buf ( n348429 , n348428 );
buf ( n348430 , n348429 );
nand ( n348431 , n348425 , n348430 );
buf ( n348432 , n348431 );
buf ( n348433 , n348432 );
xor ( n348434 , n348412 , n348433 );
buf ( n348435 , n348434 );
buf ( n348436 , n348435 );
xor ( n28404 , n348286 , n348436 );
buf ( n348438 , n348408 );
not ( n348439 , n348438 );
buf ( n348440 , n348374 );
not ( n348441 , n348440 );
and ( n28409 , n348439 , n348441 );
buf ( n348443 , n348408 );
buf ( n348444 , n348374 );
and ( n348445 , n348443 , n348444 );
nor ( n28413 , n28409 , n348445 );
buf ( n348447 , n28413 );
buf ( n348448 , n348447 );
not ( n28416 , n348448 );
buf ( n348450 , n348369 );
not ( n28418 , n348450 );
or ( n28419 , n28416 , n28418 );
buf ( n348453 , n348369 );
buf ( n348454 , n348447 );
or ( n348455 , n348453 , n348454 );
nand ( n28423 , n28419 , n348455 );
buf ( n348457 , n28423 );
buf ( n348458 , n348457 );
buf ( n348459 , n343530 );
not ( n28427 , n348459 );
buf ( n348461 , n28245 );
not ( n28429 , n348461 );
or ( n28430 , n28427 , n28429 );
and ( n348464 , n602 , n346202 );
not ( n28432 , n602 );
and ( n28433 , n28432 , n346199 );
or ( n348467 , n348464 , n28433 );
buf ( n348468 , n348467 );
buf ( n348469 , n343592 );
nand ( n28437 , n348468 , n348469 );
buf ( n348471 , n28437 );
buf ( n348472 , n348471 );
nand ( n348473 , n28430 , n348472 );
buf ( n348474 , n348473 );
buf ( n348475 , n348474 );
xor ( n28443 , n348458 , n348475 );
xor ( n28444 , n348405 , n348388 );
buf ( n348478 , n28444 );
buf ( n348479 , n344014 );
buf ( n348480 , n347074 );
nor ( n28448 , n348479 , n348480 );
buf ( n348482 , n28448 );
buf ( n348483 , n348482 );
and ( n348484 , n14749 , n343553 );
not ( n28452 , n14749 );
and ( n348486 , n28452 , n602 );
or ( n348487 , n348484 , n348486 );
buf ( n348488 , n348487 );
buf ( n348489 , n343530 );
and ( n348490 , n348488 , n348489 );
and ( n28458 , n602 , n347074 );
not ( n28459 , n602 );
and ( n28460 , n28459 , n26233 );
nor ( n28461 , n28458 , n28460 );
buf ( n348495 , n28461 );
buf ( n28463 , n343592 );
not ( n28464 , n28463 );
buf ( n348498 , n28464 );
buf ( n348499 , n348498 );
nor ( n28467 , n348495 , n348499 );
buf ( n348501 , n28467 );
buf ( n348502 , n348501 );
nor ( n348503 , n348490 , n348502 );
buf ( n348504 , n348503 );
buf ( n348505 , n348504 );
buf ( n348506 , n603 );
buf ( n348507 , n604 );
or ( n28475 , n348506 , n348507 );
buf ( n348509 , n26233 );
nand ( n28477 , n28475 , n348509 );
buf ( n348511 , n28477 );
buf ( n28479 , n348511 );
buf ( n348513 , n603 );
buf ( n348514 , n604 );
nand ( n348515 , n348513 , n348514 );
buf ( n348516 , n348515 );
buf ( n348517 , n348516 );
buf ( n348518 , n602 );
nand ( n348519 , n28479 , n348517 , n348518 );
buf ( n348520 , n348519 );
buf ( n348521 , n348520 );
nor ( n28489 , n348505 , n348521 );
buf ( n348523 , n28489 );
buf ( n348524 , n348523 );
xor ( n28492 , n348483 , n348524 );
not ( n348526 , n348487 );
not ( n28494 , n343592 );
or ( n28495 , n348526 , n28494 );
buf ( n348529 , n602 );
buf ( n348530 , n346231 );
and ( n28498 , n348529 , n348530 );
not ( n28499 , n348529 );
buf ( n348533 , n346179 );
and ( n28501 , n28499 , n348533 );
nor ( n348535 , n28498 , n28501 );
buf ( n348536 , n348535 );
buf ( n348537 , n343530 );
not ( n348538 , n348537 );
buf ( n348539 , n348538 );
or ( n28507 , n348536 , n348539 );
nand ( n348541 , n28495 , n28507 );
buf ( n348542 , n348541 );
and ( n348543 , n28492 , n348542 );
and ( n28511 , n348483 , n348524 );
or ( n28512 , n348543 , n28511 );
buf ( n348546 , n28512 );
buf ( n28514 , n348546 );
xor ( n28515 , n348478 , n28514 );
buf ( n348549 , n343530 );
not ( n348550 , n348549 );
buf ( n348551 , n348467 );
not ( n348552 , n348551 );
or ( n28520 , n348550 , n348552 );
buf ( n348554 , n348536 );
not ( n28522 , n348554 );
buf ( n348556 , n343592 );
nand ( n28524 , n28522 , n348556 );
buf ( n348558 , n28524 );
buf ( n348559 , n348558 );
nand ( n348560 , n28520 , n348559 );
buf ( n348561 , n348560 );
buf ( n348562 , n348561 );
and ( n348563 , n28515 , n348562 );
and ( n348564 , n348478 , n28514 );
or ( n348565 , n348563 , n348564 );
buf ( n348566 , n348565 );
buf ( n348567 , n348566 );
and ( n348568 , n28443 , n348567 );
and ( n28536 , n348458 , n348475 );
or ( n348570 , n348568 , n28536 );
buf ( n348571 , n348570 );
buf ( n348572 , n348571 );
and ( n28540 , n28404 , n348572 );
and ( n348574 , n348286 , n348436 );
or ( n348575 , n28540 , n348574 );
buf ( n348576 , n348575 );
buf ( n348577 , n348576 );
buf ( n348578 , n607 );
not ( n28546 , n348578 );
buf ( n348580 , n606 );
buf ( n348581 , n344185 );
and ( n28549 , n348580 , n348581 );
not ( n348583 , n348580 );
buf ( n348584 , n344185 );
not ( n28552 , n348584 );
buf ( n348586 , n28552 );
buf ( n348587 , n348586 );
and ( n28555 , n348583 , n348587 );
nor ( n28556 , n28549 , n28555 );
buf ( n348590 , n28556 );
buf ( n348591 , n348590 );
not ( n28559 , n348591 );
or ( n348593 , n28546 , n28559 );
buf ( n348594 , n606 );
buf ( n348595 , n24059 );
not ( n28563 , n348595 );
buf ( n348597 , n28563 );
buf ( n28565 , n348597 );
and ( n28566 , n348594 , n28565 );
not ( n348600 , n348594 );
buf ( n348601 , n26331 );
and ( n28569 , n348600 , n348601 );
nor ( n28570 , n28566 , n28569 );
buf ( n348604 , n28570 );
buf ( n348605 , n348604 );
buf ( n348606 , n344454 );
nand ( n28574 , n348605 , n348606 );
buf ( n348608 , n28574 );
buf ( n348609 , n348608 );
nand ( n28577 , n348593 , n348609 );
buf ( n348611 , n28577 );
buf ( n28579 , n348611 );
xor ( n28580 , n348577 , n28579 );
buf ( n348614 , n343531 );
not ( n348615 , n348614 );
not ( n28583 , n602 );
not ( n348617 , n345175 );
or ( n348618 , n28583 , n348617 );
buf ( n348619 , n25403 );
buf ( n348620 , n343553 );
nand ( n348621 , n348619 , n348620 );
buf ( n348622 , n348621 );
nand ( n348623 , n348618 , n348622 );
buf ( n348624 , n348623 );
not ( n28592 , n348624 );
or ( n28593 , n348615 , n28592 );
buf ( n348627 , n28235 );
buf ( n348628 , n343592 );
nand ( n348629 , n348627 , n348628 );
buf ( n348630 , n348629 );
buf ( n348631 , n348630 );
nand ( n28599 , n28593 , n348631 );
buf ( n348633 , n28599 );
buf ( n348634 , n348633 );
buf ( n348635 , n23911 );
not ( n348636 , n348635 );
buf ( n348637 , n598 );
not ( n348638 , n348637 );
buf ( n348639 , n348347 );
not ( n348640 , n348639 );
or ( n28608 , n348638 , n348640 );
buf ( n28609 , n14746 );
buf ( n348643 , n343953 );
nand ( n348644 , n28609 , n348643 );
buf ( n348645 , n348644 );
buf ( n348646 , n348645 );
nand ( n28614 , n28608 , n348646 );
buf ( n348648 , n28614 );
buf ( n348649 , n348648 );
not ( n28617 , n348649 );
or ( n348651 , n348636 , n28617 );
buf ( n348652 , n348310 );
buf ( n348653 , n343945 );
nand ( n348654 , n348652 , n348653 );
buf ( n348655 , n348654 );
buf ( n348656 , n348655 );
nand ( n28624 , n348651 , n348656 );
buf ( n348658 , n28624 );
buf ( n348659 , n26233 );
buf ( n348660 , n343863 );
nand ( n348661 , n348659 , n348660 );
buf ( n348662 , n348661 );
buf ( n348663 , n348662 );
not ( n348664 , n348663 );
buf ( n348665 , n348328 );
not ( n28633 , n348665 );
buf ( n348667 , n348302 );
nor ( n348668 , n28633 , n348667 );
buf ( n348669 , n348668 );
buf ( n348670 , n348669 );
nor ( n348671 , n348664 , n348670 );
buf ( n348672 , n348671 );
xor ( n28640 , n348658 , n348672 );
buf ( n348674 , n28640 );
not ( n28642 , n28389 );
not ( n348676 , n28642 );
not ( n348677 , n344017 );
and ( n28645 , n348676 , n348677 );
buf ( n28646 , n600 );
not ( n28647 , n28646 );
buf ( n28648 , n25665 );
not ( n28649 , n28648 );
or ( n28650 , n28647 , n28649 );
buf ( n348684 , n348276 );
buf ( n348685 , n23906 );
nand ( n28653 , n348684 , n348685 );
buf ( n348687 , n28653 );
buf ( n348688 , n348687 );
nand ( n28656 , n28650 , n348688 );
buf ( n348690 , n28656 );
and ( n28658 , n348690 , n344015 );
nor ( n348692 , n28645 , n28658 );
buf ( n348693 , n348692 );
xor ( n348694 , n348674 , n348693 );
xor ( n28662 , n348337 , n348411 );
and ( n28663 , n28662 , n348433 );
and ( n28664 , n348337 , n348411 );
or ( n348698 , n28663 , n28664 );
buf ( n348699 , n348698 );
buf ( n348700 , n348699 );
xor ( n348701 , n348694 , n348700 );
buf ( n348702 , n348701 );
buf ( n348703 , n348702 );
xor ( n348704 , n348634 , n348703 );
buf ( n348705 , n344338 );
not ( n28673 , n348705 );
buf ( n348707 , n604 );
not ( n348708 , n348707 );
buf ( n348709 , n24091 );
not ( n348710 , n348709 );
or ( n348711 , n348708 , n348710 );
buf ( n348712 , n344155 );
buf ( n348713 , n23530 );
nand ( n348714 , n348712 , n348713 );
buf ( n348715 , n348714 );
buf ( n348716 , n348715 );
nand ( n348717 , n348711 , n348716 );
buf ( n348718 , n348717 );
buf ( n348719 , n348718 );
not ( n348720 , n348719 );
or ( n348721 , n28673 , n348720 );
buf ( n348722 , n604 );
not ( n28690 , n348722 );
buf ( n348724 , n24109 );
not ( n28692 , n348724 );
or ( n28693 , n28690 , n28692 );
buf ( n348727 , n23530 );
buf ( n348728 , n24108 );
nand ( n28696 , n348727 , n348728 );
buf ( n348730 , n28696 );
buf ( n348731 , n348730 );
nand ( n28699 , n28693 , n348731 );
buf ( n348733 , n28699 );
buf ( n28701 , n348733 );
buf ( n348735 , n344397 );
nand ( n348736 , n28701 , n348735 );
buf ( n348737 , n348736 );
buf ( n348738 , n348737 );
nand ( n348739 , n348721 , n348738 );
buf ( n348740 , n348739 );
buf ( n348741 , n348740 );
xor ( n348742 , n348704 , n348741 );
buf ( n348743 , n348742 );
buf ( n348744 , n348743 );
xnor ( n28712 , n28580 , n348744 );
buf ( n28713 , n28712 );
buf ( n348747 , n28713 );
and ( n28715 , n607 , n348604 );
buf ( n348749 , n344445 );
not ( n28717 , n348749 );
buf ( n348751 , n344155 );
not ( n28719 , n348751 );
or ( n28720 , n28717 , n28719 );
buf ( n348754 , n24091 );
buf ( n348755 , n606 );
nand ( n28723 , n348754 , n348755 );
buf ( n348757 , n28723 );
buf ( n348758 , n348757 );
nand ( n28726 , n28720 , n348758 );
buf ( n348760 , n28726 );
and ( n28728 , n348760 , n344454 );
nor ( n28729 , n28715 , n28728 );
buf ( n348763 , n28729 );
buf ( n348764 , n604 );
buf ( n348765 , n25403 );
and ( n348766 , n348764 , n348765 );
not ( n348767 , n348764 );
buf ( n348768 , n25403 );
not ( n348769 , n348768 );
buf ( n348770 , n348769 );
buf ( n348771 , n348770 );
and ( n348772 , n348767 , n348771 );
nor ( n348773 , n348766 , n348772 );
buf ( n348774 , n348773 );
buf ( n348775 , n348774 );
not ( n348776 , n348775 );
buf ( n348777 , n348776 );
buf ( n348778 , n348777 );
not ( n28746 , n348778 );
buf ( n348780 , n344397 );
not ( n28748 , n348780 );
buf ( n348782 , n28748 );
buf ( n348783 , n348782 );
not ( n28751 , n348783 );
and ( n28752 , n28746 , n28751 );
buf ( n348786 , n348733 );
buf ( n348787 , n344338 );
and ( n28755 , n348786 , n348787 );
nor ( n28756 , n28752 , n28755 );
buf ( n348790 , n28756 );
buf ( n348791 , n348790 );
nand ( n348792 , n348763 , n348791 );
buf ( n348793 , n348792 );
buf ( n348794 , n348793 );
xor ( n348795 , n348286 , n348436 );
xor ( n348796 , n348795 , n348572 );
buf ( n348797 , n348796 );
buf ( n348798 , n348797 );
and ( n348799 , n348794 , n348798 );
buf ( n348800 , n28729 );
buf ( n348801 , n348790 );
nor ( n348802 , n348800 , n348801 );
buf ( n348803 , n348802 );
buf ( n348804 , n348803 );
nor ( n28772 , n348799 , n348804 );
buf ( n28773 , n28772 );
buf ( n348807 , n28773 );
nand ( n348808 , n348747 , n348807 );
buf ( n348809 , n348808 );
buf ( n348810 , n348809 );
buf ( n348811 , n24108 );
not ( n348812 , n348811 );
buf ( n348813 , n344445 );
not ( n348814 , n348813 );
and ( n348815 , n348812 , n348814 );
buf ( n348816 , n24108 );
buf ( n348817 , n344445 );
and ( n28785 , n348816 , n348817 );
nor ( n28786 , n348815 , n28785 );
buf ( n348820 , n28786 );
buf ( n348821 , n348820 );
not ( n28789 , n348821 );
buf ( n348823 , n344631 );
not ( n28791 , n348823 );
and ( n28792 , n28789 , n28791 );
buf ( n348826 , n348760 );
buf ( n348827 , n607 );
and ( n348828 , n348826 , n348827 );
nor ( n348829 , n28792 , n348828 );
buf ( n348830 , n348829 );
not ( n28798 , n348830 );
buf ( n348832 , n344338 );
not ( n28800 , n348832 );
buf ( n348834 , n348774 );
not ( n348835 , n348834 );
or ( n28803 , n28800 , n348835 );
and ( n348837 , n604 , n345454 );
not ( n28805 , n604 );
and ( n348839 , n28805 , n345451 );
or ( n28807 , n348837 , n348839 );
buf ( n348841 , n28807 );
buf ( n348842 , n344397 );
nand ( n348843 , n348841 , n348842 );
buf ( n348844 , n348843 );
buf ( n348845 , n348844 );
nand ( n348846 , n28803 , n348845 );
buf ( n348847 , n348846 );
buf ( n348848 , n348847 );
not ( n28816 , n348848 );
buf ( n28817 , n28816 );
not ( n28818 , n28817 );
or ( n28819 , n28798 , n28818 );
xor ( n348853 , n348458 , n348475 );
xor ( n28821 , n348853 , n348567 );
buf ( n348855 , n28821 );
nand ( n28823 , n28819 , n348855 );
buf ( n348857 , n348830 );
not ( n348858 , n348857 );
buf ( n28826 , n348847 );
nand ( n28827 , n348858 , n28826 );
buf ( n348861 , n28827 );
nand ( n348862 , n28823 , n348861 );
buf ( n348863 , n348862 );
not ( n348864 , n348863 );
xor ( n348865 , n348797 , n348790 );
xnor ( n348866 , n348865 , n28729 );
buf ( n348867 , n348866 );
nand ( n348868 , n348864 , n348867 );
buf ( n348869 , n348868 );
not ( n348870 , n348869 );
xor ( n28838 , n348478 , n28514 );
xor ( n28839 , n28838 , n348562 );
buf ( n348873 , n28839 );
buf ( n348874 , n348873 );
buf ( n348875 , n344338 );
not ( n348876 , n348875 );
buf ( n348877 , n28807 );
not ( n28845 , n348877 );
or ( n348879 , n348876 , n28845 );
buf ( n348880 , n344397 );
buf ( n348881 , n604 );
not ( n28849 , n348881 );
buf ( n348883 , n25665 );
not ( n348884 , n348883 );
or ( n28852 , n28849 , n348884 );
buf ( n348886 , n348276 );
buf ( n348887 , n23530 );
nand ( n28855 , n348886 , n348887 );
buf ( n28856 , n28855 );
buf ( n348890 , n28856 );
nand ( n28858 , n28852 , n348890 );
buf ( n348892 , n28858 );
buf ( n348893 , n348892 );
nand ( n28861 , n348880 , n348893 );
buf ( n348895 , n28861 );
buf ( n348896 , n348895 );
nand ( n28864 , n348879 , n348896 );
buf ( n348898 , n28864 );
buf ( n348899 , n348898 );
xor ( n28867 , n348874 , n348899 );
xor ( n28868 , n348483 , n348524 );
xor ( n348902 , n28868 , n348542 );
buf ( n348903 , n348902 );
buf ( n348904 , n348903 );
not ( n348905 , n348904 );
buf ( n348906 , n604 );
not ( n28874 , n348906 );
buf ( n348908 , n346202 );
not ( n348909 , n348908 );
or ( n28877 , n28874 , n348909 );
buf ( n348911 , n346199 );
buf ( n348912 , n23530 );
nand ( n28880 , n348911 , n348912 );
buf ( n28881 , n28880 );
buf ( n348915 , n28881 );
nand ( n28883 , n28877 , n348915 );
buf ( n348917 , n28883 );
buf ( n348918 , n348917 );
not ( n28886 , n348918 );
buf ( n348920 , n28886 );
buf ( n348921 , n348920 );
not ( n28889 , n348921 );
buf ( n348923 , n348782 );
not ( n348924 , n348923 );
and ( n28892 , n28889 , n348924 );
buf ( n348926 , n348892 );
buf ( n348927 , n344338 );
and ( n28895 , n348926 , n348927 );
nor ( n348929 , n28892 , n28895 );
buf ( n348930 , n348929 );
buf ( n348931 , n348930 );
not ( n28899 , n348931 );
buf ( n348933 , n28899 );
buf ( n348934 , n348933 );
not ( n28902 , n348934 );
or ( n348936 , n348905 , n28902 );
buf ( n348937 , n604 );
not ( n348938 , n348937 );
buf ( n348939 , n346231 );
not ( n28907 , n348939 );
or ( n348941 , n348938 , n28907 );
buf ( n348942 , n346179 );
buf ( n348943 , n23530 );
nand ( n28911 , n348942 , n348943 );
buf ( n348945 , n28911 );
buf ( n28913 , n348945 );
nand ( n28914 , n348941 , n28913 );
buf ( n28915 , n28914 );
buf ( n348949 , n28915 );
not ( n28917 , n348949 );
buf ( n348951 , n28917 );
buf ( n348952 , n348951 );
not ( n28920 , n348952 );
buf ( n348954 , n348782 );
not ( n28922 , n348954 );
and ( n28923 , n28920 , n28922 );
buf ( n348957 , n348917 );
buf ( n348958 , n344338 );
and ( n348959 , n348957 , n348958 );
nor ( n348960 , n28923 , n348959 );
buf ( n348961 , n348960 );
buf ( n348962 , n348961 );
not ( n28930 , n348962 );
buf ( n348964 , n28930 );
buf ( n348965 , n348964 );
not ( n28933 , n348965 );
buf ( n348967 , n348504 );
buf ( n348968 , n348520 );
xor ( n28936 , n348967 , n348968 );
buf ( n348970 , n28936 );
buf ( n348971 , n348970 );
not ( n348972 , n348971 );
or ( n28940 , n28933 , n348972 );
buf ( n348974 , n348970 );
not ( n348975 , n348974 );
buf ( n348976 , n348975 );
buf ( n348977 , n348976 );
not ( n348978 , n348977 );
buf ( n348979 , n348961 );
not ( n348980 , n348979 );
or ( n348981 , n348978 , n348980 );
buf ( n348982 , n347074 );
buf ( n348983 , n348539 );
nor ( n348984 , n348982 , n348983 );
buf ( n348985 , n348984 );
buf ( n348986 , n348985 );
buf ( n348987 , n604 );
not ( n348988 , n348987 );
buf ( n348989 , n346254 );
not ( n28957 , n348989 );
or ( n348991 , n348988 , n28957 );
buf ( n348992 , n14749 );
buf ( n348993 , n23530 );
nand ( n348994 , n348992 , n348993 );
buf ( n348995 , n348994 );
buf ( n348996 , n348995 );
nand ( n348997 , n348991 , n348996 );
buf ( n348998 , n348997 );
buf ( n348999 , n348998 );
buf ( n349000 , n344338 );
and ( n349001 , n348999 , n349000 );
buf ( n349002 , n347074 );
buf ( n349003 , n604 );
and ( n28971 , n349002 , n349003 );
buf ( n349005 , n26233 );
buf ( n349006 , n23530 );
and ( n349007 , n349005 , n349006 );
nor ( n349008 , n28971 , n349007 );
buf ( n349009 , n349008 );
buf ( n349010 , n349009 );
buf ( n349011 , n348782 );
nor ( n28979 , n349010 , n349011 );
buf ( n349013 , n28979 );
buf ( n349014 , n349013 );
nor ( n28982 , n349001 , n349014 );
buf ( n349016 , n28982 );
buf ( n349017 , n349016 );
buf ( n349018 , n605 );
buf ( n349019 , n606 );
or ( n28987 , n349018 , n349019 );
buf ( n349021 , n26233 );
nand ( n28989 , n28987 , n349021 );
buf ( n349023 , n28989 );
buf ( n349024 , n349023 );
buf ( n349025 , n605 );
buf ( n349026 , n606 );
and ( n28994 , n349025 , n349026 );
buf ( n349028 , n23530 );
nor ( n28996 , n28994 , n349028 );
buf ( n349030 , n28996 );
buf ( n349031 , n349030 );
and ( n28999 , n349024 , n349031 );
buf ( n349033 , n28999 );
buf ( n349034 , n349033 );
not ( n29002 , n349034 );
buf ( n29003 , n29002 );
buf ( n349037 , n29003 );
nor ( n29005 , n349017 , n349037 );
buf ( n349039 , n29005 );
buf ( n349040 , n349039 );
xor ( n29008 , n348986 , n349040 );
buf ( n349042 , n344338 );
not ( n29010 , n349042 );
buf ( n349044 , n28915 );
not ( n29012 , n349044 );
or ( n29013 , n29010 , n29012 );
buf ( n349047 , n348998 );
buf ( n349048 , n344397 );
nand ( n29016 , n349047 , n349048 );
buf ( n349050 , n29016 );
buf ( n349051 , n349050 );
nand ( n29019 , n29013 , n349051 );
buf ( n349053 , n29019 );
buf ( n349054 , n349053 );
and ( n29022 , n29008 , n349054 );
and ( n29023 , n348986 , n349040 );
or ( n29024 , n29022 , n29023 );
buf ( n349058 , n29024 );
buf ( n349059 , n349058 );
nand ( n29027 , n348981 , n349059 );
buf ( n349061 , n29027 );
buf ( n349062 , n349061 );
nand ( n29030 , n28940 , n349062 );
buf ( n349064 , n29030 );
buf ( n349065 , n349064 );
buf ( n349066 , n348903 );
not ( n349067 , n349066 );
buf ( n349068 , n348930 );
nand ( n349069 , n349067 , n349068 );
buf ( n349070 , n349069 );
buf ( n349071 , n349070 );
nand ( n349072 , n349065 , n349071 );
buf ( n349073 , n349072 );
buf ( n349074 , n349073 );
nand ( n29042 , n348936 , n349074 );
buf ( n29043 , n29042 );
buf ( n349077 , n29043 );
and ( n29045 , n28867 , n349077 );
and ( n349079 , n348874 , n348899 );
or ( n349080 , n29045 , n349079 );
buf ( n349081 , n349080 );
buf ( n349082 , n349081 );
buf ( n349083 , n607 );
not ( n349084 , n349083 );
and ( n349085 , n606 , n25665 );
not ( n29053 , n606 );
and ( n349087 , n29053 , n348276 );
or ( n29055 , n349085 , n349087 );
buf ( n349089 , n29055 );
not ( n349090 , n349089 );
or ( n29058 , n349084 , n349090 );
buf ( n349092 , n606 );
not ( n349093 , n349092 );
buf ( n349094 , n346202 );
not ( n349095 , n349094 );
or ( n349096 , n349093 , n349095 );
buf ( n349097 , n346205 );
buf ( n349098 , n344445 );
nand ( n29066 , n349097 , n349098 );
buf ( n349100 , n29066 );
buf ( n349101 , n349100 );
nand ( n29069 , n349096 , n349101 );
buf ( n349103 , n29069 );
buf ( n349104 , n349103 );
buf ( n349105 , n344454 );
nand ( n29073 , n349104 , n349105 );
buf ( n349107 , n29073 );
buf ( n349108 , n349107 );
nand ( n29076 , n29058 , n349108 );
buf ( n349110 , n29076 );
buf ( n29078 , n349110 );
xor ( n29079 , n348986 , n349040 );
xor ( n29080 , n29079 , n349054 );
buf ( n349114 , n29080 );
buf ( n349115 , n349114 );
nor ( n349116 , n29078 , n349115 );
buf ( n349117 , n349116 );
buf ( n349118 , n349117 );
buf ( n349119 , n349016 );
buf ( n349120 , n29003 );
and ( n349121 , n349119 , n349120 );
not ( n29089 , n349119 );
buf ( n349123 , n349033 );
and ( n349124 , n29089 , n349123 );
nor ( n349125 , n349121 , n349124 );
buf ( n349126 , n349125 );
buf ( n349127 , n349126 );
buf ( n349128 , n344338 );
not ( n29096 , n349128 );
buf ( n29097 , n29096 );
buf ( n349131 , n29097 );
buf ( n349132 , n347074 );
nor ( n29100 , n349131 , n349132 );
buf ( n349134 , n29100 );
buf ( n349135 , n349134 );
not ( n29103 , n26233 );
not ( n29104 , n344631 );
and ( n29105 , n29103 , n29104 );
buf ( n349139 , n606 );
not ( n29107 , n349139 );
buf ( n349141 , n347774 );
not ( n349142 , n349141 );
or ( n349143 , n29107 , n349142 );
buf ( n349144 , n14749 );
buf ( n349145 , n344445 );
nand ( n29113 , n349144 , n349145 );
buf ( n349147 , n29113 );
buf ( n349148 , n349147 );
nand ( n349149 , n349143 , n349148 );
buf ( n349150 , n349149 );
and ( n29118 , n607 , n349150 );
nor ( n349152 , n29105 , n29118 );
buf ( n349153 , n349152 );
nor ( n29121 , n26232 , n344452 );
buf ( n349155 , n29121 );
not ( n349156 , n349155 );
buf ( n349157 , n606 );
nand ( n349158 , n349156 , n349157 );
buf ( n349159 , n349158 );
buf ( n349160 , n349159 );
nor ( n349161 , n349153 , n349160 );
buf ( n349162 , n349161 );
buf ( n349163 , n349162 );
xor ( n29131 , n349135 , n349163 );
not ( n29132 , n349150 );
not ( n349166 , n344454 );
or ( n349167 , n29132 , n349166 );
buf ( n349168 , n346231 );
buf ( n349169 , n606 );
and ( n349170 , n349168 , n349169 );
buf ( n349171 , n346179 );
buf ( n349172 , n344445 );
and ( n349173 , n349171 , n349172 );
nor ( n349174 , n349170 , n349173 );
buf ( n349175 , n349174 );
or ( n349176 , n349175 , n344452 );
nand ( n349177 , n349167 , n349176 );
buf ( n349178 , n349177 );
and ( n349179 , n29131 , n349178 );
and ( n349180 , n349135 , n349163 );
or ( n29148 , n349179 , n349180 );
buf ( n349182 , n29148 );
buf ( n349183 , n349182 );
xor ( n349184 , n349127 , n349183 );
buf ( n349185 , n607 );
not ( n29153 , n349185 );
buf ( n349187 , n349103 );
not ( n349188 , n349187 );
or ( n349189 , n29153 , n349188 );
buf ( n349190 , n349175 );
not ( n349191 , n349190 );
buf ( n349192 , n344454 );
nand ( n29160 , n349191 , n349192 );
buf ( n29161 , n29160 );
buf ( n349195 , n29161 );
nand ( n29163 , n349189 , n349195 );
buf ( n349197 , n29163 );
buf ( n29165 , n349197 );
and ( n29166 , n349184 , n29165 );
and ( n349200 , n349127 , n349183 );
or ( n349201 , n29166 , n349200 );
buf ( n349202 , n349201 );
buf ( n349203 , n349202 );
not ( n29171 , n349203 );
buf ( n349205 , n29171 );
buf ( n349206 , n349205 );
or ( n349207 , n349118 , n349206 );
buf ( n349208 , n349110 );
buf ( n349209 , n349114 );
nand ( n29177 , n349208 , n349209 );
buf ( n349211 , n29177 );
buf ( n349212 , n349211 );
nand ( n349213 , n349207 , n349212 );
buf ( n349214 , n349213 );
buf ( n349215 , n349214 );
buf ( n349216 , n348970 );
buf ( n349217 , n348964 );
xor ( n349218 , n349216 , n349217 );
buf ( n349219 , n349058 );
xnor ( n29187 , n349218 , n349219 );
buf ( n349221 , n29187 );
buf ( n349222 , n29055 );
not ( n349223 , n349222 );
buf ( n349224 , n349223 );
buf ( n349225 , n349224 );
not ( n349226 , n349225 );
buf ( n349227 , n344631 );
not ( n29195 , n349227 );
and ( n29196 , n349226 , n29195 );
buf ( n349230 , n606 );
not ( n29198 , n349230 );
buf ( n349232 , n345454 );
not ( n29200 , n349232 );
or ( n29201 , n29198 , n29200 );
buf ( n349235 , n345451 );
buf ( n349236 , n344445 );
nand ( n349237 , n349235 , n349236 );
buf ( n349238 , n349237 );
buf ( n349239 , n349238 );
nand ( n349240 , n29201 , n349239 );
buf ( n349241 , n349240 );
buf ( n349242 , n349241 );
buf ( n349243 , n607 );
and ( n349244 , n349242 , n349243 );
nor ( n29212 , n29196 , n349244 );
buf ( n29213 , n29212 );
nand ( n349247 , n349221 , n29213 );
buf ( n349248 , n349247 );
nand ( n349249 , n349215 , n349248 );
buf ( n349250 , n349249 );
buf ( n349251 , n349250 );
buf ( n349252 , n349221 );
not ( n349253 , n349252 );
buf ( n349254 , n349253 );
buf ( n349255 , n29213 );
not ( n349256 , n349255 );
buf ( n349257 , n349256 );
nand ( n29225 , n349254 , n349257 );
buf ( n349259 , n29225 );
nand ( n29227 , n349251 , n349259 );
buf ( n349261 , n29227 );
buf ( n349262 , n349261 );
buf ( n349263 , n348903 );
buf ( n349264 , n348933 );
xor ( n349265 , n349263 , n349264 );
buf ( n349266 , n349064 );
xnor ( n29234 , n349265 , n349266 );
buf ( n349268 , n29234 );
buf ( n349269 , n349268 );
buf ( n349270 , n606 );
not ( n29238 , n349270 );
buf ( n349272 , n348770 );
not ( n349273 , n349272 );
or ( n29241 , n29238 , n349273 );
buf ( n349275 , n25403 );
buf ( n349276 , n344445 );
nand ( n29244 , n349275 , n349276 );
buf ( n349278 , n29244 );
buf ( n349279 , n349278 );
nand ( n29247 , n29241 , n349279 );
buf ( n349281 , n29247 );
buf ( n349282 , n349281 );
buf ( n349283 , n607 );
and ( n349284 , n349282 , n349283 );
buf ( n349285 , n349241 );
not ( n29253 , n349285 );
buf ( n349287 , n344631 );
nor ( n29255 , n29253 , n349287 );
buf ( n349289 , n29255 );
buf ( n349290 , n349289 );
nor ( n349291 , n349284 , n349290 );
buf ( n349292 , n349291 );
buf ( n29260 , n349292 );
nand ( n29261 , n349269 , n29260 );
buf ( n29262 , n29261 );
buf ( n349296 , n29262 );
nand ( n29264 , n349262 , n349296 );
buf ( n349298 , n29264 );
buf ( n349299 , n349298 );
buf ( n349300 , n349292 );
not ( n29268 , n349300 );
buf ( n349302 , n29268 );
buf ( n349303 , n349302 );
buf ( n349304 , n349268 );
not ( n29272 , n349304 );
buf ( n349306 , n29272 );
buf ( n349307 , n349306 );
nand ( n349308 , n349303 , n349307 );
buf ( n349309 , n349308 );
buf ( n349310 , n349309 );
and ( n29278 , n349299 , n349310 );
buf ( n349312 , n29278 );
buf ( n349313 , n349312 );
buf ( n349314 , n348820 );
buf ( n349315 , n344452 );
or ( n29283 , n349314 , n349315 );
buf ( n349317 , n349281 );
buf ( n349318 , n344454 );
nand ( n29286 , n349317 , n349318 );
buf ( n29287 , n29286 );
buf ( n349321 , n29287 );
nand ( n29289 , n29283 , n349321 );
buf ( n29290 , n29289 );
buf ( n349324 , n29290 );
xor ( n349325 , n348874 , n348899 );
xor ( n29293 , n349325 , n349077 );
buf ( n349327 , n29293 );
buf ( n349328 , n349327 );
nor ( n349329 , n349324 , n349328 );
buf ( n349330 , n349329 );
buf ( n349331 , n349330 );
or ( n349332 , n349313 , n349331 );
buf ( n349333 , n349327 );
buf ( n349334 , n29290 );
nand ( n349335 , n349333 , n349334 );
buf ( n349336 , n349335 );
buf ( n349337 , n349336 );
nand ( n349338 , n349332 , n349337 );
buf ( n349339 , n349338 );
buf ( n349340 , n349339 );
xor ( n29308 , n349082 , n349340 );
buf ( n349342 , n348830 );
not ( n349343 , n349342 );
buf ( n349344 , n348855 );
buf ( n349345 , n348847 );
and ( n29313 , n349344 , n349345 );
not ( n29314 , n349344 );
buf ( n349348 , n28817 );
and ( n29316 , n29314 , n349348 );
nor ( n29317 , n29313 , n29316 );
buf ( n349351 , n29317 );
buf ( n349352 , n349351 );
not ( n29320 , n349352 );
or ( n29321 , n349343 , n29320 );
buf ( n349355 , n349351 );
buf ( n349356 , n348830 );
or ( n29324 , n349355 , n349356 );
nand ( n29325 , n29321 , n29324 );
buf ( n349359 , n29325 );
buf ( n349360 , n349359 );
and ( n349361 , n29308 , n349360 );
and ( n29329 , n349082 , n349340 );
or ( n29330 , n349361 , n29329 );
buf ( n349364 , n29330 );
not ( n349365 , n349364 );
or ( n349366 , n348870 , n349365 );
buf ( n349367 , n348866 );
not ( n349368 , n349367 );
buf ( n349369 , n349368 );
buf ( n349370 , n349369 );
buf ( n349371 , n348862 );
nand ( n349372 , n349370 , n349371 );
buf ( n349373 , n349372 );
nand ( n349374 , n349366 , n349373 );
buf ( n349375 , n349374 );
nand ( n29343 , n348810 , n349375 );
buf ( n29344 , n29343 );
buf ( n349378 , n29344 );
buf ( n29346 , n28713 );
not ( n29347 , n29346 );
buf ( n29348 , n29347 );
buf ( n29349 , n29348 );
buf ( n349383 , n28773 );
not ( n349384 , n349383 );
buf ( n349385 , n349384 );
buf ( n349386 , n349385 );
nand ( n349387 , n29349 , n349386 );
buf ( n349388 , n349387 );
buf ( n349389 , n349388 );
nand ( n349390 , n349378 , n349389 );
buf ( n349391 , n349390 );
not ( n29359 , n349391 );
xor ( n29360 , n348634 , n348703 );
and ( n349394 , n29360 , n348741 );
and ( n29362 , n348634 , n348703 );
or ( n29363 , n349394 , n29362 );
buf ( n349397 , n29363 );
not ( n349398 , n349397 );
not ( n349399 , n349398 );
buf ( n349400 , n607 );
not ( n29368 , n349400 );
buf ( n349402 , n606 );
buf ( n349403 , n346493 );
and ( n29371 , n349402 , n349403 );
not ( n349405 , n349402 );
buf ( n349406 , n344484 );
and ( n349407 , n349405 , n349406 );
nor ( n29375 , n29371 , n349407 );
buf ( n349409 , n29375 );
buf ( n349410 , n349409 );
not ( n29378 , n349410 );
or ( n29379 , n29368 , n29378 );
buf ( n349413 , n348590 );
buf ( n349414 , n344454 );
nand ( n29382 , n349413 , n349414 );
buf ( n349416 , n29382 );
buf ( n349417 , n349416 );
nand ( n29385 , n29379 , n349417 );
buf ( n349419 , n29385 );
not ( n349420 , n349419 );
not ( n349421 , n349420 );
or ( n29389 , n349399 , n349421 );
nand ( n349423 , n349419 , n349397 );
nand ( n29391 , n29389 , n349423 );
buf ( n349425 , n343531 );
not ( n29393 , n349425 );
buf ( n349427 , n24108 );
not ( n29395 , n349427 );
buf ( n349429 , n343553 );
not ( n29397 , n349429 );
and ( n29398 , n29395 , n29397 );
buf ( n349432 , n24108 );
buf ( n349433 , n343553 );
and ( n29401 , n349432 , n349433 );
nor ( n29402 , n29398 , n29401 );
buf ( n349436 , n29402 );
buf ( n349437 , n349436 );
not ( n29405 , n349437 );
buf ( n349439 , n29405 );
buf ( n349440 , n349439 );
not ( n29408 , n349440 );
or ( n29409 , n29393 , n29408 );
buf ( n349443 , n348623 );
buf ( n349444 , n343592 );
nand ( n29412 , n349443 , n349444 );
buf ( n29413 , n29412 );
buf ( n349447 , n29413 );
nand ( n29415 , n29409 , n349447 );
buf ( n29416 , n29415 );
buf ( n349450 , n29416 );
not ( n29418 , n28640 );
not ( n29419 , n348692 );
and ( n29420 , n29418 , n29419 );
buf ( n349454 , n348692 );
buf ( n349455 , n28640 );
nand ( n349456 , n349454 , n349455 );
buf ( n349457 , n349456 );
and ( n349458 , n349457 , n348699 );
nor ( n349459 , n29420 , n349458 );
buf ( n349460 , n347812 );
not ( n349461 , n349460 );
buf ( n349462 , n347834 );
not ( n29430 , n349462 );
or ( n349464 , n349461 , n29430 );
buf ( n349465 , n347834 );
buf ( n349466 , n347812 );
or ( n29434 , n349465 , n349466 );
nand ( n349468 , n349464 , n29434 );
buf ( n349469 , n349468 );
buf ( n349470 , n349469 );
buf ( n349471 , n348662 );
not ( n29439 , n349471 );
buf ( n349473 , n29439 );
buf ( n349474 , n349473 );
not ( n29442 , n349474 );
buf ( n349476 , n348658 );
not ( n29444 , n349476 );
or ( n29445 , n29442 , n29444 );
buf ( n29446 , n348658 );
buf ( n349480 , n348669 );
nand ( n29448 , n29446 , n349480 );
buf ( n349482 , n29448 );
buf ( n349483 , n349482 );
nand ( n29451 , n29445 , n349483 );
buf ( n349485 , n29451 );
buf ( n349486 , n349485 );
xor ( n29454 , n349470 , n349486 );
buf ( n349488 , n23911 );
not ( n29456 , n349488 );
buf ( n349490 , n598 );
not ( n29458 , n349490 );
buf ( n349492 , n346202 );
not ( n29460 , n349492 );
or ( n29461 , n29458 , n29460 );
buf ( n349495 , n343953 );
buf ( n349496 , n346199 );
nand ( n349497 , n349495 , n349496 );
buf ( n349498 , n349497 );
buf ( n349499 , n349498 );
nand ( n349500 , n29461 , n349499 );
buf ( n349501 , n349500 );
buf ( n349502 , n349501 );
not ( n29470 , n349502 );
or ( n349504 , n29456 , n29470 );
buf ( n349505 , n348648 );
buf ( n349506 , n343945 );
nand ( n349507 , n349505 , n349506 );
buf ( n349508 , n349507 );
buf ( n349509 , n349508 );
nand ( n349510 , n349504 , n349509 );
buf ( n349511 , n349510 );
buf ( n349512 , n349511 );
xor ( n29480 , n29454 , n349512 );
buf ( n349514 , n29480 );
buf ( n349515 , n344015 );
not ( n349516 , n349515 );
buf ( n349517 , n600 );
not ( n349518 , n349517 );
buf ( n349519 , n345454 );
not ( n349520 , n349519 );
or ( n29488 , n349518 , n349520 );
buf ( n349522 , n23906 );
buf ( n349523 , n345451 );
nand ( n29491 , n349522 , n349523 );
buf ( n29492 , n29491 );
buf ( n349526 , n29492 );
nand ( n29494 , n29488 , n349526 );
buf ( n349528 , n29494 );
buf ( n349529 , n349528 );
not ( n29497 , n349529 );
or ( n29498 , n349516 , n29497 );
buf ( n349532 , n348690 );
buf ( n349533 , n344018 );
nand ( n349534 , n349532 , n349533 );
buf ( n349535 , n349534 );
buf ( n349536 , n349535 );
nand ( n29504 , n29498 , n349536 );
buf ( n349538 , n29504 );
xor ( n349539 , n349514 , n349538 );
not ( n29507 , n349539 );
xor ( n29508 , n349459 , n29507 );
buf ( n349542 , n29508 );
xor ( n349543 , n349450 , n349542 );
buf ( n349544 , n344338 );
not ( n349545 , n349544 );
buf ( n349546 , n348597 );
not ( n29514 , n349546 );
buf ( n349548 , n23530 );
not ( n29516 , n349548 );
and ( n349550 , n29514 , n29516 );
buf ( n349551 , n348597 );
buf ( n349552 , n23530 );
and ( n349553 , n349551 , n349552 );
nor ( n29521 , n349550 , n349553 );
buf ( n349555 , n29521 );
buf ( n349556 , n349555 );
not ( n29524 , n349556 );
buf ( n29525 , n29524 );
buf ( n349559 , n29525 );
not ( n29527 , n349559 );
or ( n29528 , n349545 , n29527 );
buf ( n349562 , n348718 );
buf ( n349563 , n344397 );
nand ( n29531 , n349562 , n349563 );
buf ( n349565 , n29531 );
buf ( n349566 , n349565 );
nand ( n29534 , n29528 , n349566 );
buf ( n29535 , n29534 );
buf ( n29536 , n29535 );
xor ( n29537 , n349543 , n29536 );
buf ( n29538 , n29537 );
and ( n349572 , n29391 , n29538 );
not ( n349573 , n29391 );
not ( n29541 , n29538 );
and ( n349575 , n349573 , n29541 );
nor ( n349576 , n349572 , n349575 );
buf ( n349577 , n349576 );
buf ( n349578 , n348576 );
not ( n349579 , n349578 );
buf ( n349580 , n348611 );
not ( n349581 , n349580 );
buf ( n349582 , n349581 );
buf ( n349583 , n349582 );
nand ( n29551 , n349579 , n349583 );
buf ( n349585 , n29551 );
buf ( n29553 , n349585 );
buf ( n29554 , n348743 );
and ( n29555 , n29553 , n29554 );
buf ( n349589 , n348576 );
not ( n349590 , n349589 );
buf ( n349591 , n349582 );
nor ( n349592 , n349590 , n349591 );
buf ( n349593 , n349592 );
buf ( n349594 , n349593 );
nor ( n349595 , n29555 , n349594 );
buf ( n349596 , n349595 );
buf ( n349597 , n349596 );
nand ( n349598 , n349577 , n349597 );
buf ( n349599 , n349598 );
not ( n349600 , n349599 );
or ( n349601 , n29359 , n349600 );
not ( n29569 , n349576 );
buf ( n29570 , n349596 );
not ( n349604 , n29570 );
buf ( n349605 , n349604 );
nand ( n349606 , n29569 , n349605 );
nand ( n29574 , n349601 , n349606 );
not ( n29575 , n29574 );
buf ( n349609 , n349409 );
not ( n349610 , n349609 );
buf ( n349611 , n349610 );
buf ( n349612 , n349611 );
not ( n29580 , n349612 );
buf ( n349614 , n344631 );
not ( n349615 , n349614 );
and ( n349616 , n29580 , n349615 );
buf ( n349617 , n606 );
not ( n349618 , n349617 );
buf ( n349619 , n346918 );
not ( n29587 , n349619 );
or ( n29588 , n349618 , n29587 );
buf ( n349622 , n23758 );
buf ( n29590 , n344445 );
nand ( n29591 , n349622 , n29590 );
buf ( n349625 , n29591 );
buf ( n349626 , n349625 );
nand ( n29594 , n29588 , n349626 );
buf ( n349628 , n29594 );
buf ( n349629 , n349628 );
buf ( n349630 , n607 );
and ( n29598 , n349629 , n349630 );
nor ( n349632 , n349616 , n29598 );
buf ( n349633 , n349632 );
buf ( n349634 , n349633 );
not ( n29602 , n349634 );
xor ( n349636 , n349450 , n349542 );
and ( n349637 , n349636 , n29536 );
and ( n29605 , n349450 , n349542 );
or ( n349639 , n349637 , n29605 );
buf ( n349640 , n349639 );
buf ( n349641 , n349640 );
not ( n349642 , n349641 );
buf ( n349643 , n349436 );
not ( n349644 , n349643 );
buf ( n349645 , n348498 );
not ( n29613 , n349645 );
and ( n349647 , n349644 , n29613 );
buf ( n349648 , n602 );
not ( n29616 , n349648 );
buf ( n349650 , n24091 );
not ( n349651 , n349650 );
or ( n29619 , n29616 , n349651 );
buf ( n349653 , n344155 );
buf ( n349654 , n343553 );
nand ( n29622 , n349653 , n349654 );
buf ( n29623 , n29622 );
buf ( n349657 , n29623 );
nand ( n349658 , n29619 , n349657 );
buf ( n349659 , n349658 );
buf ( n349660 , n349659 );
buf ( n349661 , n343530 );
and ( n349662 , n349660 , n349661 );
nor ( n29630 , n349647 , n349662 );
buf ( n29631 , n29630 );
buf ( n349665 , n344015 );
not ( n29633 , n349665 );
buf ( n349667 , n600 );
not ( n349668 , n349667 );
buf ( n349669 , n25141 );
not ( n349670 , n349669 );
or ( n29638 , n349668 , n349670 );
not ( n349672 , n600 );
nand ( n349673 , n349672 , n25140 );
buf ( n349674 , n349673 );
nand ( n349675 , n29638 , n349674 );
buf ( n349676 , n349675 );
buf ( n349677 , n349676 );
not ( n349678 , n349677 );
or ( n349679 , n29633 , n349678 );
buf ( n349680 , n349528 );
buf ( n349681 , n344018 );
nand ( n349682 , n349680 , n349681 );
buf ( n349683 , n349682 );
buf ( n349684 , n349683 );
nand ( n29652 , n349679 , n349684 );
buf ( n349686 , n29652 );
buf ( n29654 , n349686 );
buf ( n349688 , n347837 );
buf ( n349689 , n27763 );
nand ( n349690 , n349688 , n349689 );
buf ( n349691 , n349690 );
xor ( n29659 , n349691 , n347791 );
buf ( n349693 , n29659 );
buf ( n349694 , n23911 );
not ( n349695 , n349694 );
buf ( n349696 , n598 );
not ( n29664 , n349696 );
buf ( n349698 , n25665 );
not ( n29666 , n349698 );
or ( n349700 , n29664 , n29666 );
buf ( n349701 , n598 );
not ( n29669 , n349701 );
buf ( n349703 , n348276 );
nand ( n349704 , n29669 , n349703 );
buf ( n349705 , n349704 );
buf ( n349706 , n349705 );
nand ( n349707 , n349700 , n349706 );
buf ( n349708 , n349707 );
buf ( n349709 , n349708 );
not ( n29677 , n349709 );
or ( n29678 , n349695 , n29677 );
buf ( n349712 , n349501 );
buf ( n349713 , n343945 );
nand ( n349714 , n349712 , n349713 );
buf ( n349715 , n349714 );
buf ( n349716 , n349715 );
nand ( n29684 , n29678 , n349716 );
buf ( n349718 , n29684 );
buf ( n349719 , n349718 );
xor ( n349720 , n349693 , n349719 );
xor ( n29688 , n349470 , n349486 );
and ( n349722 , n29688 , n349512 );
and ( n349723 , n349470 , n349486 );
or ( n349724 , n349722 , n349723 );
buf ( n349725 , n349724 );
buf ( n349726 , n349725 );
xor ( n349727 , n349720 , n349726 );
buf ( n349728 , n349727 );
buf ( n349729 , n349728 );
xor ( n349730 , n29654 , n349729 );
not ( n349731 , n349538 );
not ( n29699 , n349514 );
or ( n29700 , n349731 , n29699 );
buf ( n29701 , n349538 );
buf ( n29702 , n349514 );
nor ( n29703 , n29701 , n29702 );
buf ( n29704 , n29703 );
or ( n349738 , n349459 , n29704 );
nand ( n29706 , n29700 , n349738 );
buf ( n349740 , n29706 );
xor ( n349741 , n349730 , n349740 );
buf ( n349742 , n349741 );
xor ( n349743 , n29631 , n349742 );
buf ( n349744 , n349555 );
not ( n349745 , n349744 );
buf ( n349746 , n348782 );
not ( n29714 , n349746 );
and ( n29715 , n349745 , n29714 );
buf ( n349749 , n604 );
not ( n349750 , n349749 );
buf ( n349751 , n343672 );
not ( n29719 , n349751 );
or ( n349753 , n349750 , n29719 );
buf ( n349754 , n344185 );
buf ( n349755 , n23530 );
nand ( n349756 , n349754 , n349755 );
buf ( n349757 , n349756 );
buf ( n349758 , n349757 );
nand ( n349759 , n349753 , n349758 );
buf ( n349760 , n349759 );
buf ( n349761 , n349760 );
buf ( n349762 , n344338 );
and ( n29730 , n349761 , n349762 );
nor ( n29731 , n29715 , n29730 );
buf ( n349765 , n29731 );
xnor ( n349766 , n349743 , n349765 );
buf ( n349767 , n349766 );
not ( n349768 , n349767 );
or ( n29736 , n349642 , n349768 );
buf ( n349770 , n349640 );
buf ( n349771 , n349766 );
or ( n29739 , n349770 , n349771 );
nand ( n29740 , n29736 , n29739 );
buf ( n349774 , n29740 );
buf ( n349775 , n349774 );
not ( n29743 , n349775 );
or ( n29744 , n29602 , n29743 );
buf ( n349778 , n349633 );
buf ( n349779 , n349774 );
or ( n29747 , n349778 , n349779 );
nand ( n29748 , n29744 , n29747 );
buf ( n349782 , n29748 );
not ( n29750 , n349782 );
buf ( n349784 , n349397 );
buf ( n349785 , n349419 );
or ( n29753 , n349784 , n349785 );
buf ( n349787 , n29538 );
nand ( n29755 , n29753 , n349787 );
buf ( n349789 , n29755 );
buf ( n349790 , n349789 );
buf ( n29758 , n349419 );
buf ( n349792 , n349397 );
nand ( n349793 , n29758 , n349792 );
buf ( n349794 , n349793 );
buf ( n349795 , n349794 );
nand ( n349796 , n349790 , n349795 );
buf ( n349797 , n349796 );
not ( n29765 , n349797 );
nand ( n29766 , n29750 , n29765 );
not ( n29767 , n29766 );
or ( n29768 , n29575 , n29767 );
nand ( n29769 , n349797 , n349782 );
nand ( n29770 , n29768 , n29769 );
not ( n29771 , n29770 );
buf ( n349805 , n29631 );
not ( n29773 , n349805 );
buf ( n349807 , n349765 );
not ( n29775 , n349807 );
or ( n29776 , n29773 , n29775 );
buf ( n349810 , n349742 );
nand ( n29778 , n29776 , n349810 );
buf ( n349812 , n29778 );
buf ( n349813 , n349812 );
buf ( n349814 , n349765 );
buf ( n349815 , n29631 );
or ( n29783 , n349814 , n349815 );
buf ( n29784 , n29783 );
buf ( n349818 , n29784 );
nand ( n29786 , n349813 , n349818 );
buf ( n349820 , n29786 );
buf ( n349821 , n349820 );
buf ( n349822 , n607 );
not ( n29790 , n349822 );
not ( n349824 , n347904 );
xor ( n349825 , n606 , n349824 );
buf ( n349826 , n349825 );
not ( n349827 , n349826 );
or ( n349828 , n29790 , n349827 );
buf ( n349829 , n349628 );
buf ( n349830 , n344454 );
nand ( n349831 , n349829 , n349830 );
buf ( n349832 , n349831 );
buf ( n349833 , n349832 );
nand ( n349834 , n349828 , n349833 );
buf ( n349835 , n349834 );
buf ( n349836 , n349835 );
xor ( n349837 , n349821 , n349836 );
xor ( n349838 , n29654 , n349729 );
and ( n29806 , n349838 , n349740 );
and ( n349840 , n29654 , n349729 );
or ( n349841 , n29806 , n349840 );
buf ( n349842 , n349841 );
buf ( n349843 , n349842 );
buf ( n29811 , n344338 );
not ( n29812 , n29811 );
buf ( n349846 , n604 );
not ( n29814 , n349846 );
buf ( n349848 , n344484 );
not ( n29816 , n349848 );
or ( n349850 , n29814 , n29816 );
buf ( n349851 , n24452 );
buf ( n349852 , n23530 );
nand ( n349853 , n349851 , n349852 );
buf ( n349854 , n349853 );
buf ( n349855 , n349854 );
nand ( n349856 , n349850 , n349855 );
buf ( n349857 , n349856 );
buf ( n349858 , n349857 );
not ( n349859 , n349858 );
or ( n349860 , n29812 , n349859 );
buf ( n349861 , n344397 );
buf ( n349862 , n349760 );
nand ( n349863 , n349861 , n349862 );
buf ( n349864 , n349863 );
buf ( n349865 , n349864 );
nand ( n349866 , n349860 , n349865 );
buf ( n349867 , n349866 );
buf ( n349868 , n349867 );
xor ( n29836 , n349843 , n349868 );
buf ( n349870 , n344015 );
not ( n349871 , n349870 );
buf ( n349872 , n600 );
not ( n29840 , n349872 );
buf ( n349874 , n24109 );
not ( n349875 , n349874 );
or ( n29843 , n29840 , n349875 );
buf ( n349877 , n347595 );
buf ( n349878 , n23906 );
nand ( n349879 , n349877 , n349878 );
buf ( n349880 , n349879 );
buf ( n349881 , n349880 );
nand ( n29849 , n29843 , n349881 );
buf ( n349883 , n29849 );
buf ( n349884 , n349883 );
not ( n349885 , n349884 );
or ( n29853 , n349871 , n349885 );
buf ( n349887 , n349676 );
buf ( n349888 , n344018 );
nand ( n349889 , n349887 , n349888 );
buf ( n349890 , n349889 );
buf ( n349891 , n349890 );
nand ( n29859 , n29853 , n349891 );
buf ( n349893 , n29859 );
buf ( n349894 , n349893 );
xor ( n349895 , n347752 , n347840 );
xor ( n29863 , n349895 , n347854 );
buf ( n349897 , n29863 );
buf ( n349898 , n349897 );
buf ( n349899 , n23911 );
not ( n349900 , n349899 );
and ( n349901 , n346695 , n598 );
not ( n349902 , n346695 );
and ( n29870 , n349902 , n343953 );
or ( n349904 , n349901 , n29870 );
buf ( n349905 , n349904 );
not ( n349906 , n349905 );
or ( n29874 , n349900 , n349906 );
buf ( n349908 , n349708 );
buf ( n29876 , n343945 );
nand ( n29877 , n349908 , n29876 );
buf ( n29878 , n29877 );
buf ( n349912 , n29878 );
nand ( n29880 , n29874 , n349912 );
buf ( n29881 , n29880 );
buf ( n349915 , n29881 );
xor ( n29883 , n349898 , n349915 );
xor ( n29884 , n349693 , n349719 );
and ( n349918 , n29884 , n349726 );
and ( n29886 , n349693 , n349719 );
or ( n349920 , n349918 , n29886 );
buf ( n349921 , n349920 );
buf ( n349922 , n349921 );
xor ( n349923 , n29883 , n349922 );
buf ( n349924 , n349923 );
buf ( n349925 , n349924 );
xor ( n349926 , n349894 , n349925 );
buf ( n349927 , n343531 );
not ( n349928 , n349927 );
buf ( n349929 , n602 );
not ( n29897 , n349929 );
buf ( n349931 , n26331 );
not ( n29899 , n349931 );
or ( n29900 , n29897 , n29899 );
buf ( n349934 , n23606 );
buf ( n349935 , n343553 );
nand ( n29903 , n349934 , n349935 );
buf ( n349937 , n29903 );
buf ( n349938 , n349937 );
nand ( n29906 , n29900 , n349938 );
buf ( n349940 , n29906 );
buf ( n349941 , n349940 );
not ( n29909 , n349941 );
or ( n349943 , n349928 , n29909 );
buf ( n349944 , n349659 );
buf ( n349945 , n343592 );
nand ( n29913 , n349944 , n349945 );
buf ( n349947 , n29913 );
buf ( n349948 , n349947 );
nand ( n349949 , n349943 , n349948 );
buf ( n349950 , n349949 );
buf ( n349951 , n349950 );
xor ( n349952 , n349926 , n349951 );
buf ( n349953 , n349952 );
buf ( n349954 , n349953 );
xor ( n349955 , n29836 , n349954 );
buf ( n349956 , n349955 );
buf ( n349957 , n349956 );
xnor ( n29925 , n349837 , n349957 );
buf ( n349959 , n29925 );
buf ( n349960 , n349959 );
buf ( n349961 , n349640 );
not ( n349962 , n349961 );
buf ( n349963 , n349633 );
nand ( n349964 , n349962 , n349963 );
buf ( n349965 , n349964 );
buf ( n349966 , n349965 );
buf ( n349967 , n349766 );
not ( n29935 , n349967 );
buf ( n349969 , n29935 );
buf ( n349970 , n349969 );
and ( n349971 , n349966 , n349970 );
buf ( n349972 , n349640 );
not ( n29940 , n349972 );
buf ( n349974 , n349633 );
nor ( n29942 , n29940 , n349974 );
buf ( n349976 , n29942 );
buf ( n349977 , n349976 );
nor ( n29945 , n349971 , n349977 );
buf ( n349979 , n29945 );
buf ( n29947 , n349979 );
nand ( n29948 , n349960 , n29947 );
buf ( n29949 , n29948 );
not ( n349983 , n29949 );
or ( n29951 , n29771 , n349983 );
buf ( n349985 , n349959 );
not ( n349986 , n349985 );
buf ( n349987 , n349986 );
buf ( n349988 , n349987 );
buf ( n349989 , n349979 );
not ( n349990 , n349989 );
buf ( n349991 , n349990 );
buf ( n349992 , n349991 );
nand ( n349993 , n349988 , n349992 );
buf ( n349994 , n349993 );
nand ( n349995 , n29951 , n349994 );
buf ( n29963 , n349995 );
buf ( n349997 , n349820 );
not ( n29965 , n349997 );
buf ( n349999 , n349835 );
not ( n29967 , n349999 );
buf ( n350001 , n29967 );
buf ( n350002 , n350001 );
not ( n29970 , n350002 );
buf ( n350004 , n29970 );
buf ( n350005 , n350004 );
not ( n350006 , n350005 );
or ( n350007 , n29965 , n350006 );
buf ( n350008 , n349820 );
not ( n29976 , n350008 );
buf ( n350010 , n29976 );
buf ( n350011 , n350010 );
not ( n29979 , n350011 );
buf ( n350013 , n350001 );
not ( n350014 , n350013 );
or ( n29982 , n29979 , n350014 );
buf ( n350016 , n349956 );
nand ( n350017 , n29982 , n350016 );
buf ( n350018 , n350017 );
buf ( n350019 , n350018 );
nand ( n350020 , n350007 , n350019 );
buf ( n350021 , n350020 );
buf ( n350022 , n350021 );
not ( n29990 , n350022 );
buf ( n350024 , n606 );
not ( n350025 , n350024 );
buf ( n350026 , n347358 );
not ( n350027 , n350026 );
or ( n350028 , n350025 , n350027 );
buf ( n350029 , n344230 );
not ( n29997 , n350029 );
buf ( n350031 , n344445 );
nand ( n29999 , n29997 , n350031 );
buf ( n350033 , n29999 );
buf ( n350034 , n350033 );
nand ( n30002 , n350028 , n350034 );
buf ( n350036 , n30002 );
buf ( n350037 , n350036 );
buf ( n350038 , n607 );
and ( n30006 , n350037 , n350038 );
buf ( n350040 , n349825 );
not ( n30008 , n350040 );
buf ( n350042 , n344631 );
nor ( n30010 , n30008 , n350042 );
buf ( n350044 , n30010 );
buf ( n350045 , n350044 );
nor ( n30013 , n30006 , n350045 );
buf ( n350047 , n30013 );
buf ( n350048 , n350047 );
not ( n30016 , n350048 );
xor ( n30017 , n349843 , n349868 );
and ( n30018 , n30017 , n349954 );
and ( n30019 , n349843 , n349868 );
or ( n30020 , n30018 , n30019 );
buf ( n350054 , n30020 );
buf ( n350055 , n350054 );
not ( n30023 , n350055 );
and ( n350057 , n30016 , n30023 );
buf ( n350058 , n350047 );
buf ( n350059 , n350054 );
and ( n350060 , n350058 , n350059 );
nor ( n30028 , n350057 , n350060 );
buf ( n350062 , n30028 );
buf ( n350063 , n350062 );
not ( n30031 , n350063 );
xor ( n350065 , n349894 , n349925 );
and ( n350066 , n350065 , n349951 );
and ( n30034 , n349894 , n349925 );
or ( n30035 , n350066 , n30034 );
buf ( n350069 , n30035 );
buf ( n350070 , n350069 );
buf ( n350071 , n344338 );
not ( n30039 , n350071 );
buf ( n350073 , n604 );
not ( n350074 , n350073 );
buf ( n350075 , n346918 );
not ( n350076 , n350075 );
or ( n350077 , n350074 , n350076 );
buf ( n350078 , n23758 );
buf ( n350079 , n23530 );
nand ( n350080 , n350078 , n350079 );
buf ( n350081 , n350080 );
buf ( n350082 , n350081 );
nand ( n350083 , n350077 , n350082 );
buf ( n350084 , n350083 );
buf ( n350085 , n350084 );
not ( n350086 , n350085 );
or ( n30054 , n30039 , n350086 );
buf ( n350088 , n349857 );
buf ( n350089 , n344397 );
nand ( n30057 , n350088 , n350089 );
buf ( n350091 , n30057 );
buf ( n350092 , n350091 );
nand ( n30060 , n30054 , n350092 );
buf ( n350094 , n30060 );
buf ( n350095 , n350094 );
xor ( n30063 , n350070 , n350095 );
xor ( n30064 , n349898 , n349915 );
and ( n350098 , n30064 , n349922 );
and ( n350099 , n349898 , n349915 );
or ( n350100 , n350098 , n350099 );
buf ( n350101 , n350100 );
buf ( n350102 , n350101 );
buf ( n350103 , n343531 );
not ( n350104 , n350103 );
buf ( n350105 , n602 );
not ( n350106 , n350105 );
buf ( n350107 , n343678 );
not ( n30075 , n350107 );
or ( n350109 , n350106 , n30075 );
buf ( n350110 , n343675 );
buf ( n350111 , n343553 );
nand ( n350112 , n350110 , n350111 );
buf ( n350113 , n350112 );
buf ( n350114 , n350113 );
nand ( n350115 , n350109 , n350114 );
buf ( n350116 , n350115 );
buf ( n350117 , n350116 );
not ( n350118 , n350117 );
or ( n350119 , n350104 , n350118 );
buf ( n30087 , n349940 );
buf ( n30088 , n343592 );
nand ( n30089 , n30087 , n30088 );
buf ( n30090 , n30089 );
buf ( n350124 , n30090 );
nand ( n350125 , n350119 , n350124 );
buf ( n350126 , n350125 );
buf ( n350127 , n350126 );
xor ( n30095 , n350102 , n350127 );
buf ( n350129 , n23911 );
not ( n30097 , n350129 );
buf ( n350131 , n28134 );
not ( n350132 , n350131 );
or ( n350133 , n30097 , n350132 );
buf ( n350134 , n349904 );
buf ( n350135 , n343945 );
nand ( n350136 , n350134 , n350135 );
buf ( n350137 , n350136 );
buf ( n350138 , n350137 );
nand ( n350139 , n350133 , n350138 );
buf ( n350140 , n350139 );
buf ( n350141 , n350140 );
buf ( n30109 , n347743 );
buf ( n30110 , n347728 );
xor ( n30111 , n30109 , n30110 );
buf ( n350145 , n347861 );
xnor ( n350146 , n30111 , n350145 );
buf ( n350147 , n350146 );
buf ( n350148 , n350147 );
xor ( n350149 , n350141 , n350148 );
buf ( n350150 , n344015 );
not ( n350151 , n350150 );
buf ( n350152 , n348191 );
not ( n30120 , n350152 );
or ( n30121 , n350151 , n30120 );
buf ( n350155 , n349883 );
buf ( n350156 , n344018 );
nand ( n350157 , n350155 , n350156 );
buf ( n350158 , n350157 );
buf ( n350159 , n350158 );
nand ( n30127 , n30121 , n350159 );
buf ( n350161 , n30127 );
buf ( n350162 , n350161 );
xor ( n30130 , n350149 , n350162 );
buf ( n350164 , n30130 );
buf ( n350165 , n350164 );
xor ( n30133 , n30095 , n350165 );
buf ( n350167 , n30133 );
buf ( n30135 , n350167 );
xor ( n30136 , n30063 , n30135 );
buf ( n30137 , n30136 );
buf ( n350171 , n30137 );
not ( n30139 , n350171 );
and ( n30140 , n30031 , n30139 );
buf ( n350174 , n30137 );
buf ( n350175 , n350062 );
and ( n30143 , n350174 , n350175 );
nor ( n350177 , n30140 , n30143 );
buf ( n350178 , n350177 );
buf ( n350179 , n350178 );
nand ( n350180 , n29990 , n350179 );
buf ( n350181 , n350180 );
buf ( n350182 , n350181 );
and ( n30150 , n29963 , n350182 );
buf ( n350184 , n30150 );
buf ( n350185 , n350184 );
not ( n30153 , n30137 );
buf ( n350187 , n350054 );
not ( n350188 , n350187 );
buf ( n350189 , n350047 );
nand ( n350190 , n350188 , n350189 );
buf ( n350191 , n350190 );
not ( n30159 , n350191 );
or ( n350193 , n30153 , n30159 );
buf ( n30161 , n350047 );
not ( n30162 , n30161 );
buf ( n350196 , n350054 );
nand ( n30164 , n30162 , n350196 );
buf ( n350198 , n30164 );
nand ( n30166 , n350193 , n350198 );
not ( n350200 , n30166 );
buf ( n350201 , n607 );
not ( n30169 , n350201 );
buf ( n350203 , n606 );
not ( n350204 , n350203 );
buf ( n350205 , n343911 );
not ( n350206 , n350205 );
or ( n350207 , n350204 , n350206 );
buf ( n350208 , n347209 );
buf ( n350209 , n344445 );
nand ( n350210 , n350208 , n350209 );
buf ( n350211 , n350210 );
buf ( n350212 , n350211 );
nand ( n350213 , n350207 , n350212 );
buf ( n350214 , n350213 );
buf ( n350215 , n350214 );
not ( n30183 , n350215 );
or ( n30184 , n30169 , n30183 );
buf ( n350218 , n350036 );
buf ( n350219 , n344454 );
nand ( n30187 , n350218 , n350219 );
buf ( n350221 , n30187 );
buf ( n350222 , n350221 );
nand ( n30190 , n30184 , n350222 );
buf ( n350224 , n30190 );
xor ( n350225 , n350070 , n350095 );
and ( n30193 , n350225 , n30135 );
and ( n350227 , n350070 , n350095 );
or ( n350228 , n30193 , n350227 );
buf ( n350229 , n350228 );
xnor ( n30197 , n350224 , n350229 );
xor ( n30198 , n350102 , n350127 );
and ( n30199 , n30198 , n350165 );
and ( n350233 , n350102 , n350127 );
or ( n350234 , n30199 , n350233 );
buf ( n350235 , n350234 );
buf ( n350236 , n350235 );
buf ( n350237 , n344338 );
not ( n30205 , n350237 );
and ( n350239 , n604 , n347904 );
not ( n350240 , n604 );
and ( n30208 , n350240 , n343723 );
or ( n350242 , n350239 , n30208 );
buf ( n350243 , n350242 );
not ( n30211 , n350243 );
or ( n350245 , n30205 , n30211 );
buf ( n350246 , n350084 );
buf ( n350247 , n344400 );
nand ( n350248 , n350246 , n350247 );
buf ( n350249 , n350248 );
buf ( n350250 , n350249 );
nand ( n350251 , n350245 , n350250 );
buf ( n350252 , n350251 );
buf ( n350253 , n350252 );
xor ( n30221 , n350236 , n350253 );
xor ( n350255 , n350141 , n350148 );
and ( n350256 , n350255 , n350162 );
and ( n30224 , n350141 , n350148 );
or ( n350258 , n350256 , n30224 );
buf ( n350259 , n350258 );
buf ( n350260 , n350259 );
buf ( n350261 , n343531 );
not ( n30229 , n350261 );
buf ( n350263 , n28193 );
not ( n350264 , n350263 );
or ( n350265 , n30229 , n350264 );
buf ( n350266 , n350116 );
buf ( n350267 , n343592 );
nand ( n350268 , n350266 , n350267 );
buf ( n350269 , n350268 );
buf ( n350270 , n350269 );
nand ( n30238 , n350265 , n350270 );
buf ( n350272 , n30238 );
buf ( n350273 , n350272 );
xor ( n350274 , n350260 , n350273 );
xor ( n350275 , n348160 , n348173 );
xor ( n350276 , n350275 , n348199 );
buf ( n350277 , n350276 );
buf ( n350278 , n350277 );
xor ( n350279 , n350274 , n350278 );
buf ( n350280 , n350279 );
buf ( n350281 , n350280 );
xor ( n350282 , n30221 , n350281 );
buf ( n350283 , n350282 );
and ( n350284 , n30197 , n350283 );
not ( n350285 , n30197 );
buf ( n350286 , n350283 );
not ( n30254 , n350286 );
buf ( n350288 , n30254 );
and ( n30256 , n350285 , n350288 );
nor ( n30257 , n350284 , n30256 );
nand ( n30258 , n350200 , n30257 );
buf ( n350292 , n30258 );
nand ( n30260 , n350185 , n350292 );
buf ( n350294 , n30260 );
buf ( n350295 , n350294 );
buf ( n350296 , n30258 );
not ( n30264 , n350178 );
nand ( n350298 , n30264 , n350021 );
buf ( n350299 , n350298 );
not ( n30267 , n350299 );
buf ( n350301 , n30267 );
buf ( n350302 , n350301 );
nand ( n30270 , n350296 , n350302 );
buf ( n350304 , n30270 );
buf ( n350305 , n350304 );
buf ( n350306 , n30257 );
not ( n350307 , n350306 );
buf ( n350308 , n30166 );
nand ( n30276 , n350307 , n350308 );
buf ( n350310 , n30276 );
buf ( n350311 , n350310 );
nand ( n30279 , n350295 , n350305 , n350311 );
buf ( n30280 , n30279 );
not ( n350314 , n30280 );
xor ( n350315 , n350236 , n350253 );
and ( n350316 , n350315 , n350281 );
and ( n30284 , n350236 , n350253 );
or ( n30285 , n350316 , n30284 );
buf ( n350319 , n30285 );
buf ( n350320 , n350319 );
buf ( n350321 , n607 );
not ( n350322 , n350321 );
buf ( n350323 , n606 );
not ( n350324 , n350323 );
buf ( n350325 , n347525 );
not ( n350326 , n350325 );
or ( n30294 , n350324 , n350326 );
buf ( n350328 , n343872 );
not ( n350329 , n350328 );
buf ( n350330 , n344445 );
nand ( n30298 , n350329 , n350330 );
buf ( n350332 , n30298 );
buf ( n350333 , n350332 );
nand ( n350334 , n30294 , n350333 );
buf ( n350335 , n350334 );
buf ( n350336 , n350335 );
not ( n30304 , n350336 );
or ( n30305 , n350322 , n30304 );
buf ( n30306 , n350214 );
buf ( n350340 , n344454 );
nand ( n30308 , n30306 , n350340 );
buf ( n30309 , n30308 );
buf ( n350343 , n30309 );
nand ( n350344 , n30305 , n350343 );
buf ( n350345 , n350344 );
buf ( n350346 , n350345 );
xor ( n30314 , n350320 , n350346 );
xor ( n30315 , n350260 , n350273 );
and ( n30316 , n30315 , n350278 );
and ( n30317 , n350260 , n350273 );
or ( n30318 , n30316 , n30317 );
buf ( n350352 , n30318 );
buf ( n350353 , n350352 );
buf ( n350354 , n344338 );
not ( n350355 , n350354 );
buf ( n350356 , n28116 );
not ( n350357 , n350356 );
or ( n350358 , n350355 , n350357 );
buf ( n350359 , n350242 );
buf ( n350360 , n344400 );
nand ( n30328 , n350359 , n350360 );
buf ( n350362 , n30328 );
buf ( n350363 , n350362 );
nand ( n30331 , n350358 , n350363 );
buf ( n350365 , n30331 );
buf ( n350366 , n350365 );
xor ( n350367 , n350353 , n350366 );
xor ( n350368 , n348204 , n348216 );
xor ( n30336 , n350368 , n348234 );
buf ( n350370 , n30336 );
buf ( n350371 , n350370 );
xnor ( n350372 , n350367 , n350371 );
buf ( n350373 , n350372 );
buf ( n350374 , n350373 );
xor ( n30342 , n30314 , n350374 );
buf ( n350376 , n30342 );
buf ( n350377 , n350224 );
not ( n30345 , n350377 );
buf ( n350379 , n350288 );
nand ( n350380 , n30345 , n350379 );
buf ( n350381 , n350380 );
and ( n350382 , n350381 , n350229 );
buf ( n350383 , n350224 );
not ( n350384 , n350383 );
buf ( n350385 , n350288 );
nor ( n350386 , n350384 , n350385 );
buf ( n350387 , n350386 );
nor ( n30355 , n350382 , n350387 );
nand ( n30356 , n350376 , n30355 );
not ( n30357 , n30356 );
or ( n30358 , n350314 , n30357 );
not ( n350392 , n30355 );
buf ( n350393 , n350376 );
not ( n30361 , n350393 );
buf ( n350395 , n30361 );
nand ( n350396 , n350392 , n350395 );
nand ( n350397 , n30358 , n350396 );
not ( n30365 , n350397 );
not ( n350399 , n348104 );
buf ( n350400 , n350399 );
not ( n350401 , n350400 );
not ( n30369 , n348126 );
not ( n350403 , n28210 );
or ( n350404 , n30369 , n350403 );
or ( n350405 , n28210 , n348126 );
nand ( n30373 , n350404 , n350405 );
not ( n350407 , n30373 );
buf ( n350408 , n350407 );
not ( n350409 , n350408 );
or ( n30377 , n350401 , n350409 );
buf ( n350411 , n30373 );
buf ( n350412 , n348104 );
nand ( n350413 , n350411 , n350412 );
buf ( n350414 , n350413 );
buf ( n350415 , n350414 );
nand ( n350416 , n30377 , n350415 );
buf ( n350417 , n350416 );
buf ( n350418 , n350417 );
buf ( n350419 , n350365 );
not ( n350420 , n350419 );
buf ( n350421 , n350420 );
buf ( n350422 , n350421 );
not ( n350423 , n350422 );
buf ( n350424 , n350352 );
not ( n350425 , n350424 );
buf ( n350426 , n350425 );
buf ( n350427 , n350426 );
not ( n30395 , n350427 );
or ( n30396 , n350423 , n30395 );
buf ( n350430 , n350370 );
nand ( n350431 , n30396 , n350430 );
buf ( n350432 , n350431 );
buf ( n350433 , n350432 );
buf ( n350434 , n350426 );
not ( n30402 , n350434 );
buf ( n350436 , n350365 );
nand ( n350437 , n30402 , n350436 );
buf ( n350438 , n350437 );
buf ( n350439 , n350438 );
nand ( n350440 , n350433 , n350439 );
buf ( n350441 , n350440 );
buf ( n350442 , n350441 );
buf ( n350443 , n607 );
not ( n350444 , n350443 );
buf ( n350445 , n347575 );
not ( n350446 , n350445 );
or ( n30414 , n350444 , n350446 );
buf ( n350448 , n350335 );
buf ( n350449 , n344454 );
nand ( n30417 , n350448 , n350449 );
buf ( n30418 , n30417 );
buf ( n350452 , n30418 );
nand ( n350453 , n30414 , n350452 );
buf ( n350454 , n350453 );
buf ( n350455 , n350454 );
xor ( n30423 , n350442 , n350455 );
buf ( n350457 , n348238 );
buf ( n350458 , n348156 );
xor ( n350459 , n350457 , n350458 );
buf ( n350460 , n348131 );
xor ( n350461 , n350459 , n350460 );
buf ( n350462 , n350461 );
buf ( n350463 , n350462 );
and ( n30431 , n30423 , n350463 );
and ( n30432 , n350442 , n350455 );
or ( n30433 , n30431 , n30432 );
buf ( n350467 , n30433 );
buf ( n350468 , n350467 );
nor ( n350469 , n350418 , n350468 );
buf ( n350470 , n350469 );
buf ( n350471 , n350470 );
xor ( n30439 , n350442 , n350455 );
xor ( n30440 , n30439 , n350463 );
buf ( n350474 , n30440 );
buf ( n350475 , n350474 );
xor ( n350476 , n350319 , n350345 );
not ( n350477 , n350373 );
and ( n350478 , n350476 , n350477 );
and ( n30446 , n350319 , n350345 );
or ( n30447 , n350478 , n30446 );
buf ( n350481 , n30447 );
nor ( n30449 , n350475 , n350481 );
buf ( n30450 , n30449 );
buf ( n350484 , n30450 );
nor ( n350485 , n350471 , n350484 );
buf ( n350486 , n350485 );
not ( n30454 , n350486 );
or ( n30455 , n30365 , n30454 );
buf ( n350489 , n350467 );
not ( n30457 , n350489 );
buf ( n350491 , n350417 );
not ( n30459 , n350491 );
buf ( n350493 , n30459 );
buf ( n350494 , n350493 );
nand ( n30462 , n30457 , n350494 );
buf ( n350496 , n30462 );
buf ( n350497 , n350496 );
buf ( n350498 , n350474 );
buf ( n350499 , n30447 );
and ( n350500 , n350498 , n350499 );
buf ( n350501 , n350500 );
buf ( n350502 , n350501 );
and ( n350503 , n350497 , n350502 );
buf ( n350504 , n350467 );
not ( n30472 , n350504 );
buf ( n350506 , n350493 );
nor ( n30474 , n30472 , n350506 );
buf ( n350508 , n30474 );
buf ( n350509 , n350508 );
nor ( n30477 , n350503 , n350509 );
buf ( n30478 , n30477 );
nand ( n350512 , n30455 , n30478 );
or ( n350513 , n347489 , n347296 );
not ( n30481 , n347342 );
not ( n350515 , n347316 );
or ( n350516 , n30481 , n350515 );
nor ( n350517 , n347316 , n347342 );
buf ( n350518 , n347483 );
not ( n350519 , n350518 );
buf ( n350520 , n350519 );
or ( n350521 , n350517 , n350520 );
nand ( n30489 , n350516 , n350521 );
nand ( n350523 , n347296 , n30489 );
nand ( n350524 , n350513 , n350523 );
buf ( n350525 , n350524 );
buf ( n350526 , n347305 );
and ( n30494 , n350525 , n350526 );
not ( n350528 , n350525 );
buf ( n350529 , n347495 );
and ( n350530 , n350528 , n350529 );
nor ( n350531 , n30494 , n350530 );
buf ( n350532 , n350531 );
xor ( n350533 , n348041 , n348059 );
and ( n350534 , n350533 , n348075 );
and ( n30502 , n348041 , n348059 );
or ( n30503 , n350534 , n30502 );
buf ( n350537 , n30503 );
nand ( n350538 , n350532 , n350537 );
nand ( n30506 , n348262 , n350512 , n350538 );
buf ( n350540 , n30506 );
buf ( n350541 , n348077 );
not ( n30509 , n350541 );
buf ( n30510 , n30509 );
buf ( n350544 , n348036 );
not ( n30512 , n350544 );
buf ( n350546 , n30512 );
nand ( n350547 , n30510 , n350546 );
not ( n30515 , n350547 );
not ( n350549 , n348036 );
not ( n30517 , n348077 );
or ( n30518 , n350549 , n30517 );
buf ( n30519 , n348082 );
buf ( n30520 , n348257 );
nor ( n30521 , n30519 , n30520 );
buf ( n30522 , n30521 );
nand ( n350556 , n30518 , n30522 );
not ( n30524 , n350556 );
or ( n350558 , n30515 , n30524 );
nand ( n350559 , n350558 , n350538 );
buf ( n350560 , n350559 );
not ( n30528 , n350532 );
not ( n350562 , n350537 );
nand ( n350563 , n30528 , n350562 );
buf ( n350564 , n350563 );
nand ( n350565 , n350540 , n350560 , n350564 );
buf ( n350566 , n350565 );
not ( n30534 , n350566 );
or ( n350568 , n347511 , n30534 );
not ( n350569 , n27251 );
nand ( n350570 , n347504 , n347499 );
nand ( n350571 , n346873 , n27250 );
nand ( n30539 , n350570 , n350571 );
nand ( n350573 , n350569 , n30539 );
buf ( n350574 , n350573 );
not ( n350575 , n350574 );
buf ( n350576 , n350575 );
buf ( n350577 , n346861 );
buf ( n30545 , n350577 );
buf ( n350579 , n30545 );
and ( n30547 , n350576 , n350579 );
buf ( n350581 , n345981 );
buf ( n350582 , n346427 );
nand ( n350583 , n350581 , n350582 );
buf ( n350584 , n350583 );
buf ( n350585 , n350584 );
not ( n350586 , n26403 );
buf ( n350587 , n26827 );
not ( n350588 , n350587 );
buf ( n350589 , n350588 );
nand ( n30557 , n350586 , n350589 );
buf ( n350591 , n30557 );
nand ( n30559 , n350585 , n350591 );
buf ( n350593 , n30559 );
nor ( n30561 , n30547 , n350593 );
nand ( n350595 , n350568 , n30561 );
not ( n350596 , n350595 );
or ( n30564 , n26401 , n350596 );
xor ( n350598 , n345081 , n345381 );
xor ( n30566 , n350598 , n345389 );
buf ( n350600 , n30566 );
buf ( n30568 , n350600 );
buf ( n350602 , n345639 );
buf ( n350603 , n25592 );
buf ( n350604 , n350603 );
buf ( n350605 , n350604 );
buf ( n350606 , n350605 );
or ( n30574 , n350602 , n350606 );
buf ( n350608 , n345403 );
nand ( n30576 , n30574 , n350608 );
buf ( n350610 , n30576 );
buf ( n350611 , n350610 );
buf ( n350612 , n350605 );
buf ( n350613 , n345639 );
nand ( n30581 , n350612 , n350613 );
buf ( n30582 , n30581 );
buf ( n350616 , n30582 );
nand ( n30584 , n350611 , n350616 );
buf ( n350618 , n30584 );
buf ( n350619 , n350618 );
nand ( n350620 , n30568 , n350619 );
buf ( n350621 , n350620 );
buf ( n350622 , n350621 );
buf ( n350623 , n345643 );
buf ( n350624 , n345967 );
nand ( n350625 , n350623 , n350624 );
buf ( n350626 , n350625 );
buf ( n350627 , n350626 );
and ( n30595 , n350622 , n350627 );
buf ( n350629 , n30595 );
nand ( n30597 , n30564 , n350629 );
buf ( n350631 , n350600 );
buf ( n350632 , n350631 );
buf ( n350633 , n350632 );
buf ( n350634 , n350633 );
not ( n350635 , n350634 );
buf ( n350636 , n350635 );
buf ( n350637 , n350636 );
buf ( n350638 , n350618 );
not ( n350639 , n350638 );
buf ( n350640 , n350639 );
nand ( n350641 , n350637 , n350640 );
buf ( n350642 , n350641 );
nand ( n30610 , n30597 , n350642 );
not ( n30611 , n30610 );
not ( n350645 , n30611 );
or ( n30613 , n25365 , n350645 );
nor ( n350647 , n25034 , n345396 );
not ( n30615 , n350647 );
buf ( n30616 , n30615 );
nand ( n350650 , n30613 , n30616 );
buf ( n350651 , n23889 );
not ( n30619 , n350651 );
buf ( n350653 , n344577 );
not ( n350654 , n350653 );
or ( n30622 , n30619 , n350654 );
xor ( n350656 , n596 , n23993 );
buf ( n30624 , n350656 );
buf ( n30625 , n343863 );
nand ( n30626 , n30624 , n30625 );
buf ( n30627 , n30626 );
buf ( n30628 , n30627 );
nand ( n30629 , n30622 , n30628 );
buf ( n30630 , n30629 );
buf ( n30631 , n30630 );
not ( n350665 , n23911 );
buf ( n350666 , n598 );
not ( n350667 , n350666 );
buf ( n350668 , n344308 );
not ( n30636 , n350668 );
or ( n30637 , n350667 , n30636 );
buf ( n350671 , n345322 );
buf ( n350672 , n343953 );
nand ( n30640 , n350671 , n350672 );
buf ( n350674 , n30640 );
buf ( n350675 , n350674 );
nand ( n30643 , n30637 , n350675 );
buf ( n30644 , n30643 );
not ( n350678 , n30644 );
or ( n30646 , n350665 , n350678 );
nand ( n350680 , n344595 , n343948 );
nand ( n350681 , n30646 , n350680 );
buf ( n350682 , n350681 );
xor ( n350683 , n30631 , n350682 );
not ( n30651 , n343531 );
not ( n350685 , n602 );
not ( n350686 , n344353 );
or ( n30654 , n350685 , n350686 );
nand ( n30655 , n343553 , n344361 );
nand ( n350689 , n30654 , n30655 );
not ( n30657 , n350689 );
or ( n350691 , n30651 , n30657 );
nand ( n30659 , n344738 , n343595 );
nand ( n30660 , n350691 , n30659 );
buf ( n350694 , n30660 );
xnor ( n350695 , n350683 , n350694 );
buf ( n350696 , n350695 );
not ( n350697 , n344751 );
not ( n350698 , n344655 );
not ( n30666 , n350698 );
and ( n350700 , n350697 , n30666 );
nand ( n30668 , n344751 , n350698 );
buf ( n350702 , n344722 );
not ( n30670 , n350702 );
buf ( n350704 , n30670 );
and ( n30672 , n30668 , n350704 );
nor ( n350706 , n350700 , n30672 );
not ( n350707 , n350706 );
xor ( n30675 , n350696 , n350707 );
not ( n350709 , n344018 );
not ( n30677 , n24612 );
or ( n350711 , n350709 , n30677 );
buf ( n350712 , n600 );
not ( n30680 , n350712 );
buf ( n350714 , n24800 );
not ( n30682 , n350714 );
or ( n350716 , n30680 , n30682 );
buf ( n350717 , n343545 );
buf ( n350718 , n23906 );
nand ( n350719 , n350717 , n350718 );
buf ( n350720 , n350719 );
buf ( n350721 , n350720 );
nand ( n350722 , n350716 , n350721 );
buf ( n350723 , n350722 );
buf ( n350724 , n350723 );
buf ( n350725 , n344015 );
nand ( n350726 , n350724 , n350725 );
buf ( n350727 , n350726 );
nand ( n30695 , n350711 , n350727 );
buf ( n350729 , n344686 );
not ( n350730 , n350729 );
buf ( n350731 , n344717 );
nand ( n350732 , n350730 , n350731 );
buf ( n350733 , n350732 );
buf ( n30701 , n350733 );
not ( n30702 , n30701 );
buf ( n350736 , n344684 );
not ( n30704 , n350736 );
buf ( n350738 , n30704 );
buf ( n350739 , n350738 );
not ( n30707 , n350739 );
or ( n350741 , n30702 , n30707 );
buf ( n350742 , n344717 );
not ( n30710 , n350742 );
buf ( n350744 , n344686 );
nand ( n350745 , n30710 , n350744 );
buf ( n350746 , n350745 );
buf ( n350747 , n350746 );
nand ( n350748 , n350741 , n350747 );
buf ( n350749 , n350748 );
xor ( n350750 , n30695 , n350749 );
and ( n350751 , n343908 , n343624 );
not ( n350752 , n343908 );
and ( n30720 , n350752 , n592 );
or ( n350754 , n350751 , n30720 );
buf ( n350755 , n350754 );
buf ( n350756 , n23613 );
and ( n350757 , n350755 , n350756 );
buf ( n350758 , n343699 );
not ( n30726 , n350758 );
buf ( n350760 , n344697 );
nor ( n30728 , n30726 , n350760 );
buf ( n350762 , n30728 );
buf ( n350763 , n350762 );
nor ( n350764 , n350757 , n350763 );
buf ( n350765 , n350764 );
buf ( n350766 , n347904 );
not ( n30734 , n350766 );
buf ( n350768 , n592 );
nand ( n350769 , n30734 , n350768 );
buf ( n350770 , n350769 );
xor ( n30738 , n350765 , n350770 );
buf ( n350772 , n343765 );
not ( n350773 , n350772 );
buf ( n350774 , n344679 );
not ( n30742 , n350774 );
or ( n30743 , n350773 , n30742 );
buf ( n350777 , n343632 );
not ( n350778 , n350777 );
buf ( n350779 , n343966 );
not ( n30747 , n350779 );
or ( n350781 , n350778 , n30747 );
buf ( n350782 , n343966 );
buf ( n350783 , n343632 );
or ( n30751 , n350782 , n350783 );
nand ( n30752 , n350781 , n30751 );
buf ( n350786 , n30752 );
buf ( n350787 , n350786 );
buf ( n350788 , n23681 );
nand ( n350789 , n350787 , n350788 );
buf ( n350790 , n350789 );
buf ( n350791 , n350790 );
nand ( n350792 , n30743 , n350791 );
buf ( n350793 , n350792 );
xor ( n30761 , n30738 , n350793 );
xor ( n30762 , n350750 , n30761 );
xnor ( n350796 , n30675 , n30762 );
buf ( n350797 , n344271 );
not ( n30765 , n350797 );
buf ( n350799 , n24512 );
not ( n350800 , n350799 );
or ( n30768 , n30765 , n350800 );
buf ( n350802 , n344271 );
buf ( n350803 , n24512 );
or ( n350804 , n350802 , n350803 );
buf ( n350805 , n344636 );
nand ( n350806 , n350804 , n350805 );
buf ( n350807 , n350806 );
buf ( n350808 , n350807 );
nand ( n350809 , n30768 , n350808 );
buf ( n350810 , n350809 );
xor ( n350811 , n350796 , n350810 );
not ( n30779 , n344338 );
buf ( n350813 , n604 );
not ( n350814 , n350813 );
not ( n350815 , n24391 );
buf ( n350816 , n350815 );
not ( n350817 , n350816 );
or ( n350818 , n350814 , n350817 );
buf ( n350819 , n24392 );
not ( n350820 , n350819 );
buf ( n350821 , n350820 );
buf ( n350822 , n350821 );
buf ( n350823 , n23530 );
nand ( n350824 , n350822 , n350823 );
buf ( n350825 , n350824 );
buf ( n350826 , n350825 );
nand ( n350827 , n350818 , n350826 );
buf ( n350828 , n350827 );
not ( n30796 , n350828 );
or ( n350830 , n30779 , n30796 );
buf ( n350831 , n24729 );
buf ( n350832 , n344400 );
nand ( n30800 , n350831 , n350832 );
buf ( n350834 , n30800 );
nand ( n30802 , n350830 , n350834 );
not ( n30803 , n30802 );
not ( n350837 , n344454 );
not ( n350838 , n344626 );
or ( n30806 , n350837 , n350838 );
not ( n350840 , n606 );
not ( n350841 , n22150 );
not ( n30809 , n350841 );
nand ( n350843 , n334232 , n14213 , n14387 );
nand ( n350844 , n334617 , n14771 );
nor ( n30812 , n350843 , n350844 );
nand ( n30813 , n30812 , n14668 );
not ( n350847 , n30813 );
or ( n350848 , n30809 , n350847 );
nand ( n30816 , n30812 , n14668 , n22150 );
nand ( n350850 , n350848 , n30816 );
buf ( n350851 , n350850 );
not ( n30819 , n350851 );
buf ( n30820 , n30819 );
not ( n350854 , n30820 );
or ( n30822 , n350840 , n350854 );
buf ( n350856 , n344445 );
buf ( n350857 , n350850 );
nand ( n350858 , n350856 , n350857 );
buf ( n350859 , n350858 );
nand ( n30827 , n30822 , n350859 );
nand ( n350861 , n30827 , n607 );
nand ( n30829 , n30806 , n350861 );
not ( n350863 , n30829 );
xor ( n30831 , n344570 , n24546 );
and ( n30832 , n30831 , n344605 );
and ( n350866 , n344570 , n24546 );
or ( n30834 , n30832 , n350866 );
buf ( n350868 , n30834 );
not ( n30836 , n350868 );
buf ( n350870 , n30836 );
and ( n350871 , n350863 , n350870 );
not ( n350872 , n350863 );
and ( n30840 , n350872 , n30834 );
nor ( n350874 , n350871 , n30840 );
nand ( n350875 , n30803 , n350874 );
not ( n30843 , n350863 );
or ( n350877 , n30843 , n350870 );
or ( n350878 , n350863 , n30834 );
nand ( n350879 , n350877 , n350878 , n30802 );
nand ( n30847 , n350875 , n350879 );
not ( n350881 , n24601 );
not ( n350882 , n24573 );
not ( n30850 , n344551 );
nand ( n350884 , n350882 , n30850 );
not ( n350885 , n350884 );
or ( n350886 , n350881 , n350885 );
nand ( n30854 , n344551 , n24574 );
nand ( n350888 , n350886 , n30854 );
and ( n350889 , n30847 , n350888 );
not ( n30857 , n30847 );
not ( n350891 , n350888 );
and ( n350892 , n30857 , n350891 );
nor ( n350893 , n350889 , n350892 );
buf ( n350894 , n344772 );
buf ( n350895 , n344787 );
or ( n350896 , n350894 , n350895 );
buf ( n350897 , n344754 );
nand ( n30865 , n350896 , n350897 );
buf ( n30866 , n30865 );
buf ( n350900 , n344772 );
buf ( n350901 , n344787 );
nand ( n350902 , n350900 , n350901 );
buf ( n350903 , n350902 );
nand ( n350904 , n30866 , n350903 );
buf ( n30872 , n350904 );
and ( n30873 , n350893 , n30872 );
not ( n350907 , n350893 );
not ( n30875 , n30872 );
and ( n350909 , n350907 , n30875 );
nor ( n30877 , n30873 , n350909 );
xnor ( n30878 , n350811 , n30877 );
buf ( n350912 , n345061 );
not ( n350913 , n350912 );
buf ( n350914 , n25025 );
nand ( n350915 , n350913 , n350914 );
buf ( n350916 , n350915 );
nand ( n30884 , n350916 , n344638 );
buf ( n350918 , n25024 );
buf ( n350919 , n345061 );
nand ( n350920 , n350918 , n350919 );
buf ( n350921 , n350920 );
nand ( n350922 , n30884 , n350921 );
buf ( n350923 , n350922 );
not ( n30891 , n350923 );
buf ( n30892 , n30891 );
nand ( n350926 , n30878 , n30892 );
buf ( n350927 , n350926 );
buf ( n30895 , n350927 );
buf ( n350929 , n30895 );
buf ( n350930 , n30892 );
not ( n350931 , n350930 );
buf ( n350932 , n30878 );
not ( n30900 , n350932 );
buf ( n350934 , n30900 );
buf ( n350935 , n350934 );
nand ( n350936 , n350931 , n350935 );
buf ( n350937 , n350936 );
nand ( n30905 , n350929 , n350937 );
not ( n30906 , n30905 );
and ( n350940 , n350650 , n30906 );
not ( n350941 , n350650 );
and ( n30909 , n350941 , n30905 );
nor ( n350943 , n350940 , n30909 );
buf ( n30911 , n350943 );
buf ( n30912 , n30911 );
buf ( n350946 , n30912 );
xor ( n350947 , n343521 , n23525 );
xor ( n350948 , n350947 , n350946 );
buf ( n350949 , n350948 );
xor ( n30917 , n343521 , n23525 );
and ( n350951 , n30917 , n350946 );
and ( n350952 , n343521 , n23525 );
or ( n30920 , n350951 , n350952 );
buf ( n350954 , n30920 );
buf ( n350955 , n320951 );
buf ( n350956 , n320946 );
not ( n30924 , n349257 );
not ( n350958 , n349254 );
or ( n30926 , n30924 , n350958 );
nand ( n30927 , n30926 , n349247 );
buf ( n350961 , n30927 );
buf ( n350962 , n349214 );
xnor ( n30930 , n350961 , n350962 );
buf ( n30931 , n30930 );
buf ( n350965 , n30931 );
xor ( n30933 , n350955 , n350956 );
xor ( n30934 , n30933 , n350965 );
buf ( n350968 , n30934 );
xor ( n350969 , n350955 , n350956 );
and ( n30937 , n350969 , n350965 );
and ( n350971 , n350955 , n350956 );
or ( n350972 , n30937 , n350971 );
buf ( n350973 , n350972 );
buf ( n350974 , n320658 );
buf ( n350975 , n320752 );
buf ( n350976 , n349309 );
buf ( n30944 , n350976 );
buf ( n350978 , n30944 );
buf ( n350979 , n29262 );
not ( n350980 , n350979 );
buf ( n350981 , n350980 );
not ( n30949 , n350981 );
nand ( n350983 , n350978 , n30949 );
not ( n30951 , n349261 );
and ( n350985 , n350983 , n30951 );
not ( n30953 , n350983 );
and ( n350987 , n30953 , n349261 );
nor ( n350988 , n350985 , n350987 );
buf ( n350989 , n350988 );
xor ( n350990 , n350974 , n350975 );
xor ( n350991 , n350990 , n350989 );
buf ( n350992 , n350991 );
xor ( n30960 , n350974 , n350975 );
and ( n350994 , n30960 , n350989 );
and ( n350995 , n350974 , n350975 );
or ( n30963 , n350994 , n350995 );
buf ( n350997 , n30963 );
buf ( n350998 , n320803 );
buf ( n350999 , n14144 );
buf ( n351000 , n349330 );
not ( n351001 , n351000 );
buf ( n351002 , n349336 );
nand ( n30970 , n351001 , n351002 );
buf ( n351004 , n30970 );
buf ( n351005 , n351004 );
buf ( n351006 , n349312 );
and ( n351007 , n351005 , n351006 );
not ( n30975 , n351005 );
not ( n351009 , n349312 );
buf ( n351010 , n351009 );
and ( n30978 , n30975 , n351010 );
nor ( n30979 , n351007 , n30978 );
buf ( n351013 , n30979 );
buf ( n30981 , n351013 );
xor ( n30982 , n350998 , n350999 );
xor ( n30983 , n30982 , n30981 );
buf ( n351017 , n30983 );
xor ( n351018 , n350998 , n350999 );
and ( n351019 , n351018 , n30981 );
and ( n30987 , n350998 , n350999 );
or ( n30988 , n351019 , n30987 );
buf ( n351022 , n30988 );
buf ( n351023 , n321111 );
buf ( n351024 , n14156 );
xor ( n351025 , n349082 , n349340 );
xor ( n30993 , n351025 , n349360 );
buf ( n351027 , n30993 );
buf ( n351028 , n351027 );
xor ( n351029 , n351023 , n351024 );
xor ( n30997 , n351029 , n351028 );
buf ( n351031 , n30997 );
xor ( n351032 , n351023 , n351024 );
and ( n31000 , n351032 , n351028 );
and ( n351034 , n351023 , n351024 );
or ( n31002 , n31000 , n351034 );
buf ( n351036 , n31002 );
buf ( n351037 , n322438 );
buf ( n351038 , n334015 );
not ( n351039 , n349797 );
xor ( n351040 , n351039 , n29750 );
not ( n31008 , n29574 );
xor ( n31009 , n351040 , n31008 );
not ( n351043 , n31009 );
buf ( n351044 , n351043 );
buf ( n351045 , n351044 );
xor ( n351046 , n351037 , n351038 );
xor ( n351047 , n351046 , n351045 );
buf ( n351048 , n351047 );
xor ( n351049 , n351037 , n351038 );
and ( n351050 , n351049 , n351045 );
and ( n351051 , n351037 , n351038 );
or ( n351052 , n351050 , n351051 );
buf ( n351053 , n351052 );
buf ( n351054 , n324344 );
buf ( n351055 , n334005 );
and ( n351056 , n350298 , n350181 );
buf ( n31024 , n349995 );
and ( n31025 , n351056 , n31024 );
not ( n351059 , n351056 );
not ( n351060 , n31024 );
and ( n31028 , n351059 , n351060 );
nor ( n351062 , n31025 , n31028 );
buf ( n351063 , n351062 );
buf ( n351064 , n351063 );
xor ( n351065 , n351054 , n351055 );
xor ( n351066 , n351065 , n351064 );
buf ( n351067 , n351066 );
xor ( n31035 , n351054 , n351055 );
and ( n351069 , n31035 , n351064 );
and ( n351070 , n351054 , n351055 );
or ( n31038 , n351069 , n351070 );
buf ( n351072 , n31038 );
buf ( n351073 , n331910 );
buf ( n351074 , n331824 );
buf ( n351075 , n350595 );
buf ( n351076 , n351075 );
buf ( n351077 , n351076 );
not ( n351078 , n351077 );
buf ( n351079 , n346430 );
not ( n351080 , n351079 );
buf ( n351081 , n351080 );
not ( n31049 , n351081 );
buf ( n351083 , n345970 );
buf ( n31051 , n351083 );
buf ( n351085 , n31051 );
nor ( n31053 , n31049 , n351085 );
not ( n31054 , n31053 );
or ( n351088 , n351078 , n31054 );
buf ( n351089 , n350626 );
buf ( n31057 , n351089 );
buf ( n31058 , n31057 );
nand ( n351092 , n351088 , n31058 );
buf ( n351093 , n350642 );
buf ( n351094 , n350621 );
buf ( n351095 , n351094 );
nand ( n351096 , n351093 , n351095 );
buf ( n351097 , n351096 );
buf ( n351098 , n351097 );
not ( n351099 , n351098 );
buf ( n351100 , n351099 );
and ( n31068 , n351092 , n351100 );
not ( n351102 , n351092 );
and ( n351103 , n351102 , n351097 );
nor ( n31071 , n31068 , n351103 );
buf ( n31072 , n31071 );
not ( n31073 , n31072 );
not ( n351107 , n31073 );
buf ( n351108 , n351107 );
xor ( n31076 , n351073 , n351074 );
xor ( n31077 , n31076 , n351108 );
buf ( n351111 , n31077 );
xor ( n351112 , n351073 , n351074 );
and ( n351113 , n351112 , n351108 );
and ( n31081 , n351073 , n351074 );
or ( n31082 , n351113 , n31081 );
buf ( n351116 , n31082 );
buf ( n351117 , n324056 );
buf ( n351118 , n334014 );
buf ( n351119 , n350396 );
buf ( n351120 , n30356 );
nand ( n31088 , n351119 , n351120 );
buf ( n351122 , n31088 );
buf ( n351123 , n30280 );
buf ( n31091 , n351123 );
buf ( n351125 , n31091 );
xnor ( n31093 , n351122 , n351125 );
buf ( n351127 , n31093 );
xor ( n31095 , n351117 , n351118 );
xor ( n31096 , n31095 , n351127 );
buf ( n351130 , n31096 );
xor ( n31098 , n351117 , n351118 );
and ( n351132 , n31098 , n351127 );
and ( n351133 , n351117 , n351118 );
or ( n31101 , n351132 , n351133 );
buf ( n351135 , n31101 );
buf ( n351136 , n327542 );
buf ( n31104 , n334010 );
buf ( n351138 , n350508 );
not ( n31106 , n351138 );
buf ( n351140 , n350496 );
nand ( n31108 , n31106 , n351140 );
buf ( n351142 , n31108 );
buf ( n351143 , n30450 );
not ( n351144 , n351143 );
buf ( n351145 , n351144 );
buf ( n351146 , n351145 );
not ( n31114 , n351146 );
buf ( n351148 , n350397 );
not ( n351149 , n351148 );
or ( n351150 , n31114 , n351149 );
buf ( n351151 , n350501 );
not ( n351152 , n351151 );
buf ( n351153 , n351152 );
buf ( n351154 , n351153 );
nand ( n351155 , n351150 , n351154 );
buf ( n351156 , n351155 );
xnor ( n31124 , n351142 , n351156 );
buf ( n351158 , n31124 );
buf ( n31126 , n351158 );
buf ( n351160 , n31126 );
buf ( n351161 , n351160 );
xor ( n351162 , n351136 , n31104 );
xor ( n31130 , n351162 , n351161 );
buf ( n351164 , n31130 );
xor ( n351165 , n351136 , n31104 );
and ( n31133 , n351165 , n351161 );
and ( n351167 , n351136 , n31104 );
or ( n351168 , n31133 , n351167 );
buf ( n351169 , n351168 );
buf ( n351170 , n327374 );
buf ( n351171 , n7530 );
buf ( n351172 , n350512 );
buf ( n351173 , n351172 );
buf ( n351174 , n351173 );
buf ( n351175 , n351174 );
buf ( n351176 , n30522 );
not ( n31144 , n351176 );
buf ( n351178 , n31144 );
buf ( n351179 , n351178 );
buf ( n351180 , n348260 );
nand ( n31148 , n351179 , n351180 );
buf ( n351182 , n31148 );
buf ( n351183 , n351182 );
not ( n31151 , n351183 );
buf ( n31152 , n31151 );
buf ( n351186 , n31152 );
and ( n351187 , n351175 , n351186 );
not ( n351188 , n351175 );
buf ( n351189 , n351182 );
and ( n351190 , n351188 , n351189 );
nor ( n351191 , n351187 , n351190 );
buf ( n351192 , n351191 );
buf ( n351193 , n351192 );
buf ( n351194 , n351193 );
buf ( n351195 , n351194 );
buf ( n351196 , n351195 );
xor ( n31164 , n351170 , n351171 );
xor ( n31165 , n31164 , n351196 );
buf ( n351199 , n31165 );
xor ( n31167 , n351170 , n351171 );
and ( n31168 , n31167 , n351196 );
and ( n31169 , n351170 , n351171 );
or ( n31170 , n31168 , n31169 );
buf ( n351204 , n31170 );
buf ( n351205 , n326633 );
buf ( n351206 , n351205 );
buf ( n351207 , n326638 );
not ( n351208 , n348036 );
not ( n31176 , n348077 );
or ( n351210 , n351208 , n31176 );
nand ( n31178 , n351210 , n350547 );
not ( n31179 , n31178 );
not ( n31180 , n31179 );
buf ( n351214 , n348260 );
not ( n351215 , n351214 );
buf ( n351216 , n350512 );
not ( n31184 , n351216 );
or ( n351218 , n351215 , n31184 );
buf ( n351219 , n351178 );
nand ( n31187 , n351218 , n351219 );
buf ( n351221 , n31187 );
not ( n31189 , n351221 );
not ( n351223 , n31189 );
or ( n351224 , n31180 , n351223 );
nand ( n31192 , n351221 , n31178 );
nand ( n31193 , n351224 , n31192 );
not ( n31194 , n31193 );
buf ( n351228 , n31194 );
buf ( n351229 , n351228 );
not ( n31197 , n351229 );
buf ( n351231 , n31197 );
xor ( n31199 , n351206 , n351207 );
xor ( n351233 , n31199 , n351231 );
buf ( n351234 , n351233 );
xor ( n31202 , n351206 , n351207 );
and ( n351236 , n31202 , n351231 );
and ( n31204 , n351206 , n351207 );
or ( n31205 , n351236 , n31204 );
buf ( n351239 , n31205 );
buf ( n351240 , n326370 );
buf ( n351241 , n326478 );
buf ( n351242 , n348262 );
not ( n31210 , n351242 );
buf ( n351244 , n351174 );
not ( n351245 , n351244 );
or ( n31213 , n31210 , n351245 );
and ( n351247 , n350547 , n350556 );
buf ( n351248 , n351247 );
nand ( n31216 , n31213 , n351248 );
buf ( n351250 , n31216 );
buf ( n351251 , n350563 );
not ( n31219 , n350562 );
nand ( n351253 , n31219 , n350532 );
buf ( n351254 , n351253 );
nand ( n351255 , n351251 , n351254 );
buf ( n351256 , n351255 );
buf ( n351257 , n351256 );
not ( n31225 , n351257 );
buf ( n351259 , n31225 );
and ( n351260 , n351250 , n351259 );
not ( n31228 , n351250 );
and ( n351262 , n31228 , n351256 );
nor ( n31230 , n351260 , n351262 );
buf ( n31231 , n31230 );
buf ( n351265 , n31231 );
xor ( n351266 , n351240 , n351241 );
xor ( n351267 , n351266 , n351265 );
buf ( n351268 , n351267 );
xor ( n351269 , n351240 , n351241 );
and ( n351270 , n351269 , n351265 );
and ( n31238 , n351240 , n351241 );
or ( n351272 , n351270 , n31238 );
buf ( n351273 , n351272 );
buf ( n351274 , n326959 );
buf ( n351275 , n327094 );
nand ( n351276 , n347502 , n27472 );
not ( n351277 , n351276 );
nand ( n31245 , n30506 , n350559 , n350563 );
not ( n351279 , n31245 );
or ( n351280 , n351277 , n351279 );
buf ( n31248 , n350570 );
buf ( n31249 , n31248 );
buf ( n31250 , n31249 );
nand ( n351284 , n351280 , n31250 );
nand ( n31252 , n350569 , n350571 );
not ( n31253 , n31252 );
and ( n351287 , n351284 , n31253 );
not ( n351288 , n351284 );
and ( n31256 , n351288 , n31252 );
nor ( n351290 , n351287 , n31256 );
buf ( n351291 , n351290 );
not ( n351292 , n351291 );
not ( n31260 , n351292 );
buf ( n351294 , n31260 );
buf ( n351295 , n351294 );
xor ( n351296 , n351274 , n351275 );
xor ( n351297 , n351296 , n351295 );
buf ( n351298 , n351297 );
xor ( n31266 , n351274 , n351275 );
and ( n351300 , n31266 , n351295 );
and ( n31268 , n351274 , n351275 );
or ( n351302 , n351300 , n31268 );
buf ( n351303 , n351302 );
buf ( n351304 , n331459 );
buf ( n351305 , n14151 );
nand ( n31273 , n351077 , n351081 );
not ( n351307 , n31273 );
not ( n351308 , n31058 );
nor ( n31276 , n351308 , n351085 );
nand ( n351310 , n351307 , n31276 );
not ( n351311 , n351085 );
not ( n31279 , n351311 );
not ( n31280 , n31058 );
or ( n351314 , n31279 , n31280 );
nand ( n351315 , n351314 , n31273 );
nand ( n31283 , n351310 , n351315 );
not ( n351317 , n31283 );
not ( n351318 , n351317 );
buf ( n31286 , n351318 );
not ( n351320 , n31286 );
buf ( n31288 , n351320 );
xor ( n31289 , n351304 , n351305 );
xor ( n351323 , n31289 , n31288 );
buf ( n351324 , n351323 );
xor ( n31292 , n351304 , n351305 );
and ( n351326 , n31292 , n31288 );
and ( n351327 , n351304 , n351305 );
or ( n31295 , n351326 , n351327 );
buf ( n351329 , n31295 );
buf ( n351330 , n323822 );
buf ( n351331 , n324005 );
buf ( n351332 , n350184 );
not ( n351333 , n351332 );
buf ( n351334 , n351333 );
buf ( n351335 , n350301 );
not ( n351336 , n351335 );
buf ( n351337 , n351336 );
nand ( n31305 , n351334 , n351337 );
nand ( n351339 , n350310 , n30258 );
not ( n351340 , n351339 );
and ( n31308 , n31305 , n351340 );
not ( n351342 , n31305 );
and ( n351343 , n351342 , n351339 );
nor ( n31311 , n31308 , n351343 );
buf ( n351345 , n31311 );
buf ( n351346 , n351345 );
xor ( n31314 , n351330 , n351331 );
xor ( n351348 , n31314 , n351346 );
buf ( n351349 , n351348 );
xor ( n351350 , n351330 , n351331 );
and ( n31318 , n351350 , n351346 );
and ( n351352 , n351330 , n351331 );
or ( n31320 , n31318 , n351352 );
buf ( n351354 , n31320 );
buf ( n351355 , n332112 );
buf ( n351356 , n332119 );
nand ( n351357 , n30615 , n345397 );
not ( n31325 , n351357 );
not ( n31326 , n30611 );
or ( n351360 , n31325 , n31326 );
not ( n351361 , n351357 );
nand ( n31329 , n350642 , n30597 );
nand ( n351363 , n351361 , n31329 );
nand ( n351364 , n351360 , n351363 );
buf ( n351365 , n351364 );
buf ( n351366 , n351365 );
buf ( n351367 , n351366 );
buf ( n351368 , n351367 );
xor ( n31336 , n351355 , n351356 );
xor ( n351370 , n31336 , n351368 );
buf ( n351371 , n351370 );
xor ( n31339 , n351355 , n351356 );
and ( n351373 , n31339 , n351368 );
and ( n351374 , n351355 , n351356 );
or ( n351375 , n351373 , n351374 );
buf ( n351376 , n351375 );
buf ( n351377 , n321253 );
buf ( n351378 , n14143 );
xor ( n31346 , n351377 , n351378 );
buf ( n351380 , n31346 );
and ( n351381 , n351377 , n351378 );
buf ( n351382 , n351381 );
buf ( n351383 , n332801 );
buf ( n351384 , n332794 );
xor ( n31352 , n351383 , n351384 );
buf ( n351386 , n31352 );
buf ( n351387 , n332589 );
buf ( n351388 , n332582 );
xor ( n351389 , n351387 , n351388 );
nand ( n31357 , n345397 , n350926 );
buf ( n351391 , n350633 );
buf ( n351392 , n350638 );
nor ( n351393 , n351391 , n351392 );
buf ( n351394 , n351393 );
nor ( n351395 , n31357 , n351394 );
not ( n31363 , n351395 );
not ( n351397 , n30597 );
or ( n31365 , n31363 , n351397 );
nand ( n31366 , n350926 , n350647 );
buf ( n351400 , n31366 );
buf ( n351401 , n350937 );
nand ( n351402 , n351400 , n351401 );
buf ( n351403 , n351402 );
buf ( n351404 , n351403 );
not ( n351405 , n351404 );
buf ( n351406 , n351405 );
nand ( n351407 , n31365 , n351406 );
buf ( n351408 , n607 );
not ( n31376 , n351408 );
buf ( n351410 , n606 );
not ( n351411 , n351410 );
not ( n351412 , n15992 );
not ( n31380 , n351412 );
not ( n351414 , n334058 );
nor ( n351415 , n351414 , n14667 );
nand ( n31383 , n351415 , n30812 );
not ( n351417 , n31383 );
not ( n351418 , n351417 );
or ( n31386 , n31380 , n351418 );
not ( n351420 , n14349 );
not ( n31388 , n351420 );
nand ( n351422 , n31388 , n31383 );
nand ( n31390 , n31386 , n351422 );
not ( n351424 , n31390 );
buf ( n351425 , n351424 );
not ( n31393 , n351425 );
buf ( n351427 , n31393 );
buf ( n351428 , n351427 );
not ( n351429 , n351428 );
or ( n31397 , n351411 , n351429 );
buf ( n351431 , n31390 );
not ( n351432 , n351431 );
buf ( n351433 , n351432 );
buf ( n351434 , n351433 );
buf ( n351435 , n344445 );
nand ( n31403 , n351434 , n351435 );
buf ( n351437 , n31403 );
buf ( n351438 , n351437 );
nand ( n351439 , n31397 , n351438 );
buf ( n351440 , n351439 );
buf ( n351441 , n351440 );
not ( n351442 , n351441 );
or ( n31410 , n31376 , n351442 );
nand ( n351444 , n30827 , n344454 );
buf ( n351445 , n351444 );
nand ( n31413 , n31410 , n351445 );
buf ( n351447 , n31413 );
buf ( n351448 , n23613 );
buf ( n351449 , n350754 );
and ( n351450 , n351448 , n351449 );
buf ( n351451 , n350762 );
nor ( n31419 , n351450 , n351451 );
buf ( n351453 , n31419 );
buf ( n351454 , n351453 );
not ( n351455 , n351454 );
buf ( n351456 , n350770 );
not ( n351457 , n351456 );
and ( n351458 , n351455 , n351457 );
buf ( n351459 , n350793 );
buf ( n351460 , n351453 );
buf ( n351461 , n350770 );
nand ( n31429 , n351460 , n351461 );
buf ( n351463 , n31429 );
buf ( n351464 , n351463 );
and ( n351465 , n351459 , n351464 );
nor ( n31433 , n351458 , n351465 );
buf ( n31434 , n31433 );
buf ( n351468 , n31434 );
not ( n31436 , n351468 );
buf ( n351470 , n343837 );
buf ( n351471 , n592 );
and ( n31439 , n351470 , n351471 );
buf ( n351473 , n31439 );
buf ( n351474 , n351473 );
buf ( n351475 , n23613 );
not ( n31443 , n351475 );
and ( n31444 , n592 , n343872 );
not ( n31445 , n592 );
and ( n351479 , n31445 , n343869 );
or ( n351480 , n31444 , n351479 );
buf ( n351481 , n351480 );
not ( n351482 , n351481 );
or ( n31450 , n31443 , n351482 );
buf ( n351484 , n350754 );
buf ( n351485 , n344705 );
nand ( n31453 , n351484 , n351485 );
buf ( n351487 , n31453 );
buf ( n351488 , n351487 );
nand ( n31456 , n31450 , n351488 );
buf ( n31457 , n31456 );
buf ( n351491 , n31457 );
xor ( n31459 , n351474 , n351491 );
buf ( n351493 , n23681 );
not ( n351494 , n351493 );
buf ( n351495 , n594 );
not ( n31463 , n351495 );
buf ( n351497 , n343985 );
not ( n351498 , n351497 );
or ( n351499 , n31463 , n351498 );
buf ( n351500 , n343982 );
buf ( n351501 , n343632 );
nand ( n31469 , n351500 , n351501 );
buf ( n351503 , n31469 );
buf ( n351504 , n351503 );
nand ( n31472 , n351499 , n351504 );
buf ( n351506 , n31472 );
buf ( n351507 , n351506 );
not ( n351508 , n351507 );
or ( n31476 , n351494 , n351508 );
buf ( n351510 , n350786 );
buf ( n351511 , n343765 );
nand ( n351512 , n351510 , n351511 );
buf ( n351513 , n351512 );
buf ( n351514 , n351513 );
nand ( n31482 , n31476 , n351514 );
buf ( n351516 , n31482 );
buf ( n351517 , n351516 );
xor ( n31485 , n31459 , n351517 );
buf ( n351519 , n31485 );
buf ( n351520 , n351519 );
not ( n351521 , n351520 );
or ( n31489 , n31436 , n351521 );
buf ( n351523 , n351519 );
buf ( n351524 , n31434 );
or ( n351525 , n351523 , n351524 );
nand ( n31493 , n31489 , n351525 );
buf ( n31494 , n31493 );
xor ( n351528 , n351447 , n31494 );
buf ( n351529 , n351528 );
not ( n31497 , n351529 );
buf ( n31498 , n31497 );
xor ( n31499 , n30695 , n350749 );
and ( n351533 , n31499 , n30761 );
and ( n351534 , n30695 , n350749 );
or ( n31502 , n351533 , n351534 );
not ( n351536 , n31502 );
buf ( n351537 , n343863 );
not ( n31505 , n351537 );
buf ( n351539 , n596 );
not ( n31507 , n351539 );
buf ( n351541 , n344055 );
not ( n31509 , n351541 );
or ( n351543 , n31507 , n31509 );
buf ( n351544 , n344588 );
buf ( n351545 , n343882 );
nand ( n351546 , n351544 , n351545 );
buf ( n351547 , n351546 );
buf ( n351548 , n351547 );
nand ( n351549 , n351543 , n351548 );
buf ( n351550 , n351549 );
buf ( n351551 , n351550 );
not ( n31519 , n351551 );
or ( n31520 , n31505 , n31519 );
buf ( n351554 , n350656 );
buf ( n351555 , n23889 );
nand ( n31523 , n351554 , n351555 );
buf ( n351557 , n31523 );
buf ( n351558 , n351557 );
nand ( n351559 , n31520 , n351558 );
buf ( n351560 , n351559 );
buf ( n351561 , n343948 );
not ( n31529 , n351561 );
buf ( n351563 , n30644 );
not ( n351564 , n351563 );
or ( n31532 , n31529 , n351564 );
and ( n351566 , n14695 , n343953 );
not ( n31534 , n14695 );
and ( n351568 , n31534 , n598 );
or ( n31536 , n351566 , n351568 );
buf ( n351570 , n31536 );
buf ( n351571 , n23911 );
nand ( n31539 , n351570 , n351571 );
buf ( n351573 , n31539 );
buf ( n351574 , n351573 );
nand ( n31542 , n31532 , n351574 );
buf ( n31543 , n31542 );
xor ( n351577 , n351560 , n31543 );
buf ( n351578 , n351577 );
buf ( n351579 , n344015 );
not ( n351580 , n351579 );
and ( n31548 , n600 , n344383 );
not ( n31549 , n600 );
and ( n351583 , n31549 , n24346 );
or ( n31551 , n31548 , n351583 );
buf ( n31552 , n31551 );
not ( n31553 , n31552 );
or ( n31554 , n351580 , n31553 );
buf ( n351588 , n350723 );
buf ( n351589 , n344018 );
nand ( n351590 , n351588 , n351589 );
buf ( n351591 , n351590 );
buf ( n351592 , n351591 );
nand ( n31560 , n31554 , n351592 );
buf ( n31561 , n31560 );
buf ( n351595 , n31561 );
buf ( n31563 , n351595 );
buf ( n31564 , n31563 );
buf ( n31565 , n31564 );
not ( n351599 , n31565 );
buf ( n351600 , n351599 );
buf ( n351601 , n351600 );
and ( n31569 , n351578 , n351601 );
not ( n31570 , n351578 );
buf ( n351604 , n31564 );
and ( n31572 , n31570 , n351604 );
nor ( n351606 , n31569 , n31572 );
buf ( n351607 , n351606 );
and ( n31575 , n351536 , n351607 );
not ( n351609 , n351536 );
buf ( n351610 , n351607 );
not ( n31578 , n351610 );
buf ( n31579 , n31578 );
and ( n351613 , n351609 , n31579 );
nor ( n31581 , n31575 , n351613 );
or ( n351615 , n31498 , n31581 );
nand ( n351616 , n31581 , n31498 );
nand ( n351617 , n351615 , n351616 );
buf ( n351618 , n351617 );
not ( n351619 , n350904 );
nand ( n351620 , n351619 , n350891 );
not ( n31588 , n351620 );
buf ( n351622 , n30847 );
buf ( n351623 , n351622 );
buf ( n351624 , n351623 );
not ( n351625 , n351624 );
or ( n31593 , n31588 , n351625 );
not ( n351627 , n350891 );
nand ( n31595 , n351627 , n350904 );
nand ( n351629 , n31593 , n31595 );
buf ( n351630 , n351629 );
xor ( n31598 , n351618 , n351630 );
buf ( n31599 , n350696 );
not ( n351633 , n31599 );
buf ( n351634 , n351633 );
buf ( n351635 , n351634 );
not ( n351636 , n351635 );
buf ( n351637 , n350707 );
not ( n351638 , n351637 );
or ( n351639 , n351636 , n351638 );
buf ( n351640 , n350696 );
not ( n31608 , n351640 );
buf ( n351642 , n350706 );
not ( n351643 , n351642 );
or ( n31611 , n31608 , n351643 );
buf ( n351645 , n30762 );
nand ( n351646 , n31611 , n351645 );
buf ( n351647 , n351646 );
buf ( n351648 , n351647 );
nand ( n351649 , n351639 , n351648 );
buf ( n351650 , n351649 );
not ( n31618 , n30802 );
nand ( n31619 , n31618 , n350863 );
buf ( n351653 , n30834 );
buf ( n351654 , n351653 );
buf ( n351655 , n351654 );
and ( n31623 , n31619 , n351655 );
buf ( n351657 , n30802 );
buf ( n351658 , n30829 );
and ( n351659 , n351657 , n351658 );
buf ( n351660 , n351659 );
nor ( n351661 , n31623 , n351660 );
not ( n351662 , n351661 );
xor ( n31630 , n351650 , n351662 );
xor ( n31631 , n344618 , n23530 );
buf ( n351665 , n31631 );
not ( n351666 , n351665 );
buf ( n351667 , n29097 );
not ( n351668 , n351667 );
and ( n31636 , n351666 , n351668 );
buf ( n351670 , n350828 );
buf ( n351671 , n344400 );
and ( n351672 , n351670 , n351671 );
nor ( n31640 , n31636 , n351672 );
buf ( n351674 , n31640 );
not ( n351675 , n351674 );
not ( n351676 , n351675 );
buf ( n351677 , n30630 );
not ( n351678 , n351677 );
buf ( n351679 , n351678 );
not ( n31647 , n351679 );
buf ( n351681 , n350681 );
not ( n351682 , n351681 );
buf ( n351683 , n351682 );
not ( n31651 , n351683 );
or ( n351685 , n31647 , n31651 );
nand ( n351686 , n351685 , n30660 );
nand ( n31654 , n350681 , n30630 );
nand ( n351688 , n351686 , n31654 );
not ( n351689 , n343531 );
buf ( n351690 , n602 );
not ( n351691 , n351690 );
buf ( n351692 , n344435 );
not ( n351693 , n351692 );
or ( n31661 , n351691 , n351693 );
buf ( n351695 , n344435 );
not ( n31663 , n351695 );
buf ( n351697 , n31663 );
buf ( n351698 , n351697 );
buf ( n351699 , n343553 );
nand ( n351700 , n351698 , n351699 );
buf ( n351701 , n351700 );
buf ( n351702 , n351701 );
nand ( n351703 , n31661 , n351702 );
buf ( n351704 , n351703 );
not ( n31672 , n351704 );
or ( n351706 , n351689 , n31672 );
buf ( n351707 , n350689 );
buf ( n351708 , n343595 );
nand ( n351709 , n351707 , n351708 );
buf ( n351710 , n351709 );
nand ( n351711 , n351706 , n351710 );
and ( n31679 , n351688 , n351711 );
not ( n351713 , n351688 );
not ( n351714 , n351711 );
and ( n31682 , n351713 , n351714 );
nor ( n351716 , n31679 , n31682 );
not ( n351717 , n351716 );
or ( n31685 , n351676 , n351717 );
or ( n351719 , n351716 , n351675 );
nand ( n31687 , n31685 , n351719 );
buf ( n351721 , n31687 );
not ( n31689 , n351721 );
buf ( n351723 , n31689 );
xor ( n351724 , n31630 , n351723 );
buf ( n351725 , n351724 );
xnor ( n351726 , n31598 , n351725 );
buf ( n351727 , n351726 );
not ( n31695 , n30877 );
buf ( n31696 , n350796 );
buf ( n351730 , n31696 );
buf ( n351731 , n351730 );
not ( n351732 , n351731 );
nand ( n351733 , n31695 , n351732 );
buf ( n31701 , n350810 );
and ( n351735 , n351733 , n31701 );
buf ( n351736 , n351731 );
not ( n351737 , n351736 );
buf ( n351738 , n31695 );
nor ( n351739 , n351737 , n351738 );
buf ( n351740 , n351739 );
nor ( n31708 , n351735 , n351740 );
nand ( n351742 , n351727 , n31708 );
buf ( n351743 , n351742 );
not ( n351744 , n351743 );
nor ( n31712 , n351727 , n31708 );
buf ( n351746 , n31712 );
not ( n31714 , n351746 );
buf ( n351748 , n31714 );
buf ( n351749 , n351748 );
not ( n351750 , n351749 );
buf ( n351751 , n351750 );
buf ( n351752 , n351751 );
nor ( n351753 , n351744 , n351752 );
buf ( n351754 , n351753 );
and ( n31722 , n351407 , n351754 );
not ( n351756 , n351407 );
buf ( n351757 , n351754 );
not ( n31725 , n351757 );
buf ( n31726 , n31725 );
and ( n351760 , n351756 , n31726 );
nor ( n31728 , n31722 , n351760 );
buf ( n351762 , n31728 );
buf ( n31730 , n351762 );
buf ( n351764 , n31730 );
buf ( n351765 , n351764 );
and ( n31733 , n351389 , n351765 );
and ( n351767 , n351387 , n351388 );
or ( n31735 , n31733 , n351767 );
buf ( n351769 , n31735 );
buf ( n351770 , n351769 );
buf ( n351771 , n332686 );
buf ( n351772 , n332693 );
xor ( n351773 , n351771 , n351772 );
not ( n351774 , n351742 );
nor ( n31742 , n351774 , n31357 );
not ( n351776 , n31742 );
not ( n351777 , n30611 );
or ( n31745 , n351776 , n351777 );
buf ( n351779 , n351742 );
not ( n351780 , n351779 );
buf ( n351781 , n351403 );
not ( n31749 , n351781 );
or ( n351783 , n351780 , n31749 );
buf ( n31751 , n351748 );
nand ( n31752 , n351783 , n31751 );
buf ( n31753 , n31752 );
buf ( n351787 , n31753 );
not ( n31755 , n351787 );
buf ( n351789 , n31755 );
nand ( n31757 , n31745 , n351789 );
not ( n351791 , n344015 );
buf ( n351792 , n600 );
not ( n31760 , n351792 );
buf ( n351794 , n344353 );
not ( n31762 , n351794 );
or ( n351796 , n31760 , n31762 );
buf ( n351797 , n344361 );
buf ( n351798 , n23906 );
nand ( n31766 , n351797 , n351798 );
buf ( n351800 , n31766 );
buf ( n351801 , n351800 );
nand ( n351802 , n351796 , n351801 );
buf ( n351803 , n351802 );
not ( n31771 , n351803 );
or ( n31772 , n351791 , n31771 );
buf ( n351806 , n31551 );
buf ( n351807 , n344018 );
nand ( n31775 , n351806 , n351807 );
buf ( n351809 , n31775 );
nand ( n31777 , n31772 , n351809 );
buf ( n351811 , n31777 );
not ( n31779 , n351811 );
buf ( n351813 , n23681 );
not ( n31781 , n351813 );
buf ( n351815 , n594 );
not ( n351816 , n351815 );
buf ( n351817 , n23996 );
not ( n31785 , n351817 );
or ( n351819 , n351816 , n31785 );
buf ( n351820 , n344035 );
buf ( n351821 , n343632 );
nand ( n351822 , n351820 , n351821 );
buf ( n351823 , n351822 );
buf ( n351824 , n351823 );
nand ( n31792 , n351819 , n351824 );
buf ( n351826 , n31792 );
buf ( n351827 , n351826 );
not ( n31795 , n351827 );
or ( n351829 , n31781 , n31795 );
buf ( n351830 , n351506 );
buf ( n351831 , n343765 );
nand ( n31799 , n351830 , n351831 );
buf ( n351833 , n31799 );
buf ( n351834 , n351833 );
nand ( n31802 , n351829 , n351834 );
buf ( n351836 , n31802 );
not ( n351837 , n351836 );
buf ( n351838 , n23911 );
not ( n31806 , n351838 );
buf ( n31807 , n598 );
not ( n31808 , n31807 );
buf ( n31809 , n24800 );
not ( n31810 , n31809 );
or ( n31811 , n31808 , n31810 );
buf ( n351845 , n343545 );
buf ( n351846 , n343953 );
nand ( n31814 , n351845 , n351846 );
buf ( n351848 , n31814 );
buf ( n351849 , n351848 );
nand ( n351850 , n31811 , n351849 );
buf ( n351851 , n351850 );
buf ( n351852 , n351851 );
not ( n351853 , n351852 );
or ( n31821 , n31806 , n351853 );
buf ( n351855 , n31536 );
buf ( n351856 , n343948 );
nand ( n31824 , n351855 , n351856 );
buf ( n351858 , n31824 );
buf ( n351859 , n351858 );
nand ( n351860 , n31821 , n351859 );
buf ( n351861 , n351860 );
not ( n31829 , n351861 );
not ( n31830 , n31829 );
or ( n31831 , n351837 , n31830 );
not ( n351865 , n351836 );
nand ( n351866 , n351865 , n351861 );
nand ( n31834 , n31831 , n351866 );
not ( n31835 , n31834 );
or ( n31836 , n31779 , n31835 );
or ( n351870 , n31834 , n351811 );
nand ( n351871 , n31836 , n351870 );
buf ( n351872 , n351871 );
buf ( n351873 , n31434 );
not ( n31841 , n351873 );
buf ( n351875 , n31841 );
nor ( n351876 , n351447 , n351875 );
not ( n31844 , n351876 );
not ( n351878 , n351519 );
not ( n31846 , n351878 );
and ( n31847 , n31844 , n31846 );
buf ( n351881 , n607 );
not ( n351882 , n351881 );
buf ( n351883 , n351440 );
not ( n31851 , n351883 );
or ( n31852 , n351882 , n31851 );
buf ( n351886 , n351444 );
nand ( n351887 , n31852 , n351886 );
buf ( n351888 , n351887 );
and ( n31856 , n351888 , n351875 );
nor ( n31857 , n31847 , n31856 );
buf ( n351891 , n31857 );
xor ( n351892 , n351872 , n351891 );
xor ( n351893 , n351474 , n351491 );
and ( n31861 , n351893 , n351517 );
and ( n351895 , n351474 , n351491 );
or ( n31863 , n31861 , n351895 );
buf ( n351897 , n31863 );
not ( n351898 , n344338 );
and ( n31866 , n604 , n30820 );
not ( n351900 , n604 );
and ( n31868 , n351900 , n350850 );
or ( n31869 , n31866 , n31868 );
not ( n351903 , n31869 );
or ( n31871 , n351898 , n351903 );
buf ( n351905 , n31631 );
not ( n31873 , n351905 );
buf ( n351907 , n344400 );
nand ( n351908 , n31873 , n351907 );
buf ( n351909 , n351908 );
nand ( n351910 , n31871 , n351909 );
xor ( n351911 , n351897 , n351910 );
and ( n31879 , n347209 , n592 );
buf ( n351913 , n23613 );
not ( n351914 , n351913 );
nand ( n351915 , n343969 , n592 );
buf ( n351916 , n343966 );
buf ( n351917 , n343624 );
nand ( n31885 , n351916 , n351917 );
buf ( n351919 , n31885 );
nand ( n31887 , n351915 , n351919 );
buf ( n351921 , n31887 );
not ( n351922 , n351921 );
or ( n351923 , n351914 , n351922 );
buf ( n351924 , n351480 );
buf ( n351925 , n344705 );
nand ( n351926 , n351924 , n351925 );
buf ( n351927 , n351926 );
buf ( n351928 , n351927 );
nand ( n351929 , n351923 , n351928 );
buf ( n351930 , n351929 );
xor ( n31898 , n31879 , n351930 );
buf ( n351932 , n343863 );
not ( n351933 , n351932 );
buf ( n351934 , n596 );
not ( n351935 , n351934 );
buf ( n351936 , n344301 );
not ( n31904 , n351936 );
or ( n351938 , n351935 , n31904 );
buf ( n351939 , n345322 );
buf ( n351940 , n343882 );
nand ( n351941 , n351939 , n351940 );
buf ( n351942 , n351941 );
buf ( n351943 , n351942 );
nand ( n31911 , n351938 , n351943 );
buf ( n351945 , n31911 );
buf ( n351946 , n351945 );
not ( n31914 , n351946 );
or ( n31915 , n351933 , n31914 );
buf ( n351949 , n351550 );
buf ( n351950 , n23889 );
nand ( n351951 , n351949 , n351950 );
buf ( n351952 , n351951 );
buf ( n351953 , n351952 );
nand ( n351954 , n31915 , n351953 );
buf ( n351955 , n351954 );
xor ( n351956 , n31898 , n351955 );
xnor ( n351957 , n351911 , n351956 );
buf ( n351958 , n351957 );
xor ( n31926 , n351892 , n351958 );
buf ( n351960 , n31926 );
not ( n31928 , n351661 );
not ( n31929 , n31687 );
or ( n351963 , n31928 , n31929 );
nand ( n31931 , n351963 , n351650 );
buf ( n351965 , n31931 );
nand ( n31933 , n351723 , n351662 );
buf ( n351967 , n31933 );
and ( n351968 , n351965 , n351967 );
buf ( n351969 , n351968 );
xor ( n31937 , n351960 , n351969 );
not ( n351971 , n351714 );
not ( n351972 , n351674 );
or ( n31940 , n351971 , n351972 );
nand ( n351974 , n31940 , n351688 );
buf ( n31942 , n351974 );
nand ( n351976 , n351675 , n351711 );
buf ( n351977 , n351976 );
nand ( n351978 , n31942 , n351977 );
buf ( n351979 , n351978 );
buf ( n351980 , n351979 );
not ( n351981 , n351980 );
buf ( n351982 , n351981 );
buf ( n351983 , n351982 );
not ( n351984 , n351983 );
buf ( n351985 , n351560 );
not ( n31953 , n351985 );
buf ( n351987 , n31543 );
not ( n351988 , n351987 );
or ( n31956 , n31953 , n351988 );
buf ( n351990 , n351560 );
buf ( n351991 , n31543 );
or ( n351992 , n351990 , n351991 );
buf ( n351993 , n31561 );
nand ( n351994 , n351992 , n351993 );
buf ( n351995 , n351994 );
buf ( n351996 , n351995 );
nand ( n351997 , n31956 , n351996 );
buf ( n351998 , n351997 );
buf ( n351999 , n351998 );
buf ( n352000 , n343531 );
not ( n31968 , n352000 );
not ( n352002 , n602 );
not ( n352003 , n24392 );
or ( n31971 , n352002 , n352003 );
or ( n352005 , n24392 , n602 );
nand ( n352006 , n31971 , n352005 );
buf ( n352007 , n352006 );
not ( n352008 , n352007 );
or ( n352009 , n31968 , n352008 );
buf ( n352010 , n351704 );
buf ( n352011 , n343595 );
nand ( n352012 , n352010 , n352011 );
buf ( n352013 , n352012 );
buf ( n352014 , n352013 );
nand ( n352015 , n352009 , n352014 );
buf ( n352016 , n352015 );
buf ( n352017 , n352016 );
xor ( n31985 , n351999 , n352017 );
buf ( n352019 , n344454 );
not ( n352020 , n352019 );
buf ( n352021 , n351440 );
not ( n31989 , n352021 );
or ( n31990 , n352020 , n31989 );
not ( n31991 , n14349 );
nand ( n352025 , n15289 , n14329 );
not ( n352026 , n352025 );
nand ( n31994 , n31991 , n14199 , n352026 );
not ( n31995 , n334248 );
nand ( n31996 , n31995 , n334633 , n14720 );
nor ( n352030 , n31994 , n31996 );
not ( n352031 , n342097 );
or ( n31999 , n352030 , n352031 );
not ( n32000 , n31994 );
not ( n352034 , n31996 );
nand ( n32002 , n32000 , n352031 , n352034 );
nand ( n352036 , n31999 , n32002 );
and ( n32004 , n352036 , n344445 );
not ( n32005 , n352036 );
and ( n352039 , n32005 , n606 );
or ( n352040 , n32004 , n352039 );
buf ( n352041 , n352040 );
buf ( n352042 , n607 );
nand ( n352043 , n352041 , n352042 );
buf ( n352044 , n352043 );
buf ( n352045 , n352044 );
nand ( n32013 , n31990 , n352045 );
buf ( n352047 , n32013 );
not ( n32015 , n352047 );
buf ( n352049 , n32015 );
xor ( n32017 , n31985 , n352049 );
buf ( n352051 , n32017 );
buf ( n352052 , n352051 );
not ( n32020 , n352052 );
buf ( n352054 , n32020 );
buf ( n352055 , n352054 );
not ( n32023 , n352055 );
or ( n352057 , n351984 , n32023 );
buf ( n352058 , n352051 );
buf ( n352059 , n351979 );
nand ( n352060 , n352058 , n352059 );
buf ( n352061 , n352060 );
buf ( n352062 , n352061 );
nand ( n32030 , n352057 , n352062 );
buf ( n352064 , n32030 );
buf ( n352065 , n352064 );
not ( n32033 , n351528 );
buf ( n352067 , n351536 );
buf ( n352068 , n351607 );
nand ( n352069 , n352067 , n352068 );
buf ( n352070 , n352069 );
not ( n32038 , n352070 );
or ( n352072 , n32033 , n32038 );
buf ( n352073 , n31579 );
buf ( n32041 , n31502 );
nand ( n32042 , n352073 , n32041 );
buf ( n32043 , n32042 );
nand ( n352077 , n352072 , n32043 );
buf ( n352078 , n352077 );
not ( n32046 , n352078 );
buf ( n352080 , n32046 );
buf ( n352081 , n352080 );
and ( n352082 , n352065 , n352081 );
not ( n352083 , n352065 );
buf ( n352084 , n352077 );
and ( n352085 , n352083 , n352084 );
nor ( n352086 , n352082 , n352085 );
buf ( n352087 , n352086 );
xor ( n32055 , n31937 , n352087 );
buf ( n352089 , n351617 );
buf ( n352090 , n352089 );
buf ( n352091 , n352090 );
buf ( n352092 , n352091 );
not ( n32060 , n352092 );
buf ( n352094 , n351629 );
not ( n352095 , n352094 );
buf ( n352096 , n352095 );
buf ( n352097 , n352096 );
nand ( n32065 , n32060 , n352097 );
buf ( n352099 , n32065 );
and ( n352100 , n352099 , n351724 );
buf ( n352101 , n352091 );
not ( n32069 , n352101 );
buf ( n352103 , n352096 );
nor ( n352104 , n32069 , n352103 );
buf ( n352105 , n352104 );
nor ( n32073 , n352100 , n352105 );
nor ( n32074 , n32055 , n32073 );
not ( n32075 , n32074 );
nand ( n352109 , n32055 , n32073 );
buf ( n352110 , n352109 );
and ( n32078 , n32075 , n352110 );
and ( n32079 , n31757 , n32078 );
not ( n32080 , n31757 );
not ( n352114 , n32078 );
and ( n32082 , n32080 , n352114 );
nor ( n32083 , n32079 , n32082 );
buf ( n32084 , n32083 );
not ( n32085 , n32084 );
buf ( n352119 , n32085 );
not ( n32087 , n352119 );
buf ( n32088 , n32087 );
buf ( n352122 , n32088 );
xor ( n352123 , n351773 , n352122 );
buf ( n352124 , n352123 );
buf ( n352125 , n352124 );
xor ( n352126 , n351387 , n351388 );
xor ( n352127 , n352126 , n351765 );
buf ( n352128 , n352127 );
buf ( n352129 , n352128 );
buf ( n352130 , n350954 );
xor ( n352131 , n352129 , n352130 );
buf ( n32099 , n350949 );
not ( n352133 , n32099 );
buf ( n352134 , n352133 );
buf ( n352135 , n352134 );
buf ( n352136 , n351376 );
not ( n32104 , n352136 );
buf ( n352138 , n32104 );
buf ( n352139 , n352138 );
nand ( n32107 , n352135 , n352139 );
buf ( n352141 , n32107 );
buf ( n32109 , n352141 );
buf ( n352143 , n351111 );
not ( n32111 , n352143 );
buf ( n352145 , n351329 );
not ( n352146 , n352145 );
buf ( n352147 , n352146 );
buf ( n352148 , n352147 );
nand ( n352149 , n32111 , n352148 );
buf ( n352150 , n352149 );
buf ( n352151 , n352150 );
nand ( n352152 , n32109 , n352151 );
buf ( n352153 , n352152 );
buf ( n352154 , n352153 );
buf ( n352155 , n351116 );
buf ( n352156 , n351371 );
nor ( n352157 , n352155 , n352156 );
buf ( n352158 , n352157 );
buf ( n352159 , n352158 );
nor ( n352160 , n352154 , n352159 );
buf ( n352161 , n352160 );
buf ( n352162 , n352161 );
not ( n352163 , n352162 );
buf ( n352164 , n327911 );
buf ( n352165 , n352164 );
buf ( n352166 , n327916 );
xor ( n352167 , n352165 , n352166 );
buf ( n352168 , n350579 );
not ( n32136 , n352168 );
not ( n352170 , n350576 );
not ( n32138 , n347507 );
nand ( n352172 , n31245 , n32138 );
nand ( n352173 , n352170 , n352172 );
buf ( n352174 , n352173 );
not ( n352175 , n352174 );
or ( n352176 , n32136 , n352175 );
buf ( n352177 , n30557 );
buf ( n352178 , n352177 );
buf ( n352179 , n352178 );
buf ( n352180 , n352179 );
nand ( n32148 , n352176 , n352180 );
buf ( n352182 , n32148 );
buf ( n352183 , n350584 );
buf ( n32151 , n352183 );
buf ( n352185 , n32151 );
nand ( n32153 , n351081 , n352185 );
not ( n32154 , n32153 );
and ( n352188 , n352182 , n32154 );
not ( n352189 , n352182 );
and ( n32157 , n352189 , n32153 );
nor ( n352191 , n352188 , n32157 );
buf ( n352192 , n352191 );
not ( n32160 , n352192 );
buf ( n352194 , n32160 );
not ( n352195 , n352194 );
buf ( n352196 , n352195 );
and ( n32164 , n352167 , n352196 );
and ( n352198 , n352165 , n352166 );
or ( n352199 , n32164 , n352198 );
buf ( n352200 , n352199 );
buf ( n352201 , n352200 );
buf ( n352202 , n351324 );
xor ( n352203 , n352201 , n352202 );
buf ( n352204 , n327223 );
buf ( n352205 , n327229 );
xor ( n32173 , n352204 , n352205 );
and ( n32174 , n350579 , n352179 );
xor ( n32175 , n32174 , n352173 );
buf ( n352209 , n32175 );
buf ( n352210 , n352209 );
buf ( n352211 , n352210 );
buf ( n352212 , n352211 );
buf ( n352213 , n352212 );
and ( n352214 , n32173 , n352213 );
and ( n352215 , n352204 , n352205 );
or ( n32183 , n352214 , n352215 );
buf ( n352217 , n32183 );
buf ( n352218 , n352217 );
xor ( n352219 , n352165 , n352166 );
xor ( n32187 , n352219 , n352196 );
buf ( n352221 , n32187 );
buf ( n352222 , n352221 );
xor ( n32190 , n352218 , n352222 );
buf ( n352224 , n351303 );
xor ( n32192 , n352204 , n352205 );
xor ( n352226 , n32192 , n352213 );
buf ( n352227 , n352226 );
buf ( n352228 , n352227 );
xor ( n352229 , n352224 , n352228 );
buf ( n32197 , n325919 );
xor ( n32198 , n326250 , n32197 );
nand ( n32199 , n30506 , n350559 , n350563 );
nand ( n352233 , n31250 , n351276 );
xnor ( n352234 , n32199 , n352233 );
buf ( n32202 , n352234 );
and ( n352236 , n32198 , n32202 );
and ( n32204 , n326250 , n32197 );
or ( n32205 , n352236 , n32204 );
buf ( n32206 , n32205 );
buf ( n32207 , n351298 );
xor ( n32208 , n32206 , n32207 );
buf ( n352242 , n351273 );
xor ( n32210 , n326250 , n32197 );
xor ( n352244 , n32210 , n32202 );
buf ( n352245 , n352244 );
xor ( n32213 , n352242 , n352245 );
buf ( n32214 , n351239 );
buf ( n32215 , n351268 );
xor ( n32216 , n32214 , n32215 );
buf ( n352250 , n351169 );
buf ( n352251 , n351199 );
xor ( n32219 , n352250 , n352251 );
buf ( n352253 , n327464 );
buf ( n352254 , n327508 );
xor ( n32222 , n352253 , n352254 );
not ( n32223 , n350397 );
not ( n32224 , n32223 );
buf ( n352258 , n351153 );
buf ( n352259 , n351145 );
nand ( n32227 , n352258 , n352259 );
buf ( n352261 , n32227 );
not ( n32229 , n352261 );
not ( n352263 , n32229 );
or ( n352264 , n32224 , n352263 );
nand ( n32232 , n352261 , n350397 );
nand ( n352266 , n352264 , n32232 );
not ( n32234 , n352266 );
not ( n352268 , n32234 );
buf ( n352269 , n352268 );
and ( n352270 , n32222 , n352269 );
and ( n352271 , n352253 , n352254 );
or ( n352272 , n352270 , n352271 );
buf ( n352273 , n352272 );
buf ( n352274 , n352273 );
buf ( n352275 , n351164 );
xor ( n352276 , n352274 , n352275 );
xor ( n352277 , n352253 , n352254 );
xor ( n352278 , n352277 , n352269 );
buf ( n352279 , n352278 );
buf ( n352280 , n352279 );
buf ( n352281 , n351135 );
nor ( n352282 , n352280 , n352281 );
buf ( n352283 , n352282 );
buf ( n352284 , n352283 );
or ( n32252 , n351130 , n351354 );
not ( n352286 , n32252 );
buf ( n352287 , n351072 );
buf ( n352288 , n351349 );
xor ( n352289 , n352287 , n352288 );
buf ( n32257 , n324377 );
buf ( n32258 , n324388 );
buf ( n352292 , n32258 );
xor ( n352293 , n32257 , n352292 );
buf ( n352294 , n29949 );
buf ( n32262 , n352294 );
buf ( n352296 , n32262 );
buf ( n352297 , n352296 );
buf ( n352298 , n349994 );
nand ( n352299 , n352297 , n352298 );
buf ( n352300 , n352299 );
buf ( n352301 , n352300 );
buf ( n32269 , n29770 );
buf ( n32270 , n32269 );
buf ( n352304 , n32270 );
buf ( n352305 , n352304 );
not ( n352306 , n352305 );
buf ( n352307 , n352306 );
buf ( n352308 , n352307 );
and ( n352309 , n352301 , n352308 );
not ( n352310 , n352301 );
buf ( n352311 , n352304 );
and ( n32279 , n352310 , n352311 );
nor ( n352313 , n352309 , n32279 );
buf ( n352314 , n352313 );
buf ( n352315 , n352314 );
and ( n32283 , n352293 , n352315 );
and ( n32284 , n32257 , n352292 );
or ( n352318 , n32283 , n32284 );
buf ( n352319 , n352318 );
buf ( n352320 , n352319 );
buf ( n352321 , n351067 );
xor ( n352322 , n352320 , n352321 );
xor ( n352323 , n32257 , n352292 );
xor ( n32291 , n352323 , n352315 );
buf ( n352325 , n32291 );
buf ( n352326 , n352325 );
buf ( n352327 , n351053 );
or ( n352328 , n352326 , n352327 );
buf ( n352329 , n352328 );
buf ( n352330 , n352329 );
not ( n32298 , n352330 );
buf ( n352332 , n322279 );
buf ( n352333 , n334007 );
xor ( n32301 , n352332 , n352333 );
buf ( n352335 , n349391 );
buf ( n32303 , n352335 );
buf ( n352337 , n32303 );
buf ( n352338 , n352337 );
not ( n32306 , n352338 );
buf ( n352340 , n32306 );
not ( n32308 , n352340 );
not ( n352342 , n349605 );
not ( n32310 , n29569 );
or ( n32311 , n352342 , n32310 );
nand ( n32312 , n32311 , n349599 );
not ( n32313 , n32312 );
not ( n32314 , n32313 );
or ( n32315 , n32308 , n32314 );
buf ( n352349 , n352337 );
buf ( n352350 , n32312 );
nand ( n32318 , n352349 , n352350 );
buf ( n352352 , n32318 );
nand ( n352353 , n32315 , n352352 );
buf ( n352354 , n352353 );
xor ( n32322 , n32301 , n352354 );
buf ( n352356 , n32322 );
buf ( n352357 , n352356 );
buf ( n352358 , n322648 );
buf ( n352359 , n14146 );
xor ( n352360 , n352358 , n352359 );
buf ( n352361 , n349388 );
buf ( n352362 , n348809 );
nand ( n352363 , n352361 , n352362 );
buf ( n352364 , n352363 );
buf ( n352365 , n352364 );
buf ( n352366 , n349374 );
buf ( n32334 , n352366 );
buf ( n352368 , n32334 );
buf ( n352369 , n352368 );
or ( n32337 , n352365 , n352369 );
buf ( n352371 , n352368 );
buf ( n352372 , n348809 );
buf ( n352373 , n349388 );
nand ( n352374 , n352372 , n352373 );
buf ( n352375 , n352374 );
buf ( n352376 , n352375 );
nand ( n32344 , n352371 , n352376 );
buf ( n352378 , n32344 );
buf ( n352379 , n352378 );
nand ( n352380 , n32337 , n352379 );
buf ( n352381 , n352380 );
buf ( n352382 , n352381 );
and ( n32350 , n352360 , n352382 );
and ( n32351 , n352358 , n352359 );
or ( n352385 , n32350 , n32351 );
buf ( n352386 , n352385 );
buf ( n352387 , n352386 );
or ( n32355 , n352357 , n352387 );
xor ( n32356 , n352358 , n352359 );
xor ( n32357 , n32356 , n352382 );
buf ( n32358 , n32357 );
buf ( n352392 , n32358 );
buf ( n352393 , n322701 );
buf ( n352394 , n14159 );
xor ( n352395 , n352393 , n352394 );
buf ( n352396 , n349373 );
buf ( n352397 , n348869 );
nand ( n352398 , n352396 , n352397 );
buf ( n352399 , n352398 );
not ( n32367 , n349364 );
and ( n352401 , n352399 , n32367 );
not ( n352402 , n352399 );
and ( n32370 , n352402 , n349364 );
nor ( n352404 , n352401 , n32370 );
buf ( n352405 , n352404 );
and ( n352406 , n352395 , n352405 );
and ( n32374 , n352393 , n352394 );
or ( n32375 , n352406 , n32374 );
buf ( n352409 , n32375 );
buf ( n352410 , n352409 );
or ( n32378 , n352392 , n352410 );
buf ( n352412 , n351036 );
xor ( n352413 , n352393 , n352394 );
xor ( n32381 , n352413 , n352405 );
buf ( n352415 , n32381 );
buf ( n352416 , n352415 );
or ( n32384 , n352412 , n352416 );
buf ( n352418 , n350973 );
buf ( n352419 , n351382 );
buf ( n352420 , n351380 );
buf ( n352421 , n321437 );
xor ( n32389 , n352420 , n352421 );
buf ( n352423 , n1699 );
buf ( n352424 , n321335 );
xor ( n32392 , n352423 , n352424 );
buf ( n352426 , n321458 );
not ( n352427 , n321499 );
not ( n352428 , n352427 );
buf ( n352429 , n352428 );
xor ( n352430 , n352426 , n352429 );
buf ( n352431 , n1738 );
and ( n32399 , n352430 , n352431 );
or ( n352433 , n32399 , C0 );
buf ( n352434 , n352433 );
buf ( n352435 , n352434 );
and ( n32403 , n32392 , n352435 );
and ( n32404 , n352423 , n352424 );
or ( n352438 , n32403 , n32404 );
buf ( n352439 , n352438 );
buf ( n352440 , n352439 );
and ( n32408 , n32389 , n352440 );
and ( n352442 , n352420 , n352421 );
or ( n32410 , n32408 , n352442 );
buf ( n352444 , n32410 );
buf ( n352445 , n352444 );
xor ( n32413 , n352419 , n352445 );
buf ( n352447 , n350968 );
and ( n352448 , n32413 , n352447 );
and ( n352449 , n352419 , n352445 );
or ( n32417 , n352448 , n352449 );
buf ( n352451 , n32417 );
buf ( n352452 , n352451 );
xor ( n32420 , n352418 , n352452 );
buf ( n352454 , n350992 );
and ( n352455 , n32420 , n352454 );
and ( n32423 , n352418 , n352452 );
or ( n352457 , n352455 , n32423 );
buf ( n352458 , n352457 );
buf ( n352459 , n351017 );
not ( n352460 , n352459 );
buf ( n352461 , n352460 );
buf ( n352462 , n352461 );
buf ( n352463 , n350997 );
not ( n32431 , n352463 );
buf ( n352465 , n32431 );
buf ( n352466 , n352465 );
nand ( n352467 , n352462 , n352466 );
buf ( n352468 , n352467 );
and ( n32436 , n352458 , n352468 );
buf ( n352470 , n352461 );
buf ( n352471 , n352465 );
nor ( n352472 , n352470 , n352471 );
buf ( n352473 , n352472 );
nor ( n32441 , n32436 , n352473 );
buf ( n352475 , n32441 );
buf ( n352476 , n351031 );
buf ( n32444 , n351022 );
nor ( n32445 , n352476 , n32444 );
buf ( n352479 , n32445 );
buf ( n352480 , n352479 );
or ( n352481 , n352475 , n352480 );
buf ( n352482 , n351031 );
buf ( n352483 , n351022 );
nand ( n352484 , n352482 , n352483 );
buf ( n352485 , n352484 );
buf ( n352486 , n352485 );
nand ( n352487 , n352481 , n352486 );
buf ( n352488 , n352487 );
buf ( n352489 , n352488 );
nand ( n352490 , n32384 , n352489 );
buf ( n352491 , n352490 );
buf ( n352492 , n352491 );
buf ( n352493 , n351036 );
buf ( n32461 , n352415 );
nand ( n32462 , n352493 , n32461 );
buf ( n352496 , n32462 );
buf ( n352497 , n352496 );
nand ( n352498 , n352492 , n352497 );
buf ( n352499 , n352498 );
buf ( n352500 , n352499 );
nand ( n32468 , n32378 , n352500 );
buf ( n352502 , n32468 );
buf ( n352503 , n352502 );
buf ( n352504 , n32358 );
buf ( n32472 , n352409 );
nand ( n32473 , n352504 , n32472 );
buf ( n352507 , n32473 );
buf ( n352508 , n352507 );
nand ( n352509 , n352503 , n352508 );
buf ( n352510 , n352509 );
buf ( n352511 , n352510 );
nand ( n32479 , n32355 , n352511 );
buf ( n352513 , n32479 );
buf ( n352514 , n352513 );
buf ( n352515 , n352356 );
buf ( n352516 , n352386 );
nand ( n352517 , n352515 , n352516 );
buf ( n352518 , n352517 );
buf ( n352519 , n352518 );
nand ( n352520 , n352514 , n352519 );
buf ( n352521 , n352520 );
buf ( n352522 , n352521 );
not ( n32490 , n352522 );
buf ( n352524 , n32490 );
buf ( n352525 , n352524 );
buf ( n352526 , n351048 );
xor ( n32494 , n352332 , n352333 );
and ( n352528 , n32494 , n352354 );
and ( n352529 , n352332 , n352333 );
or ( n32497 , n352528 , n352529 );
buf ( n352531 , n32497 );
buf ( n352532 , n352531 );
nor ( n352533 , n352526 , n352532 );
buf ( n352534 , n352533 );
buf ( n352535 , n352534 );
or ( n352536 , n352525 , n352535 );
buf ( n352537 , n351048 );
buf ( n352538 , n352531 );
nand ( n352539 , n352537 , n352538 );
buf ( n352540 , n352539 );
buf ( n352541 , n352540 );
nand ( n32509 , n352536 , n352541 );
buf ( n352543 , n32509 );
buf ( n352544 , n352543 );
not ( n32512 , n352544 );
or ( n32513 , n32298 , n32512 );
buf ( n352547 , n352325 );
buf ( n352548 , n351053 );
nand ( n352549 , n352547 , n352548 );
buf ( n352550 , n352549 );
buf ( n352551 , n352550 );
nand ( n32519 , n32513 , n352551 );
buf ( n352553 , n32519 );
buf ( n352554 , n352553 );
and ( n352555 , n352322 , n352554 );
and ( n352556 , n352320 , n352321 );
or ( n32524 , n352555 , n352556 );
buf ( n352558 , n32524 );
buf ( n32526 , n352558 );
and ( n32527 , n352289 , n32526 );
and ( n32528 , n352287 , n352288 );
or ( n32529 , n32527 , n32528 );
buf ( n32530 , n32529 );
not ( n352564 , n32530 );
or ( n32532 , n352286 , n352564 );
nand ( n32533 , n351130 , n351354 );
nand ( n32534 , n32532 , n32533 );
buf ( n352568 , n32534 );
not ( n352569 , n352568 );
buf ( n352570 , n352569 );
buf ( n352571 , n352570 );
or ( n32539 , n352284 , n352571 );
buf ( n352573 , n352279 );
buf ( n352574 , n351135 );
nand ( n352575 , n352573 , n352574 );
buf ( n352576 , n352575 );
buf ( n352577 , n352576 );
nand ( n32545 , n32539 , n352577 );
buf ( n352579 , n32545 );
buf ( n352580 , n352579 );
and ( n32548 , n352276 , n352580 );
and ( n32549 , n352274 , n352275 );
or ( n32550 , n32548 , n32549 );
buf ( n352584 , n32550 );
buf ( n352585 , n352584 );
and ( n32553 , n32219 , n352585 );
and ( n32554 , n352250 , n352251 );
or ( n32555 , n32553 , n32554 );
buf ( n352589 , n32555 );
buf ( n352590 , n352589 );
buf ( n32558 , n351204 );
xor ( n32559 , n352590 , n32558 );
buf ( n352593 , n351234 );
and ( n32561 , n32559 , n352593 );
and ( n352595 , n352590 , n32558 );
or ( n352596 , n32561 , n352595 );
buf ( n352597 , n352596 );
buf ( n352598 , n352597 );
and ( n32566 , n32216 , n352598 );
and ( n352600 , n32214 , n32215 );
or ( n352601 , n32566 , n352600 );
buf ( n352602 , n352601 );
buf ( n352603 , n352602 );
and ( n352604 , n32213 , n352603 );
and ( n32572 , n352242 , n352245 );
or ( n352606 , n352604 , n32572 );
buf ( n352607 , n352606 );
buf ( n352608 , n352607 );
and ( n32576 , n32208 , n352608 );
and ( n352610 , n32206 , n32207 );
or ( n352611 , n32576 , n352610 );
buf ( n352612 , n352611 );
buf ( n352613 , n352612 );
and ( n352614 , n352229 , n352613 );
and ( n352615 , n352224 , n352228 );
or ( n32583 , n352614 , n352615 );
buf ( n352617 , n32583 );
buf ( n352618 , n352617 );
and ( n32586 , n32190 , n352618 );
and ( n32587 , n352218 , n352222 );
or ( n352621 , n32586 , n32587 );
buf ( n352622 , n352621 );
buf ( n352623 , n352622 );
and ( n32591 , n352203 , n352623 );
and ( n352625 , n352201 , n352202 );
or ( n352626 , n32591 , n352625 );
buf ( n352627 , n352626 );
buf ( n352628 , n352627 );
not ( n32596 , n352628 );
or ( n32597 , n352163 , n32596 );
buf ( n352631 , n352158 );
buf ( n352632 , n351111 );
buf ( n352633 , n351329 );
nand ( n32601 , n352632 , n352633 );
buf ( n352635 , n32601 );
buf ( n352636 , n352635 );
or ( n352637 , n352631 , n352636 );
buf ( n352638 , n351116 );
buf ( n352639 , n351371 );
nand ( n32607 , n352638 , n352639 );
buf ( n352641 , n32607 );
buf ( n352642 , n352641 );
nand ( n352643 , n352637 , n352642 );
buf ( n352644 , n352643 );
buf ( n352645 , n352644 );
buf ( n352646 , n352141 );
and ( n32614 , n352645 , n352646 );
buf ( n352648 , n352134 );
buf ( n352649 , n352138 );
nor ( n32617 , n352648 , n352649 );
buf ( n352651 , n32617 );
buf ( n352652 , n352651 );
nor ( n352653 , n32614 , n352652 );
buf ( n352654 , n352653 );
buf ( n352655 , n352654 );
nand ( n352656 , n32597 , n352655 );
buf ( n352657 , n352656 );
buf ( n352658 , n352657 );
and ( n32626 , n352131 , n352658 );
and ( n32627 , n352129 , n352130 );
or ( n32628 , n32626 , n32627 );
buf ( n352662 , n32628 );
buf ( n352663 , n352662 );
xor ( n352664 , n351770 , n352125 );
xor ( n32632 , n352664 , n352663 );
buf ( n352666 , n32632 );
xor ( n32634 , n351770 , n352125 );
and ( n352668 , n32634 , n352663 );
and ( n352669 , n351770 , n352125 );
or ( n32637 , n352668 , n352669 );
buf ( n352671 , n32637 );
xor ( n32639 , n352129 , n352130 );
xor ( n352673 , n32639 , n352658 );
buf ( n352674 , n352673 );
buf ( n352675 , n352158 );
not ( n352676 , n352675 );
buf ( n352677 , n352676 );
buf ( n352678 , n352677 );
not ( n32646 , n352150 );
not ( n352680 , n352627 );
or ( n352681 , n32646 , n352680 );
nand ( n32649 , n352681 , n352635 );
buf ( n352683 , n32649 );
buf ( n352684 , n352641 );
not ( n352685 , n352678 );
not ( n32653 , n352683 );
or ( n32654 , n352685 , n32653 );
nand ( n32655 , n32654 , n352684 );
buf ( n352689 , n32655 );
xor ( n32657 , n352201 , n352202 );
xor ( n352691 , n32657 , n352623 );
buf ( n352692 , n352691 );
xor ( n32660 , n352218 , n352222 );
xor ( n352694 , n32660 , n352618 );
buf ( n352695 , n352694 );
xor ( n32663 , n352224 , n352228 );
xor ( n32664 , n32663 , n352613 );
buf ( n352698 , n32664 );
xor ( n32666 , n32206 , n32207 );
xor ( n352700 , n32666 , n352608 );
buf ( n352701 , n352700 );
xor ( n32669 , n352242 , n352245 );
xor ( n352703 , n32669 , n352603 );
buf ( n352704 , n352703 );
xor ( n32672 , n32214 , n32215 );
xor ( n32673 , n32672 , n352598 );
buf ( n32674 , n32673 );
xor ( n32675 , n352590 , n32558 );
xor ( n32676 , n32675 , n352593 );
buf ( n352710 , n32676 );
xor ( n32678 , n352250 , n352251 );
xor ( n32679 , n32678 , n352585 );
buf ( n352713 , n32679 );
xor ( n32681 , n352274 , n352275 );
xor ( n32682 , n32681 , n352580 );
buf ( n352716 , n32682 );
buf ( n352717 , n352570 );
buf ( n352718 , n32534 );
buf ( n352719 , n352279 );
buf ( n352720 , n351135 );
xor ( n32688 , n352719 , n352720 );
buf ( n352722 , n32688 );
buf ( n352723 , n352722 );
and ( n352724 , n352723 , n352718 );
not ( n32692 , n352723 );
and ( n32693 , n32692 , n352717 );
nor ( n32694 , n352724 , n32693 );
buf ( n352728 , n32694 );
xor ( n32696 , n352320 , n352321 );
xor ( n32697 , n32696 , n352554 );
buf ( n352731 , n32697 );
buf ( n352732 , n352325 );
buf ( n352733 , n351053 );
xor ( n32701 , n352732 , n352733 );
buf ( n352735 , n32701 );
buf ( n352736 , n352735 );
buf ( n352737 , n352543 );
xor ( n32705 , n352736 , n352737 );
buf ( n352739 , n32705 );
buf ( n352740 , n352524 );
buf ( n352741 , n352521 );
buf ( n352742 , n351048 );
buf ( n352743 , n352531 );
xor ( n32711 , n352742 , n352743 );
buf ( n352745 , n32711 );
buf ( n352746 , n352745 );
and ( n32714 , n352746 , n352741 );
not ( n352748 , n352746 );
and ( n352749 , n352748 , n352740 );
nor ( n32717 , n32714 , n352749 );
buf ( n352751 , n32717 );
buf ( n352752 , n352356 );
buf ( n352753 , n352386 );
xor ( n352754 , n352752 , n352753 );
buf ( n352755 , n352754 );
buf ( n352756 , n352755 );
buf ( n352757 , n352510 );
xor ( n32725 , n352756 , n352757 );
buf ( n352759 , n32725 );
buf ( n352760 , n32358 );
buf ( n352761 , n352409 );
xor ( n352762 , n352760 , n352761 );
buf ( n352763 , n352762 );
buf ( n352764 , n352763 );
buf ( n352765 , n352499 );
xor ( n32733 , n352764 , n352765 );
buf ( n352767 , n32733 );
buf ( n352768 , n352415 );
buf ( n352769 , n351036 );
xor ( n352770 , n352768 , n352769 );
buf ( n352771 , n352770 );
buf ( n352772 , n352771 );
buf ( n352773 , n352488 );
xor ( n32741 , n352772 , n352773 );
buf ( n352775 , n32741 );
buf ( n352776 , n351017 );
buf ( n352777 , n352465 );
xnor ( n32745 , n352776 , n352777 );
buf ( n32746 , n32745 );
buf ( n32747 , n32746 );
buf ( n352781 , n352458 );
xor ( n352782 , n32747 , n352781 );
buf ( n352783 , n352782 );
xor ( n352784 , n352418 , n352452 );
xor ( n352785 , n352784 , n352454 );
buf ( n352786 , n352785 );
xor ( n32754 , n352419 , n352445 );
xor ( n352788 , n32754 , n352447 );
buf ( n352789 , n352788 );
xor ( n32757 , n352420 , n352421 );
xor ( n352791 , n32757 , n352440 );
buf ( n352792 , n352791 );
xor ( n32760 , n352423 , n352424 );
xor ( n352794 , n32760 , n352435 );
buf ( n352795 , n352794 );
xor ( n32763 , n352426 , n352429 );
xor ( n352797 , n32763 , n352431 );
buf ( n352798 , n352797 );
buf ( n352799 , n352138 );
buf ( n352800 , n351376 );
buf ( n352801 , n350949 );
and ( n32769 , n352801 , n352800 );
not ( n32770 , n352801 );
and ( n352804 , n32770 , n352799 );
nor ( n32772 , n32769 , n352804 );
buf ( n32773 , n32772 );
buf ( n32774 , n352147 );
buf ( n352808 , n351329 );
buf ( n352809 , n351111 );
and ( n32777 , n352809 , n352808 );
not ( n352811 , n352809 );
and ( n32779 , n352811 , n32774 );
nor ( n352813 , n32777 , n32779 );
buf ( n352814 , n352813 );
buf ( n352815 , n352689 );
buf ( n352816 , n32773 );
xor ( n32784 , n352815 , n352816 );
buf ( n352818 , n32784 );
buf ( n32786 , n352627 );
buf ( n352820 , n352814 );
xor ( n352821 , n32786 , n352820 );
buf ( n352822 , n352821 );
xor ( n32790 , n351771 , n351772 );
and ( n352824 , n32790 , n352122 );
and ( n32792 , n351771 , n351772 );
or ( n352826 , n352824 , n32792 );
buf ( n352827 , n352826 );
buf ( n352828 , n352827 );
buf ( n352829 , n351386 );
xor ( n352830 , n352828 , n352829 );
buf ( n352831 , n352830 );
buf ( n352832 , n576 );
buf ( n352833 , n24388 );
and ( n32801 , n352832 , n352833 );
buf ( n352835 , n32801 );
buf ( n352836 , n336167 );
not ( n352837 , n352836 );
buf ( n352838 , n576 );
nand ( n352839 , n352837 , n352838 );
buf ( n352840 , n352839 );
buf ( n352841 , n352840 );
not ( n352842 , n352841 );
buf ( n352843 , n352842 );
xor ( n32811 , n352835 , n352843 );
buf ( n32812 , n334643 );
not ( n352846 , n32812 );
buf ( n352847 , n352846 );
buf ( n352848 , n352847 );
not ( n352849 , n352848 );
buf ( n352850 , n335406 );
not ( n352851 , n352850 );
or ( n352852 , n352849 , n352851 );
buf ( n352853 , n580 );
not ( n352854 , n352853 );
buf ( n32822 , n14099 );
not ( n352856 , n32822 );
buf ( n352857 , n352856 );
buf ( n352858 , n352857 );
not ( n32826 , n352858 );
or ( n352860 , n352854 , n32826 );
buf ( n352861 , n352857 );
not ( n32829 , n352861 );
buf ( n32830 , n32829 );
buf ( n352864 , n32830 );
buf ( n352865 , n334650 );
nand ( n32833 , n352864 , n352865 );
buf ( n352867 , n32833 );
buf ( n352868 , n352867 );
nand ( n32836 , n352860 , n352868 );
buf ( n352870 , n32836 );
buf ( n352871 , n352870 );
nand ( n352872 , n352852 , n352871 );
buf ( n352873 , n352872 );
xor ( n32841 , n32811 , n352873 );
buf ( n352875 , n14822 );
not ( n352876 , n352875 );
buf ( n352877 , n580 );
not ( n352878 , n352877 );
buf ( n32846 , n342097 );
not ( n32847 , n32846 );
buf ( n352881 , n32847 );
not ( n32849 , n352881 );
or ( n32850 , n352878 , n32849 );
buf ( n352884 , n32846 );
buf ( n352885 , n334650 );
nand ( n32853 , n352884 , n352885 );
buf ( n352887 , n32853 );
buf ( n352888 , n352887 );
nand ( n32856 , n32850 , n352888 );
buf ( n352890 , n32856 );
buf ( n352891 , n352890 );
not ( n352892 , n352891 );
or ( n32860 , n352876 , n352892 );
buf ( n352894 , n352870 );
buf ( n352895 , n334643 );
nand ( n352896 , n352894 , n352895 );
buf ( n352897 , n352896 );
buf ( n352898 , n352897 );
nand ( n352899 , n32860 , n352898 );
buf ( n352900 , n352899 );
buf ( n352901 , n352900 );
not ( n352902 , n352901 );
buf ( n352903 , n337902 );
buf ( n352904 , n576 );
nand ( n352905 , n352903 , n352904 );
buf ( n352906 , n352905 );
buf ( n352907 , n352906 );
buf ( n352908 , n337085 );
buf ( n352909 , n576 );
nand ( n352910 , n352908 , n352909 );
buf ( n352911 , n352910 );
buf ( n352912 , n352911 );
nand ( n352913 , n352907 , n352912 );
buf ( n352914 , n352913 );
buf ( n352915 , n352914 );
not ( n352916 , n352915 );
buf ( n32884 , n14891 );
not ( n32885 , n32884 );
xor ( n352919 , n352832 , n352833 );
buf ( n352920 , n352919 );
buf ( n352921 , n352920 );
not ( n352922 , n352921 );
or ( n32890 , n32885 , n352922 );
buf ( n352924 , n576 );
not ( n32892 , n352924 );
buf ( n352926 , n336167 );
not ( n352927 , n352926 );
or ( n352928 , n32892 , n352927 );
buf ( n352929 , n15217 );
buf ( n352930 , n332672 );
nand ( n352931 , n352929 , n352930 );
buf ( n352932 , n352931 );
buf ( n352933 , n352932 );
nand ( n352934 , n352928 , n352933 );
buf ( n352935 , n352934 );
buf ( n352936 , n352935 );
buf ( n352937 , n334786 );
nand ( n352938 , n352936 , n352937 );
buf ( n352939 , n352938 );
buf ( n352940 , n352939 );
nand ( n352941 , n32890 , n352940 );
buf ( n352942 , n352941 );
buf ( n352943 , n352942 );
not ( n352944 , n352943 );
or ( n32912 , n352916 , n352944 );
buf ( n352946 , n352911 );
not ( n352947 , n352946 );
buf ( n352948 , n352906 );
not ( n352949 , n352948 );
buf ( n352950 , n352949 );
buf ( n352951 , n352950 );
nand ( n32919 , n352947 , n352951 );
buf ( n352953 , n32919 );
buf ( n352954 , n352953 );
nand ( n32922 , n32912 , n352954 );
buf ( n352956 , n32922 );
not ( n352957 , n352956 );
buf ( n352958 , n352957 );
nand ( n352959 , n352902 , n352958 );
buf ( n352960 , n352959 );
buf ( n352961 , n352960 );
not ( n352962 , n352961 );
buf ( n32930 , n334694 );
not ( n32931 , n32930 );
buf ( n32932 , n32931 );
not ( n32933 , n32932 );
not ( n352967 , n336910 );
or ( n352968 , n32933 , n352967 );
buf ( n352969 , n352857 );
buf ( n352970 , n334702 );
xnor ( n32938 , n352969 , n352970 );
buf ( n352972 , n32938 );
buf ( n352973 , n352972 );
not ( n32941 , n352973 );
buf ( n352975 , n32941 );
nand ( n32943 , n352968 , n352975 );
not ( n32944 , n32943 );
not ( n32945 , n334850 );
buf ( n352979 , n578 );
not ( n32947 , n352979 );
buf ( n352981 , n22150 );
not ( n32949 , n352981 );
or ( n32950 , n32947 , n32949 );
not ( n32951 , n15975 );
buf ( n352985 , n32951 );
buf ( n352986 , n334748 );
nand ( n32954 , n352985 , n352986 );
buf ( n352988 , n32954 );
buf ( n352989 , n352988 );
nand ( n32957 , n32950 , n352989 );
buf ( n352991 , n32957 );
not ( n32959 , n352991 );
or ( n32960 , n32945 , n32959 );
buf ( n352994 , n578 );
not ( n32962 , n352994 );
buf ( n352996 , n335808 );
not ( n352997 , n352996 );
or ( n32965 , n32962 , n352997 );
buf ( n352999 , n15290 );
buf ( n353000 , n334748 );
nand ( n32968 , n352999 , n353000 );
buf ( n32969 , n32968 );
buf ( n353003 , n32969 );
nand ( n32971 , n32965 , n353003 );
buf ( n32972 , n32971 );
buf ( n353006 , n32972 );
buf ( n353007 , n14949 );
buf ( n353008 , n353007 );
buf ( n353009 , n353008 );
buf ( n353010 , n353009 );
nand ( n353011 , n353006 , n353010 );
buf ( n353012 , n353011 );
nand ( n32980 , n32960 , n353012 );
not ( n353014 , n32980 );
or ( n353015 , n32944 , n353014 );
not ( n32983 , n334727 );
not ( n353017 , n334694 );
and ( n32985 , n32983 , n353017 );
nor ( n32986 , n32985 , n352972 );
not ( n353020 , n32986 );
not ( n32988 , n32980 );
not ( n353022 , n32988 );
or ( n353023 , n353020 , n353022 );
not ( n32991 , n334643 );
not ( n353025 , n352890 );
or ( n353026 , n32991 , n353025 );
buf ( n353027 , n580 );
not ( n353028 , n353027 );
buf ( n353029 , n335851 );
not ( n353030 , n353029 );
buf ( n353031 , n353030 );
buf ( n353032 , n353031 );
not ( n353033 , n353032 );
buf ( n353034 , n353033 );
buf ( n353035 , n353034 );
not ( n33003 , n353035 );
buf ( n353037 , n33003 );
buf ( n353038 , n353037 );
not ( n33006 , n353038 );
or ( n353040 , n353028 , n33006 );
buf ( n353041 , n353034 );
buf ( n353042 , n334650 );
nand ( n353043 , n353041 , n353042 );
buf ( n353044 , n353043 );
buf ( n353045 , n353044 );
nand ( n353046 , n353040 , n353045 );
buf ( n353047 , n353046 );
buf ( n353048 , n353047 );
buf ( n353049 , n14822 );
nand ( n33017 , n353048 , n353049 );
buf ( n353051 , n33017 );
nand ( n33019 , n353026 , n353051 );
nand ( n353053 , n353023 , n33019 );
nand ( n353054 , n353015 , n353053 );
buf ( n353055 , n353054 );
not ( n353056 , n353055 );
or ( n33024 , n352962 , n353056 );
buf ( n353058 , n352956 );
buf ( n33026 , n352900 );
buf ( n353060 , n33026 );
nand ( n353061 , n353058 , n353060 );
buf ( n353062 , n353061 );
buf ( n353063 , n353062 );
nand ( n353064 , n33024 , n353063 );
buf ( n353065 , n353064 );
xor ( n353066 , n32841 , n353065 );
buf ( n353067 , n352840 );
buf ( n353068 , n14891 );
not ( n33036 , n353068 );
buf ( n353070 , n576 );
not ( n33038 , n353070 );
buf ( n353072 , n335808 );
not ( n353073 , n353072 );
or ( n33041 , n33038 , n353073 );
buf ( n33042 , n335808 );
not ( n353076 , n33042 );
buf ( n353077 , n353076 );
buf ( n353078 , n353077 );
buf ( n353079 , n332672 );
nand ( n33047 , n353078 , n353079 );
buf ( n33048 , n33047 );
buf ( n33049 , n33048 );
nand ( n33050 , n33041 , n33049 );
buf ( n33051 , n33050 );
buf ( n353085 , n33051 );
not ( n353086 , n353085 );
or ( n353087 , n33036 , n353086 );
buf ( n353088 , n352920 );
buf ( n353089 , n334786 );
nand ( n33057 , n353088 , n353089 );
buf ( n33058 , n33057 );
buf ( n353092 , n33058 );
nand ( n33060 , n353087 , n353092 );
buf ( n33061 , n33060 );
buf ( n33062 , n33061 );
xor ( n33063 , n353067 , n33062 );
buf ( n353097 , n353009 );
not ( n353098 , n353097 );
buf ( n353099 , n352991 );
not ( n353100 , n353099 );
or ( n33068 , n353098 , n353100 );
buf ( n353102 , n578 );
not ( n353103 , n353102 );
buf ( n353104 , n353037 );
not ( n33072 , n353104 );
or ( n353106 , n353103 , n33072 );
buf ( n353107 , n353037 );
not ( n33075 , n353107 );
buf ( n353109 , n33075 );
buf ( n353110 , n353109 );
buf ( n353111 , n334748 );
nand ( n33079 , n353110 , n353111 );
buf ( n33080 , n33079 );
buf ( n353114 , n33080 );
nand ( n33082 , n353106 , n353114 );
buf ( n33083 , n33082 );
buf ( n353117 , n33083 );
buf ( n353118 , n334850 );
nand ( n353119 , n353117 , n353118 );
buf ( n353120 , n353119 );
buf ( n353121 , n353120 );
nand ( n33089 , n33068 , n353121 );
buf ( n353123 , n33089 );
buf ( n353124 , n353123 );
and ( n353125 , n33063 , n353124 );
and ( n353126 , n353067 , n33062 );
or ( n33094 , n353125 , n353126 );
buf ( n353128 , n33094 );
buf ( n353129 , n578 );
not ( n353130 , n353129 );
buf ( n353131 , n32847 );
not ( n353132 , n353131 );
or ( n353133 , n353130 , n353132 );
buf ( n353134 , n32846 );
buf ( n353135 , n334748 );
nand ( n353136 , n353134 , n353135 );
buf ( n353137 , n353136 );
buf ( n353138 , n353137 );
nand ( n353139 , n353133 , n353138 );
buf ( n353140 , n353139 );
and ( n353141 , n353140 , n334850 );
not ( n33109 , n33083 );
buf ( n353143 , n353009 );
not ( n353144 , n353143 );
buf ( n353145 , n353144 );
nor ( n353146 , n33109 , n353145 );
nor ( n353147 , n353141 , n353146 );
not ( n33115 , n33051 );
not ( n33116 , n334786 );
or ( n353150 , n33115 , n33116 );
buf ( n353151 , n576 );
not ( n33119 , n353151 );
buf ( n353153 , n15975 );
not ( n353154 , n353153 );
or ( n33122 , n33119 , n353154 );
buf ( n353156 , n32951 );
buf ( n353157 , n332672 );
nand ( n353158 , n353156 , n353157 );
buf ( n353159 , n353158 );
buf ( n353160 , n353159 );
nand ( n353161 , n33122 , n353160 );
buf ( n353162 , n353161 );
nand ( n353163 , n353162 , n14891 );
nand ( n353164 , n353150 , n353163 );
not ( n353165 , n353164 );
and ( n33133 , n353147 , n353165 );
not ( n353167 , n353147 );
and ( n33135 , n353167 , n353164 );
nor ( n353169 , n33133 , n33135 );
xor ( n33137 , n353128 , n353169 );
xor ( n33138 , n353066 , n33137 );
not ( n353172 , n33138 );
xor ( n353173 , n353067 , n33062 );
xor ( n33141 , n353173 , n353124 );
buf ( n353175 , n33141 );
and ( n353176 , n352911 , n352950 );
not ( n33144 , n352911 );
and ( n353178 , n33144 , n352906 );
or ( n353179 , n353176 , n353178 );
and ( n33147 , n353179 , n352942 );
not ( n33148 , n353179 );
not ( n353182 , n352942 );
and ( n33150 , n33148 , n353182 );
nor ( n353184 , n33147 , n33150 );
buf ( n353185 , n353184 );
buf ( n353186 , n352911 );
buf ( n353187 , n334786 );
not ( n33155 , n353187 );
and ( n33156 , n335121 , n332672 );
not ( n353190 , n335121 );
and ( n353191 , n353190 , n576 );
or ( n33159 , n33156 , n353191 );
buf ( n353193 , n33159 );
not ( n353194 , n353193 );
or ( n33162 , n33155 , n353194 );
buf ( n353196 , n352935 );
buf ( n353197 , n14891 );
nand ( n353198 , n353196 , n353197 );
buf ( n353199 , n353198 );
buf ( n353200 , n353199 );
nand ( n353201 , n33162 , n353200 );
buf ( n353202 , n353201 );
buf ( n353203 , n353202 );
xor ( n353204 , n353186 , n353203 );
buf ( n353205 , n334850 );
not ( n353206 , n353205 );
buf ( n353207 , n32972 );
not ( n353208 , n353207 );
or ( n353209 , n353206 , n353208 );
buf ( n353210 , n578 );
not ( n353211 , n353210 );
buf ( n353212 , n24387 );
not ( n33180 , n353212 );
or ( n353214 , n353211 , n33180 );
buf ( n353215 , n15300 );
buf ( n353216 , n334748 );
nand ( n33184 , n353215 , n353216 );
buf ( n33185 , n33184 );
buf ( n353219 , n33185 );
nand ( n33187 , n353214 , n353219 );
buf ( n353221 , n33187 );
buf ( n33189 , n353221 );
buf ( n33190 , n353009 );
nand ( n33191 , n33189 , n33190 );
buf ( n33192 , n33191 );
buf ( n33193 , n33192 );
nand ( n33194 , n353209 , n33193 );
buf ( n33195 , n33194 );
buf ( n353229 , n33195 );
and ( n353230 , n353204 , n353229 );
and ( n33198 , n353186 , n353203 );
or ( n353232 , n353230 , n33198 );
buf ( n353233 , n353232 );
buf ( n353234 , n353233 );
xor ( n353235 , n353185 , n353234 );
buf ( n353236 , n17240 );
buf ( n353237 , n576 );
nand ( n353238 , n353236 , n353237 );
buf ( n353239 , n353238 );
buf ( n353240 , n353239 );
buf ( n353241 , n336886 );
not ( n353242 , n353241 );
buf ( n33210 , n576 );
nand ( n33211 , n353242 , n33210 );
buf ( n353245 , n33211 );
buf ( n353246 , n353245 );
nand ( n33214 , n353240 , n353246 );
buf ( n353248 , n33214 );
buf ( n353249 , n353248 );
not ( n33217 , n353249 );
buf ( n353251 , n335432 );
not ( n33219 , n353251 );
buf ( n353253 , n353221 );
not ( n353254 , n353253 );
or ( n353255 , n33219 , n353254 );
buf ( n353256 , n578 );
not ( n353257 , n353256 );
buf ( n353258 , n336167 );
not ( n33226 , n353258 );
or ( n353260 , n353257 , n33226 );
buf ( n353261 , n15217 );
buf ( n353262 , n334748 );
nand ( n353263 , n353261 , n353262 );
buf ( n353264 , n353263 );
buf ( n353265 , n353264 );
nand ( n33233 , n353260 , n353265 );
buf ( n353267 , n33233 );
buf ( n33235 , n353267 );
buf ( n353269 , n353009 );
nand ( n353270 , n33235 , n353269 );
buf ( n353271 , n353270 );
buf ( n353272 , n353271 );
nand ( n33240 , n353255 , n353272 );
buf ( n33241 , n33240 );
buf ( n353275 , n33241 );
not ( n33243 , n353275 );
or ( n353277 , n33217 , n33243 );
buf ( n353278 , n353239 );
not ( n33246 , n353278 );
buf ( n33247 , n353245 );
not ( n353281 , n33247 );
buf ( n353282 , n353281 );
buf ( n353283 , n353282 );
nand ( n33251 , n33246 , n353283 );
buf ( n353285 , n33251 );
buf ( n353286 , n353285 );
nand ( n353287 , n353277 , n353286 );
buf ( n353288 , n353287 );
not ( n33256 , n353288 );
buf ( n353290 , n580 );
not ( n353291 , n353290 );
buf ( n353292 , n15975 );
not ( n33260 , n353292 );
or ( n353294 , n353291 , n33260 );
not ( n353295 , n22150 );
nand ( n33263 , n353295 , n334650 );
buf ( n353297 , n33263 );
nand ( n353298 , n353294 , n353297 );
buf ( n353299 , n353298 );
buf ( n353300 , n353299 );
not ( n33268 , n353300 );
buf ( n353302 , n33268 );
not ( n33270 , n353302 );
not ( n353304 , n335406 );
and ( n353305 , n33270 , n353304 );
and ( n33273 , n353047 , n334643 );
nor ( n353307 , n353305 , n33273 );
buf ( n353308 , n352972 );
not ( n33276 , n353308 );
buf ( n353310 , n32932 );
not ( n33278 , n353310 );
and ( n353312 , n33276 , n33278 );
buf ( n353313 , n582 );
not ( n33281 , n353313 );
buf ( n353315 , n352031 );
not ( n353316 , n353315 );
or ( n33284 , n33281 , n353316 );
buf ( n353318 , n342097 );
buf ( n353319 , n334702 );
nand ( n33287 , n353318 , n353319 );
buf ( n353321 , n33287 );
buf ( n353322 , n353321 );
nand ( n33290 , n33284 , n353322 );
buf ( n353324 , n33290 );
buf ( n353325 , n353324 );
buf ( n353326 , n334727 );
and ( n33294 , n353325 , n353326 );
nor ( n353328 , n353312 , n33294 );
buf ( n353329 , n353328 );
nand ( n353330 , n353307 , n353329 );
not ( n33298 , n353330 );
or ( n353332 , n33256 , n33298 );
not ( n353333 , n353329 );
buf ( n353334 , n334643 );
not ( n33302 , n353334 );
buf ( n353336 , n353047 );
not ( n33304 , n353336 );
or ( n353338 , n33302 , n33304 );
buf ( n353339 , n353302 );
not ( n353340 , n353339 );
buf ( n353341 , n14822 );
nand ( n353342 , n353340 , n353341 );
buf ( n353343 , n353342 );
buf ( n353344 , n353343 );
nand ( n353345 , n353338 , n353344 );
buf ( n353346 , n353345 );
nand ( n33314 , n353333 , n353346 );
nand ( n33315 , n353332 , n33314 );
buf ( n353349 , n33315 );
and ( n33317 , n353235 , n353349 );
and ( n33318 , n353185 , n353234 );
or ( n353352 , n33317 , n33318 );
buf ( n353353 , n353352 );
xor ( n33321 , n353175 , n353353 );
xnor ( n353355 , n352900 , n352957 );
buf ( n353356 , n353355 );
buf ( n353357 , n353054 );
xor ( n353358 , n353356 , n353357 );
buf ( n353359 , n353358 );
and ( n33327 , n33321 , n353359 );
and ( n353361 , n353175 , n353353 );
or ( n353362 , n33327 , n353361 );
not ( n353363 , n353362 );
nand ( n33331 , n353172 , n353363 );
nand ( n353365 , n33138 , n353362 );
nand ( n353366 , n33331 , n353365 );
not ( n33334 , n353366 );
buf ( n353368 , n337183 );
buf ( n353369 , n576 );
and ( n33337 , n353368 , n353369 );
buf ( n353371 , n33337 );
not ( n33339 , n353371 );
buf ( n353373 , n334786 );
not ( n33341 , n353373 );
and ( n33342 , n337163 , n332672 );
not ( n353376 , n337163 );
and ( n353377 , n353376 , n576 );
or ( n33345 , n33342 , n353377 );
buf ( n353379 , n33345 );
not ( n33347 , n353379 );
or ( n353381 , n33341 , n33347 );
buf ( n353382 , n14890 );
not ( n353383 , n353382 );
buf ( n353384 , n576 );
not ( n33352 , n353384 );
buf ( n353386 , n334890 );
not ( n353387 , n353386 );
or ( n353388 , n33352 , n353387 );
buf ( n353389 , n334896 );
buf ( n353390 , n332672 );
nand ( n33358 , n353389 , n353390 );
buf ( n353392 , n33358 );
buf ( n353393 , n353392 );
nand ( n33361 , n353388 , n353393 );
buf ( n353395 , n33361 );
buf ( n353396 , n353395 );
nand ( n33364 , n353383 , n353396 );
buf ( n353398 , n33364 );
buf ( n353399 , n353398 );
nand ( n33367 , n353381 , n353399 );
buf ( n33368 , n33367 );
not ( n353402 , n33368 );
not ( n33370 , n353402 );
or ( n353404 , n33339 , n33370 );
buf ( n33372 , n353371 );
not ( n353406 , n33372 );
buf ( n353407 , n353406 );
nand ( n353408 , n33368 , n353407 );
nand ( n353409 , n353404 , n353408 );
not ( n33377 , n353409 );
not ( n353411 , n33377 );
buf ( n353412 , n335432 );
not ( n33380 , n353412 );
buf ( n33381 , n578 );
not ( n33382 , n33381 );
buf ( n33383 , n337088 );
not ( n33384 , n33383 );
or ( n33385 , n33382 , n33384 );
buf ( n353419 , n337085 );
buf ( n353420 , n334748 );
nand ( n353421 , n353419 , n353420 );
buf ( n353422 , n353421 );
buf ( n353423 , n353422 );
nand ( n353424 , n33385 , n353423 );
buf ( n353425 , n353424 );
buf ( n353426 , n353425 );
not ( n353427 , n353426 );
or ( n353428 , n33380 , n353427 );
buf ( n353429 , n578 );
not ( n353430 , n353429 );
buf ( n353431 , n17937 );
not ( n33399 , n353431 );
or ( n353433 , n353430 , n33399 );
buf ( n33401 , n15012 );
buf ( n33402 , n334748 );
nand ( n33403 , n33401 , n33402 );
buf ( n33404 , n33403 );
buf ( n33405 , n33404 );
nand ( n33406 , n353433 , n33405 );
buf ( n33407 , n33406 );
buf ( n353441 , n33407 );
buf ( n353442 , n353009 );
nand ( n33410 , n353441 , n353442 );
buf ( n353444 , n33410 );
buf ( n353445 , n353444 );
nand ( n353446 , n353428 , n353445 );
buf ( n353447 , n353446 );
not ( n353448 , n353447 );
not ( n353449 , n353448 );
or ( n353450 , n353411 , n353449 );
nand ( n33418 , n353409 , n353447 );
nand ( n353452 , n353450 , n33418 );
not ( n33420 , n353009 );
not ( n33421 , n578 );
not ( n353455 , n336868 );
or ( n33423 , n33421 , n353455 );
buf ( n353457 , n336865 );
buf ( n353458 , n334748 );
nand ( n33426 , n353457 , n353458 );
buf ( n353460 , n33426 );
nand ( n353461 , n33423 , n353460 );
not ( n33429 , n353461 );
or ( n353463 , n33420 , n33429 );
buf ( n353464 , n578 );
not ( n33432 , n353464 );
buf ( n353466 , n14837 );
not ( n353467 , n353466 );
or ( n353468 , n33432 , n353467 );
buf ( n353469 , n334896 );
buf ( n353470 , n334748 );
nand ( n353471 , n353469 , n353470 );
buf ( n353472 , n353471 );
buf ( n353473 , n353472 );
nand ( n353474 , n353468 , n353473 );
buf ( n353475 , n353474 );
buf ( n353476 , n353475 );
buf ( n353477 , n335432 );
nand ( n33445 , n353476 , n353477 );
buf ( n353479 , n33445 );
nand ( n353480 , n353463 , n353479 );
not ( n33448 , n353480 );
and ( n353482 , n576 , n334662 );
not ( n353483 , n576 );
and ( n353484 , n353483 , n334561 );
or ( n33452 , n353482 , n353484 );
buf ( n33453 , n33452 );
not ( n33454 , n33453 );
buf ( n33455 , n33454 );
buf ( n353489 , n33455 );
not ( n353490 , n353489 );
buf ( n353491 , n15711 );
not ( n33459 , n353491 );
and ( n353493 , n353490 , n33459 );
buf ( n353494 , n576 );
not ( n33462 , n353494 );
buf ( n353496 , n335237 );
not ( n353497 , n353496 );
or ( n33465 , n33462 , n353497 );
buf ( n353499 , n334647 );
buf ( n353500 , n332672 );
nand ( n33468 , n353499 , n353500 );
buf ( n353502 , n33468 );
buf ( n353503 , n353502 );
nand ( n353504 , n33465 , n353503 );
buf ( n353505 , n353504 );
buf ( n353506 , n353505 );
buf ( n353507 , n14891 );
and ( n353508 , n353506 , n353507 );
nor ( n33476 , n353493 , n353508 );
buf ( n33477 , n33476 );
buf ( n353511 , n33477 );
not ( n33479 , n14891 );
not ( n353513 , n33452 );
or ( n353514 , n33479 , n353513 );
not ( n353515 , n576 );
not ( n33483 , n334837 );
or ( n353517 , n353515 , n33483 );
nand ( n33485 , n14698 , n332672 );
nand ( n353519 , n353517 , n33485 );
nand ( n353520 , n334786 , n353519 );
nand ( n33488 , n353514 , n353520 );
buf ( n353522 , n33488 );
not ( n33490 , n353522 );
buf ( n353524 , n33490 );
buf ( n353525 , n353524 );
nand ( n33493 , n353511 , n353525 );
buf ( n353527 , n33493 );
not ( n353528 , n353527 );
or ( n33496 , n33448 , n353528 );
buf ( n353530 , n33477 );
not ( n353531 , n353530 );
buf ( n353532 , n33488 );
nand ( n353533 , n353531 , n353532 );
buf ( n353534 , n353533 );
nand ( n33502 , n33496 , n353534 );
buf ( n353536 , n33502 );
buf ( n353537 , n15239 );
not ( n353538 , n353537 );
buf ( n353539 , n335111 );
not ( n353540 , n353539 );
or ( n353541 , n353538 , n353540 );
buf ( n353542 , n588 );
not ( n353543 , n353542 );
buf ( n353544 , n352857 );
not ( n33512 , n353544 );
or ( n353546 , n353543 , n33512 );
buf ( n353547 , n14099 );
buf ( n353548 , n334972 );
nand ( n33516 , n353547 , n353548 );
buf ( n353550 , n33516 );
buf ( n353551 , n353550 );
nand ( n33519 , n353546 , n353551 );
buf ( n353553 , n33519 );
buf ( n353554 , n353553 );
nand ( n33522 , n353541 , n353554 );
buf ( n33523 , n33522 );
buf ( n353557 , n33523 );
nor ( n33525 , n353536 , n353557 );
buf ( n33526 , n33525 );
buf ( n353560 , n33526 );
not ( n33528 , n353560 );
buf ( n353562 , n336030 );
buf ( n353563 , n576 );
and ( n353564 , n353562 , n353563 );
buf ( n353565 , n353564 );
buf ( n353566 , n353565 );
buf ( n353567 , n353505 );
not ( n33535 , n353567 );
buf ( n33536 , n33535 );
buf ( n353570 , n33536 );
not ( n33538 , n353570 );
buf ( n353572 , n15711 );
not ( n33540 , n353572 );
and ( n353574 , n33538 , n33540 );
buf ( n353575 , n33345 );
buf ( n353576 , n14891 );
and ( n33544 , n353575 , n353576 );
nor ( n33545 , n353574 , n33544 );
buf ( n353579 , n33545 );
buf ( n353580 , n353579 );
not ( n33548 , n353580 );
buf ( n353582 , n33548 );
buf ( n353583 , n353582 );
xor ( n353584 , n353566 , n353583 );
buf ( n353585 , n335432 );
not ( n33553 , n353585 );
buf ( n353587 , n33407 );
not ( n353588 , n353587 );
or ( n353589 , n33553 , n353588 );
buf ( n353590 , n353475 );
buf ( n353591 , n353009 );
nand ( n353592 , n353590 , n353591 );
buf ( n353593 , n353592 );
buf ( n353594 , n353593 );
nand ( n33562 , n353589 , n353594 );
buf ( n353596 , n33562 );
buf ( n353597 , n353596 );
xor ( n33565 , n353584 , n353597 );
buf ( n353599 , n33565 );
buf ( n353600 , n353599 );
nand ( n353601 , n33528 , n353600 );
buf ( n353602 , n353601 );
buf ( n353603 , n33502 );
buf ( n353604 , n33523 );
nand ( n353605 , n353603 , n353604 );
buf ( n353606 , n353605 );
nand ( n33574 , n353602 , n353606 );
xor ( n353608 , n353452 , n33574 );
not ( n353609 , n14822 );
not ( n353610 , n334650 );
not ( n353611 , n337894 );
or ( n33579 , n353610 , n353611 );
buf ( n353613 , n15264 );
buf ( n33581 , n580 );
nand ( n353615 , n353613 , n33581 );
buf ( n353616 , n353615 );
nand ( n33584 , n33579 , n353616 );
not ( n353618 , n33584 );
or ( n353619 , n353609 , n353618 );
buf ( n353620 , n580 );
not ( n353621 , n353620 );
buf ( n353622 , n336167 );
not ( n33590 , n353622 );
or ( n353624 , n353621 , n33590 );
buf ( n353625 , n15217 );
buf ( n353626 , n334650 );
nand ( n33594 , n353625 , n353626 );
buf ( n353628 , n33594 );
buf ( n353629 , n353628 );
nand ( n33597 , n353624 , n353629 );
buf ( n353631 , n33597 );
nand ( n33599 , n353631 , n15528 );
nand ( n33600 , n353619 , n33599 );
not ( n353634 , n33600 );
buf ( n353635 , n334694 );
not ( n33603 , n353635 );
buf ( n353637 , n582 );
not ( n353638 , n353637 );
buf ( n353639 , n15290 );
not ( n353640 , n353639 );
buf ( n353641 , n353640 );
buf ( n353642 , n353641 );
not ( n33610 , n353642 );
or ( n353644 , n353638 , n33610 );
buf ( n353645 , n15290 );
buf ( n353646 , n334702 );
nand ( n353647 , n353645 , n353646 );
buf ( n353648 , n353647 );
buf ( n353649 , n353648 );
nand ( n33617 , n353644 , n353649 );
buf ( n353651 , n33617 );
buf ( n353652 , n353651 );
not ( n353653 , n353652 );
or ( n33621 , n33603 , n353653 );
buf ( n353655 , n582 );
not ( n33623 , n353655 );
buf ( n353657 , n335163 );
not ( n353658 , n353657 );
or ( n33626 , n33623 , n353658 );
nand ( n353660 , n15300 , n334702 );
buf ( n353661 , n353660 );
nand ( n33629 , n33626 , n353661 );
buf ( n353663 , n33629 );
buf ( n353664 , n353663 );
buf ( n353665 , n334727 );
nand ( n353666 , n353664 , n353665 );
buf ( n353667 , n353666 );
buf ( n353668 , n353667 );
nand ( n33636 , n33621 , n353668 );
buf ( n353670 , n33636 );
buf ( n353671 , n353670 );
not ( n33639 , n353671 );
buf ( n353673 , n33639 );
not ( n33641 , n353673 );
or ( n353675 , n353634 , n33641 );
not ( n353676 , n353670 );
or ( n33644 , n353676 , n33600 );
nand ( n353678 , n353675 , n33644 );
not ( n33646 , n353678 );
buf ( n353680 , n353565 );
not ( n33648 , n353680 );
buf ( n353682 , n353582 );
not ( n33650 , n353682 );
or ( n353684 , n33648 , n33650 );
buf ( n353685 , n353565 );
not ( n33653 , n353685 );
buf ( n33654 , n33653 );
buf ( n353688 , n33654 );
not ( n353689 , n353688 );
buf ( n353690 , n353579 );
not ( n33658 , n353690 );
or ( n353692 , n353689 , n33658 );
buf ( n33660 , n353596 );
nand ( n33661 , n353692 , n33660 );
buf ( n33662 , n33661 );
buf ( n353696 , n33662 );
nand ( n353697 , n353684 , n353696 );
buf ( n353698 , n353697 );
nand ( n33666 , n33646 , n353698 );
not ( n353700 , n353698 );
nand ( n353701 , n353700 , n353678 );
nand ( n33669 , n33666 , n353701 );
xnor ( n353703 , n353608 , n33669 );
buf ( n353704 , n15164 );
not ( n353705 , n353704 );
buf ( n353706 , n586 );
not ( n33674 , n353706 );
buf ( n353708 , n15975 );
not ( n33676 , n353708 );
or ( n353710 , n33674 , n33676 );
buf ( n353711 , n14199 );
buf ( n353712 , n334982 );
nand ( n353713 , n353711 , n353712 );
buf ( n353714 , n353713 );
buf ( n353715 , n353714 );
nand ( n353716 , n353710 , n353715 );
buf ( n353717 , n353716 );
buf ( n353718 , n353717 );
not ( n353719 , n353718 );
or ( n353720 , n353705 , n353719 );
buf ( n353721 , n586 );
not ( n33689 , n353721 );
buf ( n353723 , n15992 );
not ( n353724 , n353723 );
or ( n33692 , n33689 , n353724 );
buf ( n353726 , n335851 );
buf ( n353727 , n334982 );
nand ( n33695 , n353726 , n353727 );
buf ( n353729 , n33695 );
buf ( n353730 , n353729 );
nand ( n353731 , n33692 , n353730 );
buf ( n353732 , n353731 );
buf ( n353733 , n353732 );
buf ( n353734 , n334978 );
nand ( n33702 , n353733 , n353734 );
buf ( n353736 , n33702 );
buf ( n353737 , n353736 );
nand ( n33705 , n353720 , n353737 );
buf ( n353739 , n33705 );
not ( n33707 , n353739 );
not ( n353741 , n335114 );
not ( n33709 , n588 );
not ( n33710 , n342097 );
not ( n353744 , n33710 );
or ( n353745 , n33709 , n353744 );
buf ( n353746 , n342097 );
buf ( n353747 , n334972 );
nand ( n353748 , n353746 , n353747 );
buf ( n353749 , n353748 );
nand ( n353750 , n353745 , n353749 );
not ( n353751 , n353750 );
or ( n353752 , n353741 , n353751 );
buf ( n353753 , n353553 );
buf ( n353754 , n15275 );
nand ( n353755 , n353753 , n353754 );
buf ( n353756 , n353755 );
nand ( n353757 , n353752 , n353756 );
not ( n353758 , n353757 );
or ( n33726 , n33707 , n353758 );
buf ( n353760 , n353739 );
not ( n33728 , n353760 );
buf ( n353762 , n33728 );
not ( n353763 , n353762 );
not ( n353764 , n335114 );
not ( n33732 , n353750 );
or ( n353766 , n353764 , n33732 );
nand ( n33734 , n353766 , n353756 );
not ( n33735 , n33734 );
not ( n33736 , n33735 );
or ( n353770 , n353763 , n33736 );
buf ( n353771 , n582 );
buf ( n353772 , n333978 );
and ( n353773 , n353771 , n353772 );
not ( n33741 , n353771 );
buf ( n353775 , n335003 );
and ( n33743 , n33741 , n353775 );
nor ( n33744 , n353773 , n33743 );
buf ( n353778 , n33744 );
buf ( n353779 , n353778 );
not ( n353780 , n353779 );
buf ( n353781 , n353780 );
not ( n33749 , n353781 );
not ( n353783 , n336910 );
and ( n33751 , n33749 , n353783 );
not ( n33752 , n334702 );
not ( n33753 , n337894 );
or ( n33754 , n33752 , n33753 );
nand ( n353788 , n15264 , n582 );
nand ( n33756 , n33754 , n353788 );
and ( n33757 , n33756 , n334694 );
nor ( n33758 , n33751 , n33757 );
not ( n353792 , n33758 );
not ( n353793 , n353792 );
not ( n33761 , n353524 );
or ( n33762 , n353793 , n33761 );
buf ( n353796 , n33488 );
not ( n353797 , n353796 );
buf ( n353798 , n33758 );
not ( n33766 , n353798 );
or ( n33767 , n353797 , n33766 );
buf ( n353801 , n14897 );
buf ( n353802 , n576 );
nand ( n353803 , n353801 , n353802 );
buf ( n353804 , n353803 );
buf ( n353805 , n353804 );
not ( n353806 , n353805 );
buf ( n353807 , n353806 );
buf ( n353808 , n353807 );
not ( n353809 , n353808 );
not ( n33777 , n15528 );
not ( n33778 , n580 );
not ( n33779 , n14837 );
or ( n33780 , n33778 , n33779 );
buf ( n353814 , n14688 );
buf ( n353815 , n334650 );
nand ( n33783 , n353814 , n353815 );
buf ( n353817 , n33783 );
nand ( n33785 , n33780 , n353817 );
not ( n33786 , n33785 );
or ( n33787 , n33777 , n33786 );
buf ( n353821 , n342151 );
buf ( n353822 , n14822 );
nand ( n33790 , n353821 , n353822 );
buf ( n33791 , n33790 );
nand ( n353825 , n33787 , n33791 );
buf ( n353826 , n353825 );
not ( n353827 , n353826 );
or ( n353828 , n353809 , n353827 );
buf ( n353829 , n353825 );
buf ( n353830 , n353807 );
or ( n33798 , n353829 , n353830 );
buf ( n353832 , n14891 );
not ( n353833 , n353832 );
buf ( n353834 , n353519 );
not ( n353835 , n353834 );
or ( n353836 , n353833 , n353835 );
buf ( n353837 , n342211 );
buf ( n353838 , n334786 );
nand ( n33806 , n353837 , n353838 );
buf ( n353840 , n33806 );
buf ( n353841 , n353840 );
nand ( n33809 , n353836 , n353841 );
buf ( n353843 , n33809 );
buf ( n353844 , n353843 );
nand ( n353845 , n33798 , n353844 );
buf ( n353846 , n353845 );
buf ( n353847 , n353846 );
nand ( n33815 , n353828 , n353847 );
buf ( n353849 , n33815 );
buf ( n353850 , n353849 );
nand ( n353851 , n33767 , n353850 );
buf ( n353852 , n353851 );
nand ( n33820 , n33762 , n353852 );
nand ( n33821 , n353770 , n33820 );
nand ( n353855 , n33726 , n33821 );
not ( n353856 , n353855 );
not ( n33824 , n353856 );
not ( n353858 , n334917 );
and ( n33826 , n15290 , n334879 );
not ( n33827 , n15290 );
and ( n33828 , n33827 , n584 );
or ( n353862 , n33826 , n33828 );
not ( n353863 , n353862 );
or ( n33831 , n353858 , n353863 );
not ( n33832 , n334868 );
not ( n353866 , n33832 );
not ( n353867 , n584 );
not ( n33835 , n15975 );
or ( n33836 , n353867 , n33835 );
buf ( n353870 , n14199 );
buf ( n353871 , n334879 );
nand ( n353872 , n353870 , n353871 );
buf ( n353873 , n353872 );
nand ( n33841 , n33836 , n353873 );
nand ( n353875 , n353866 , n33841 );
nand ( n33843 , n33831 , n353875 );
buf ( n353877 , n33843 );
not ( n353878 , n353877 );
buf ( n353879 , n353878 );
not ( n33847 , n353879 );
not ( n353881 , n15164 );
not ( n353882 , n353732 );
or ( n33850 , n353881 , n353882 );
nand ( n353884 , n586 , n33710 );
not ( n353885 , n353884 );
buf ( n353886 , n342097 );
buf ( n353887 , n334982 );
nand ( n353888 , n353886 , n353887 );
buf ( n353889 , n353888 );
not ( n353890 , n353889 );
or ( n33858 , n353885 , n353890 );
nand ( n353892 , n33858 , n334978 );
nand ( n353893 , n33850 , n353892 );
not ( n353894 , n353893 );
or ( n33862 , n33847 , n353894 );
not ( n353896 , n353893 );
nand ( n353897 , n353896 , n33843 );
nand ( n353898 , n33862 , n353897 );
not ( n33866 , n335261 );
nand ( n353900 , n33866 , n576 );
not ( n353901 , n353900 );
not ( n33869 , n334727 );
not ( n353903 , n33756 );
or ( n353904 , n33869 , n353903 );
buf ( n353905 , n582 );
not ( n33873 , n353905 );
buf ( n353907 , n336167 );
not ( n353908 , n353907 );
or ( n33876 , n33873 , n353908 );
buf ( n353910 , n15217 );
buf ( n353911 , n334702 );
nand ( n353912 , n353910 , n353911 );
buf ( n353913 , n353912 );
buf ( n353914 , n353913 );
nand ( n353915 , n33876 , n353914 );
buf ( n353916 , n353915 );
nand ( n33884 , n353916 , n334694 );
nand ( n33885 , n353904 , n33884 );
not ( n353919 , n33885 );
or ( n353920 , n353901 , n353919 );
buf ( n353921 , n33885 );
buf ( n353922 , n353900 );
nor ( n353923 , n353921 , n353922 );
buf ( n353924 , n353923 );
not ( n353925 , n15528 );
buf ( n353926 , n580 );
not ( n353927 , n353926 );
buf ( n353928 , n335003 );
not ( n33896 , n353928 );
or ( n353930 , n353927 , n33896 );
buf ( n353931 , n333978 );
buf ( n353932 , n334650 );
nand ( n353933 , n353931 , n353932 );
buf ( n353934 , n353933 );
buf ( n353935 , n353934 );
nand ( n33903 , n353930 , n353935 );
buf ( n353937 , n33903 );
not ( n33905 , n353937 );
or ( n353939 , n353925 , n33905 );
not ( n33907 , n580 );
not ( n33908 , n33907 );
not ( n353942 , n15012 );
not ( n353943 , n353942 );
or ( n33911 , n33908 , n353943 );
or ( n353945 , n353942 , n33907 );
nand ( n353946 , n33911 , n353945 );
not ( n33914 , n353946 );
nand ( n353948 , n33914 , n14822 );
nand ( n353949 , n353939 , n353948 );
buf ( n353950 , n353949 );
not ( n33918 , n353950 );
buf ( n353952 , n33918 );
or ( n353953 , n353924 , n353952 );
nand ( n353954 , n353920 , n353953 );
not ( n33922 , n353954 );
and ( n33923 , n353898 , n33922 );
not ( n33924 , n353898 );
and ( n353958 , n33924 , n353954 );
nor ( n33926 , n33923 , n353958 );
not ( n353960 , n33926 );
or ( n353961 , n33824 , n353960 );
buf ( n33929 , n353900 );
buf ( n353963 , n353949 );
xor ( n353964 , n33929 , n353963 );
buf ( n353965 , n33885 );
xnor ( n33933 , n353964 , n353965 );
buf ( n353967 , n33933 );
buf ( n353968 , n353967 );
not ( n353969 , n353968 );
buf ( n353970 , n335177 );
not ( n33938 , n353970 );
buf ( n353972 , n338457 );
not ( n33940 , n353972 );
or ( n353974 , n33938 , n33940 );
and ( n33942 , n14099 , n335097 );
not ( n33943 , n14099 );
and ( n353977 , n33943 , n590 );
or ( n353978 , n33942 , n353977 );
buf ( n353979 , n353978 );
nand ( n353980 , n353974 , n353979 );
buf ( n353981 , n353980 );
buf ( n353982 , n334868 );
not ( n353983 , n353982 );
and ( n353984 , n15300 , n334879 );
not ( n353985 , n15300 );
and ( n33953 , n353985 , n584 );
or ( n353987 , n353984 , n33953 );
buf ( n353988 , n353987 );
not ( n33956 , n353988 );
or ( n353990 , n353983 , n33956 );
and ( n353991 , n15217 , n334879 );
not ( n33959 , n15217 );
and ( n33960 , n33959 , n584 );
or ( n33961 , n353991 , n33960 );
buf ( n353995 , n33961 );
buf ( n353996 , n334917 );
nand ( n33964 , n353995 , n353996 );
buf ( n353998 , n33964 );
buf ( n353999 , n353998 );
nand ( n354000 , n353990 , n353999 );
buf ( n354001 , n354000 );
nor ( n33969 , n353981 , n354001 );
buf ( n354003 , n33969 );
not ( n33971 , n354003 );
not ( n354005 , n16686 );
nand ( n354006 , n354005 , n576 );
not ( n33974 , n334643 );
xor ( n33975 , n33907 , n353942 );
not ( n354009 , n33975 );
or ( n354010 , n33974 , n354009 );
nand ( n33978 , n33785 , n14822 );
nand ( n354012 , n354010 , n33978 );
xor ( n33980 , n354006 , n354012 );
not ( n354014 , n14941 );
not ( n33982 , n353461 );
or ( n33983 , n354014 , n33982 );
and ( n354017 , n15381 , n334748 );
not ( n33985 , n15381 );
and ( n354019 , n33985 , n578 );
or ( n33987 , n354017 , n354019 );
nand ( n33988 , n33987 , n353009 );
nand ( n354022 , n33983 , n33988 );
xnor ( n354023 , n33980 , n354022 );
buf ( n354024 , n354023 );
nand ( n354025 , n33971 , n354024 );
buf ( n354026 , n354025 );
buf ( n354027 , n334868 );
not ( n354028 , n354027 );
buf ( n354029 , n353987 );
not ( n354030 , n354029 );
or ( n33998 , n354028 , n354030 );
buf ( n354032 , n353998 );
nand ( n354033 , n33998 , n354032 );
buf ( n354034 , n354033 );
buf ( n354035 , n354034 );
buf ( n354036 , n353981 );
nand ( n354037 , n354035 , n354036 );
buf ( n354038 , n354037 );
and ( n354039 , n354026 , n354038 );
buf ( n354040 , n354039 );
not ( n34008 , n354040 );
or ( n354042 , n353969 , n34008 );
and ( n34010 , n33477 , n353524 );
not ( n354044 , n33477 );
and ( n34012 , n354044 , n33488 );
nor ( n34013 , n34010 , n34012 );
not ( n354047 , n353480 );
and ( n354048 , n34013 , n354047 );
not ( n34016 , n34013 );
and ( n354050 , n34016 , n353480 );
nor ( n354051 , n354048 , n354050 );
not ( n34019 , n354051 );
not ( n354053 , n33975 );
not ( n354054 , n334643 );
or ( n354055 , n354053 , n354054 );
and ( n34023 , n33785 , n14822 );
not ( n354057 , n354006 );
nor ( n354058 , n34023 , n354057 );
nand ( n34026 , n354055 , n354058 );
not ( n354060 , n34026 );
not ( n354061 , n354022 );
or ( n34029 , n354060 , n354061 );
nand ( n34030 , n354012 , n354057 );
nand ( n34031 , n34029 , n34030 );
not ( n354065 , n34031 );
or ( n354066 , n34019 , n354065 );
not ( n34034 , n354051 );
not ( n34035 , n34031 );
nand ( n34036 , n34034 , n34035 );
nand ( n354070 , n354066 , n34036 );
not ( n354071 , n334917 );
not ( n34039 , n353987 );
or ( n34040 , n354071 , n34039 );
buf ( n354074 , n353862 );
buf ( n354075 , n334868 );
nand ( n354076 , n354074 , n354075 );
buf ( n354077 , n354076 );
nand ( n34045 , n34040 , n354077 );
and ( n34046 , n354070 , n34045 );
not ( n354080 , n354070 );
not ( n354081 , n34045 );
and ( n34049 , n354080 , n354081 );
nor ( n34050 , n34046 , n34049 );
buf ( n354084 , n34050 );
nand ( n354085 , n354042 , n354084 );
buf ( n354086 , n354085 );
buf ( n354087 , n353967 );
not ( n34055 , n354087 );
buf ( n354089 , n354026 );
buf ( n354090 , n354038 );
nand ( n354091 , n354089 , n354090 );
buf ( n354092 , n354091 );
buf ( n354093 , n354092 );
nand ( n354094 , n34055 , n354093 );
buf ( n354095 , n354094 );
nand ( n34063 , n354086 , n354095 );
nand ( n34064 , n353961 , n34063 );
buf ( n354098 , n34064 );
buf ( n354099 , n33926 );
not ( n354100 , n354099 );
buf ( n354101 , n354100 );
buf ( n354102 , n354101 );
buf ( n354103 , n353855 );
nand ( n354104 , n354102 , n354103 );
buf ( n354105 , n354104 );
buf ( n354106 , n354105 );
and ( n354107 , n354098 , n354106 );
buf ( n354108 , n354107 );
xor ( n34076 , n353703 , n354108 );
buf ( n354110 , n353954 );
not ( n354111 , n354110 );
buf ( n354112 , n353896 );
buf ( n354113 , n353879 );
nand ( n354114 , n354112 , n354113 );
buf ( n354115 , n354114 );
buf ( n354116 , n354115 );
not ( n354117 , n354116 );
or ( n354118 , n354111 , n354117 );
buf ( n354119 , n353896 );
not ( n354120 , n354119 );
buf ( n354121 , n33843 );
nand ( n354122 , n354120 , n354121 );
buf ( n354123 , n354122 );
buf ( n354124 , n354123 );
nand ( n34092 , n354118 , n354124 );
buf ( n354126 , n34092 );
buf ( n354127 , n354126 );
buf ( n354128 , n353900 );
not ( n354129 , n354128 );
buf ( n354130 , n354129 );
buf ( n354131 , n354130 );
buf ( n354132 , n334694 );
not ( n354133 , n354132 );
buf ( n354134 , n353663 );
not ( n354135 , n354134 );
or ( n354136 , n354133 , n354135 );
buf ( n354137 , n353916 );
buf ( n354138 , n334727 );
nand ( n34106 , n354137 , n354138 );
buf ( n354140 , n34106 );
buf ( n354141 , n354140 );
nand ( n354142 , n354136 , n354141 );
buf ( n354143 , n354142 );
buf ( n354144 , n354143 );
xor ( n34112 , n354131 , n354144 );
not ( n354146 , n15528 );
not ( n34114 , n33584 );
or ( n34115 , n354146 , n34114 );
buf ( n354149 , n14822 );
buf ( n354150 , n353937 );
nand ( n354151 , n354149 , n354150 );
buf ( n354152 , n354151 );
nand ( n34120 , n34115 , n354152 );
buf ( n354154 , n34120 );
and ( n354155 , n34112 , n354154 );
and ( n34123 , n354131 , n354144 );
or ( n354157 , n354155 , n34123 );
buf ( n354158 , n354157 );
not ( n34126 , n354158 );
not ( n354160 , n34126 );
not ( n34128 , n334917 );
not ( n354162 , n33841 );
or ( n34130 , n34128 , n354162 );
buf ( n354164 , n584 );
not ( n354165 , n354164 );
buf ( n354166 , n15992 );
not ( n354167 , n354166 );
or ( n34135 , n354165 , n354167 );
buf ( n354169 , n335851 );
buf ( n354170 , n334879 );
nand ( n354171 , n354169 , n354170 );
buf ( n354172 , n354171 );
buf ( n354173 , n354172 );
nand ( n354174 , n34135 , n354173 );
buf ( n354175 , n354174 );
nand ( n354176 , n354175 , n334868 );
nand ( n354177 , n34130 , n354176 );
not ( n354178 , n354177 );
not ( n34146 , n586 );
not ( n354180 , n33710 );
or ( n354181 , n34146 , n354180 );
nand ( n34149 , n354181 , n353889 );
and ( n354183 , n34149 , n15163 );
not ( n354184 , n325557 );
not ( n34152 , n14099 );
or ( n34153 , n354184 , n34152 );
buf ( n34154 , n325557 );
or ( n354188 , n34154 , n14099 );
nand ( n354189 , n34153 , n354188 );
nand ( n34157 , n354189 , n334978 );
not ( n354191 , n34157 );
nor ( n354192 , n354183 , n354191 );
not ( n34160 , n354192 );
or ( n354194 , n354178 , n34160 );
and ( n34162 , n34149 , n15163 );
nor ( n34163 , n34162 , n354191 );
or ( n354197 , n34163 , n354177 );
nand ( n34165 , n354194 , n354197 );
not ( n354199 , n34165 );
or ( n34167 , n354160 , n354199 );
not ( n34168 , n34165 );
nand ( n354202 , n34168 , n354158 );
nand ( n354203 , n34167 , n354202 );
buf ( n354204 , n354203 );
xor ( n354205 , n354127 , n354204 );
xor ( n354206 , n354131 , n354144 );
xor ( n34174 , n354206 , n354154 );
buf ( n354208 , n34174 );
not ( n354209 , n354208 );
nand ( n354210 , n34035 , n354081 );
not ( n34178 , n354051 );
and ( n354212 , n354210 , n34178 );
not ( n354213 , n334917 );
not ( n34181 , n353987 );
or ( n354215 , n354213 , n34181 );
nand ( n354216 , n354215 , n354077 );
and ( n34184 , n34031 , n354216 );
nor ( n354218 , n354212 , n34184 );
nand ( n34186 , n354209 , n354218 );
not ( n34187 , n34186 );
buf ( n354221 , n33526 );
not ( n34189 , n354221 );
buf ( n354223 , n353606 );
nand ( n354224 , n34189 , n354223 );
buf ( n354225 , n354224 );
buf ( n354226 , n354225 );
buf ( n34194 , n353599 );
not ( n354228 , n34194 );
buf ( n354229 , n354228 );
buf ( n354230 , n354229 );
and ( n354231 , n354226 , n354230 );
not ( n34199 , n354226 );
buf ( n354233 , n353599 );
and ( n354234 , n34199 , n354233 );
nor ( n34202 , n354231 , n354234 );
buf ( n354236 , n34202 );
not ( n34204 , n354236 );
or ( n354238 , n34187 , n34204 );
buf ( n354239 , n354218 );
not ( n34207 , n354239 );
buf ( n354241 , n34207 );
buf ( n354242 , n354241 );
buf ( n354243 , n354208 );
nand ( n354244 , n354242 , n354243 );
buf ( n354245 , n354244 );
nand ( n34213 , n354238 , n354245 );
buf ( n354247 , n34213 );
xnor ( n354248 , n354205 , n354247 );
buf ( n354249 , n354248 );
xor ( n354250 , n34076 , n354249 );
buf ( n354251 , n354208 );
buf ( n354252 , n354241 );
xor ( n354253 , n354251 , n354252 );
buf ( n354254 , n354236 );
xnor ( n34222 , n354253 , n354254 );
buf ( n354256 , n34222 );
buf ( n354257 , n334978 );
not ( n354258 , n354257 );
buf ( n354259 , n353717 );
not ( n34227 , n354259 );
or ( n354261 , n354258 , n34227 );
buf ( n354262 , n586 );
not ( n354263 , n354262 );
buf ( n34231 , n15290 );
not ( n354265 , n34231 );
buf ( n354266 , n354265 );
buf ( n354267 , n354266 );
not ( n354268 , n354267 );
or ( n34236 , n354263 , n354268 );
buf ( n354270 , n15290 );
buf ( n354271 , n334982 );
nand ( n354272 , n354270 , n354271 );
buf ( n354273 , n354272 );
buf ( n354274 , n354273 );
nand ( n354275 , n34236 , n354274 );
buf ( n354276 , n354275 );
buf ( n354277 , n354276 );
buf ( n354278 , n15164 );
nand ( n354279 , n354277 , n354278 );
buf ( n354280 , n354279 );
buf ( n354281 , n354280 );
nand ( n34249 , n354261 , n354281 );
buf ( n354283 , n34249 );
nand ( n354284 , n334694 , n353778 );
buf ( n354285 , n342175 );
buf ( n354286 , n334727 );
nand ( n354287 , n354285 , n354286 );
buf ( n354288 , n354287 );
and ( n34256 , n33987 , n334850 );
and ( n354290 , n342240 , n14949 );
nor ( n354291 , n34256 , n354290 );
nand ( n34259 , n354284 , n354288 , n354291 );
not ( n34260 , n34259 );
xor ( n354294 , n342197 , n342222 );
and ( n354295 , n354294 , n342248 );
and ( n34263 , n342197 , n342222 );
or ( n354297 , n354295 , n34263 );
buf ( n354298 , n354297 );
not ( n34266 , n354298 );
or ( n354300 , n34260 , n34266 );
not ( n354301 , n354291 );
nand ( n34269 , n354284 , n354288 );
nand ( n354303 , n354301 , n34269 );
nand ( n34271 , n354300 , n354303 );
xor ( n354305 , n354283 , n34271 );
buf ( n354306 , n15275 );
not ( n34274 , n354306 );
buf ( n354308 , n353750 );
not ( n34276 , n354308 );
or ( n354310 , n34274 , n34276 );
not ( n34278 , n588 );
not ( n34279 , n353031 );
or ( n354313 , n34278 , n34279 );
buf ( n354314 , n335851 );
buf ( n354315 , n334972 );
nand ( n354316 , n354314 , n354315 );
buf ( n354317 , n354316 );
nand ( n34285 , n354313 , n354317 );
buf ( n354319 , n34285 );
buf ( n354320 , n335114 );
nand ( n354321 , n354319 , n354320 );
buf ( n354322 , n354321 );
buf ( n354323 , n354322 );
nand ( n354324 , n354310 , n354323 );
buf ( n354325 , n354324 );
and ( n354326 , n354305 , n354325 );
and ( n354327 , n354283 , n34271 );
or ( n34295 , n354326 , n354327 );
buf ( n354329 , n34295 );
not ( n34297 , n354329 );
not ( n354331 , n353739 );
not ( n354332 , n33735 );
or ( n34300 , n354331 , n354332 );
buf ( n354334 , n353757 );
buf ( n354335 , n353762 );
nand ( n354336 , n354334 , n354335 );
buf ( n354337 , n354336 );
nand ( n34305 , n34300 , n354337 );
xor ( n354339 , n33820 , n34305 );
buf ( n354340 , n354339 );
not ( n34308 , n354340 );
buf ( n34309 , n34308 );
buf ( n354343 , n34309 );
nand ( n34311 , n34297 , n354343 );
buf ( n34312 , n34311 );
not ( n354346 , n334917 );
not ( n354347 , n22356 );
or ( n34315 , n354346 , n354347 );
buf ( n354349 , n33961 );
buf ( n354350 , n334868 );
nand ( n354351 , n354349 , n354350 );
buf ( n354352 , n354351 );
nand ( n34320 , n34315 , n354352 );
not ( n354354 , n34320 );
not ( n354355 , n354354 );
buf ( n354356 , n334978 );
not ( n34324 , n354356 );
buf ( n354358 , n354276 );
not ( n354359 , n354358 );
or ( n354360 , n34324 , n354359 );
buf ( n354361 , n342263 );
buf ( n354362 , n15164 );
nand ( n34330 , n354361 , n354362 );
buf ( n354364 , n34330 );
buf ( n354365 , n354364 );
nand ( n34333 , n354360 , n354365 );
buf ( n354367 , n34333 );
buf ( n354368 , n354367 );
not ( n354369 , n354368 );
buf ( n354370 , n354369 );
not ( n34338 , n354370 );
or ( n34339 , n354355 , n34338 );
not ( n34340 , n334643 );
not ( n354374 , n33785 );
or ( n354375 , n34340 , n354374 );
nand ( n34343 , n354375 , n33791 );
buf ( n354377 , n353843 );
not ( n34345 , n354377 );
buf ( n354379 , n353804 );
not ( n354380 , n354379 );
and ( n34348 , n34345 , n354380 );
buf ( n354382 , n14891 );
not ( n354383 , n354382 );
buf ( n354384 , n353519 );
not ( n34352 , n354384 );
or ( n354386 , n354383 , n34352 );
buf ( n354387 , n353840 );
nand ( n34355 , n354386 , n354387 );
buf ( n354389 , n34355 );
buf ( n354390 , n354389 );
buf ( n354391 , n353804 );
and ( n354392 , n354390 , n354391 );
nor ( n354393 , n34348 , n354392 );
buf ( n354394 , n354393 );
xor ( n34362 , n34343 , n354394 );
not ( n34363 , n34362 );
nand ( n34364 , n34339 , n34363 );
buf ( n354398 , n34364 );
not ( n354399 , n354370 );
nand ( n354400 , n354399 , n34320 );
buf ( n354401 , n354400 );
nand ( n354402 , n354398 , n354401 );
buf ( n354403 , n354402 );
buf ( n354404 , n354403 );
not ( n34372 , n354404 );
not ( n34373 , n354001 );
not ( n354407 , n34373 );
not ( n354408 , n353981 );
not ( n34376 , n354408 );
or ( n354410 , n354407 , n34376 );
nand ( n354411 , n354410 , n354038 );
and ( n34379 , n354411 , n354023 );
not ( n354413 , n354411 );
buf ( n354414 , n354023 );
not ( n34382 , n354414 );
buf ( n354416 , n34382 );
and ( n34384 , n354413 , n354416 );
nor ( n354418 , n34379 , n34384 );
not ( n34386 , n354418 );
buf ( n354420 , n34386 );
not ( n354421 , n354420 );
or ( n354422 , n34372 , n354421 );
buf ( n354423 , n354403 );
not ( n354424 , n354423 );
buf ( n354425 , n354424 );
buf ( n354426 , n354425 );
not ( n354427 , n354426 );
buf ( n354428 , n354418 );
not ( n34396 , n354428 );
or ( n354430 , n354427 , n34396 );
xor ( n34398 , n33488 , n353849 );
xnor ( n354432 , n34398 , n33758 );
not ( n354433 , n354432 );
buf ( n354434 , n354433 );
nand ( n354435 , n354430 , n354434 );
buf ( n354436 , n354435 );
buf ( n354437 , n354436 );
nand ( n34405 , n354422 , n354437 );
buf ( n354439 , n34405 );
and ( n354440 , n34312 , n354439 );
buf ( n354441 , n34295 );
buf ( n354442 , n354339 );
and ( n34410 , n354441 , n354442 );
buf ( n354444 , n34410 );
nor ( n34412 , n354440 , n354444 );
xor ( n354446 , n354256 , n34412 );
buf ( n354447 , n353855 );
buf ( n354448 , n354101 );
xor ( n354449 , n354447 , n354448 );
buf ( n354450 , n34063 );
xnor ( n34418 , n354449 , n354450 );
buf ( n34419 , n34418 );
and ( n354453 , n354446 , n34419 );
and ( n354454 , n354256 , n34412 );
or ( n34422 , n354453 , n354454 );
nand ( n354456 , n354250 , n34422 );
buf ( n354457 , n354456 );
or ( n34425 , n342182 , n342161 );
nand ( n354459 , n34425 , n342188 );
buf ( n354460 , n342182 );
buf ( n354461 , n342161 );
nand ( n354462 , n354460 , n354461 );
buf ( n354463 , n354462 );
nand ( n34431 , n354459 , n354463 );
buf ( n354465 , n34431 );
buf ( n354466 , n335114 );
not ( n354467 , n354466 );
buf ( n354468 , n342081 );
not ( n354469 , n354468 );
or ( n34437 , n354467 , n354469 );
nand ( n34438 , n34285 , n15275 );
buf ( n354472 , n34438 );
nand ( n354473 , n34437 , n354472 );
buf ( n354474 , n354473 );
buf ( n354475 , n354474 );
xor ( n354476 , n354465 , n354475 );
buf ( n354477 , n335181 );
not ( n354478 , n354477 );
buf ( n34446 , n22180 );
not ( n34447 , n34446 );
or ( n34448 , n354478 , n34447 );
buf ( n34449 , n353978 );
buf ( n34450 , n591 );
nand ( n34451 , n34449 , n34450 );
buf ( n34452 , n34451 );
buf ( n34453 , n34452 );
nand ( n34454 , n34448 , n34453 );
buf ( n34455 , n34454 );
buf ( n354489 , n34455 );
xor ( n34457 , n354476 , n354489 );
buf ( n354491 , n34457 );
not ( n34459 , n354491 );
not ( n34460 , n34459 );
not ( n354494 , n22167 );
not ( n354495 , n342108 );
or ( n34463 , n354494 , n354495 );
or ( n354497 , n342108 , n22167 );
nand ( n34465 , n354497 , n342066 );
nand ( n354499 , n34463 , n34465 );
not ( n354500 , n354499 );
not ( n34468 , n354500 );
or ( n354502 , n34460 , n34468 );
not ( n354503 , n22361 );
nand ( n34471 , n342192 , n342136 );
not ( n354505 , n34471 );
or ( n354506 , n354503 , n354505 );
nand ( n34474 , n342189 , n342135 );
nand ( n34475 , n354506 , n34474 );
nand ( n354509 , n354502 , n34475 );
nand ( n354510 , n354491 , n354499 );
and ( n34478 , n354509 , n354510 );
not ( n354512 , n34478 );
buf ( n354513 , n354433 );
not ( n34481 , n354513 );
buf ( n354515 , n354425 );
not ( n354516 , n354515 );
or ( n354517 , n34481 , n354516 );
buf ( n354518 , n354432 );
buf ( n354519 , n354403 );
nand ( n354520 , n354518 , n354519 );
buf ( n354521 , n354520 );
buf ( n354522 , n354521 );
nand ( n354523 , n354517 , n354522 );
buf ( n354524 , n354523 );
buf ( n354525 , n354524 );
buf ( n354526 , n354418 );
not ( n34494 , n354526 );
buf ( n354528 , n34494 );
and ( n354529 , n354525 , n354528 );
not ( n34497 , n354525 );
buf ( n354531 , n354526 );
and ( n354532 , n34497 , n354531 );
nor ( n34500 , n354529 , n354532 );
buf ( n354534 , n34500 );
buf ( n354535 , n354534 );
not ( n34503 , n354535 );
not ( n34504 , n34503 );
and ( n34505 , n354512 , n34504 );
buf ( n354539 , n34478 );
buf ( n354540 , n34503 );
nand ( n354541 , n354539 , n354540 );
buf ( n354542 , n354541 );
xor ( n34510 , n354465 , n354475 );
and ( n354544 , n34510 , n354489 );
and ( n34512 , n354465 , n354475 );
or ( n34513 , n354544 , n34512 );
buf ( n354547 , n34513 );
buf ( n354548 , n354547 );
xor ( n34516 , n354283 , n34271 );
xor ( n354550 , n34516 , n354325 );
buf ( n354551 , n354550 );
xor ( n34519 , n354548 , n354551 );
not ( n34520 , n354291 );
not ( n354554 , n354298 );
xor ( n34522 , n34520 , n354554 );
not ( n354556 , n34269 );
xnor ( n34524 , n34522 , n354556 );
not ( n354558 , n34524 );
xor ( n34526 , n342250 , n22346 );
and ( n34527 , n34526 , n22360 );
and ( n354561 , n342250 , n22346 );
or ( n34529 , n34527 , n354561 );
buf ( n354563 , n34529 );
not ( n354564 , n354563 );
buf ( n354565 , n354564 );
not ( n34533 , n354565 );
or ( n354567 , n354558 , n34533 );
not ( n354568 , n354354 );
not ( n34536 , n354367 );
nand ( n354570 , n34536 , n34363 );
nand ( n354571 , n354367 , n34362 );
nand ( n34539 , n354570 , n354571 );
not ( n34540 , n34539 );
or ( n354574 , n354568 , n34540 );
nand ( n354575 , n354570 , n34320 , n354571 );
nand ( n34543 , n354574 , n354575 );
nand ( n354577 , n354567 , n34543 );
buf ( n354578 , n354565 );
not ( n34546 , n354578 );
xor ( n354580 , n34520 , n354554 );
buf ( n354581 , n34269 );
xnor ( n354582 , n354580 , n354581 );
buf ( n354583 , n354582 );
nand ( n354584 , n34546 , n354583 );
buf ( n354585 , n354584 );
nand ( n34553 , n354577 , n354585 );
buf ( n354587 , n34553 );
xor ( n34555 , n34519 , n354587 );
buf ( n354589 , n34555 );
buf ( n354590 , n354589 );
buf ( n34558 , n354590 );
buf ( n354592 , n34558 );
and ( n354593 , n354542 , n354592 );
nor ( n34561 , n34505 , n354593 );
buf ( n354595 , n353967 );
buf ( n354596 , n354092 );
xor ( n34564 , n354595 , n354596 );
buf ( n354598 , n34050 );
xnor ( n354599 , n34564 , n354598 );
buf ( n354600 , n354599 );
buf ( n354601 , n354600 );
xor ( n354602 , n354548 , n354551 );
and ( n354603 , n354602 , n354587 );
and ( n34571 , n354548 , n354551 );
or ( n354605 , n354603 , n34571 );
buf ( n354606 , n354605 );
buf ( n354607 , n354606 );
xor ( n34575 , n354601 , n354607 );
xor ( n34576 , n354441 , n354442 );
buf ( n354610 , n34576 );
xor ( n34578 , n354610 , n354439 );
buf ( n354612 , n34578 );
xnor ( n354613 , n34575 , n354612 );
buf ( n354614 , n354613 );
nand ( n354615 , n34561 , n354614 );
buf ( n354616 , n354615 );
nand ( n34584 , n354457 , n354616 );
buf ( n354618 , n34584 );
not ( n34586 , n354618 );
buf ( n354620 , n34586 );
not ( n354621 , n354620 );
xor ( n354622 , n354256 , n34412 );
xor ( n354623 , n354622 , n34419 );
buf ( n354624 , n354600 );
buf ( n354625 , n354624 );
buf ( n354626 , n354625 );
buf ( n354627 , n354626 );
not ( n34595 , n354627 );
buf ( n354629 , n354606 );
not ( n354630 , n354629 );
buf ( n354631 , n354630 );
buf ( n354632 , n354631 );
nand ( n354633 , n34595 , n354632 );
buf ( n354634 , n354633 );
buf ( n34602 , n34578 );
and ( n354636 , n354634 , n34602 );
buf ( n354637 , n354626 );
not ( n34605 , n354637 );
buf ( n354639 , n354631 );
nor ( n354640 , n34605 , n354639 );
buf ( n354641 , n354640 );
nor ( n34609 , n354636 , n354641 );
nand ( n354643 , n354623 , n34609 );
buf ( n354644 , n354643 );
buf ( n354645 , n34561 );
not ( n354646 , n354645 );
buf ( n354647 , n354646 );
buf ( n354648 , n354614 );
not ( n354649 , n354648 );
buf ( n354650 , n354649 );
nand ( n354651 , n354647 , n354650 );
buf ( n354652 , n354534 );
buf ( n354653 , n354589 );
xor ( n34621 , n354652 , n354653 );
buf ( n354655 , n34478 );
xnor ( n34623 , n34621 , n354655 );
buf ( n354657 , n34623 );
buf ( n354658 , n34529 );
buf ( n354659 , n354582 );
and ( n354660 , n354658 , n354659 );
not ( n34628 , n354658 );
buf ( n34629 , n34524 );
and ( n354663 , n34628 , n34629 );
nor ( n34631 , n354660 , n354663 );
buf ( n34632 , n34631 );
and ( n354666 , n34543 , n34632 );
not ( n34634 , n34543 );
not ( n354668 , n34632 );
and ( n354669 , n34634 , n354668 );
or ( n34637 , n354666 , n354669 );
not ( n354671 , n34637 );
buf ( n354672 , n342035 );
buf ( n354673 , n354672 );
not ( n34641 , n354673 );
buf ( n354675 , n342050 );
not ( n34643 , n354675 );
or ( n34644 , n34641 , n34643 );
buf ( n354678 , n342035 );
not ( n354679 , n354678 );
buf ( n354680 , n354679 );
buf ( n354681 , n354680 );
not ( n354682 , n354681 );
buf ( n354683 , n342056 );
not ( n34651 , n354683 );
or ( n34652 , n354682 , n34651 );
buf ( n354686 , n342111 );
nand ( n34654 , n34652 , n354686 );
buf ( n354688 , n34654 );
buf ( n354689 , n354688 );
nand ( n34657 , n34644 , n354689 );
buf ( n354691 , n34657 );
not ( n34659 , n354691 );
not ( n34660 , n34659 );
or ( n34661 , n354671 , n34660 );
not ( n34662 , n354499 );
not ( n354696 , n34459 );
or ( n34664 , n34662 , n354696 );
nand ( n34665 , n354500 , n354491 );
nand ( n34666 , n34664 , n34665 );
and ( n34667 , n34666 , n34475 );
not ( n354701 , n34666 );
not ( n354702 , n34475 );
and ( n34670 , n354701 , n354702 );
nor ( n354704 , n34667 , n34670 );
nand ( n354705 , n34661 , n354704 );
buf ( n354706 , n354705 );
not ( n34674 , n34637 );
nand ( n354708 , n34674 , n354691 );
buf ( n354709 , n354708 );
nand ( n354710 , n354706 , n354709 );
buf ( n354711 , n354710 );
nand ( n34679 , n354657 , n354711 );
nand ( n34680 , n354651 , n34679 );
buf ( n354714 , n34680 );
nand ( n34682 , n354644 , n354714 );
buf ( n354716 , n34682 );
not ( n34684 , n354716 );
buf ( n354718 , n34684 );
not ( n354719 , n354718 );
or ( n354720 , n354621 , n354719 );
not ( n34688 , n354456 );
buf ( n354722 , n354623 );
not ( n354723 , n354722 );
buf ( n354724 , n354723 );
not ( n354725 , n34609 );
nand ( n354726 , n354724 , n354725 );
not ( n34694 , n354726 );
not ( n354728 , n34694 );
or ( n354729 , n34688 , n354728 );
not ( n34697 , n34422 );
not ( n354731 , n354250 );
nand ( n34699 , n34697 , n354731 );
buf ( n354733 , n34699 );
nand ( n354734 , n354729 , n354733 );
buf ( n354735 , n354734 );
not ( n354736 , n354735 );
buf ( n354737 , n354736 );
buf ( n354738 , n354737 );
nand ( n34706 , n354720 , n354738 );
buf ( n354740 , n34706 );
xor ( n34708 , n353175 , n353353 );
xor ( n354742 , n34708 , n353359 );
buf ( n354743 , n354742 );
not ( n34711 , n354743 );
buf ( n354745 , n34711 );
xor ( n354746 , n353186 , n353203 );
xor ( n34714 , n354746 , n353229 );
buf ( n354748 , n34714 );
buf ( n354749 , n354748 );
not ( n34717 , n354749 );
buf ( n354751 , n584 );
not ( n354752 , n354751 );
buf ( n354753 , n352857 );
not ( n34721 , n354753 );
or ( n354755 , n354752 , n34721 );
buf ( n354756 , n14099 );
buf ( n354757 , n334879 );
nand ( n354758 , n354756 , n354757 );
buf ( n354759 , n354758 );
buf ( n354760 , n354759 );
nand ( n34728 , n354755 , n354760 );
buf ( n354762 , n34728 );
buf ( n354763 , n354762 );
buf ( n34731 , n336786 );
buf ( n354765 , n33832 );
nand ( n34733 , n34731 , n354765 );
buf ( n354767 , n34733 );
buf ( n354768 , n354767 );
nand ( n34736 , n354763 , n354768 );
buf ( n354770 , n34736 );
buf ( n354771 , n354770 );
buf ( n354772 , n14891 );
not ( n34740 , n354772 );
buf ( n354774 , n33159 );
not ( n354775 , n354774 );
or ( n34743 , n34740 , n354775 );
not ( n354777 , n576 );
not ( n354778 , n337088 );
or ( n34746 , n354777 , n354778 );
buf ( n354780 , n337085 );
buf ( n354781 , n332672 );
nand ( n354782 , n354780 , n354781 );
buf ( n354783 , n354782 );
nand ( n354784 , n34746 , n354783 );
buf ( n354785 , n354784 );
buf ( n354786 , n334786 );
nand ( n34754 , n354785 , n354786 );
buf ( n354788 , n34754 );
buf ( n354789 , n354788 );
nand ( n34757 , n34743 , n354789 );
buf ( n34758 , n34757 );
buf ( n354792 , n34758 );
xor ( n354793 , n354771 , n354792 );
buf ( n354794 , n334643 );
not ( n354795 , n354794 );
buf ( n354796 , n353299 );
not ( n34764 , n354796 );
or ( n354798 , n354795 , n34764 );
buf ( n354799 , n580 );
not ( n34767 , n354799 );
buf ( n354801 , n335808 );
not ( n354802 , n354801 );
or ( n34770 , n34767 , n354802 );
buf ( n354804 , n15290 );
buf ( n354805 , n334650 );
nand ( n34773 , n354804 , n354805 );
buf ( n354807 , n34773 );
buf ( n354808 , n354807 );
nand ( n34776 , n34770 , n354808 );
buf ( n34777 , n34776 );
buf ( n354811 , n34777 );
buf ( n354812 , n14822 );
nand ( n354813 , n354811 , n354812 );
buf ( n354814 , n354813 );
buf ( n354815 , n354814 );
nand ( n34783 , n354798 , n354815 );
buf ( n34784 , n34783 );
buf ( n354818 , n34784 );
and ( n34786 , n354793 , n354818 );
and ( n354820 , n354771 , n354792 );
or ( n354821 , n34786 , n354820 );
buf ( n354822 , n354821 );
buf ( n354823 , n354822 );
not ( n354824 , n354823 );
or ( n34792 , n34717 , n354824 );
buf ( n354826 , n354748 );
not ( n354827 , n354826 );
buf ( n354828 , n354827 );
buf ( n354829 , n354828 );
not ( n354830 , n354829 );
buf ( n354831 , n354822 );
not ( n354832 , n354831 );
buf ( n354833 , n354832 );
buf ( n34801 , n354833 );
not ( n34802 , n34801 );
or ( n34803 , n354830 , n34802 );
buf ( n354837 , n334694 );
not ( n34805 , n354837 );
buf ( n354839 , n353324 );
not ( n354840 , n354839 );
or ( n354841 , n34805 , n354840 );
buf ( n354842 , n582 );
not ( n354843 , n354842 );
buf ( n354844 , n353031 );
not ( n34812 , n354844 );
or ( n354846 , n354843 , n34812 );
buf ( n354847 , n353034 );
buf ( n354848 , n334702 );
nand ( n354849 , n354847 , n354848 );
buf ( n354850 , n354849 );
buf ( n354851 , n354850 );
nand ( n34819 , n354846 , n354851 );
buf ( n34820 , n34819 );
buf ( n34821 , n34820 );
buf ( n354855 , n334727 );
nand ( n354856 , n34821 , n354855 );
buf ( n354857 , n354856 );
buf ( n354858 , n354857 );
nand ( n34826 , n354841 , n354858 );
buf ( n354860 , n34826 );
buf ( n354861 , n354860 );
not ( n354862 , n354861 );
buf ( n354863 , n33241 );
not ( n34831 , n354863 );
buf ( n354865 , n353239 );
not ( n354866 , n354865 );
buf ( n354867 , n353282 );
not ( n34835 , n354867 );
and ( n354869 , n354866 , n34835 );
buf ( n354870 , n353282 );
buf ( n354871 , n353239 );
and ( n34839 , n354870 , n354871 );
nor ( n354873 , n354869 , n34839 );
buf ( n354874 , n354873 );
buf ( n354875 , n354874 );
not ( n34843 , n354875 );
and ( n354877 , n34831 , n34843 );
buf ( n354878 , n33241 );
buf ( n354879 , n354874 );
and ( n34847 , n354878 , n354879 );
nor ( n354881 , n354877 , n34847 );
buf ( n354882 , n354881 );
buf ( n354883 , n354882 );
nand ( n354884 , n354862 , n354883 );
buf ( n354885 , n354884 );
buf ( n354886 , n354885 );
buf ( n354887 , n353245 );
not ( n354888 , n354887 );
buf ( n354889 , n334643 );
not ( n34857 , n354889 );
buf ( n354891 , n34777 );
not ( n354892 , n354891 );
or ( n34860 , n34857 , n354892 );
buf ( n354894 , n580 );
not ( n354895 , n354894 );
buf ( n354896 , n24387 );
not ( n354897 , n354896 );
or ( n34865 , n354895 , n354897 );
buf ( n354899 , n15300 );
buf ( n354900 , n334650 );
nand ( n34868 , n354899 , n354900 );
buf ( n354902 , n34868 );
buf ( n354903 , n354902 );
nand ( n354904 , n34865 , n354903 );
buf ( n354905 , n354904 );
buf ( n354906 , n354905 );
buf ( n354907 , n14822 );
nand ( n354908 , n354906 , n354907 );
buf ( n354909 , n354908 );
buf ( n354910 , n354909 );
nand ( n34878 , n34860 , n354910 );
buf ( n354912 , n34878 );
buf ( n354913 , n354912 );
not ( n354914 , n354913 );
or ( n34882 , n354888 , n354914 );
buf ( n354916 , n354912 );
buf ( n354917 , n353245 );
or ( n34885 , n354916 , n354917 );
not ( n354919 , n14891 );
not ( n354920 , n354784 );
or ( n34888 , n354919 , n354920 );
xor ( n34889 , n576 , n15341 );
buf ( n34890 , n34889 );
buf ( n34891 , n334786 );
nand ( n34892 , n34890 , n34891 );
buf ( n34893 , n34892 );
nand ( n354927 , n34888 , n34893 );
buf ( n354928 , n354927 );
nand ( n354929 , n34885 , n354928 );
buf ( n354930 , n354929 );
buf ( n354931 , n354930 );
nand ( n34899 , n34882 , n354931 );
buf ( n354933 , n34899 );
buf ( n354934 , n354933 );
and ( n354935 , n354886 , n354934 );
buf ( n354936 , n354860 );
not ( n34904 , n354936 );
buf ( n354938 , n354882 );
nor ( n354939 , n34904 , n354938 );
buf ( n354940 , n354939 );
buf ( n354941 , n354940 );
nor ( n34909 , n354935 , n354941 );
buf ( n354943 , n34909 );
buf ( n34911 , n354943 );
not ( n354945 , n34911 );
buf ( n354946 , n354945 );
buf ( n354947 , n354946 );
nand ( n34915 , n34803 , n354947 );
buf ( n354949 , n34915 );
buf ( n354950 , n354949 );
nand ( n354951 , n34792 , n354950 );
buf ( n354952 , n354951 );
buf ( n354953 , n354952 );
and ( n354954 , n32980 , n32986 );
not ( n34922 , n32980 );
and ( n354956 , n34922 , n32943 );
or ( n354957 , n354954 , n354956 );
and ( n34925 , n354957 , n33019 );
not ( n354959 , n354957 );
not ( n354960 , n33019 );
and ( n34928 , n354959 , n354960 );
nor ( n354962 , n34925 , n34928 );
buf ( n354963 , n354962 );
or ( n354964 , n354953 , n354963 );
xor ( n354965 , n353185 , n353234 );
xor ( n34933 , n354965 , n353349 );
buf ( n354967 , n34933 );
buf ( n354968 , n354967 );
nand ( n34936 , n354964 , n354968 );
buf ( n354970 , n34936 );
buf ( n354971 , n354952 );
buf ( n354972 , n354962 );
nand ( n354973 , n354971 , n354972 );
buf ( n354974 , n354973 );
nand ( n34942 , n354970 , n354974 );
not ( n34943 , n34942 );
nand ( n354977 , n354745 , n34943 );
xor ( n354978 , n353329 , n353288 );
xor ( n34946 , n354978 , n353346 );
xor ( n34947 , n354748 , n354833 );
xnor ( n34948 , n34947 , n354943 );
xor ( n354982 , n34946 , n34948 );
xor ( n354983 , n354771 , n354792 );
xor ( n34951 , n354983 , n354818 );
buf ( n354985 , n34951 );
not ( n34953 , n354985 );
buf ( n354987 , n336865 );
buf ( n354988 , n576 );
nand ( n34956 , n354987 , n354988 );
buf ( n354990 , n34956 );
buf ( n354991 , n354990 );
buf ( n354992 , n353407 );
nand ( n34960 , n354991 , n354992 );
buf ( n354994 , n34960 );
buf ( n354995 , n354994 );
not ( n34963 , n354995 );
buf ( n354997 , n334786 );
not ( n34965 , n354997 );
buf ( n354999 , n353395 );
not ( n355000 , n354999 );
or ( n34968 , n34965 , n355000 );
buf ( n355002 , n34889 );
buf ( n355003 , n14891 );
nand ( n355004 , n355002 , n355003 );
buf ( n355005 , n355004 );
buf ( n355006 , n355005 );
nand ( n34974 , n34968 , n355006 );
buf ( n355008 , n34974 );
buf ( n355009 , n355008 );
not ( n355010 , n355009 );
or ( n34978 , n34963 , n355010 );
buf ( n355012 , n354990 );
not ( n34980 , n355012 );
buf ( n355014 , n353371 );
nand ( n34982 , n34980 , n355014 );
buf ( n355016 , n34982 );
buf ( n355017 , n355016 );
nand ( n34985 , n34978 , n355017 );
buf ( n34986 , n34985 );
not ( n34987 , n353009 );
buf ( n355021 , n334748 );
not ( n34989 , n355021 );
buf ( n355023 , n337902 );
not ( n34991 , n355023 );
or ( n355025 , n34989 , n34991 );
buf ( n355026 , n337894 );
not ( n34994 , n355026 );
buf ( n355028 , n578 );
nand ( n355029 , n34994 , n355028 );
buf ( n355030 , n355029 );
buf ( n355031 , n355030 );
nand ( n355032 , n355025 , n355031 );
buf ( n355033 , n355032 );
not ( n355034 , n355033 );
or ( n355035 , n34987 , n355034 );
buf ( n355036 , n353267 );
buf ( n355037 , n334850 );
nand ( n355038 , n355036 , n355037 );
buf ( n355039 , n355038 );
nand ( n355040 , n355035 , n355039 );
xor ( n355041 , n34986 , n355040 );
buf ( n355042 , n334917 );
not ( n35010 , n355042 );
not ( n35011 , n584 );
not ( n35012 , n352031 );
or ( n35013 , n35011 , n35012 );
buf ( n355047 , n342097 );
buf ( n355048 , n334879 );
nand ( n35016 , n355047 , n355048 );
buf ( n355050 , n35016 );
nand ( n35018 , n35013 , n355050 );
buf ( n355052 , n35018 );
not ( n35020 , n355052 );
or ( n35021 , n35010 , n35020 );
buf ( n355055 , n354762 );
buf ( n355056 , n334868 );
nand ( n355057 , n355055 , n355056 );
buf ( n355058 , n355057 );
buf ( n355059 , n355058 );
nand ( n35027 , n35021 , n355059 );
buf ( n355061 , n35027 );
and ( n35029 , n355041 , n355061 );
and ( n355063 , n34986 , n355040 );
or ( n355064 , n35029 , n355063 );
not ( n35032 , n355064 );
and ( n35033 , n34953 , n35032 );
xor ( n355067 , n354860 , n354933 );
and ( n355068 , n355067 , n354882 );
not ( n35036 , n355067 );
buf ( n355070 , n354882 );
not ( n35038 , n355070 );
buf ( n355072 , n35038 );
and ( n35040 , n35036 , n355072 );
nor ( n355074 , n355068 , n35040 );
nor ( n355075 , n35033 , n355074 );
buf ( n355076 , n355064 );
buf ( n355077 , n354985 );
and ( n355078 , n355076 , n355077 );
buf ( n355079 , n355078 );
nor ( n355080 , n355075 , n355079 );
and ( n355081 , n354982 , n355080 );
and ( n35049 , n34946 , n34948 );
or ( n355083 , n355081 , n35049 );
buf ( n35051 , n355083 );
buf ( n355085 , n354962 );
buf ( n355086 , n354967 );
xor ( n35054 , n355085 , n355086 );
buf ( n355088 , n354952 );
xnor ( n355089 , n35054 , n355088 );
buf ( n355090 , n355089 );
buf ( n355091 , n355090 );
nand ( n355092 , n35051 , n355091 );
buf ( n355093 , n355092 );
nand ( n355094 , n354977 , n355093 );
not ( n35062 , n355094 );
not ( n355096 , n35062 );
not ( n35064 , n353452 );
nand ( n355098 , n35064 , n353701 , n33666 );
not ( n35066 , n355098 );
not ( n355100 , n33574 );
or ( n35068 , n35066 , n355100 );
not ( n35069 , n353701 );
not ( n35070 , n33666 );
or ( n355104 , n35069 , n35070 );
nand ( n355105 , n355104 , n353452 );
nand ( n35073 , n35068 , n355105 );
not ( n35074 , n35073 );
not ( n355108 , n354158 );
buf ( n355109 , n334917 );
not ( n35077 , n355109 );
buf ( n355111 , n33841 );
not ( n355112 , n355111 );
or ( n355113 , n35077 , n355112 );
buf ( n355114 , n354176 );
nand ( n35082 , n355113 , n355114 );
buf ( n355116 , n35082 );
not ( n355117 , n355116 );
nand ( n355118 , n355117 , n34163 );
not ( n35086 , n355118 );
or ( n35087 , n355108 , n35086 );
not ( n355121 , n354192 );
nand ( n355122 , n355121 , n355116 );
nand ( n355123 , n35087 , n355122 );
not ( n35091 , n355123 );
not ( n355125 , n355008 );
not ( n35093 , n354990 );
and ( n35094 , n353371 , n35093 );
not ( n355128 , n353371 );
and ( n35096 , n355128 , n354990 );
nor ( n355130 , n35094 , n35096 );
not ( n35098 , n355130 );
and ( n35099 , n355125 , n35098 );
and ( n355133 , n355008 , n355130 );
nor ( n355134 , n35099 , n355133 );
buf ( n355135 , n353651 );
not ( n355136 , n355135 );
buf ( n355137 , n355136 );
not ( n35105 , n355137 );
not ( n355139 , n336910 );
and ( n355140 , n35105 , n355139 );
buf ( n355141 , n582 );
not ( n35109 , n355141 );
buf ( n355143 , n15975 );
not ( n355144 , n355143 );
or ( n35112 , n35109 , n355144 );
buf ( n355146 , n14199 );
buf ( n35114 , n334702 );
nand ( n35115 , n355146 , n35114 );
buf ( n355149 , n35115 );
buf ( n355150 , n355149 );
nand ( n355151 , n35112 , n355150 );
buf ( n355152 , n355151 );
and ( n355153 , n355152 , n334694 );
nor ( n35121 , n355140 , n355153 );
and ( n35122 , n355134 , n35121 );
not ( n355156 , n355134 );
not ( n355157 , n35121 );
and ( n35125 , n355156 , n355157 );
or ( n355159 , n35122 , n35125 );
not ( n355160 , n334868 );
not ( n35128 , n35018 );
or ( n355162 , n355160 , n35128 );
nand ( n355163 , n354175 , n334917 );
nand ( n35131 , n355162 , n355163 );
buf ( n35132 , n35131 );
and ( n355166 , n355159 , n35132 );
not ( n355167 , n355159 );
not ( n35135 , n35131 );
and ( n355169 , n355167 , n35135 );
nor ( n355170 , n355166 , n355169 );
not ( n35138 , n355170 );
nand ( n355172 , n35091 , n35138 );
not ( n355173 , n355172 );
or ( n355174 , n35074 , n355173 );
not ( n35142 , n35091 );
nand ( n35143 , n35142 , n355170 );
nand ( n35144 , n355174 , n35143 );
buf ( n355178 , n35144 );
not ( n35146 , n355178 );
buf ( n355180 , n334694 );
not ( n35148 , n355180 );
buf ( n355182 , n34820 );
not ( n355183 , n355182 );
or ( n355184 , n35148 , n355183 );
buf ( n355185 , n355152 );
buf ( n355186 , n334727 );
nand ( n355187 , n355185 , n355186 );
buf ( n355188 , n355187 );
buf ( n355189 , n355188 );
nand ( n355190 , n355184 , n355189 );
buf ( n355191 , n355190 );
buf ( n355192 , n355191 );
or ( n35160 , n15164 , n334978 );
nand ( n355194 , n354189 , n35160 );
buf ( n355195 , n355194 );
buf ( n355196 , n334643 );
not ( n35164 , n355196 );
buf ( n355198 , n354905 );
not ( n355199 , n355198 );
or ( n355200 , n35164 , n355199 );
buf ( n355201 , n353631 );
buf ( n355202 , n14822 );
nand ( n355203 , n355201 , n355202 );
buf ( n355204 , n355203 );
buf ( n355205 , n355204 );
nand ( n355206 , n355200 , n355205 );
buf ( n355207 , n355206 );
buf ( n355208 , n355207 );
xor ( n355209 , n355195 , n355208 );
buf ( n355210 , n335432 );
not ( n35178 , n355210 );
buf ( n355212 , n355033 );
not ( n355213 , n355212 );
or ( n35181 , n35178 , n355213 );
buf ( n355215 , n353425 );
buf ( n355216 , n353009 );
nand ( n35184 , n355215 , n355216 );
buf ( n355218 , n35184 );
buf ( n355219 , n355218 );
nand ( n355220 , n35181 , n355219 );
buf ( n355221 , n355220 );
buf ( n355222 , n355221 );
and ( n35190 , n355209 , n355222 );
and ( n35191 , n355195 , n355208 );
or ( n355225 , n35190 , n35191 );
buf ( n355226 , n355225 );
buf ( n355227 , n355226 );
xor ( n35195 , n355192 , n355227 );
buf ( n355229 , n353282 );
buf ( n355230 , n354927 );
xor ( n355231 , n355229 , n355230 );
buf ( n355232 , n354912 );
xnor ( n355233 , n355231 , n355232 );
buf ( n355234 , n355233 );
buf ( n355235 , n355234 );
xor ( n355236 , n35195 , n355235 );
buf ( n355237 , n355236 );
buf ( n355238 , n355237 );
not ( n355239 , n355238 );
buf ( n355240 , n355239 );
buf ( n355241 , n355240 );
nand ( n35209 , n35146 , n355241 );
buf ( n355243 , n35209 );
buf ( n355244 , n355243 );
or ( n35212 , n35131 , n355157 );
nand ( n35213 , n35212 , n355134 );
buf ( n355247 , n35213 );
nand ( n35215 , n35131 , n355157 );
buf ( n355249 , n35215 );
nand ( n355250 , n355247 , n355249 );
buf ( n355251 , n355250 );
buf ( n355252 , n355251 );
xor ( n35220 , n34986 , n355040 );
xor ( n35221 , n35220 , n355061 );
buf ( n355255 , n35221 );
xor ( n35223 , n355252 , n355255 );
not ( n355257 , n33368 );
nand ( n35225 , n355257 , n353371 );
not ( n35226 , n35225 );
not ( n35227 , n353447 );
or ( n355261 , n35226 , n35227 );
buf ( n35229 , n33368 );
buf ( n355263 , n353407 );
nand ( n35231 , n35229 , n355263 );
buf ( n355265 , n35231 );
nand ( n35233 , n355261 , n355265 );
buf ( n355267 , n35233 );
not ( n35235 , n355267 );
buf ( n355269 , n35235 );
buf ( n355270 , n355269 );
not ( n35238 , n355270 );
not ( n355272 , n353673 );
not ( n355273 , n33600 );
not ( n35241 , n355273 );
and ( n355275 , n355272 , n35241 );
nand ( n355276 , n353673 , n355273 );
and ( n35244 , n355276 , n353698 );
nor ( n355278 , n355275 , n35244 );
buf ( n355279 , n355278 );
not ( n35247 , n355279 );
or ( n355281 , n35238 , n35247 );
xor ( n35249 , n355195 , n355208 );
xor ( n355283 , n35249 , n355222 );
buf ( n355284 , n355283 );
buf ( n355285 , n355284 );
nand ( n355286 , n355281 , n355285 );
buf ( n355287 , n355286 );
buf ( n355288 , n355287 );
buf ( n355289 , n355278 );
not ( n35257 , n355289 );
buf ( n355291 , n35233 );
buf ( n355292 , n355291 );
nand ( n35260 , n35257 , n355292 );
buf ( n355294 , n35260 );
buf ( n355295 , n355294 );
nand ( n355296 , n355288 , n355295 );
buf ( n355297 , n355296 );
buf ( n355298 , n355297 );
xor ( n355299 , n35223 , n355298 );
buf ( n355300 , n355299 );
buf ( n355301 , n355300 );
buf ( n35269 , n355301 );
buf ( n355303 , n35269 );
buf ( n355304 , n355303 );
and ( n35272 , n355244 , n355304 );
buf ( n355306 , n35144 );
not ( n35274 , n355306 );
buf ( n355308 , n355240 );
nor ( n355309 , n35274 , n355308 );
buf ( n355310 , n355309 );
buf ( n355311 , n355310 );
nor ( n35279 , n35272 , n355311 );
buf ( n355313 , n35279 );
buf ( n355314 , n355313 );
xor ( n35282 , n355192 , n355227 );
and ( n35283 , n35282 , n355235 );
and ( n35284 , n355192 , n355227 );
or ( n355318 , n35283 , n35284 );
buf ( n355319 , n355318 );
buf ( n355320 , n355319 );
xor ( n35288 , n355252 , n355255 );
and ( n35289 , n35288 , n355298 );
and ( n355323 , n355252 , n355255 );
or ( n355324 , n35289 , n355323 );
buf ( n355325 , n355324 );
buf ( n355326 , n355325 );
xor ( n355327 , n355320 , n355326 );
xor ( n35295 , n355076 , n355077 );
buf ( n355329 , n35295 );
not ( n355330 , n355329 );
and ( n355331 , n355074 , n355330 );
not ( n35299 , n355074 );
and ( n35300 , n35299 , n355329 );
nor ( n355334 , n355331 , n35300 );
buf ( n355335 , n355334 );
xnor ( n35303 , n355327 , n355335 );
buf ( n355337 , n35303 );
buf ( n355338 , n355337 );
nand ( n355339 , n355314 , n355338 );
buf ( n355340 , n355339 );
buf ( n355341 , n355340 );
xor ( n35309 , n34946 , n34948 );
xor ( n355343 , n35309 , n355080 );
buf ( n35311 , n355343 );
buf ( n355345 , n355319 );
buf ( n355346 , n355334 );
or ( n355347 , n355345 , n355346 );
buf ( n355348 , n355325 );
nand ( n35316 , n355347 , n355348 );
buf ( n355350 , n35316 );
buf ( n35318 , n355334 );
buf ( n355352 , n355319 );
nand ( n35320 , n35318 , n355352 );
buf ( n35321 , n35320 );
and ( n355355 , n355350 , n35321 );
buf ( n355356 , n355355 );
nand ( n35324 , n35311 , n355356 );
buf ( n355358 , n35324 );
buf ( n35326 , n355358 );
and ( n35327 , n355341 , n35326 );
buf ( n35328 , n35327 );
not ( n355362 , n354108 );
not ( n35330 , n353703 );
nand ( n355364 , n355362 , n35330 );
and ( n355365 , n354249 , n355364 );
and ( n35333 , n353703 , n354108 );
nor ( n355367 , n355365 , n35333 );
not ( n35335 , n355367 );
buf ( n355369 , n355284 );
buf ( n355370 , n355269 );
and ( n35338 , n355369 , n355370 );
not ( n355372 , n355369 );
buf ( n355373 , n355291 );
and ( n35341 , n355372 , n355373 );
nor ( n355375 , n35338 , n35341 );
buf ( n355376 , n355375 );
buf ( n355377 , n355278 );
buf ( n355378 , n355377 );
buf ( n355379 , n355378 );
xnor ( n355380 , n355376 , n355379 );
buf ( n355381 , n355380 );
buf ( n355382 , n34213 );
buf ( n355383 , n354126 );
not ( n35351 , n355383 );
buf ( n355385 , n354203 );
not ( n355386 , n355385 );
buf ( n355387 , n355386 );
buf ( n355388 , n355387 );
nand ( n355389 , n35351 , n355388 );
buf ( n355390 , n355389 );
buf ( n355391 , n355390 );
and ( n35359 , n355382 , n355391 );
not ( n355393 , n354126 );
nor ( n35361 , n355393 , n355387 );
buf ( n355395 , n35361 );
nor ( n355396 , n35359 , n355395 );
buf ( n355397 , n355396 );
buf ( n355398 , n355397 );
xor ( n355399 , n355381 , n355398 );
and ( n355400 , n355170 , n355123 );
not ( n35368 , n355170 );
and ( n355402 , n35368 , n35091 );
nor ( n355403 , n355400 , n355402 );
not ( n35371 , n35073 );
and ( n35372 , n355403 , n35371 );
not ( n35373 , n355403 );
and ( n355407 , n35373 , n35073 );
nor ( n355408 , n35372 , n355407 );
buf ( n355409 , n355408 );
xor ( n35377 , n355399 , n355409 );
buf ( n355411 , n35377 );
nand ( n355412 , n35335 , n355411 );
buf ( n35380 , n355237 );
buf ( n355414 , n355300 );
xor ( n35382 , n35380 , n355414 );
buf ( n355416 , n35144 );
xnor ( n355417 , n35382 , n355416 );
buf ( n355418 , n355417 );
buf ( n355419 , n355418 );
xor ( n35387 , n355381 , n355398 );
and ( n355421 , n35387 , n355409 );
and ( n355422 , n355381 , n355398 );
or ( n355423 , n355421 , n355422 );
buf ( n355424 , n355423 );
buf ( n355425 , n355424 );
nand ( n355426 , n355419 , n355425 );
buf ( n355427 , n355426 );
nand ( n35395 , n355412 , n355427 );
not ( n355429 , n35395 );
nand ( n35397 , n35328 , n355429 );
nor ( n35398 , n355096 , n35397 );
and ( n355432 , n354740 , n35398 );
buf ( n355433 , n354657 );
not ( n35401 , n355433 );
buf ( n355435 , n35401 );
buf ( n355436 , n354711 );
not ( n355437 , n355436 );
buf ( n355438 , n355437 );
nand ( n355439 , n355435 , n355438 );
buf ( n355440 , n355439 );
buf ( n355441 , n355427 );
and ( n35409 , n34637 , n354691 );
not ( n355443 , n34637 );
and ( n355444 , n355443 , n34659 );
nor ( n35412 , n35409 , n355444 );
xor ( n355446 , n354704 , n35412 );
not ( n355447 , n342111 );
not ( n35415 , n342060 );
or ( n35416 , n355447 , n35415 );
nand ( n355450 , n35416 , n342116 );
not ( n355451 , n355450 );
not ( n35419 , n22366 );
and ( n355453 , n355451 , n35419 );
buf ( n355454 , n355450 );
buf ( n355455 , n22366 );
nand ( n35423 , n355454 , n355455 );
buf ( n355457 , n35423 );
buf ( n355458 , n342130 );
and ( n355459 , n355457 , n355458 );
nor ( n35427 , n355453 , n355459 );
nor ( n355461 , n355446 , n35427 );
buf ( n355462 , n355461 );
and ( n35430 , n355440 , n355441 , n355462 );
buf ( n35431 , n35430 );
buf ( n355465 , n354643 );
buf ( n355466 , n354615 );
and ( n35434 , n355465 , n355466 );
buf ( n355468 , n35434 );
buf ( n355469 , n354456 );
buf ( n35437 , n355412 );
and ( n35438 , n355469 , n35437 );
buf ( n355472 , n35438 );
nand ( n35440 , n35431 , n355468 , n355472 , n35328 );
not ( n355474 , n35440 );
buf ( n355475 , n35062 );
and ( n35443 , n355474 , n355475 );
nor ( n35444 , n355432 , n35443 );
nand ( n35445 , n355343 , n355355 );
nand ( n355479 , n354643 , n35445 , n355340 );
nor ( n355480 , n355479 , n354618 );
not ( n35448 , n355439 );
nor ( n35449 , n35448 , n35395 );
nand ( n35450 , n355480 , n35449 );
not ( n355484 , n35450 );
buf ( n355485 , n355484 );
buf ( n355486 , n341900 );
not ( n35454 , n355486 );
buf ( n355488 , n341998 );
not ( n355489 , n355488 );
or ( n355490 , n35454 , n355489 );
nand ( n35458 , n355446 , n35427 );
buf ( n355492 , n35458 );
not ( n355493 , n355492 );
buf ( n355494 , n16358 );
buf ( n355495 , n342304 );
nand ( n35463 , n355494 , n355495 );
buf ( n355497 , n35463 );
buf ( n355498 , n355497 );
nor ( n355499 , n355493 , n355498 );
buf ( n355500 , n355499 );
buf ( n355501 , n355500 );
nand ( n35469 , n355490 , n355501 );
buf ( n355503 , n35469 );
buf ( n35471 , n355503 );
not ( n35472 , n342304 );
buf ( n355506 , n16361 );
not ( n355507 , n355506 );
buf ( n355508 , n355507 );
not ( n35476 , n355508 );
or ( n35477 , n35472 , n35476 );
nand ( n35478 , n35477 , n342315 );
buf ( n355512 , n35458 );
not ( n35480 , n355512 );
buf ( n355514 , n35480 );
not ( n355515 , n355514 );
nand ( n35483 , n35478 , n355515 );
buf ( n355517 , n35483 );
nand ( n35485 , n35471 , n355517 );
buf ( n355519 , n35485 );
not ( n355520 , n35478 );
not ( n355521 , n22078 );
nand ( n35489 , n355520 , n22728 , n355521 );
and ( n355523 , n355519 , n35489 , n35062 );
buf ( n355524 , n355523 );
nand ( n355525 , n355485 , n355524 );
buf ( n355526 , n355525 );
or ( n35494 , n355424 , n355418 );
not ( n355528 , n355411 );
nand ( n35496 , n355528 , n355367 );
nand ( n355530 , n35494 , n35496 );
not ( n35498 , n355530 );
buf ( n355532 , n355427 );
buf ( n355533 , n355340 );
nand ( n35501 , n355532 , n355533 );
buf ( n35502 , n35501 );
nand ( n355536 , n355343 , n355355 );
not ( n35504 , n355536 );
nor ( n35505 , n35502 , n35504 );
not ( n35506 , n35505 );
or ( n355540 , n35498 , n35506 );
or ( n355541 , n355337 , n355313 );
not ( n35509 , n355343 );
not ( n35510 , n355355 );
nand ( n355544 , n35509 , n35510 );
and ( n355545 , n355541 , n355544 );
nor ( n35513 , n355545 , n35504 );
not ( n35514 , n35513 );
nand ( n35515 , n355540 , n35514 );
nand ( n355549 , n35515 , n355475 );
buf ( n35517 , n355090 );
not ( n35518 , n35517 );
buf ( n355552 , n35518 );
buf ( n355553 , n355552 );
buf ( n355554 , n355083 );
not ( n355555 , n355554 );
buf ( n355556 , n355555 );
buf ( n355557 , n355556 );
nand ( n35525 , n355553 , n355557 );
buf ( n355559 , n35525 );
buf ( n355560 , n355559 );
nor ( n355561 , n354742 , n34942 );
buf ( n355562 , n355561 );
or ( n35530 , n355560 , n355562 );
nand ( n35531 , n354742 , n34942 );
buf ( n355565 , n35531 );
nand ( n355566 , n35530 , n355565 );
buf ( n355567 , n355566 );
buf ( n355568 , n355567 );
not ( n35536 , n355568 );
buf ( n355570 , n35536 );
nand ( n355571 , n35444 , n355526 , n355549 , n355570 );
not ( n35539 , n355571 );
or ( n35540 , n33334 , n35539 );
not ( n35541 , n355570 );
nor ( n355575 , n35541 , n353366 );
nand ( n355576 , n35444 , n355526 , n355549 , n355575 );
nand ( n35544 , n35540 , n355576 );
buf ( n355578 , n35544 );
not ( n355579 , n355578 );
buf ( n35547 , n355579 );
not ( n35548 , n35547 );
buf ( n355582 , n35548 );
buf ( n35550 , n592 );
buf ( n355584 , n334531 );
buf ( n35552 , n355584 );
buf ( n355586 , n35552 );
buf ( n355587 , n355586 );
and ( n35555 , n35550 , n355587 );
buf ( n355589 , n35555 );
not ( n35557 , n355589 );
buf ( n355591 , n352036 );
buf ( n355592 , n355591 );
buf ( n355593 , n355592 );
buf ( n355594 , n355593 );
not ( n35562 , n355594 );
buf ( n355596 , n35562 );
buf ( n355597 , n355596 );
not ( n35565 , n355597 );
buf ( n355599 , n35565 );
buf ( n355600 , n355599 );
buf ( n355601 , n592 );
nand ( n35569 , n355600 , n355601 );
buf ( n355603 , n35569 );
buf ( n355604 , n355603 );
not ( n35572 , n355604 );
buf ( n355606 , n35572 );
buf ( n355607 , n355606 );
not ( n355608 , n355607 );
buf ( n355609 , n592 );
buf ( n355610 , n334537 );
not ( n35578 , n355610 );
buf ( n355612 , n35578 );
buf ( n355613 , n355612 );
not ( n355614 , n355613 );
buf ( n355615 , n355614 );
buf ( n355616 , n355615 );
and ( n35584 , n355609 , n355616 );
buf ( n35585 , n35584 );
buf ( n355619 , n35585 );
not ( n35587 , n355619 );
or ( n355621 , n355608 , n35587 );
buf ( n355622 , n355603 );
not ( n35590 , n355622 );
buf ( n35591 , n35585 );
not ( n355625 , n35591 );
buf ( n355626 , n355625 );
buf ( n355627 , n355626 );
not ( n355628 , n355627 );
or ( n35596 , n35590 , n355628 );
xor ( n355630 , n35550 , n355587 );
buf ( n355631 , n355630 );
buf ( n355632 , n355631 );
buf ( n355633 , n23613 );
not ( n355634 , n355633 );
buf ( n355635 , n344705 );
not ( n355636 , n355635 );
buf ( n355637 , n355636 );
buf ( n355638 , n355637 );
nand ( n35606 , n355634 , n355638 );
buf ( n355640 , n35606 );
buf ( n355641 , n355640 );
and ( n35609 , n355632 , n355641 );
buf ( n355643 , n35609 );
buf ( n355644 , n355643 );
not ( n35612 , n355644 );
buf ( n35613 , n35612 );
buf ( n35614 , n35613 );
nand ( n35615 , n35596 , n35614 );
buf ( n35616 , n35615 );
buf ( n355650 , n35616 );
nand ( n35618 , n355621 , n355650 );
buf ( n355652 , n35618 );
not ( n355653 , n355652 );
not ( n355654 , n355653 );
or ( n35622 , n35557 , n355654 );
buf ( n355656 , n592 );
buf ( n355657 , n344618 );
and ( n35625 , n355656 , n355657 );
buf ( n355659 , n35625 );
buf ( n355660 , n355659 );
buf ( n355661 , n343863 );
buf ( n355662 , n23889 );
or ( n35630 , n355661 , n355662 );
buf ( n355664 , n596 );
not ( n355665 , n355664 );
buf ( n355666 , n355586 );
not ( n35634 , n355666 );
buf ( n355668 , n35634 );
buf ( n355669 , n355668 );
not ( n35637 , n355669 );
or ( n35638 , n355665 , n35637 );
buf ( n355672 , n355586 );
buf ( n355673 , n343882 );
nand ( n35641 , n355672 , n355673 );
buf ( n355675 , n35641 );
buf ( n355676 , n355675 );
nand ( n35644 , n35638 , n355676 );
buf ( n35645 , n35644 );
buf ( n355679 , n35645 );
nand ( n35647 , n35630 , n355679 );
buf ( n355681 , n35647 );
buf ( n355682 , n355681 );
xor ( n35650 , n355660 , n355682 );
buf ( n355684 , n23613 );
not ( n355685 , n355684 );
buf ( n355686 , n351424 );
buf ( n355687 , n592 );
xor ( n355688 , n355686 , n355687 );
buf ( n355689 , n355688 );
buf ( n355690 , n355689 );
not ( n35658 , n355690 );
or ( n35659 , n355685 , n35658 );
buf ( n355693 , n592 );
not ( n355694 , n355693 );
buf ( n355695 , n350850 );
not ( n35663 , n355695 );
buf ( n355697 , n35663 );
buf ( n355698 , n355697 );
not ( n35666 , n355698 );
or ( n355700 , n355694 , n35666 );
buf ( n35668 , n355697 );
not ( n35669 , n35668 );
buf ( n35670 , n35669 );
buf ( n355704 , n35670 );
buf ( n355705 , n343624 );
nand ( n355706 , n355704 , n355705 );
buf ( n355707 , n355706 );
buf ( n355708 , n355707 );
nand ( n35676 , n355700 , n355708 );
buf ( n355710 , n35676 );
buf ( n355711 , n355710 );
buf ( n355712 , n344705 );
nand ( n355713 , n355711 , n355712 );
buf ( n355714 , n355713 );
buf ( n355715 , n355714 );
nand ( n35683 , n35659 , n355715 );
buf ( n355717 , n35683 );
buf ( n355718 , n355717 );
and ( n355719 , n35650 , n355718 );
and ( n35687 , n355660 , n355682 );
or ( n355721 , n355719 , n35687 );
buf ( n355722 , n355721 );
buf ( n355723 , n355722 );
not ( n35691 , n355723 );
buf ( n355725 , n343765 );
not ( n35693 , n355725 );
buf ( n355727 , n343632 );
buf ( n35695 , n355615 );
not ( n355729 , n35695 );
buf ( n355730 , n355729 );
buf ( n355731 , n355730 );
and ( n355732 , n355727 , n355731 );
not ( n355733 , n355727 );
buf ( n355734 , n355615 );
and ( n35702 , n355733 , n355734 );
nor ( n355736 , n355732 , n35702 );
buf ( n355737 , n355736 );
buf ( n355738 , n355737 );
not ( n355739 , n355738 );
or ( n35707 , n35693 , n355739 );
buf ( n355741 , n594 );
not ( n35709 , n355741 );
buf ( n355743 , n355668 );
not ( n35711 , n355743 );
or ( n35712 , n35709 , n35711 );
buf ( n35713 , n355586 );
buf ( n355747 , n343632 );
nand ( n355748 , n35713 , n355747 );
buf ( n355749 , n355748 );
buf ( n355750 , n355749 );
nand ( n35718 , n35712 , n355750 );
buf ( n355752 , n35718 );
buf ( n355753 , n355752 );
buf ( n355754 , n23681 );
nand ( n355755 , n355753 , n355754 );
buf ( n355756 , n355755 );
buf ( n355757 , n355756 );
nand ( n355758 , n35707 , n355757 );
buf ( n355759 , n355758 );
buf ( n35727 , n35670 );
buf ( n35728 , n592 );
nand ( n35729 , n35727 , n35728 );
buf ( n35730 , n35729 );
buf ( n355764 , n35730 );
not ( n35732 , n355764 );
buf ( n355766 , n23613 );
not ( n355767 , n355766 );
buf ( n355768 , n592 );
not ( n355769 , n355768 );
buf ( n355770 , n355596 );
not ( n35738 , n355770 );
or ( n35739 , n355769 , n35738 );
buf ( n355773 , n355599 );
buf ( n355774 , n343624 );
nand ( n35742 , n355773 , n355774 );
buf ( n355776 , n35742 );
buf ( n355777 , n355776 );
nand ( n35745 , n35739 , n355777 );
buf ( n355779 , n35745 );
buf ( n355780 , n355779 );
not ( n35748 , n355780 );
or ( n35749 , n355767 , n35748 );
buf ( n355783 , n344705 );
buf ( n355784 , n355689 );
nand ( n35752 , n355783 , n355784 );
buf ( n355786 , n35752 );
buf ( n355787 , n355786 );
nand ( n35755 , n35749 , n355787 );
buf ( n35756 , n35755 );
buf ( n355790 , n35756 );
not ( n35758 , n355790 );
buf ( n355792 , n35758 );
buf ( n355793 , n355792 );
not ( n35761 , n355793 );
or ( n35762 , n35732 , n35761 );
buf ( n355796 , n35756 );
buf ( n355797 , n35730 );
not ( n35765 , n355797 );
buf ( n355799 , n35765 );
buf ( n355800 , n355799 );
nand ( n35768 , n355796 , n355800 );
buf ( n355802 , n35768 );
buf ( n355803 , n355802 );
nand ( n355804 , n35762 , n355803 );
buf ( n355805 , n355804 );
xnor ( n355806 , n355759 , n355805 );
not ( n35774 , n355806 );
buf ( n355808 , n35774 );
not ( n355809 , n355808 );
or ( n35777 , n35691 , n355809 );
buf ( n355811 , n23613 );
not ( n355812 , n355811 );
buf ( n355813 , n355710 );
not ( n35781 , n355813 );
or ( n355815 , n355812 , n35781 );
xor ( n35783 , n355656 , n355657 );
buf ( n355817 , n35783 );
buf ( n355818 , n355817 );
buf ( n355819 , n344705 );
nand ( n355820 , n355818 , n355819 );
buf ( n355821 , n355820 );
buf ( n355822 , n355821 );
nand ( n355823 , n355815 , n355822 );
buf ( n355824 , n355823 );
buf ( n355825 , n355824 );
buf ( n355826 , n23681 );
not ( n355827 , n355826 );
buf ( n355828 , n355737 );
not ( n35796 , n355828 );
or ( n355830 , n355827 , n35796 );
buf ( n355831 , n594 );
not ( n35799 , n355831 );
buf ( n355833 , n355596 );
not ( n355834 , n355833 );
or ( n355835 , n35799 , n355834 );
buf ( n355836 , n355593 );
buf ( n35804 , n355836 );
buf ( n35805 , n35804 );
buf ( n355839 , n35805 );
buf ( n355840 , n343632 );
nand ( n355841 , n355839 , n355840 );
buf ( n355842 , n355841 );
buf ( n355843 , n355842 );
nand ( n35811 , n355835 , n355843 );
buf ( n355845 , n35811 );
buf ( n355846 , n355845 );
buf ( n355847 , n343765 );
nand ( n355848 , n355846 , n355847 );
buf ( n355849 , n355848 );
buf ( n355850 , n355849 );
nand ( n355851 , n355830 , n355850 );
buf ( n355852 , n355851 );
buf ( n355853 , n355852 );
xor ( n355854 , n355825 , n355853 );
xor ( n35822 , n355660 , n355682 );
xor ( n355856 , n35822 , n355718 );
buf ( n355857 , n355856 );
buf ( n355858 , n355857 );
and ( n355859 , n355854 , n355858 );
and ( n355860 , n355825 , n355853 );
or ( n35828 , n355859 , n355860 );
buf ( n355862 , n35828 );
buf ( n355863 , n355862 );
buf ( n355864 , n355806 );
buf ( n355865 , n355722 );
not ( n355866 , n355865 );
buf ( n355867 , n355866 );
buf ( n355868 , n355867 );
nand ( n35836 , n355864 , n355868 );
buf ( n355870 , n35836 );
buf ( n355871 , n355870 );
nand ( n35839 , n355863 , n355871 );
buf ( n355873 , n35839 );
buf ( n355874 , n355873 );
nand ( n355875 , n35777 , n355874 );
buf ( n355876 , n355875 );
buf ( n355877 , n355799 );
buf ( n355878 , n35730 );
not ( n35846 , n355878 );
buf ( n355880 , n35756 );
not ( n355881 , n355880 );
or ( n35849 , n35846 , n355881 );
buf ( n355883 , n355799 );
not ( n355884 , n355883 );
buf ( n355885 , n355792 );
not ( n355886 , n355885 );
or ( n355887 , n355884 , n355886 );
buf ( n355888 , n355759 );
nand ( n355889 , n355887 , n355888 );
buf ( n355890 , n355889 );
buf ( n355891 , n355890 );
nand ( n355892 , n35849 , n355891 );
buf ( n355893 , n355892 );
buf ( n355894 , n355893 );
xor ( n355895 , n355877 , n355894 );
and ( n35863 , n355686 , n355687 );
buf ( n355897 , n35863 );
buf ( n355898 , n355897 );
buf ( n355899 , n23680 );
not ( n355900 , n355899 );
buf ( n355901 , n24631 );
not ( n35869 , n355901 );
or ( n35870 , n355900 , n35869 );
buf ( n355904 , n355752 );
nand ( n355905 , n35870 , n355904 );
buf ( n355906 , n355905 );
buf ( n355907 , n355906 );
xor ( n355908 , n355898 , n355907 );
buf ( n355909 , n23613 );
not ( n355910 , n355909 );
xor ( n355911 , n355609 , n355616 );
buf ( n355912 , n355911 );
buf ( n355913 , n355912 );
not ( n355914 , n355913 );
or ( n35879 , n355910 , n355914 );
buf ( n355916 , n355779 );
buf ( n355917 , n344705 );
nand ( n35882 , n355916 , n355917 );
buf ( n355919 , n35882 );
buf ( n355920 , n355919 );
nand ( n355921 , n35879 , n355920 );
buf ( n355922 , n355921 );
buf ( n355923 , n355922 );
xor ( n35888 , n355908 , n355923 );
buf ( n35889 , n35888 );
buf ( n355926 , n35889 );
xor ( n35891 , n355895 , n355926 );
buf ( n355928 , n35891 );
nor ( n35893 , n355876 , n355928 );
buf ( n355930 , n35893 );
xor ( n35895 , n355877 , n355894 );
and ( n355932 , n35895 , n355926 );
and ( n355933 , n355877 , n355894 );
or ( n35898 , n355932 , n355933 );
buf ( n355935 , n35898 );
buf ( n355936 , n355935 );
buf ( n355937 , n355603 );
buf ( n355938 , n344705 );
not ( n35903 , n355938 );
buf ( n355940 , n355912 );
not ( n35905 , n355940 );
or ( n355942 , n35903 , n35905 );
buf ( n355943 , n355631 );
buf ( n355944 , n23613 );
nand ( n35909 , n355943 , n355944 );
buf ( n355946 , n35909 );
buf ( n355947 , n355946 );
nand ( n355948 , n355942 , n355947 );
buf ( n355949 , n355948 );
buf ( n355950 , n355949 );
xor ( n355951 , n355937 , n355950 );
xor ( n355952 , n355898 , n355907 );
and ( n35917 , n355952 , n355923 );
and ( n355954 , n355898 , n355907 );
or ( n355955 , n35917 , n355954 );
buf ( n355956 , n355955 );
buf ( n355957 , n355956 );
xor ( n355958 , n355951 , n355957 );
buf ( n355959 , n355958 );
buf ( n355960 , n355959 );
nor ( n355961 , n355936 , n355960 );
buf ( n355962 , n355961 );
buf ( n355963 , n355962 );
nor ( n355964 , n355930 , n355963 );
buf ( n355965 , n355964 );
buf ( n355966 , n355965 );
not ( n35931 , n355966 );
xor ( n355968 , n355937 , n355950 );
and ( n355969 , n355968 , n355957 );
and ( n35934 , n355937 , n355950 );
or ( n355971 , n355969 , n35934 );
buf ( n355972 , n355971 );
buf ( n355973 , n355972 );
not ( n355974 , n355973 );
buf ( n355975 , n355606 );
buf ( n355976 , n35585 );
xor ( n355977 , n355975 , n355976 );
buf ( n355978 , n355643 );
xor ( n355979 , n355977 , n355978 );
buf ( n355980 , n355979 );
buf ( n355981 , n355980 );
nand ( n355982 , n355974 , n355981 );
buf ( n355983 , n355982 );
buf ( n355984 , n355983 );
not ( n355985 , n355984 );
buf ( n355986 , n355985 );
buf ( n355987 , n355986 );
nor ( n355988 , n35931 , n355987 );
buf ( n355989 , n355988 );
not ( n35954 , n355989 );
not ( n355991 , n350815 );
buf ( n355992 , n355991 );
and ( n35957 , n592 , n355992 );
buf ( n355994 , n35957 );
not ( n355995 , n355994 );
buf ( n355996 , n23889 );
not ( n35961 , n355996 );
buf ( n355998 , n596 );
not ( n35963 , n355998 );
buf ( n356000 , n355730 );
not ( n356001 , n356000 );
or ( n35966 , n35963 , n356001 );
buf ( n356003 , n355615 );
buf ( n356004 , n343882 );
nand ( n35969 , n356003 , n356004 );
buf ( n356006 , n35969 );
buf ( n356007 , n356006 );
nand ( n35972 , n35966 , n356007 );
buf ( n356009 , n35972 );
buf ( n35974 , n356009 );
not ( n35975 , n35974 );
or ( n35976 , n35961 , n35975 );
buf ( n35977 , n35645 );
buf ( n356014 , n343863 );
nand ( n356015 , n35977 , n356014 );
buf ( n356016 , n356015 );
buf ( n356017 , n356016 );
nand ( n35982 , n35976 , n356017 );
buf ( n35983 , n35982 );
buf ( n356020 , n35983 );
not ( n35985 , n356020 );
or ( n356022 , n355995 , n35985 );
buf ( n356023 , n35983 );
buf ( n356024 , n35957 );
or ( n35989 , n356023 , n356024 );
buf ( n35990 , n23681 );
not ( n35991 , n35990 );
buf ( n356028 , n355845 );
not ( n35993 , n356028 );
or ( n35994 , n35991 , n35993 );
buf ( n356031 , n594 );
not ( n35996 , n356031 );
buf ( n356033 , n351427 );
not ( n35998 , n356033 );
or ( n35999 , n35996 , n35998 );
buf ( n356036 , n351424 );
buf ( n356037 , n343632 );
nand ( n36002 , n356036 , n356037 );
buf ( n356039 , n36002 );
buf ( n356040 , n356039 );
nand ( n356041 , n35999 , n356040 );
buf ( n356042 , n356041 );
buf ( n356043 , n356042 );
buf ( n356044 , n343765 );
nand ( n36009 , n356043 , n356044 );
buf ( n356046 , n36009 );
buf ( n356047 , n356046 );
nand ( n36012 , n35994 , n356047 );
buf ( n356049 , n36012 );
buf ( n356050 , n356049 );
nand ( n36015 , n35989 , n356050 );
buf ( n356052 , n36015 );
buf ( n356053 , n356052 );
nand ( n36018 , n356022 , n356053 );
buf ( n356055 , n36018 );
buf ( n356056 , n356055 );
not ( n36021 , n356056 );
xor ( n36022 , n355825 , n355853 );
xor ( n36023 , n36022 , n355858 );
buf ( n356060 , n36023 );
buf ( n36025 , n356060 );
not ( n356062 , n36025 );
buf ( n356063 , n356062 );
buf ( n356064 , n356063 );
not ( n36029 , n356064 );
or ( n356066 , n36021 , n36029 );
buf ( n356067 , n356060 );
buf ( n356068 , n356055 );
not ( n356069 , n356068 );
buf ( n356070 , n356069 );
buf ( n356071 , n356070 );
nand ( n356072 , n356067 , n356071 );
buf ( n356073 , n356072 );
buf ( n356074 , n356073 );
nand ( n356075 , n356066 , n356074 );
buf ( n356076 , n356075 );
buf ( n356077 , n356076 );
not ( n356078 , n355824 );
buf ( n356079 , n592 );
buf ( n356080 , n345097 );
and ( n356081 , n356079 , n356080 );
buf ( n356082 , n356081 );
buf ( n356083 , n356082 );
buf ( n36048 , n23911 );
not ( n356085 , n36048 );
buf ( n356086 , n356085 );
buf ( n356087 , n356086 );
not ( n356088 , n356087 );
buf ( n356089 , n343948 );
not ( n356090 , n356089 );
buf ( n356091 , n356090 );
buf ( n356092 , n356091 );
not ( n356093 , n356092 );
or ( n356094 , n356088 , n356093 );
and ( n36059 , n355586 , n343953 );
not ( n356096 , n355586 );
and ( n356097 , n356096 , n598 );
or ( n36062 , n36059 , n356097 );
buf ( n356099 , n36062 );
nand ( n356100 , n356094 , n356099 );
buf ( n356101 , n356100 );
buf ( n356102 , n356101 );
xor ( n36067 , n356083 , n356102 );
buf ( n356104 , n23681 );
not ( n36069 , n356104 );
buf ( n356106 , n356042 );
not ( n356107 , n356106 );
or ( n36072 , n36069 , n356107 );
not ( n356109 , n594 );
not ( n356110 , n355697 );
or ( n36075 , n356109 , n356110 );
buf ( n356112 , n35670 );
buf ( n356113 , n343632 );
nand ( n36078 , n356112 , n356113 );
buf ( n356115 , n36078 );
nand ( n36080 , n36075 , n356115 );
buf ( n356117 , n36080 );
buf ( n356118 , n343765 );
nand ( n36083 , n356117 , n356118 );
buf ( n356120 , n36083 );
buf ( n356121 , n356120 );
nand ( n356122 , n36072 , n356121 );
buf ( n356123 , n356122 );
buf ( n356124 , n356123 );
and ( n356125 , n36067 , n356124 );
and ( n356126 , n356083 , n356102 );
or ( n36091 , n356125 , n356126 );
buf ( n356128 , n36091 );
buf ( n356129 , n356128 );
not ( n36094 , n356129 );
buf ( n36095 , n36094 );
not ( n356132 , n36095 );
or ( n36097 , n356078 , n356132 );
nor ( n356134 , n355824 , n36095 );
not ( n356135 , n356049 );
xor ( n36100 , n35957 , n356135 );
xnor ( n356137 , n36100 , n35983 );
or ( n356138 , n356134 , n356137 );
nand ( n36103 , n36097 , n356138 );
buf ( n356140 , n36103 );
and ( n356141 , n356077 , n356140 );
not ( n36106 , n356077 );
not ( n356143 , n36103 );
buf ( n36108 , n356143 );
and ( n36109 , n36106 , n36108 );
nor ( n356146 , n356141 , n36109 );
buf ( n356147 , n356146 );
buf ( n356148 , n356147 );
buf ( n356149 , n344436 );
not ( n356150 , n356149 );
buf ( n356151 , n592 );
nand ( n356152 , n356150 , n356151 );
buf ( n356153 , n356152 );
buf ( n356154 , n356153 );
not ( n356155 , n356154 );
buf ( n36120 , n343863 );
not ( n36121 , n36120 );
buf ( n356158 , n356009 );
not ( n36123 , n356158 );
or ( n356160 , n36121 , n36123 );
buf ( n356161 , n596 );
not ( n36126 , n356161 );
buf ( n356163 , n355596 );
not ( n36128 , n356163 );
or ( n356165 , n36126 , n36128 );
buf ( n36130 , n35805 );
buf ( n356167 , n343882 );
nand ( n36132 , n36130 , n356167 );
buf ( n356169 , n36132 );
buf ( n356170 , n356169 );
nand ( n36135 , n356165 , n356170 );
buf ( n356172 , n36135 );
buf ( n356173 , n356172 );
buf ( n356174 , n23889 );
nand ( n36139 , n356173 , n356174 );
buf ( n356176 , n36139 );
buf ( n356177 , n356176 );
nand ( n356178 , n356160 , n356177 );
buf ( n356179 , n356178 );
buf ( n356180 , n356179 );
not ( n356181 , n356180 );
buf ( n356182 , n356181 );
buf ( n356183 , n356182 );
not ( n356184 , n356183 );
or ( n356185 , n356155 , n356184 );
buf ( n356186 , n344705 );
not ( n356187 , n356186 );
xor ( n356188 , n592 , n355992 );
buf ( n356189 , n356188 );
not ( n356190 , n356189 );
or ( n356191 , n356187 , n356190 );
buf ( n36156 , n355817 );
buf ( n36157 , n23613 );
nand ( n36158 , n36156 , n36157 );
buf ( n36159 , n36158 );
buf ( n356196 , n36159 );
nand ( n36161 , n356191 , n356196 );
buf ( n356198 , n36161 );
buf ( n356199 , n356198 );
nand ( n36164 , n356185 , n356199 );
buf ( n356201 , n36164 );
buf ( n356202 , n356201 );
buf ( n356203 , n356153 );
not ( n36168 , n356203 );
buf ( n356205 , n356179 );
nand ( n356206 , n36168 , n356205 );
buf ( n356207 , n356206 );
buf ( n356208 , n356207 );
nand ( n36173 , n356202 , n356208 );
buf ( n356210 , n36173 );
buf ( n356211 , n356210 );
not ( n36176 , n356211 );
xor ( n36177 , n355824 , n36095 );
xnor ( n36178 , n36177 , n356137 );
buf ( n356215 , n36178 );
nand ( n356216 , n36176 , n356215 );
buf ( n356217 , n356216 );
buf ( n356218 , n343863 );
not ( n356219 , n356218 );
buf ( n356220 , n356172 );
not ( n356221 , n356220 );
or ( n356222 , n356219 , n356221 );
buf ( n356223 , n596 );
not ( n36188 , n356223 );
buf ( n356225 , n351427 );
not ( n36190 , n356225 );
or ( n356227 , n36188 , n36190 );
buf ( n36192 , n351424 );
buf ( n356229 , n343882 );
nand ( n356230 , n36192 , n356229 );
buf ( n356231 , n356230 );
buf ( n356232 , n356231 );
nand ( n356233 , n356227 , n356232 );
buf ( n356234 , n356233 );
buf ( n356235 , n356234 );
buf ( n356236 , n23889 );
nand ( n36201 , n356235 , n356236 );
buf ( n356238 , n36201 );
buf ( n356239 , n356238 );
nand ( n36204 , n356222 , n356239 );
buf ( n36205 , n36204 );
not ( n356242 , n36205 );
nand ( n36207 , n356242 , n356082 );
not ( n356244 , n36207 );
not ( n356245 , n343765 );
buf ( n356246 , n594 );
not ( n356247 , n356246 );
buf ( n356248 , n24586 );
not ( n36213 , n356248 );
or ( n356250 , n356247 , n36213 );
buf ( n356251 , n344618 );
buf ( n356252 , n343632 );
nand ( n36217 , n356251 , n356252 );
buf ( n356254 , n36217 );
buf ( n356255 , n356254 );
nand ( n356256 , n356250 , n356255 );
buf ( n356257 , n356256 );
not ( n36222 , n356257 );
or ( n356259 , n356245 , n36222 );
nand ( n36224 , n36080 , n23681 );
nand ( n356261 , n356259 , n36224 );
not ( n36226 , n356261 );
or ( n36227 , n356244 , n36226 );
buf ( n356264 , n36205 );
buf ( n356265 , n356082 );
not ( n36230 , n356265 );
buf ( n356267 , n36230 );
buf ( n356268 , n356267 );
nand ( n36233 , n356264 , n356268 );
buf ( n356270 , n36233 );
nand ( n36235 , n36227 , n356270 );
not ( n36236 , n36235 );
buf ( n356273 , n356153 );
buf ( n356274 , n356198 );
xor ( n356275 , n356273 , n356274 );
buf ( n356276 , n356179 );
xnor ( n356277 , n356275 , n356276 );
buf ( n356278 , n356277 );
xor ( n36243 , n356083 , n356102 );
xor ( n356280 , n36243 , n356124 );
buf ( n356281 , n356280 );
or ( n36246 , n356278 , n356281 );
not ( n356283 , n36246 );
or ( n36248 , n36236 , n356283 );
buf ( n356285 , n356278 );
buf ( n356286 , n356281 );
nand ( n356287 , n356285 , n356286 );
buf ( n356288 , n356287 );
nand ( n356289 , n36248 , n356288 );
and ( n356290 , n356217 , n356289 );
buf ( n356291 , n356210 );
not ( n356292 , n356291 );
buf ( n356293 , n36178 );
nor ( n36258 , n356292 , n356293 );
buf ( n36259 , n36258 );
nor ( n356296 , n356290 , n36259 );
buf ( n356297 , n356296 );
nand ( n356298 , n356148 , n356297 );
buf ( n356299 , n356298 );
not ( n36264 , n356299 );
not ( n356301 , n356143 );
buf ( n356302 , n356063 );
buf ( n356303 , n356070 );
nand ( n36268 , n356302 , n356303 );
buf ( n356305 , n36268 );
not ( n356306 , n356305 );
or ( n36271 , n356301 , n356306 );
nand ( n356308 , n356055 , n356060 );
nand ( n356309 , n36271 , n356308 );
not ( n36274 , n356309 );
not ( n356311 , n355867 );
not ( n36276 , n35774 );
or ( n36277 , n356311 , n36276 );
buf ( n356314 , n355806 );
buf ( n356315 , n355722 );
nand ( n356316 , n356314 , n356315 );
buf ( n356317 , n356316 );
nand ( n356318 , n36277 , n356317 );
xnor ( n36283 , n356318 , n355862 );
nand ( n356320 , n36274 , n36283 );
not ( n36285 , n356320 );
nor ( n356322 , n36264 , n36285 );
buf ( n356323 , n23613 );
not ( n36288 , n356323 );
buf ( n356325 , n356188 );
not ( n36290 , n356325 );
or ( n356327 , n36288 , n36290 );
buf ( n356328 , n592 );
not ( n36293 , n356328 );
buf ( n356330 , n344436 );
not ( n36295 , n356330 );
or ( n36296 , n36293 , n36295 );
buf ( n356333 , n344435 );
not ( n36298 , n356333 );
buf ( n356335 , n343624 );
nand ( n36300 , n36298 , n356335 );
buf ( n356337 , n36300 );
buf ( n356338 , n356337 );
nand ( n356339 , n36296 , n356338 );
buf ( n356340 , n356339 );
buf ( n356341 , n356340 );
buf ( n356342 , n344705 );
nand ( n356343 , n356341 , n356342 );
buf ( n356344 , n356343 );
buf ( n356345 , n356344 );
nand ( n356346 , n356327 , n356345 );
buf ( n356347 , n356346 );
buf ( n356348 , n356347 );
not ( n356349 , n356348 );
buf ( n356350 , n343948 );
not ( n356351 , n356350 );
buf ( n356352 , n598 );
not ( n36317 , n356352 );
buf ( n356354 , n355730 );
not ( n356355 , n356354 );
or ( n356356 , n36317 , n356355 );
buf ( n356357 , n355615 );
buf ( n356358 , n343953 );
nand ( n356359 , n356357 , n356358 );
buf ( n356360 , n356359 );
buf ( n356361 , n356360 );
nand ( n36326 , n356356 , n356361 );
buf ( n356363 , n36326 );
buf ( n356364 , n356363 );
not ( n36329 , n356364 );
or ( n356366 , n356351 , n36329 );
buf ( n356367 , n36062 );
buf ( n356368 , n23911 );
nand ( n36333 , n356367 , n356368 );
buf ( n356370 , n36333 );
buf ( n356371 , n356370 );
nand ( n36336 , n356366 , n356371 );
buf ( n356373 , n36336 );
buf ( n356374 , n356373 );
not ( n356375 , n356374 );
or ( n356376 , n356349 , n356375 );
buf ( n356377 , n356347 );
buf ( n356378 , n356373 );
or ( n36340 , n356377 , n356378 );
buf ( n356380 , n23613 );
not ( n356381 , n356380 );
xor ( n36343 , n356079 , n356080 );
buf ( n356383 , n36343 );
buf ( n356384 , n356383 );
not ( n36346 , n356384 );
or ( n356386 , n356381 , n36346 );
buf ( n356387 , n592 );
not ( n356388 , n356387 );
buf ( n356389 , n344383 );
not ( n356390 , n356389 );
or ( n36352 , n356388 , n356390 );
buf ( n356392 , n24346 );
buf ( n356393 , n343624 );
nand ( n356394 , n356392 , n356393 );
buf ( n356395 , n356394 );
buf ( n356396 , n356395 );
nand ( n356397 , n36352 , n356396 );
buf ( n356398 , n356397 );
buf ( n356399 , n356398 );
buf ( n356400 , n344705 );
nand ( n356401 , n356399 , n356400 );
buf ( n356402 , n356401 );
buf ( n356403 , n356402 );
nand ( n356404 , n356386 , n356403 );
buf ( n356405 , n356404 );
buf ( n356406 , n356405 );
buf ( n356407 , n356406 );
buf ( n356408 , n356407 );
buf ( n36358 , n356408 );
not ( n36359 , n36358 );
buf ( n36360 , n36359 );
buf ( n36361 , n36360 );
buf ( n356413 , n24346 );
buf ( n356414 , n592 );
nand ( n356415 , n356413 , n356414 );
buf ( n356416 , n356415 );
buf ( n356417 , n356416 );
nand ( n36367 , n36361 , n356417 );
buf ( n356419 , n36367 );
buf ( n356420 , n356419 );
not ( n356421 , n356420 );
buf ( n356422 , n343863 );
not ( n36372 , n356422 );
buf ( n356424 , n356234 );
not ( n36374 , n356424 );
or ( n36375 , n36372 , n36374 );
buf ( n356427 , n596 );
not ( n36377 , n356427 );
buf ( n356429 , n350850 );
buf ( n36379 , n356429 );
buf ( n356431 , n36379 );
buf ( n356432 , n356431 );
not ( n356433 , n356432 );
buf ( n356434 , n356433 );
buf ( n356435 , n356434 );
not ( n36385 , n356435 );
or ( n36386 , n36377 , n36385 );
buf ( n356438 , n35670 );
buf ( n356439 , n343882 );
nand ( n36389 , n356438 , n356439 );
buf ( n356441 , n36389 );
buf ( n356442 , n356441 );
nand ( n36392 , n36386 , n356442 );
buf ( n356444 , n36392 );
buf ( n356445 , n356444 );
buf ( n356446 , n23889 );
nand ( n36396 , n356445 , n356446 );
buf ( n356448 , n36396 );
buf ( n356449 , n356448 );
nand ( n356450 , n36375 , n356449 );
buf ( n356451 , n356450 );
buf ( n356452 , n356451 );
not ( n356453 , n356452 );
or ( n356454 , n356421 , n356453 );
buf ( n356455 , n36360 );
buf ( n356456 , n356416 );
or ( n356457 , n356455 , n356456 );
buf ( n356458 , n356457 );
buf ( n356459 , n356458 );
nand ( n356460 , n356454 , n356459 );
buf ( n356461 , n356460 );
buf ( n356462 , n356461 );
nand ( n356463 , n36340 , n356462 );
buf ( n356464 , n356463 );
buf ( n356465 , n356464 );
nand ( n356466 , n356376 , n356465 );
buf ( n356467 , n356466 );
buf ( n356468 , n356467 );
buf ( n356469 , n36235 );
buf ( n356470 , n356281 );
xor ( n36417 , n356469 , n356470 );
buf ( n356472 , n356278 );
xnor ( n36419 , n36417 , n356472 );
buf ( n356474 , n36419 );
buf ( n356475 , n356474 );
xor ( n36422 , n356468 , n356475 );
buf ( n356477 , n23613 );
not ( n36424 , n356477 );
buf ( n356479 , n356340 );
not ( n36426 , n356479 );
or ( n356481 , n36424 , n36426 );
buf ( n36428 , n356383 );
buf ( n356483 , n344705 );
nand ( n356484 , n36428 , n356483 );
buf ( n356485 , n356484 );
buf ( n356486 , n356485 );
nand ( n36433 , n356481 , n356486 );
buf ( n356488 , n36433 );
not ( n356489 , n356488 );
buf ( n356490 , n344014 );
not ( n356491 , n356490 );
buf ( n356492 , n344017 );
not ( n36439 , n356492 );
or ( n356494 , n356491 , n36439 );
buf ( n356495 , n355586 );
not ( n356496 , n356495 );
buf ( n356497 , n23906 );
not ( n356498 , n356497 );
and ( n356499 , n356496 , n356498 );
buf ( n356500 , n355586 );
buf ( n356501 , n23906 );
and ( n356502 , n356500 , n356501 );
nor ( n36449 , n356499 , n356502 );
buf ( n36450 , n36449 );
buf ( n36451 , n36450 );
not ( n36452 , n36451 );
buf ( n36453 , n36452 );
buf ( n356508 , n36453 );
nand ( n36455 , n356494 , n356508 );
buf ( n36456 , n36455 );
not ( n356511 , n36456 );
or ( n36458 , n356489 , n356511 );
not ( n356513 , n356488 );
not ( n356514 , n356513 );
not ( n36461 , n36456 );
not ( n356516 , n36461 );
or ( n356517 , n356514 , n356516 );
buf ( n356518 , n343765 );
not ( n356519 , n356518 );
buf ( n356520 , n594 );
not ( n36467 , n356520 );
buf ( n356522 , n350815 );
not ( n36469 , n356522 );
or ( n36470 , n36467 , n36469 );
buf ( n356525 , n355991 );
buf ( n356526 , n343632 );
nand ( n36473 , n356525 , n356526 );
buf ( n356528 , n36473 );
buf ( n356529 , n356528 );
nand ( n36476 , n36470 , n356529 );
buf ( n36477 , n36476 );
buf ( n356532 , n36477 );
not ( n36479 , n356532 );
or ( n356534 , n356519 , n36479 );
buf ( n356535 , n356257 );
buf ( n356536 , n23681 );
nand ( n36483 , n356535 , n356536 );
buf ( n356538 , n36483 );
buf ( n356539 , n356538 );
nand ( n36486 , n356534 , n356539 );
buf ( n36487 , n36486 );
buf ( n356542 , n36487 );
nand ( n36489 , n356517 , n356542 );
nand ( n356544 , n36458 , n36489 );
not ( n36491 , n356544 );
xor ( n36492 , n356082 , n356261 );
xnor ( n356547 , n36492 , n36205 );
not ( n36494 , n356547 );
nand ( n356549 , n36491 , n36494 );
buf ( n356550 , n356549 );
not ( n36497 , n356550 );
buf ( n36498 , n356347 );
buf ( n356553 , n356373 );
xor ( n356554 , n36498 , n356553 );
buf ( n356555 , n356461 );
xnor ( n356556 , n356554 , n356555 );
buf ( n356557 , n356556 );
buf ( n356558 , n356557 );
not ( n36505 , n356558 );
buf ( n356560 , n36505 );
buf ( n356561 , n356560 );
not ( n36508 , n356561 );
or ( n356563 , n36497 , n36508 );
nand ( n356564 , n356544 , n356547 );
buf ( n356565 , n356564 );
nand ( n36512 , n356563 , n356565 );
buf ( n356567 , n36512 );
buf ( n356568 , n356567 );
xnor ( n36515 , n36422 , n356568 );
buf ( n36516 , n36515 );
buf ( n356571 , n36516 );
not ( n356572 , n356488 );
not ( n36519 , n36461 );
or ( n356574 , n356572 , n36519 );
nand ( n356575 , n36456 , n356513 );
nand ( n36522 , n356574 , n356575 );
not ( n356577 , n356542 );
and ( n36524 , n36522 , n356577 );
not ( n356579 , n36522 );
and ( n36526 , n356579 , n356542 );
nor ( n36527 , n36524 , n36526 );
buf ( n36528 , n36527 );
buf ( n356583 , n23681 );
not ( n356584 , n356583 );
buf ( n356585 , n36477 );
not ( n36532 , n356585 );
or ( n356587 , n356584 , n36532 );
buf ( n36534 , n594 );
not ( n36535 , n36534 );
buf ( n356590 , n344435 );
not ( n36537 , n356590 );
or ( n356592 , n36535 , n36537 );
buf ( n356593 , n24408 );
buf ( n36540 , n343632 );
nand ( n36541 , n356593 , n36540 );
buf ( n36542 , n36541 );
buf ( n356597 , n36542 );
nand ( n36544 , n356592 , n356597 );
buf ( n356599 , n36544 );
buf ( n356600 , n356599 );
buf ( n356601 , n343765 );
nand ( n36548 , n356600 , n356601 );
buf ( n356603 , n36548 );
buf ( n356604 , n356603 );
nand ( n36551 , n356587 , n356604 );
buf ( n356606 , n36551 );
not ( n36553 , n356606 );
not ( n36554 , n36553 );
not ( n36555 , n36554 );
buf ( n356610 , n23911 );
not ( n356611 , n356610 );
buf ( n356612 , n598 );
not ( n356613 , n356612 );
buf ( n356614 , n355596 );
not ( n36561 , n356614 );
or ( n356616 , n356613 , n36561 );
buf ( n36563 , n355593 );
buf ( n356618 , n343953 );
nand ( n356619 , n36563 , n356618 );
buf ( n356620 , n356619 );
buf ( n356621 , n356620 );
nand ( n356622 , n356616 , n356621 );
buf ( n356623 , n356622 );
buf ( n356624 , n356623 );
not ( n36571 , n356624 );
or ( n356626 , n356611 , n36571 );
buf ( n356627 , n598 );
not ( n356628 , n356627 );
buf ( n356629 , n351427 );
not ( n356630 , n356629 );
or ( n36577 , n356628 , n356630 );
not ( n356632 , n351417 );
not ( n356633 , n351412 );
or ( n36580 , n356632 , n356633 );
nand ( n356635 , n36580 , n351422 );
not ( n356636 , n356635 );
nand ( n36583 , n356636 , n343953 );
buf ( n356638 , n36583 );
nand ( n356639 , n36577 , n356638 );
buf ( n356640 , n356639 );
buf ( n356641 , n356640 );
buf ( n356642 , n343948 );
nand ( n36589 , n356641 , n356642 );
buf ( n356644 , n36589 );
buf ( n356645 , n356644 );
nand ( n36592 , n356626 , n356645 );
buf ( n356647 , n36592 );
not ( n356648 , n356647 );
nand ( n36595 , n36555 , n356648 );
not ( n356650 , n36595 );
buf ( n356651 , n24278 );
buf ( n356652 , n592 );
nand ( n356653 , n356651 , n356652 );
buf ( n356654 , n356653 );
buf ( n356655 , n356654 );
buf ( n356656 , n343567 );
buf ( n356657 , n592 );
nand ( n36604 , n356656 , n356657 );
buf ( n356659 , n36604 );
buf ( n356660 , n356659 );
nand ( n36607 , n356655 , n356660 );
buf ( n356662 , n36607 );
buf ( n356663 , n356662 );
not ( n36610 , n356663 );
buf ( n356665 , n23613 );
not ( n356666 , n356665 );
buf ( n356667 , n356398 );
not ( n356668 , n356667 );
or ( n356669 , n356666 , n356668 );
buf ( n356670 , n592 );
not ( n356671 , n356670 );
buf ( n356672 , n24800 );
not ( n36619 , n356672 );
or ( n356674 , n356671 , n36619 );
buf ( n36621 , n343545 );
buf ( n356676 , n343624 );
nand ( n356677 , n36621 , n356676 );
buf ( n356678 , n356677 );
buf ( n356679 , n356678 );
nand ( n36626 , n356674 , n356679 );
buf ( n356681 , n36626 );
buf ( n356682 , n356681 );
buf ( n356683 , n344705 );
nand ( n356684 , n356682 , n356683 );
buf ( n356685 , n356684 );
buf ( n356686 , n356685 );
nand ( n356687 , n356669 , n356686 );
buf ( n356688 , n356687 );
buf ( n356689 , n356688 );
not ( n356690 , n356689 );
or ( n356691 , n36610 , n356690 );
buf ( n36638 , n356654 );
not ( n36639 , n36638 );
buf ( n36640 , n36639 );
buf ( n36641 , n36640 );
buf ( n356696 , n356659 );
not ( n356697 , n356696 );
buf ( n356698 , n356697 );
buf ( n356699 , n356698 );
nand ( n356700 , n36641 , n356699 );
buf ( n356701 , n356700 );
buf ( n356702 , n356701 );
nand ( n356703 , n356691 , n356702 );
buf ( n356704 , n356703 );
not ( n36651 , n356704 );
or ( n356706 , n356650 , n36651 );
buf ( n356707 , n356648 );
not ( n356708 , n356707 );
buf ( n356709 , n36554 );
buf ( n356710 , n356709 );
nand ( n356711 , n356708 , n356710 );
buf ( n356712 , n356711 );
nand ( n36659 , n356706 , n356712 );
buf ( n356714 , n36659 );
not ( n356715 , n356714 );
buf ( n356716 , n356715 );
buf ( n356717 , n356716 );
nand ( n356718 , n36528 , n356717 );
buf ( n356719 , n356718 );
not ( n356720 , n356719 );
buf ( n36667 , n356623 );
not ( n356722 , n36667 );
buf ( n356723 , n356722 );
buf ( n356724 , n356723 );
not ( n36671 , n356724 );
buf ( n356726 , n356091 );
not ( n36673 , n356726 );
and ( n356728 , n36671 , n36673 );
buf ( n356729 , n356363 );
buf ( n356730 , n23911 );
and ( n356731 , n356729 , n356730 );
nor ( n356732 , n356728 , n356731 );
buf ( n356733 , n356732 );
not ( n356734 , n343863 );
not ( n356735 , n356444 );
or ( n36682 , n356734 , n356735 );
buf ( n356737 , n596 );
not ( n356738 , n356737 );
buf ( n356739 , n24586 );
not ( n356740 , n356739 );
or ( n36687 , n356738 , n356740 );
buf ( n356742 , n344618 );
buf ( n36689 , n343882 );
nand ( n36690 , n356742 , n36689 );
buf ( n36691 , n36690 );
buf ( n356746 , n36691 );
nand ( n356747 , n36687 , n356746 );
buf ( n356748 , n356747 );
buf ( n356749 , n356748 );
buf ( n356750 , n23889 );
nand ( n36697 , n356749 , n356750 );
buf ( n356752 , n36697 );
nand ( n356753 , n36682 , n356752 );
not ( n36700 , n356753 );
not ( n36701 , n592 );
nor ( n356756 , n36701 , n343548 );
buf ( n356757 , n356756 );
not ( n356758 , n356757 );
buf ( n356759 , n356408 );
nand ( n356760 , n356758 , n356759 );
buf ( n356761 , n356760 );
not ( n36708 , n356761 );
or ( n356763 , n36700 , n36708 );
buf ( n356764 , n36360 );
buf ( n356765 , n356756 );
nand ( n356766 , n356764 , n356765 );
buf ( n356767 , n356766 );
nand ( n356768 , n356763 , n356767 );
xor ( n356769 , n356733 , n356768 );
buf ( n36714 , n356416 );
buf ( n36715 , n36360 );
xor ( n36716 , n36714 , n36715 );
buf ( n356773 , n356451 );
xnor ( n356774 , n36716 , n356773 );
buf ( n356775 , n356774 );
not ( n356776 , n356775 );
xnor ( n356777 , n356769 , n356776 );
not ( n356778 , n356777 );
or ( n356779 , n356720 , n356778 );
not ( n356780 , n36527 );
nand ( n356781 , n36659 , n356780 );
nand ( n36720 , n356779 , n356781 );
not ( n36721 , n36720 );
buf ( n356784 , n356733 );
not ( n36723 , n356784 );
buf ( n356786 , n356776 );
nand ( n356787 , n36723 , n356786 );
buf ( n356788 , n356787 );
buf ( n356789 , n356733 );
not ( n36728 , n356789 );
buf ( n356791 , n356775 );
not ( n356792 , n356791 );
or ( n36731 , n36728 , n356792 );
buf ( n356794 , n356768 );
nand ( n356795 , n36731 , n356794 );
buf ( n356796 , n356795 );
nand ( n356797 , n356788 , n356796 );
not ( n36736 , n356797 );
and ( n356799 , n356544 , n356547 );
not ( n36738 , n356544 );
and ( n36739 , n36738 , n36494 );
nor ( n356802 , n356799 , n36739 );
not ( n356803 , n356802 );
nand ( n36742 , n356560 , n356803 );
nand ( n356805 , n356557 , n356802 );
nand ( n356806 , n36736 , n36742 , n356805 );
not ( n36745 , n356806 );
or ( n356808 , n36721 , n36745 );
nand ( n356809 , n36742 , n356805 );
buf ( n356810 , n356809 );
buf ( n356811 , n356797 );
nand ( n36750 , n356810 , n356811 );
buf ( n36751 , n36750 );
nand ( n356814 , n356808 , n36751 );
buf ( n356815 , n356814 );
or ( n356816 , n356571 , n356815 );
buf ( n356817 , n356816 );
buf ( n356818 , n356289 );
not ( n356819 , n356818 );
not ( n36758 , n356210 );
not ( n356821 , n36758 );
not ( n356822 , n36178 );
or ( n36761 , n356821 , n356822 );
or ( n356824 , n36758 , n36178 );
nand ( n356825 , n36761 , n356824 );
buf ( n356826 , n356825 );
not ( n356827 , n356826 );
or ( n356828 , n356819 , n356827 );
buf ( n356829 , n356825 );
buf ( n356830 , n356289 );
or ( n36769 , n356829 , n356830 );
nand ( n356832 , n356828 , n36769 );
buf ( n356833 , n356832 );
buf ( n356834 , n356833 );
not ( n356835 , n356467 );
not ( n36774 , n356474 );
not ( n36775 , n36774 );
or ( n356838 , n356835 , n36775 );
buf ( n356839 , n356467 );
not ( n356840 , n356839 );
buf ( n356841 , n356840 );
buf ( n356842 , n356841 );
not ( n356843 , n356842 );
buf ( n356844 , n356474 );
not ( n356845 , n356844 );
or ( n356846 , n356843 , n356845 );
buf ( n356847 , n356567 );
nand ( n36783 , n356846 , n356847 );
buf ( n356849 , n36783 );
nand ( n356850 , n356838 , n356849 );
buf ( n356851 , n356850 );
nor ( n356852 , n356834 , n356851 );
buf ( n356853 , n356852 );
buf ( n356854 , n356853 );
not ( n356855 , n356854 );
buf ( n356856 , n356855 );
and ( n36792 , n356322 , n356817 , n356856 );
not ( n356858 , n36792 );
buf ( n356859 , n351955 );
buf ( n356860 , n31879 );
or ( n36796 , n356859 , n356860 );
buf ( n356862 , n351930 );
nand ( n36798 , n36796 , n356862 );
buf ( n356864 , n36798 );
buf ( n356865 , n356864 );
buf ( n356866 , n351955 );
buf ( n356867 , n31879 );
nand ( n36803 , n356866 , n356867 );
buf ( n356869 , n36803 );
buf ( n356870 , n356869 );
and ( n36806 , n356865 , n356870 );
buf ( n356872 , n36806 );
buf ( n356873 , n356872 );
not ( n36809 , n356873 );
buf ( n356875 , n36809 );
buf ( n356876 , n356875 );
not ( n356877 , n356876 );
not ( n36813 , n343595 );
not ( n36814 , n352006 );
or ( n356880 , n36813 , n36814 );
not ( n356881 , n344618 );
nand ( n36817 , n356881 , n602 );
not ( n36818 , n36817 );
buf ( n356884 , n344618 );
buf ( n356885 , n343553 );
nand ( n36821 , n356884 , n356885 );
buf ( n36822 , n36821 );
not ( n356888 , n36822 );
or ( n36824 , n36818 , n356888 );
nand ( n356890 , n36824 , n343531 );
nand ( n36826 , n356880 , n356890 );
buf ( n356892 , n36826 );
not ( n356893 , n356892 );
buf ( n356894 , n356893 );
buf ( n356895 , n356894 );
not ( n356896 , n356895 );
or ( n356897 , n356877 , n356896 );
buf ( n356898 , n36826 );
buf ( n356899 , n356872 );
nand ( n356900 , n356898 , n356899 );
buf ( n356901 , n356900 );
buf ( n356902 , n356901 );
nand ( n356903 , n356897 , n356902 );
buf ( n356904 , n356903 );
buf ( n356905 , n356904 );
buf ( n356906 , n31869 );
not ( n356907 , n356906 );
buf ( n356908 , n356907 );
buf ( n356909 , n356908 );
not ( n356910 , n356909 );
buf ( n356911 , n344400 );
not ( n36847 , n356911 );
buf ( n356913 , n36847 );
buf ( n356914 , n356913 );
not ( n356915 , n356914 );
and ( n36851 , n356910 , n356915 );
buf ( n356917 , n604 );
not ( n356918 , n356917 );
buf ( n356919 , n351427 );
not ( n36855 , n356919 );
or ( n36856 , n356918 , n36855 );
buf ( n356922 , n351433 );
buf ( n356923 , n23530 );
nand ( n36859 , n356922 , n356923 );
buf ( n356925 , n36859 );
buf ( n356926 , n356925 );
nand ( n356927 , n36856 , n356926 );
buf ( n356928 , n356927 );
buf ( n356929 , n356928 );
buf ( n356930 , n344338 );
and ( n356931 , n356929 , n356930 );
nor ( n36867 , n36851 , n356931 );
buf ( n356933 , n36867 );
buf ( n356934 , n356933 );
and ( n36870 , n356905 , n356934 );
not ( n356936 , n356905 );
buf ( n356937 , n356933 );
not ( n36873 , n356937 );
buf ( n356939 , n36873 );
buf ( n356940 , n356939 );
and ( n36876 , n356936 , n356940 );
nor ( n36877 , n36870 , n36876 );
buf ( n356943 , n36877 );
buf ( n356944 , n356943 );
not ( n36880 , n356944 );
buf ( n356946 , n36880 );
not ( n356947 , n356946 );
buf ( n356948 , n351861 );
not ( n356949 , n356948 );
buf ( n356950 , n31777 );
not ( n356951 , n356950 );
or ( n36887 , n356949 , n356951 );
buf ( n356953 , n31777 );
buf ( n356954 , n351861 );
or ( n36890 , n356953 , n356954 );
buf ( n356956 , n351836 );
nand ( n36892 , n36890 , n356956 );
buf ( n356958 , n36892 );
buf ( n36894 , n356958 );
nand ( n36895 , n36887 , n36894 );
buf ( n36896 , n36895 );
buf ( n356962 , n344015 );
not ( n36898 , n356962 );
buf ( n356964 , n600 );
not ( n36900 , n356964 );
buf ( n356966 , n344435 );
not ( n36902 , n356966 );
or ( n36903 , n36900 , n36902 );
buf ( n356969 , n23906 );
buf ( n356970 , n24408 );
nand ( n36906 , n356969 , n356970 );
buf ( n356972 , n36906 );
buf ( n356973 , n356972 );
nand ( n356974 , n36903 , n356973 );
buf ( n356975 , n356974 );
buf ( n356976 , n356975 );
not ( n356977 , n356976 );
or ( n356978 , n36898 , n356977 );
buf ( n356979 , n351803 );
buf ( n356980 , n344018 );
nand ( n356981 , n356979 , n356980 );
buf ( n356982 , n356981 );
buf ( n356983 , n356982 );
nand ( n36919 , n356978 , n356983 );
buf ( n36920 , n36919 );
xor ( n356986 , n36896 , n36920 );
buf ( n356987 , n607 );
not ( n356988 , n356987 );
buf ( n356989 , n606 );
not ( n36925 , n356989 );
buf ( n356991 , n334537 );
not ( n356992 , n356991 );
buf ( n356993 , n356992 );
buf ( n356994 , n356993 );
not ( n356995 , n356994 );
or ( n36931 , n36925 , n356995 );
buf ( n356997 , n334537 );
buf ( n356998 , n356997 );
buf ( n356999 , n356998 );
buf ( n357000 , n356999 );
buf ( n357001 , n344445 );
nand ( n36937 , n357000 , n357001 );
buf ( n357003 , n36937 );
buf ( n357004 , n357003 );
nand ( n357005 , n36931 , n357004 );
buf ( n357006 , n357005 );
buf ( n357007 , n357006 );
not ( n357008 , n357007 );
or ( n36944 , n356988 , n357008 );
buf ( n357010 , n352040 );
buf ( n357011 , n344454 );
nand ( n36947 , n357010 , n357011 );
buf ( n357013 , n36947 );
buf ( n357014 , n357013 );
nand ( n36950 , n36944 , n357014 );
buf ( n36951 , n36950 );
xor ( n357017 , n356986 , n36951 );
buf ( n357018 , n357017 );
not ( n357019 , n357018 );
buf ( n357020 , n357019 );
not ( n36956 , n357020 );
or ( n357022 , n356947 , n36956 );
buf ( n36958 , n357017 );
buf ( n357024 , n356943 );
nand ( n357025 , n36958 , n357024 );
buf ( n357026 , n357025 );
nand ( n36962 , n357022 , n357026 );
buf ( n357028 , n351897 );
not ( n357029 , n357028 );
buf ( n357030 , n31631 );
not ( n357031 , n357030 );
buf ( n357032 , n356913 );
not ( n36968 , n357032 );
and ( n36969 , n357031 , n36968 );
buf ( n357035 , n31869 );
buf ( n357036 , n344338 );
and ( n36972 , n357035 , n357036 );
nor ( n357038 , n36969 , n36972 );
buf ( n357039 , n357038 );
buf ( n357040 , n357039 );
nand ( n357041 , n357029 , n357040 );
buf ( n357042 , n357041 );
and ( n36978 , n357042 , n351956 );
buf ( n357044 , n351897 );
not ( n357045 , n357044 );
buf ( n357046 , n357039 );
nor ( n357047 , n357045 , n357046 );
buf ( n357048 , n357047 );
nor ( n36984 , n36978 , n357048 );
not ( n357050 , n36984 );
not ( n357051 , n357050 );
and ( n36987 , n31887 , n344705 );
buf ( n357053 , n592 );
not ( n357054 , n357053 );
buf ( n357055 , n343985 );
not ( n357056 , n357055 );
or ( n357057 , n357054 , n357056 );
buf ( n357058 , n343982 );
buf ( n357059 , n343624 );
nand ( n357060 , n357058 , n357059 );
buf ( n357061 , n357060 );
buf ( n357062 , n357061 );
nand ( n357063 , n357057 , n357062 );
buf ( n357064 , n357063 );
and ( n37000 , n357064 , n23613 );
nor ( n357066 , n36987 , n37000 );
not ( n357067 , n357066 );
buf ( n37003 , n344957 );
buf ( n357069 , n592 );
and ( n357070 , n37003 , n357069 );
buf ( n357071 , n357070 );
not ( n37007 , n357071 );
and ( n357073 , n357067 , n37007 );
and ( n357074 , n357066 , n357071 );
nor ( n37010 , n357073 , n357074 );
buf ( n357076 , n343863 );
not ( n357077 , n357076 );
buf ( n357078 , n596 );
not ( n357079 , n357078 );
buf ( n357080 , n14695 );
not ( n37016 , n357080 );
buf ( n37017 , n37016 );
buf ( n357083 , n37017 );
not ( n37019 , n357083 );
or ( n357085 , n357079 , n37019 );
buf ( n37021 , n14695 );
buf ( n357087 , n343882 );
nand ( n37023 , n37021 , n357087 );
buf ( n357089 , n37023 );
buf ( n357090 , n357089 );
nand ( n37026 , n357085 , n357090 );
buf ( n357092 , n37026 );
buf ( n357093 , n357092 );
not ( n37029 , n357093 );
or ( n37030 , n357077 , n37029 );
buf ( n357096 , n351945 );
buf ( n357097 , n23889 );
nand ( n37033 , n357096 , n357097 );
buf ( n357099 , n37033 );
buf ( n357100 , n357099 );
nand ( n357101 , n37030 , n357100 );
buf ( n357102 , n357101 );
not ( n357103 , n357102 );
and ( n37039 , n37010 , n357103 );
not ( n357105 , n37010 );
and ( n37041 , n357105 , n357102 );
nor ( n357107 , n37039 , n37041 );
buf ( n357108 , n343765 );
not ( n37044 , n357108 );
buf ( n357110 , n351826 );
not ( n357111 , n357110 );
or ( n37047 , n37044 , n357111 );
buf ( n357113 , n594 );
not ( n357114 , n357113 );
buf ( n357115 , n24026 );
not ( n357116 , n357115 );
or ( n357117 , n357114 , n357116 );
buf ( n357118 , n344588 );
buf ( n357119 , n343632 );
nand ( n357120 , n357118 , n357119 );
buf ( n357121 , n357120 );
buf ( n357122 , n357121 );
nand ( n357123 , n357117 , n357122 );
buf ( n357124 , n357123 );
buf ( n357125 , n357124 );
buf ( n357126 , n23681 );
nand ( n357127 , n357125 , n357126 );
buf ( n357128 , n357127 );
buf ( n357129 , n357128 );
nand ( n357130 , n37047 , n357129 );
buf ( n357131 , n357130 );
buf ( n357132 , n357131 );
not ( n37068 , n357132 );
buf ( n357134 , n23911 );
not ( n37070 , n357134 );
buf ( n357136 , n598 );
not ( n37072 , n357136 );
buf ( n357138 , n344383 );
not ( n37074 , n357138 );
or ( n37075 , n37072 , n37074 );
buf ( n357141 , n24346 );
buf ( n357142 , n343953 );
nand ( n37078 , n357141 , n357142 );
buf ( n357144 , n37078 );
buf ( n357145 , n357144 );
nand ( n357146 , n37075 , n357145 );
buf ( n357147 , n357146 );
buf ( n357148 , n357147 );
not ( n357149 , n357148 );
or ( n357150 , n37070 , n357149 );
buf ( n357151 , n351851 );
buf ( n357152 , n343948 );
nand ( n357153 , n357151 , n357152 );
buf ( n357154 , n357153 );
buf ( n357155 , n357154 );
nand ( n357156 , n357150 , n357155 );
buf ( n357157 , n357156 );
buf ( n357158 , n357157 );
not ( n357159 , n357158 );
buf ( n357160 , n357159 );
buf ( n357161 , n357160 );
not ( n357162 , n357161 );
or ( n357163 , n37068 , n357162 );
buf ( n357164 , n357160 );
buf ( n357165 , n357131 );
or ( n37100 , n357164 , n357165 );
nand ( n357167 , n357163 , n37100 );
buf ( n357168 , n357167 );
and ( n37103 , n357107 , n357168 );
not ( n37104 , n357107 );
not ( n37105 , n357168 );
and ( n37106 , n37104 , n37105 );
nor ( n357173 , n37103 , n37106 );
buf ( n357174 , n357173 );
not ( n357175 , n357174 );
buf ( n357176 , n357175 );
not ( n37111 , n357176 );
or ( n357178 , n357051 , n37111 );
buf ( n357179 , n357173 );
buf ( n357180 , n36984 );
nand ( n357181 , n357179 , n357180 );
buf ( n357182 , n357181 );
nand ( n37117 , n357178 , n357182 );
not ( n357184 , n351998 );
not ( n37119 , n352016 );
nand ( n37120 , n37119 , n32015 );
not ( n357187 , n37120 );
or ( n37122 , n357184 , n357187 );
buf ( n357189 , n352016 );
buf ( n357190 , n352047 );
nand ( n37125 , n357189 , n357190 );
buf ( n357192 , n37125 );
nand ( n37127 , n37122 , n357192 );
buf ( n357194 , n37127 );
not ( n37129 , n357194 );
buf ( n357196 , n37129 );
and ( n357197 , n37117 , n357196 );
not ( n37132 , n37117 );
buf ( n357199 , n37127 );
buf ( n37134 , n357199 );
buf ( n357201 , n37134 );
and ( n37136 , n37132 , n357201 );
nor ( n37137 , n357197 , n37136 );
not ( n37138 , n37137 );
and ( n37139 , n36962 , n37138 );
not ( n37140 , n36962 );
and ( n37141 , n37140 , n37137 );
nor ( n37142 , n37139 , n37141 );
buf ( n357209 , n37142 );
xor ( n37144 , n351872 , n351891 );
and ( n37145 , n37144 , n351958 );
and ( n37146 , n351872 , n351891 );
or ( n37147 , n37145 , n37146 );
buf ( n357214 , n37147 );
buf ( n357215 , n357214 );
not ( n357216 , n357215 );
not ( n37151 , n352054 );
not ( n37152 , n351979 );
or ( n37153 , n37151 , n37152 );
not ( n357220 , n352051 );
not ( n357221 , n351982 );
or ( n37156 , n357220 , n357221 );
nand ( n357223 , n37156 , n352077 );
nand ( n357224 , n37153 , n357223 );
buf ( n357225 , n357224 );
not ( n357226 , n357225 );
and ( n357227 , n357216 , n357226 );
buf ( n357228 , n357224 );
buf ( n357229 , n357214 );
and ( n357230 , n357228 , n357229 );
nor ( n357231 , n357227 , n357230 );
buf ( n357232 , n357231 );
buf ( n357233 , n357232 );
xor ( n357234 , n357209 , n357233 );
buf ( n357235 , n357234 );
xor ( n37167 , n351960 , n351969 );
and ( n357237 , n37167 , n352087 );
and ( n37169 , n351960 , n351969 );
or ( n357239 , n357237 , n37169 );
nand ( n357240 , n357235 , n357239 );
and ( n357241 , n31712 , n357240 , n352109 );
not ( n37173 , n357240 );
not ( n357243 , n32074 );
or ( n357244 , n37173 , n357243 );
buf ( n357245 , n357235 );
not ( n37177 , n357245 );
buf ( n357247 , n37177 );
not ( n37179 , n357239 );
nand ( n357249 , n357247 , n37179 );
nand ( n37181 , n357244 , n357249 );
or ( n37182 , n357241 , n37181 );
buf ( n357252 , n23889 );
not ( n357253 , n357252 );
buf ( n357254 , n357092 );
not ( n357255 , n357254 );
or ( n357256 , n357253 , n357255 );
buf ( n357257 , n596 );
not ( n357258 , n357257 );
buf ( n37190 , n343548 );
not ( n37191 , n37190 );
or ( n37192 , n357258 , n37191 );
buf ( n37193 , n343545 );
buf ( n37194 , n343882 );
nand ( n37195 , n37193 , n37194 );
buf ( n37196 , n37195 );
buf ( n37197 , n37196 );
nand ( n37198 , n37192 , n37197 );
buf ( n37199 , n37198 );
buf ( n357269 , n37199 );
buf ( n357270 , n343863 );
nand ( n357271 , n357269 , n357270 );
buf ( n357272 , n357271 );
buf ( n357273 , n357272 );
nand ( n357274 , n357256 , n357273 );
buf ( n357275 , n357274 );
buf ( n357276 , n357275 );
buf ( n357277 , n23911 );
not ( n357278 , n357277 );
buf ( n357279 , n598 );
not ( n357280 , n357279 );
buf ( n357281 , n345091 );
not ( n357282 , n357281 );
or ( n357283 , n357280 , n357282 );
buf ( n357284 , n344353 );
not ( n357285 , n357284 );
buf ( n357286 , n357285 );
buf ( n357287 , n357286 );
buf ( n357288 , n343953 );
nand ( n37220 , n357287 , n357288 );
buf ( n357290 , n37220 );
buf ( n357291 , n357290 );
nand ( n357292 , n357283 , n357291 );
buf ( n357293 , n357292 );
buf ( n37225 , n357293 );
not ( n37226 , n37225 );
or ( n37227 , n357278 , n37226 );
buf ( n37228 , n357147 );
buf ( n37229 , n343948 );
nand ( n37230 , n37228 , n37229 );
buf ( n37231 , n37230 );
buf ( n37232 , n37231 );
nand ( n37233 , n37227 , n37232 );
buf ( n37234 , n37233 );
buf ( n357304 , n37234 );
not ( n357305 , n357304 );
buf ( n357306 , n357305 );
buf ( n357307 , n357306 );
xor ( n357308 , n357276 , n357307 );
buf ( n357309 , n357102 );
buf ( n357310 , n357071 );
or ( n357311 , n357309 , n357310 );
buf ( n357312 , n357066 );
not ( n37244 , n357312 );
buf ( n357314 , n37244 );
buf ( n357315 , n357314 );
nand ( n37247 , n357311 , n357315 );
buf ( n37248 , n37247 );
buf ( n357318 , n37248 );
buf ( n357319 , n357102 );
buf ( n357320 , n357071 );
nand ( n357321 , n357319 , n357320 );
buf ( n357322 , n357321 );
buf ( n357323 , n357322 );
nand ( n357324 , n357318 , n357323 );
buf ( n357325 , n357324 );
buf ( n357326 , n357325 );
xnor ( n37258 , n357308 , n357326 );
buf ( n357328 , n37258 );
not ( n37260 , n36826 );
not ( n37261 , n356939 );
or ( n37262 , n37260 , n37261 );
not ( n37263 , n356894 );
not ( n37264 , n356933 );
or ( n37265 , n37263 , n37264 );
nand ( n357335 , n37265 , n356875 );
nand ( n37267 , n37262 , n357335 );
xor ( n357337 , n357328 , n37267 );
not ( n357338 , n23532 );
not ( n37270 , n356431 );
not ( n357340 , n343553 );
or ( n357341 , n37270 , n357340 );
nand ( n37273 , n355697 , n602 );
nand ( n37274 , n357341 , n37273 );
not ( n357344 , n37274 );
or ( n37276 , n357338 , n357344 );
not ( n37277 , n36817 );
not ( n357347 , n36822 );
or ( n37279 , n37277 , n357347 );
nand ( n37280 , n37279 , n343595 );
nand ( n357350 , n37276 , n37280 );
buf ( n357351 , n357350 );
not ( n357352 , n357351 );
buf ( n357353 , n357352 );
buf ( n357354 , n357353 );
not ( n37286 , n357354 );
not ( n357356 , n343969 );
nand ( n37288 , n357356 , n592 );
not ( n37289 , n23681 );
not ( n37290 , n345322 );
not ( n37291 , n343632 );
or ( n37292 , n37290 , n37291 );
nand ( n37293 , n344301 , n594 );
nand ( n37294 , n37292 , n37293 );
not ( n37295 , n37294 );
or ( n37296 , n37289 , n37295 );
nand ( n37297 , n357124 , n343765 );
nand ( n37298 , n37296 , n37297 );
xor ( n37299 , n37288 , n37298 );
not ( n37300 , n23613 );
buf ( n357370 , n592 );
not ( n37302 , n357370 );
buf ( n357372 , n23996 );
not ( n37304 , n357372 );
or ( n37305 , n37302 , n37304 );
buf ( n37306 , n23993 );
buf ( n357376 , n343624 );
nand ( n37308 , n37306 , n357376 );
buf ( n357378 , n37308 );
buf ( n357379 , n357378 );
nand ( n357380 , n37305 , n357379 );
buf ( n357381 , n357380 );
not ( n37313 , n357381 );
or ( n357383 , n37300 , n37313 );
buf ( n357384 , n357064 );
buf ( n357385 , n344705 );
nand ( n37317 , n357384 , n357385 );
buf ( n357387 , n37317 );
nand ( n37319 , n357383 , n357387 );
buf ( n357389 , n37319 );
not ( n37321 , n357389 );
buf ( n357391 , n37321 );
xnor ( n37323 , n37299 , n357391 );
buf ( n357393 , n37323 );
not ( n37325 , n357393 );
buf ( n357395 , n37325 );
buf ( n357396 , n357395 );
not ( n37328 , n357396 );
or ( n37329 , n37286 , n37328 );
buf ( n357399 , n37323 );
buf ( n357400 , n357350 );
nand ( n37332 , n357399 , n357400 );
buf ( n357402 , n37332 );
buf ( n357403 , n357402 );
nand ( n37335 , n37329 , n357403 );
buf ( n357405 , n37335 );
buf ( n357406 , n357405 );
buf ( n357407 , n344338 );
not ( n357408 , n357407 );
buf ( n357409 , n604 );
not ( n357410 , n357409 );
buf ( n37342 , n352036 );
not ( n357412 , n37342 );
buf ( n357413 , n357412 );
buf ( n357414 , n357413 );
not ( n357415 , n357414 );
or ( n37347 , n357410 , n357415 );
buf ( n357417 , n355593 );
buf ( n357418 , n23530 );
nand ( n37350 , n357417 , n357418 );
buf ( n357420 , n37350 );
buf ( n357421 , n357420 );
nand ( n357422 , n37347 , n357421 );
buf ( n357423 , n357422 );
buf ( n357424 , n357423 );
not ( n37356 , n357424 );
or ( n357426 , n357408 , n37356 );
buf ( n357427 , n356928 );
buf ( n357428 , n344400 );
nand ( n357429 , n357427 , n357428 );
buf ( n357430 , n357429 );
buf ( n357431 , n357430 );
nand ( n357432 , n357426 , n357431 );
buf ( n357433 , n357432 );
buf ( n357434 , n357433 );
buf ( n37366 , n357434 );
buf ( n357436 , n37366 );
buf ( n357437 , n357436 );
not ( n357438 , n357437 );
buf ( n357439 , n357438 );
buf ( n357440 , n357439 );
and ( n357441 , n357406 , n357440 );
not ( n37373 , n357406 );
buf ( n357443 , n357436 );
and ( n37375 , n37373 , n357443 );
nor ( n37376 , n357441 , n37375 );
buf ( n357446 , n37376 );
buf ( n357447 , n357446 );
not ( n37379 , n357447 );
buf ( n357449 , n37379 );
xor ( n37381 , n357337 , n357449 );
xor ( n37382 , n36896 , n36920 );
and ( n37383 , n37382 , n36951 );
and ( n37384 , n36896 , n36920 );
or ( n37385 , n37383 , n37384 );
not ( n37386 , n344015 );
buf ( n357456 , n600 );
not ( n357457 , n357456 );
buf ( n357458 , n24392 );
not ( n357459 , n357458 );
or ( n37391 , n357457 , n357459 );
buf ( n357461 , n350821 );
buf ( n357462 , n23906 );
nand ( n37394 , n357461 , n357462 );
buf ( n357464 , n37394 );
buf ( n357465 , n357464 );
nand ( n357466 , n37391 , n357465 );
buf ( n357467 , n357466 );
not ( n37399 , n357467 );
or ( n357469 , n37386 , n37399 );
nand ( n357470 , n356975 , n344018 );
nand ( n37402 , n357469 , n357470 );
not ( n357472 , n344454 );
not ( n357473 , n357006 );
or ( n37405 , n357472 , n357473 );
buf ( n357475 , n606 );
not ( n37407 , n357475 );
buf ( n37408 , n334531 );
not ( n37409 , n37408 );
buf ( n37410 , n37409 );
buf ( n357480 , n37410 );
not ( n37412 , n357480 );
or ( n357482 , n37407 , n37412 );
buf ( n37414 , n334531 );
buf ( n357484 , n344445 );
nand ( n357485 , n37414 , n357484 );
buf ( n357486 , n357485 );
buf ( n357487 , n357486 );
nand ( n357488 , n357482 , n357487 );
buf ( n357489 , n357488 );
buf ( n357490 , n357489 );
buf ( n357491 , n607 );
nand ( n37423 , n357490 , n357491 );
buf ( n357493 , n37423 );
nand ( n37425 , n37405 , n357493 );
xor ( n37426 , n37402 , n37425 );
buf ( n357496 , n357131 );
not ( n37428 , n357496 );
buf ( n357498 , n357160 );
nand ( n37430 , n37428 , n357498 );
buf ( n357500 , n37430 );
not ( n37432 , n357500 );
not ( n37433 , n357107 );
or ( n37434 , n37432 , n37433 );
buf ( n357504 , n357157 );
buf ( n357505 , n357131 );
nand ( n37437 , n357504 , n357505 );
buf ( n357507 , n37437 );
nand ( n37439 , n37434 , n357507 );
xor ( n37440 , n37426 , n37439 );
xor ( n357510 , n37385 , n37440 );
not ( n37442 , n357173 );
not ( n357512 , n37127 );
or ( n357513 , n37442 , n357512 );
buf ( n357514 , n37127 );
buf ( n357515 , n357173 );
or ( n357516 , n357514 , n357515 );
buf ( n357517 , n357050 );
nand ( n357518 , n357516 , n357517 );
buf ( n357519 , n357518 );
nand ( n37451 , n357513 , n357519 );
xor ( n357521 , n357510 , n37451 );
xor ( n37453 , n37381 , n357521 );
buf ( n357523 , n357017 );
not ( n357524 , n357523 );
buf ( n357525 , n356943 );
nand ( n357526 , n357524 , n357525 );
buf ( n357527 , n357526 );
not ( n357528 , n357527 );
not ( n37460 , n37138 );
or ( n357530 , n357528 , n37460 );
not ( n37462 , n356943 );
nand ( n357532 , n37462 , n357017 );
nand ( n37464 , n357530 , n357532 );
xor ( n37465 , n37453 , n37464 );
not ( n357535 , n37465 );
buf ( n357536 , n37142 );
buf ( n37468 , n357536 );
buf ( n37469 , n37468 );
buf ( n357539 , n37469 );
buf ( n357540 , n357224 );
buf ( n37472 , n357540 );
buf ( n357542 , n37472 );
buf ( n357543 , n357542 );
not ( n37475 , n357543 );
buf ( n357545 , n357214 );
nand ( n37477 , n37475 , n357545 );
buf ( n357547 , n37477 );
buf ( n357548 , n357547 );
and ( n37480 , n357539 , n357548 );
buf ( n357550 , n357542 );
buf ( n357551 , n357214 );
not ( n37483 , n357551 );
buf ( n357553 , n37483 );
buf ( n357554 , n357553 );
and ( n357555 , n357550 , n357554 );
nor ( n37487 , n37480 , n357555 );
buf ( n357557 , n37487 );
nand ( n37489 , n357535 , n357557 );
nand ( n37490 , n37182 , n37489 );
buf ( n357560 , n357557 );
not ( n357561 , n357560 );
buf ( n357562 , n37465 );
buf ( n357563 , n357562 );
buf ( n357564 , n357563 );
buf ( n357565 , n357564 );
nand ( n357566 , n357561 , n357565 );
buf ( n357567 , n357566 );
nand ( n37499 , n37490 , n357567 );
not ( n37500 , n37499 );
buf ( n357570 , n592 );
not ( n37502 , n357570 );
buf ( n357572 , n24026 );
not ( n37504 , n357572 );
or ( n37505 , n37502 , n37504 );
buf ( n357575 , n344588 );
buf ( n357576 , n343624 );
nand ( n37508 , n357575 , n357576 );
buf ( n37509 , n37508 );
buf ( n357579 , n37509 );
nand ( n37511 , n37505 , n357579 );
buf ( n357581 , n37511 );
buf ( n357582 , n357581 );
not ( n357583 , n357582 );
buf ( n357584 , n357583 );
buf ( n357585 , n357584 );
not ( n357586 , n357585 );
buf ( n357587 , n355637 );
not ( n37519 , n357587 );
and ( n357589 , n357586 , n37519 );
buf ( n357590 , n592 );
not ( n37522 , n357590 );
buf ( n357592 , n344301 );
not ( n37524 , n357592 );
or ( n37525 , n37522 , n37524 );
buf ( n357595 , n345322 );
buf ( n357596 , n343624 );
nand ( n37528 , n357595 , n357596 );
buf ( n357598 , n37528 );
buf ( n357599 , n357598 );
nand ( n37531 , n37525 , n357599 );
buf ( n357601 , n37531 );
buf ( n357602 , n357601 );
buf ( n357603 , n23613 );
and ( n37535 , n357602 , n357603 );
nor ( n357605 , n357589 , n37535 );
buf ( n357606 , n357605 );
buf ( n357607 , n357606 );
not ( n37539 , n357607 );
buf ( n357609 , n37539 );
buf ( n357610 , n344015 );
not ( n37542 , n357610 );
buf ( n357612 , n600 );
not ( n357613 , n357612 );
buf ( n357614 , n31390 );
not ( n357615 , n357614 );
or ( n37547 , n357613 , n357615 );
buf ( n357617 , n351424 );
buf ( n357618 , n23906 );
nand ( n37550 , n357617 , n357618 );
buf ( n37551 , n37550 );
buf ( n357621 , n37551 );
nand ( n37553 , n37547 , n357621 );
buf ( n357623 , n37553 );
buf ( n357624 , n357623 );
not ( n357625 , n357624 );
or ( n37557 , n37542 , n357625 );
and ( n357627 , n600 , n355697 );
not ( n357628 , n600 );
and ( n37560 , n357628 , n356431 );
or ( n357630 , n357627 , n37560 );
buf ( n37562 , n357630 );
buf ( n357632 , n344018 );
nand ( n357633 , n37562 , n357632 );
buf ( n357634 , n357633 );
buf ( n357635 , n357634 );
nand ( n357636 , n37557 , n357635 );
buf ( n357637 , n357636 );
xor ( n357638 , n357609 , n357637 );
not ( n357639 , n592 );
nor ( n37571 , n357639 , n344896 );
buf ( n37572 , n37571 );
buf ( n357642 , n344705 );
not ( n357643 , n357642 );
buf ( n357644 , n357601 );
not ( n37576 , n357644 );
or ( n357646 , n357643 , n37576 );
and ( n357647 , n592 , n37017 );
not ( n37579 , n592 );
and ( n357649 , n37579 , n14695 );
or ( n37581 , n357647 , n357649 );
buf ( n357651 , n37581 );
buf ( n357652 , n23613 );
nand ( n37584 , n357651 , n357652 );
buf ( n357654 , n37584 );
buf ( n357655 , n357654 );
nand ( n357656 , n357646 , n357655 );
buf ( n357657 , n357656 );
buf ( n357658 , n357657 );
xor ( n357659 , n37572 , n357658 );
buf ( n357660 , n23681 );
not ( n37592 , n357660 );
and ( n357662 , n594 , n344383 );
not ( n37594 , n594 );
and ( n357664 , n37594 , n24346 );
or ( n357665 , n357662 , n357664 );
buf ( n357666 , n357665 );
not ( n357667 , n357666 );
or ( n357668 , n37592 , n357667 );
buf ( n357669 , n594 );
not ( n37601 , n357669 );
buf ( n357671 , n24800 );
not ( n357672 , n357671 );
or ( n37604 , n37601 , n357672 );
buf ( n357674 , n343545 );
buf ( n357675 , n343632 );
nand ( n37607 , n357674 , n357675 );
buf ( n37608 , n37607 );
buf ( n357678 , n37608 );
nand ( n37610 , n37604 , n357678 );
buf ( n357680 , n37610 );
buf ( n357681 , n357680 );
buf ( n357682 , n343765 );
nand ( n37614 , n357681 , n357682 );
buf ( n357684 , n37614 );
buf ( n357685 , n357684 );
nand ( n357686 , n357668 , n357685 );
buf ( n357687 , n357686 );
buf ( n357688 , n357687 );
xor ( n37620 , n357659 , n357688 );
buf ( n357690 , n37620 );
xor ( n37622 , n357638 , n357690 );
buf ( n357692 , n343863 );
not ( n37624 , n357692 );
and ( n37625 , n596 , n344436 );
not ( n357695 , n596 );
and ( n357696 , n357695 , n24408 );
or ( n37628 , n37625 , n357696 );
buf ( n357698 , n37628 );
not ( n37630 , n357698 );
or ( n37631 , n37624 , n37630 );
xor ( n37632 , n596 , n344361 );
buf ( n357702 , n37632 );
buf ( n357703 , n23889 );
nand ( n37635 , n357702 , n357703 );
buf ( n357705 , n37635 );
buf ( n357706 , n357705 );
nand ( n37638 , n37631 , n357706 );
buf ( n357708 , n37638 );
xor ( n37640 , n343953 , n344618 );
buf ( n357710 , n37640 );
not ( n37642 , n357710 );
buf ( n37643 , n356086 );
not ( n37644 , n37643 );
and ( n37645 , n37642 , n37644 );
buf ( n357715 , n598 );
not ( n357716 , n357715 );
buf ( n357717 , n350815 );
not ( n357718 , n357717 );
or ( n357719 , n357716 , n357718 );
nand ( n37651 , n24390 , n24389 );
nand ( n357721 , n343953 , n37651 );
buf ( n37653 , n357721 );
nand ( n37654 , n357719 , n37653 );
buf ( n37655 , n37654 );
buf ( n357725 , n37655 );
buf ( n357726 , n343948 );
and ( n357727 , n357725 , n357726 );
nor ( n357728 , n37645 , n357727 );
buf ( n357729 , n357728 );
buf ( n357730 , n357729 );
buf ( n37659 , n29097 );
not ( n37660 , n37659 );
buf ( n357733 , n356913 );
not ( n37662 , n357733 );
or ( n37663 , n37660 , n37662 );
buf ( n357736 , n604 );
not ( n37665 , n357736 );
buf ( n357738 , n37410 );
not ( n37667 , n357738 );
or ( n37668 , n37665 , n37667 );
buf ( n357741 , n334531 );
buf ( n357742 , n23530 );
nand ( n37671 , n357741 , n357742 );
buf ( n357744 , n37671 );
buf ( n357745 , n357744 );
nand ( n37674 , n37668 , n357745 );
buf ( n357747 , n37674 );
buf ( n357748 , n357747 );
nand ( n357749 , n37663 , n357748 );
buf ( n357750 , n357749 );
buf ( n357751 , n357750 );
not ( n37680 , n357751 );
buf ( n357753 , n37680 );
buf ( n357754 , n357753 );
and ( n357755 , n357730 , n357754 );
not ( n357756 , n357730 );
buf ( n357757 , n357750 );
and ( n357758 , n357756 , n357757 );
nor ( n357759 , n357755 , n357758 );
buf ( n357760 , n357759 );
or ( n357761 , n357708 , n357760 );
nand ( n357762 , n357760 , n357708 );
nand ( n37691 , n357761 , n357762 );
not ( n357764 , n37691 );
xor ( n357765 , n37622 , n357764 );
buf ( n357766 , n343948 );
not ( n357767 , n357766 );
buf ( n357768 , n598 );
not ( n37697 , n357768 );
buf ( n357770 , n344436 );
not ( n37699 , n357770 );
or ( n37700 , n37697 , n37699 );
buf ( n357773 , n24408 );
buf ( n357774 , n343953 );
nand ( n357775 , n357773 , n357774 );
buf ( n357776 , n357775 );
buf ( n357777 , n357776 );
nand ( n357778 , n37700 , n357777 );
buf ( n357779 , n357778 );
buf ( n357780 , n357779 );
not ( n357781 , n357780 );
or ( n37710 , n357767 , n357781 );
buf ( n357783 , n37655 );
buf ( n357784 , n23911 );
nand ( n37713 , n357783 , n357784 );
buf ( n37714 , n37713 );
buf ( n357787 , n37714 );
nand ( n37716 , n37710 , n357787 );
buf ( n37717 , n37716 );
not ( n357790 , n37717 );
not ( n357791 , n343531 );
not ( n37720 , n602 );
and ( n357793 , n37720 , n355596 );
not ( n37722 , n37720 );
buf ( n357795 , n357413 );
not ( n37724 , n357795 );
buf ( n357797 , n37724 );
and ( n357798 , n37722 , n357797 );
nor ( n357799 , n357793 , n357798 );
not ( n37728 , n357799 );
or ( n37729 , n357791 , n37728 );
and ( n37730 , n356635 , n23977 );
not ( n37731 , n356635 );
and ( n37732 , n37731 , n602 );
nor ( n37733 , n37730 , n37732 );
buf ( n357806 , n37733 );
buf ( n357807 , n343595 );
nand ( n37736 , n357806 , n357807 );
buf ( n357809 , n37736 );
nand ( n37738 , n37729 , n357809 );
not ( n37739 , n37738 );
or ( n37740 , n357790 , n37739 );
buf ( n357813 , n37738 );
buf ( n357814 , n37717 );
or ( n357815 , n357813 , n357814 );
not ( n37744 , n343863 );
not ( n357817 , n343882 );
not ( n37746 , n24346 );
or ( n357819 , n357817 , n37746 );
or ( n37748 , n24346 , n343882 );
nand ( n37749 , n357819 , n37748 );
not ( n37750 , n37749 );
or ( n357823 , n37744 , n37750 );
buf ( n357824 , n37199 );
buf ( n357825 , n23889 );
nand ( n357826 , n357824 , n357825 );
buf ( n357827 , n357826 );
nand ( n37756 , n357823 , n357827 );
buf ( n357829 , n37756 );
buf ( n357830 , n23613 );
not ( n37759 , n357830 );
buf ( n357832 , n357581 );
not ( n357833 , n357832 );
or ( n37762 , n37759 , n357833 );
buf ( n357835 , n357381 );
buf ( n37764 , n344705 );
nand ( n37765 , n357835 , n37764 );
buf ( n357838 , n37765 );
buf ( n357839 , n357838 );
nand ( n37768 , n37762 , n357839 );
buf ( n357841 , n37768 );
buf ( n357842 , n357841 );
or ( n37771 , n357829 , n357842 );
buf ( n357844 , n343765 );
not ( n37773 , n357844 );
buf ( n357846 , n37294 );
not ( n37775 , n357846 );
or ( n37776 , n37773 , n37775 );
buf ( n357849 , n594 );
buf ( n357850 , n14695 );
and ( n37779 , n357849 , n357850 );
not ( n37780 , n357849 );
buf ( n357853 , n37017 );
and ( n37782 , n37780 , n357853 );
nor ( n37783 , n37779 , n37782 );
buf ( n357856 , n37783 );
buf ( n357857 , n357856 );
buf ( n357858 , n23681 );
nand ( n357859 , n357857 , n357858 );
buf ( n357860 , n357859 );
buf ( n357861 , n357860 );
nand ( n357862 , n37776 , n357861 );
buf ( n357863 , n357862 );
buf ( n357864 , n357863 );
nand ( n357865 , n37771 , n357864 );
buf ( n357866 , n357865 );
buf ( n357867 , n357866 );
buf ( n357868 , n37756 );
buf ( n357869 , n357841 );
nand ( n37798 , n357868 , n357869 );
buf ( n37799 , n37798 );
buf ( n357872 , n37799 );
nand ( n37801 , n357867 , n357872 );
buf ( n357874 , n37801 );
buf ( n357875 , n357874 );
nand ( n357876 , n357815 , n357875 );
buf ( n37802 , n357876 );
nand ( n37803 , n37740 , n37802 );
xor ( n357879 , n357765 , n37803 );
buf ( n357880 , n357353 );
not ( n37806 , n357880 );
buf ( n357882 , n357433 );
not ( n357883 , n357882 );
buf ( n357884 , n357883 );
buf ( n357885 , n357884 );
not ( n37811 , n357885 );
or ( n37812 , n37806 , n37811 );
buf ( n357888 , n357395 );
nand ( n37814 , n37812 , n357888 );
buf ( n357890 , n37814 );
buf ( n37816 , n357890 );
buf ( n357892 , n357433 );
buf ( n357893 , n357350 );
nand ( n357894 , n357892 , n357893 );
buf ( n357895 , n357894 );
buf ( n37821 , n357895 );
nand ( n37822 , n37816 , n37821 );
buf ( n37823 , n37822 );
buf ( n357899 , n37823 );
not ( n37825 , n357899 );
buf ( n357901 , n343985 );
not ( n37827 , n357901 );
buf ( n357903 , n592 );
nand ( n37829 , n37827 , n357903 );
buf ( n357905 , n37829 );
buf ( n357906 , n357905 );
not ( n357907 , n37288 );
not ( n37833 , n357907 );
not ( n357909 , n37319 );
or ( n357910 , n37833 , n357909 );
not ( n37836 , n37288 );
not ( n357912 , n357391 );
or ( n37838 , n37836 , n357912 );
buf ( n357914 , n37298 );
nand ( n37840 , n37838 , n357914 );
nand ( n37841 , n357910 , n37840 );
buf ( n357917 , n37841 );
xor ( n37843 , n357906 , n357917 );
not ( n37844 , n343595 );
not ( n37845 , n37274 );
or ( n37846 , n37844 , n37845 );
nand ( n357922 , n37733 , n343531 );
nand ( n37848 , n37846 , n357922 );
buf ( n357924 , n37848 );
xnor ( n37850 , n37843 , n357924 );
buf ( n357926 , n37850 );
buf ( n357927 , n357926 );
nand ( n37853 , n37825 , n357927 );
buf ( n357929 , n37853 );
buf ( n357930 , n344452 );
not ( n37856 , n357930 );
buf ( n357932 , n344631 );
not ( n37858 , n357932 );
or ( n37859 , n37856 , n37858 );
buf ( n357935 , n357489 );
nand ( n37861 , n37859 , n357935 );
buf ( n357937 , n37861 );
not ( n37863 , n37756 );
not ( n37864 , n37863 );
or ( n37865 , n357841 , n357863 );
nand ( n37866 , n357863 , n357841 );
nand ( n37867 , n37865 , n37866 );
not ( n37868 , n37867 );
or ( n37869 , n37864 , n37868 );
not ( n37870 , n37867 );
not ( n37871 , n37863 );
nand ( n37872 , n37870 , n37871 );
nand ( n357948 , n37869 , n37872 );
xor ( n37874 , n357937 , n357948 );
buf ( n357950 , n344018 );
not ( n357951 , n357950 );
buf ( n357952 , n357467 );
not ( n37878 , n357952 );
or ( n37879 , n357951 , n37878 );
buf ( n357955 , n344015 );
buf ( n357956 , n600 );
not ( n37882 , n357956 );
buf ( n357958 , n356881 );
not ( n37884 , n357958 );
or ( n357960 , n37882 , n37884 );
buf ( n357961 , n344618 );
buf ( n357962 , n23906 );
nand ( n357963 , n357961 , n357962 );
buf ( n357964 , n357963 );
buf ( n357965 , n357964 );
nand ( n357966 , n357960 , n357965 );
buf ( n357967 , n357966 );
buf ( n357968 , n357967 );
nand ( n357969 , n357955 , n357968 );
buf ( n357970 , n357969 );
buf ( n357971 , n357970 );
nand ( n357972 , n37879 , n357971 );
buf ( n357973 , n357972 );
buf ( n357974 , n357973 );
not ( n357975 , n357974 );
buf ( n357976 , n357975 );
xor ( n37902 , n37874 , n357976 );
and ( n357978 , n357929 , n37902 );
buf ( n357979 , n37823 );
not ( n357980 , n357979 );
buf ( n357981 , n357926 );
nor ( n37907 , n357980 , n357981 );
buf ( n357983 , n37907 );
nor ( n357984 , n357978 , n357983 );
not ( n37910 , n357984 );
not ( n357986 , n37910 );
not ( n357987 , n592 );
nor ( n37913 , n357987 , n23996 );
buf ( n357989 , n37913 );
buf ( n357990 , n357905 );
xor ( n37916 , n357989 , n357990 );
buf ( n357992 , n343863 );
not ( n37918 , n357992 );
buf ( n357994 , n37632 );
not ( n357995 , n357994 );
or ( n37921 , n37918 , n357995 );
nand ( n357997 , n37749 , n23889 );
buf ( n357998 , n357997 );
nand ( n37924 , n37921 , n357998 );
buf ( n37925 , n37924 );
buf ( n358001 , n37925 );
xnor ( n37927 , n37916 , n358001 );
buf ( n37928 , n37927 );
buf ( n358004 , n37928 );
buf ( n358005 , n344400 );
not ( n37931 , n358005 );
buf ( n358007 , n604 );
not ( n358008 , n358007 );
buf ( n358009 , n355612 );
not ( n358010 , n358009 );
or ( n37936 , n358008 , n358010 );
buf ( n358012 , n23530 );
buf ( n358013 , n334537 );
nand ( n358014 , n358012 , n358013 );
buf ( n358015 , n358014 );
buf ( n358016 , n358015 );
nand ( n358017 , n37936 , n358016 );
buf ( n358018 , n358017 );
buf ( n358019 , n358018 );
not ( n358020 , n358019 );
or ( n358021 , n37931 , n358020 );
buf ( n358022 , n357747 );
buf ( n358023 , n344338 );
nand ( n358024 , n358022 , n358023 );
buf ( n358025 , n358024 );
buf ( n358026 , n358025 );
nand ( n358027 , n358021 , n358026 );
buf ( n358028 , n358027 );
buf ( n358029 , n358028 );
xor ( n358030 , n358004 , n358029 );
not ( n37956 , n343595 );
not ( n358032 , n37274 );
or ( n358033 , n37956 , n358032 );
nand ( n37959 , n358033 , n357922 );
not ( n358035 , n37959 );
not ( n37961 , n357905 );
or ( n37962 , n358035 , n37961 );
buf ( n358038 , n37848 );
buf ( n358039 , n357905 );
or ( n358040 , n358038 , n358039 );
buf ( n358041 , n37841 );
nand ( n358042 , n358040 , n358041 );
buf ( n358043 , n358042 );
nand ( n37969 , n37962 , n358043 );
buf ( n358045 , n37969 );
xnor ( n37971 , n358030 , n358045 );
buf ( n358047 , n37971 );
buf ( n358048 , n358047 );
buf ( n37974 , n358048 );
buf ( n358050 , n37974 );
buf ( n358051 , n23911 );
not ( n358052 , n358051 );
buf ( n358053 , n357779 );
not ( n358054 , n358053 );
or ( n37980 , n358052 , n358054 );
buf ( n358056 , n357293 );
buf ( n358057 , n343948 );
nand ( n37983 , n358056 , n358057 );
buf ( n37984 , n37983 );
buf ( n358060 , n37984 );
nand ( n358061 , n37980 , n358060 );
buf ( n358062 , n358061 );
buf ( n358063 , n358062 );
not ( n358064 , n358063 );
buf ( n358065 , n357423 );
not ( n358066 , n358065 );
buf ( n358067 , n358066 );
buf ( n37993 , n358067 );
not ( n37994 , n37993 );
buf ( n37995 , n356913 );
not ( n37996 , n37995 );
and ( n37997 , n37994 , n37996 );
buf ( n358073 , n358018 );
buf ( n358074 , n344338 );
and ( n358075 , n358073 , n358074 );
nor ( n38001 , n37997 , n358075 );
buf ( n358077 , n38001 );
buf ( n38003 , n358077 );
not ( n358079 , n38003 );
buf ( n358080 , n358079 );
buf ( n358081 , n358080 );
not ( n358082 , n358081 );
or ( n38008 , n358064 , n358082 );
buf ( n358084 , n358062 );
not ( n358085 , n358084 );
buf ( n358086 , n358085 );
buf ( n358087 , n358086 );
not ( n358088 , n358087 );
buf ( n358089 , n358077 );
not ( n38015 , n358089 );
or ( n358091 , n358088 , n38015 );
buf ( n358092 , n357275 );
not ( n38018 , n358092 );
buf ( n358094 , n37234 );
not ( n38020 , n358094 );
or ( n38021 , n38018 , n38020 );
buf ( n358097 , n357325 );
buf ( n358098 , n357275 );
not ( n38024 , n358098 );
buf ( n358100 , n357306 );
nand ( n358101 , n38024 , n358100 );
buf ( n358102 , n358101 );
buf ( n38028 , n358102 );
nand ( n38029 , n358097 , n38028 );
buf ( n38030 , n38029 );
buf ( n358106 , n38030 );
nand ( n38032 , n38021 , n358106 );
buf ( n38033 , n38032 );
buf ( n358109 , n38033 );
nand ( n38035 , n358091 , n358109 );
buf ( n358111 , n38035 );
buf ( n358112 , n358111 );
nand ( n38038 , n38008 , n358112 );
buf ( n358114 , n38038 );
not ( n38040 , n358114 );
nand ( n358116 , n358050 , n38040 );
not ( n38042 , n358116 );
or ( n38043 , n357986 , n38042 );
buf ( n358119 , n358050 );
not ( n38045 , n358119 );
buf ( n358121 , n358114 );
nand ( n38047 , n38045 , n358121 );
buf ( n358123 , n38047 );
nand ( n358124 , n38043 , n358123 );
xor ( n38050 , n357879 , n358124 );
not ( n358126 , n37969 );
buf ( n38052 , n37928 );
buf ( n38053 , n38052 );
buf ( n38054 , n38053 );
or ( n358130 , n38054 , n358028 );
not ( n38056 , n358130 );
or ( n358132 , n358126 , n38056 );
buf ( n358133 , n358028 );
buf ( n358134 , n358133 );
buf ( n358135 , n38054 );
nand ( n358136 , n358134 , n358135 );
buf ( n358137 , n358136 );
nand ( n358138 , n358132 , n358137 );
buf ( n358139 , n358138 );
buf ( n358140 , n37913 );
not ( n358141 , n358140 );
buf ( n358142 , n357905 );
nand ( n358143 , n358141 , n358142 );
buf ( n358144 , n358143 );
buf ( n358145 , n358144 );
not ( n358146 , n358145 );
buf ( n358147 , n37925 );
not ( n38073 , n358147 );
or ( n358149 , n358146 , n38073 );
buf ( n358150 , n357905 );
not ( n38076 , n358150 );
buf ( n358152 , n37913 );
nand ( n38078 , n38076 , n358152 );
buf ( n358154 , n38078 );
buf ( n358155 , n358154 );
nand ( n358156 , n358149 , n358155 );
buf ( n358157 , n358156 );
buf ( n358158 , n358157 );
not ( n358159 , n343531 );
buf ( n358160 , n602 );
not ( n358161 , n358160 );
buf ( n358162 , n355612 );
not ( n38088 , n358162 );
or ( n358164 , n358161 , n38088 );
buf ( n358165 , n356993 );
not ( n38091 , n358165 );
buf ( n358167 , n343553 );
nand ( n358168 , n38091 , n358167 );
buf ( n358169 , n358168 );
buf ( n358170 , n358169 );
nand ( n38096 , n358164 , n358170 );
buf ( n358172 , n38096 );
not ( n38098 , n358172 );
or ( n358174 , n358159 , n38098 );
nand ( n38100 , n357797 , n602 );
nand ( n358176 , n355596 , n37720 );
nand ( n38102 , n38100 , n358176 , n343595 );
nand ( n358178 , n358174 , n38102 );
not ( n358179 , n358178 );
buf ( n358180 , n358179 );
not ( n358181 , n358180 );
buf ( n358182 , n358181 );
buf ( n358183 , n358182 );
xor ( n358184 , n358158 , n358183 );
buf ( n38110 , n357606 );
buf ( n358186 , n23681 );
not ( n358187 , n358186 );
buf ( n358188 , n357680 );
not ( n38114 , n358188 );
or ( n358190 , n358187 , n38114 );
buf ( n38116 , n357856 );
buf ( n38117 , n343765 );
nand ( n358193 , n38116 , n38117 );
buf ( n358194 , n358193 );
buf ( n358195 , n358194 );
nand ( n38121 , n358190 , n358195 );
buf ( n358197 , n38121 );
buf ( n358198 , n358197 );
xor ( n358199 , n38110 , n358198 );
buf ( n358200 , n344015 );
not ( n38126 , n358200 );
buf ( n358202 , n357630 );
not ( n358203 , n358202 );
or ( n38129 , n38126 , n358203 );
buf ( n358205 , n357967 );
buf ( n358206 , n344018 );
nand ( n38132 , n358205 , n358206 );
buf ( n38133 , n38132 );
buf ( n358209 , n38133 );
nand ( n38135 , n38129 , n358209 );
buf ( n38136 , n38135 );
buf ( n358212 , n38136 );
and ( n38138 , n358199 , n358212 );
and ( n358214 , n38110 , n358198 );
or ( n358215 , n38138 , n358214 );
buf ( n358216 , n358215 );
buf ( n358217 , n358216 );
xor ( n358218 , n358184 , n358217 );
buf ( n358219 , n358218 );
buf ( n358220 , n358219 );
xor ( n38146 , n358139 , n358220 );
not ( n358222 , n357948 );
not ( n358223 , n358222 );
not ( n38149 , n357937 );
nand ( n358225 , n357976 , n38149 );
not ( n358226 , n358225 );
or ( n38152 , n358223 , n358226 );
nor ( n358228 , n38149 , n357976 );
not ( n38154 , n358228 );
nand ( n358230 , n38152 , n38154 );
not ( n38156 , n358230 );
xor ( n38157 , n38110 , n358198 );
xor ( n358233 , n38157 , n358212 );
buf ( n358234 , n358233 );
not ( n38160 , n358234 );
or ( n358236 , n38156 , n38160 );
buf ( n358237 , n358234 );
not ( n38163 , n358237 );
buf ( n38164 , n38163 );
not ( n358240 , n38164 );
not ( n38166 , n358230 );
not ( n38167 , n38166 );
or ( n358243 , n358240 , n38167 );
buf ( n358244 , n357874 );
buf ( n358245 , n37717 );
xor ( n38171 , n358244 , n358245 );
buf ( n358247 , n37738 );
xor ( n38173 , n38171 , n358247 );
buf ( n358249 , n38173 );
nand ( n358250 , n358243 , n358249 );
nand ( n358251 , n358236 , n358250 );
buf ( n358252 , n358251 );
xor ( n358253 , n38146 , n358252 );
buf ( n358254 , n358253 );
xor ( n38180 , n38050 , n358254 );
xor ( n358256 , n358234 , n358230 );
xnor ( n358257 , n358256 , n358249 );
buf ( n358258 , n358257 );
not ( n358259 , n358258 );
or ( n358260 , n37425 , n37402 );
not ( n38186 , n358260 );
not ( n358262 , n37439 );
or ( n358263 , n38186 , n358262 );
nand ( n358264 , n37425 , n37402 );
nand ( n38190 , n358263 , n358264 );
not ( n358266 , n38190 );
not ( n38192 , n37267 );
not ( n358268 , n357328 );
nand ( n38194 , n38192 , n358268 );
and ( n358270 , n38194 , n357449 );
nor ( n38196 , n358268 , n38192 );
nor ( n38197 , n358270 , n38196 );
buf ( n358273 , n38197 );
not ( n358274 , n358273 );
buf ( n358275 , n358274 );
not ( n358276 , n358275 );
or ( n38202 , n358266 , n358276 );
buf ( n358278 , n38190 );
not ( n38204 , n358278 );
buf ( n358280 , n38204 );
buf ( n358281 , n358280 );
not ( n38207 , n358281 );
buf ( n358283 , n38197 );
not ( n38209 , n358283 );
or ( n38210 , n38207 , n38209 );
buf ( n358286 , n358062 );
buf ( n358287 , n358080 );
xor ( n38213 , n358286 , n358287 );
buf ( n358289 , n38033 );
xor ( n38215 , n38213 , n358289 );
buf ( n358291 , n38215 );
buf ( n358292 , n358291 );
nand ( n38218 , n38210 , n358292 );
buf ( n358294 , n38218 );
nand ( n38220 , n38202 , n358294 );
buf ( n358296 , n38220 );
nand ( n358297 , n358259 , n358296 );
buf ( n358298 , n358297 );
not ( n38224 , n358257 );
buf ( n38225 , n38220 );
not ( n38226 , n38225 );
buf ( n38227 , n38226 );
not ( n358303 , n38227 );
or ( n358304 , n38224 , n358303 );
not ( n38230 , n357984 );
not ( n358306 , n38040 );
not ( n358307 , n358047 );
not ( n38233 , n358307 );
or ( n358309 , n358306 , n38233 );
nand ( n358310 , n358047 , n358114 );
nand ( n38236 , n358309 , n358310 );
not ( n38237 , n38236 );
or ( n38238 , n38230 , n38237 );
not ( n38239 , n38236 );
nand ( n38240 , n38239 , n37910 );
nand ( n38241 , n38238 , n38240 );
buf ( n38242 , n38241 );
nand ( n38243 , n358304 , n38242 );
nand ( n38244 , n358298 , n38243 );
nor ( n358320 , n38180 , n38244 );
not ( n38246 , n358320 );
xor ( n358322 , n357609 , n357637 );
and ( n358323 , n358322 , n357690 );
and ( n38249 , n357609 , n357637 );
or ( n358325 , n358323 , n38249 );
buf ( n358326 , n357750 );
not ( n38252 , n358326 );
buf ( n358328 , n357729 );
not ( n358329 , n358328 );
buf ( n358330 , n358329 );
buf ( n358331 , n358330 );
not ( n358332 , n358331 );
or ( n358333 , n38252 , n358332 );
buf ( n358334 , n357753 );
not ( n358335 , n358334 );
buf ( n358336 , n357729 );
not ( n38262 , n358336 );
or ( n358338 , n358335 , n38262 );
buf ( n358339 , n357708 );
nand ( n358340 , n358338 , n358339 );
buf ( n358341 , n358340 );
buf ( n358342 , n358341 );
nand ( n38268 , n358333 , n358342 );
buf ( n358344 , n38268 );
xor ( n358345 , n358325 , n358344 );
buf ( n358346 , n23911 );
not ( n38272 , n358346 );
buf ( n358348 , n598 );
not ( n358349 , n358348 );
buf ( n358350 , n356434 );
not ( n358351 , n358350 );
or ( n358352 , n358349 , n358351 );
buf ( n358353 , n356431 );
buf ( n358354 , n343953 );
nand ( n358355 , n358353 , n358354 );
buf ( n358356 , n358355 );
buf ( n358357 , n358356 );
nand ( n358358 , n358352 , n358357 );
buf ( n358359 , n358358 );
buf ( n358360 , n358359 );
not ( n38286 , n358360 );
or ( n38287 , n38272 , n38286 );
buf ( n358363 , n37640 );
not ( n358364 , n358363 );
buf ( n358365 , n343948 );
nand ( n358366 , n358364 , n358365 );
buf ( n358367 , n358366 );
buf ( n358368 , n358367 );
nand ( n358369 , n38287 , n358368 );
buf ( n358370 , n358369 );
buf ( n358371 , n358370 );
xor ( n38297 , n37572 , n357658 );
and ( n358373 , n38297 , n357688 );
and ( n358374 , n37572 , n357658 );
or ( n38300 , n358373 , n358374 );
buf ( n358376 , n38300 );
buf ( n358377 , n358376 );
xor ( n38303 , n358371 , n358377 );
buf ( n358379 , n343863 );
not ( n38305 , n358379 );
and ( n358381 , n596 , n350815 );
not ( n358382 , n596 );
and ( n358383 , n358382 , n355991 );
or ( n358384 , n358381 , n358383 );
buf ( n358385 , n358384 );
not ( n358386 , n358385 );
or ( n358387 , n38305 , n358386 );
buf ( n358388 , n37628 );
buf ( n358389 , n23889 );
nand ( n358390 , n358388 , n358389 );
buf ( n358391 , n358390 );
buf ( n358392 , n358391 );
nand ( n358393 , n358387 , n358392 );
buf ( n358394 , n358393 );
buf ( n358395 , n358394 );
xor ( n358396 , n38303 , n358395 );
buf ( n358397 , n358396 );
xor ( n38318 , n358345 , n358397 );
not ( n358399 , n38318 );
not ( n38320 , n357764 );
not ( n38321 , n37622 );
or ( n358402 , n38320 , n38321 );
not ( n358403 , n37622 );
nand ( n38324 , n358403 , n37691 );
nand ( n358405 , n38324 , n37803 );
nand ( n358406 , n358402 , n358405 );
buf ( n358407 , n344015 );
not ( n358408 , n358407 );
buf ( n358409 , n600 );
not ( n38330 , n358409 );
buf ( n358411 , n357413 );
not ( n38332 , n358411 );
or ( n358413 , n38330 , n38332 );
buf ( n358414 , n355593 );
buf ( n358415 , n23906 );
nand ( n358416 , n358414 , n358415 );
buf ( n358417 , n358416 );
buf ( n358418 , n358417 );
nand ( n358419 , n358413 , n358418 );
buf ( n358420 , n358419 );
buf ( n358421 , n358420 );
not ( n358422 , n358421 );
or ( n358423 , n358408 , n358422 );
buf ( n358424 , n344018 );
buf ( n358425 , n357623 );
nand ( n358426 , n358424 , n358425 );
buf ( n358427 , n358426 );
buf ( n358428 , n358427 );
nand ( n38349 , n358423 , n358428 );
buf ( n358430 , n38349 );
buf ( n38351 , n358430 );
not ( n358432 , n23613 );
not ( n38353 , n356681 );
or ( n358434 , n358432 , n38353 );
nand ( n358435 , n37581 , n344705 );
nand ( n38356 , n358434 , n358435 );
xor ( n358437 , n36640 , n38356 );
buf ( n358438 , n23681 );
not ( n38359 , n358438 );
buf ( n358440 , n594 );
not ( n38361 , n358440 );
buf ( n358442 , n344353 );
not ( n38363 , n358442 );
or ( n38364 , n38361 , n38363 );
buf ( n358445 , n357286 );
buf ( n358446 , n343632 );
nand ( n38367 , n358445 , n358446 );
buf ( n358448 , n38367 );
buf ( n358449 , n358448 );
nand ( n38370 , n38364 , n358449 );
buf ( n358451 , n38370 );
buf ( n358452 , n358451 );
not ( n38373 , n358452 );
or ( n358454 , n38359 , n38373 );
buf ( n358455 , n357665 );
buf ( n358456 , n343765 );
nand ( n38377 , n358455 , n358456 );
buf ( n358458 , n38377 );
buf ( n358459 , n358458 );
nand ( n38380 , n358454 , n358459 );
buf ( n358461 , n38380 );
xnor ( n38382 , n358437 , n358461 );
buf ( n358463 , n38382 );
xor ( n358464 , n38351 , n358463 );
buf ( n358465 , n343595 );
not ( n358466 , n358465 );
buf ( n358467 , n358172 );
not ( n358468 , n358467 );
or ( n38389 , n358466 , n358468 );
buf ( n358470 , n602 );
not ( n358471 , n358470 );
buf ( n358472 , n37410 );
not ( n358473 , n358472 );
or ( n358474 , n358471 , n358473 );
buf ( n358475 , n334531 );
buf ( n358476 , n343553 );
nand ( n358477 , n358475 , n358476 );
buf ( n358478 , n358477 );
buf ( n358479 , n358478 );
nand ( n38400 , n358474 , n358479 );
buf ( n358481 , n38400 );
buf ( n358482 , n358481 );
buf ( n358483 , n343531 );
nand ( n38404 , n358482 , n358483 );
buf ( n358485 , n38404 );
buf ( n358486 , n358485 );
nand ( n358487 , n38389 , n358486 );
buf ( n358488 , n358487 );
buf ( n358489 , n358488 );
xor ( n38410 , n358464 , n358489 );
buf ( n358491 , n38410 );
buf ( n358492 , n358157 );
not ( n38413 , n358492 );
buf ( n358494 , n358182 );
not ( n38415 , n358494 );
or ( n358496 , n38413 , n38415 );
buf ( n358497 , n358157 );
not ( n38418 , n358497 );
buf ( n358499 , n38418 );
buf ( n358500 , n358499 );
not ( n358501 , n358500 );
buf ( n358502 , n358179 );
not ( n358503 , n358502 );
or ( n358504 , n358501 , n358503 );
buf ( n358505 , n358216 );
nand ( n358506 , n358504 , n358505 );
buf ( n358507 , n358506 );
buf ( n358508 , n358507 );
nand ( n358509 , n358496 , n358508 );
buf ( n358510 , n358509 );
not ( n358511 , n358510 );
and ( n38432 , n358491 , n358511 );
not ( n38433 , n358491 );
and ( n38434 , n38433 , n358510 );
nor ( n38435 , n38432 , n38434 );
not ( n38436 , n38435 );
and ( n38437 , n358406 , n38436 );
not ( n38438 , n358406 );
and ( n358519 , n38438 , n38435 );
nor ( n38440 , n38437 , n358519 );
not ( n38441 , n38440 );
or ( n358522 , n358399 , n38441 );
not ( n38443 , n38440 );
not ( n358524 , n38318 );
nand ( n38445 , n38443 , n358524 );
nand ( n38446 , n358522 , n38445 );
xor ( n38447 , n358139 , n358220 );
and ( n358528 , n38447 , n358252 );
and ( n358529 , n358139 , n358220 );
or ( n38450 , n358528 , n358529 );
buf ( n358531 , n38450 );
not ( n358532 , n358531 );
and ( n38453 , n38446 , n358532 );
not ( n358534 , n38446 );
and ( n358535 , n358534 , n358531 );
nor ( n358536 , n38453 , n358535 );
not ( n38457 , n358536 );
xor ( n358538 , n357879 , n358124 );
and ( n358539 , n358538 , n358254 );
and ( n38460 , n357879 , n358124 );
or ( n358541 , n358539 , n38460 );
not ( n358542 , n358541 );
nand ( n38463 , n38457 , n358542 );
nand ( n38464 , n38246 , n38463 );
buf ( n38465 , n38464 );
buf ( n358546 , n38190 );
buf ( n358547 , n358291 );
xor ( n38468 , n358546 , n358547 );
buf ( n358549 , n358275 );
xor ( n38470 , n38468 , n358549 );
buf ( n38471 , n38470 );
not ( n358552 , n38471 );
buf ( n38473 , n37823 );
xor ( n358554 , n357926 , n38473 );
not ( n38475 , n37902 );
xnor ( n38476 , n358554 , n38475 );
not ( n38477 , n38476 );
xor ( n358558 , n37385 , n37440 );
and ( n38479 , n358558 , n37451 );
and ( n358560 , n37385 , n37440 );
or ( n358561 , n38479 , n358560 );
buf ( n358562 , n358561 );
not ( n38483 , n358562 );
buf ( n38484 , n38483 );
not ( n358565 , n38484 );
or ( n38486 , n38477 , n358565 );
not ( n358567 , n38476 );
nand ( n358568 , n358567 , n358561 );
nand ( n38489 , n38486 , n358568 );
nand ( n38490 , n358552 , n38489 );
not ( n358571 , n38490 );
not ( n358572 , n358552 );
not ( n38493 , n38489 );
nand ( n358574 , n358572 , n38493 );
not ( n358575 , n358574 );
or ( n38496 , n358571 , n358575 );
buf ( n358577 , n37381 );
buf ( n358578 , n358577 );
buf ( n358579 , n358578 );
not ( n358580 , n358579 );
buf ( n358581 , n357521 );
not ( n358582 , n358581 );
buf ( n358583 , n358582 );
not ( n38504 , n358583 );
not ( n358585 , n38504 );
or ( n358586 , n358580 , n358585 );
not ( n38507 , n358579 );
not ( n38508 , n38507 );
not ( n358589 , n358583 );
or ( n38510 , n38508 , n358589 );
nand ( n38511 , n38510 , n37464 );
nand ( n358592 , n358586 , n38511 );
not ( n358593 , n358592 );
nand ( n358594 , n38496 , n358593 );
buf ( n358595 , n358594 );
not ( n358596 , n38484 );
not ( n358597 , n38476 );
or ( n38518 , n358596 , n358597 );
nand ( n358599 , n38518 , n38471 );
buf ( n358600 , n358568 );
nand ( n38521 , n358599 , n358600 );
buf ( n358602 , n38521 );
not ( n38523 , n358602 );
xor ( n358604 , n358257 , n38241 );
xnor ( n358605 , n358604 , n38227 );
buf ( n358606 , n358605 );
nand ( n38527 , n38523 , n358606 );
buf ( n358608 , n38527 );
buf ( n358609 , n358608 );
nand ( n358610 , n358595 , n358609 );
buf ( n358611 , n358610 );
buf ( n358612 , n358611 );
nor ( n38533 , n38465 , n358612 );
buf ( n358614 , n38533 );
not ( n358615 , n358614 );
or ( n38536 , n37500 , n358615 );
not ( n38537 , n358592 );
nand ( n38538 , n358574 , n38490 );
nor ( n38539 , n38537 , n38538 );
nand ( n38540 , n358608 , n38539 );
not ( n38541 , n38540 );
nand ( n358622 , n358536 , n358541 );
buf ( n358623 , n358622 );
not ( n38544 , n358623 );
buf ( n358625 , n358605 );
not ( n38546 , n358625 );
buf ( n358627 , n38546 );
buf ( n358628 , n358627 );
buf ( n358629 , n38521 );
nand ( n358630 , n358628 , n358629 );
buf ( n358631 , n358630 );
nand ( n38552 , n38180 , n38244 );
nand ( n358633 , n358631 , n38552 );
buf ( n38554 , n358633 );
nor ( n38555 , n38544 , n38554 );
buf ( n38556 , n38555 );
not ( n358637 , n38556 );
or ( n38558 , n38541 , n358637 );
buf ( n358639 , n38463 );
not ( n358640 , n358639 );
not ( n358641 , n38180 );
not ( n38562 , n38244 );
nand ( n358643 , n358641 , n38562 );
buf ( n358644 , n358643 );
not ( n38565 , n358644 );
or ( n358646 , n358640 , n38565 );
buf ( n358647 , n358622 );
buf ( n38568 , n358647 );
buf ( n358649 , n38568 );
buf ( n358650 , n358649 );
nand ( n358651 , n358646 , n358650 );
buf ( n358652 , n358651 );
nand ( n38573 , n38558 , n358652 );
nand ( n358654 , n38536 , n38573 );
not ( n358655 , n23911 );
not ( n38576 , n356640 );
or ( n358657 , n358655 , n38576 );
buf ( n358658 , n358359 );
buf ( n358659 , n343948 );
nand ( n358660 , n358658 , n358659 );
buf ( n358661 , n358660 );
nand ( n38582 , n358657 , n358661 );
not ( n38583 , n23681 );
not ( n38584 , n356599 );
or ( n358665 , n38583 , n38584 );
buf ( n358666 , n358451 );
buf ( n358667 , n343765 );
nand ( n38588 , n358666 , n358667 );
buf ( n358669 , n38588 );
nand ( n358670 , n358665 , n358669 );
buf ( n358671 , n358670 );
not ( n358672 , n23889 );
not ( n38593 , n358384 );
or ( n358674 , n358672 , n38593 );
buf ( n358675 , n356748 );
buf ( n358676 , n343863 );
nand ( n38597 , n358675 , n358676 );
buf ( n358678 , n38597 );
nand ( n358679 , n358674 , n358678 );
buf ( n38600 , n358679 );
and ( n38601 , n358671 , n38600 );
not ( n358682 , n358671 );
not ( n358683 , n358679 );
buf ( n358684 , n358683 );
and ( n358685 , n358682 , n358684 );
nor ( n358686 , n38601 , n358685 );
buf ( n358687 , n358686 );
xor ( n38608 , n38582 , n358687 );
buf ( n358689 , n38608 );
buf ( n358690 , n356698 );
buf ( n358691 , n36640 );
xor ( n358692 , n358690 , n358691 );
buf ( n358693 , n356688 );
xnor ( n38614 , n358692 , n358693 );
buf ( n38615 , n38614 );
buf ( n38616 , n38615 );
not ( n358697 , n38616 );
buf ( n358698 , n358697 );
buf ( n358699 , n358698 );
or ( n358700 , n358689 , n358699 );
xor ( n38621 , n358371 , n358377 );
and ( n358702 , n38621 , n358395 );
and ( n38623 , n358371 , n358377 );
or ( n358704 , n358702 , n38623 );
buf ( n358705 , n358704 );
buf ( n358706 , n358705 );
nand ( n38627 , n358700 , n358706 );
buf ( n358708 , n38627 );
buf ( n358709 , n358708 );
buf ( n358710 , n38608 );
buf ( n358711 , n358698 );
nand ( n358712 , n358710 , n358711 );
buf ( n38630 , n358712 );
buf ( n358714 , n38630 );
nand ( n358715 , n358709 , n358714 );
buf ( n358716 , n358715 );
buf ( n358717 , n358716 );
not ( n38635 , n356704 );
not ( n38636 , n36553 );
or ( n358720 , n38635 , n38636 );
not ( n38638 , n356704 );
nand ( n38639 , n38638 , n356606 );
nand ( n358723 , n358720 , n38639 );
and ( n38641 , n358723 , n356648 );
not ( n38642 , n358723 );
and ( n358726 , n38642 , n356647 );
nor ( n358727 , n38641 , n358726 );
buf ( n358728 , n344018 );
not ( n38646 , n358728 );
buf ( n358730 , n358420 );
not ( n358731 , n358730 );
or ( n358732 , n38646 , n358731 );
buf ( n358733 , n600 );
not ( n38651 , n358733 );
buf ( n358735 , n356993 );
not ( n358736 , n358735 );
or ( n38654 , n38651 , n358736 );
buf ( n358738 , n356999 );
buf ( n358739 , n23906 );
nand ( n358740 , n358738 , n358739 );
buf ( n358741 , n358740 );
buf ( n358742 , n358741 );
nand ( n38660 , n38654 , n358742 );
buf ( n358744 , n38660 );
buf ( n358745 , n358744 );
buf ( n358746 , n344015 );
nand ( n38664 , n358745 , n358746 );
buf ( n358748 , n38664 );
buf ( n358749 , n358748 );
nand ( n358750 , n358732 , n358749 );
buf ( n358751 , n358750 );
buf ( n358752 , n348539 );
not ( n358753 , n358752 );
buf ( n358754 , n346090 );
not ( n38672 , n358754 );
or ( n358756 , n358753 , n38672 );
buf ( n358757 , n358481 );
nand ( n358758 , n358756 , n358757 );
buf ( n358759 , n358758 );
or ( n38677 , n358751 , n358759 );
nand ( n358761 , n356654 , n38356 );
buf ( n358762 , n36640 );
not ( n38680 , n358762 );
not ( n358764 , n38356 );
buf ( n358765 , n358764 );
not ( n38683 , n358765 );
or ( n358767 , n38680 , n38683 );
buf ( n358768 , n358461 );
nand ( n38686 , n358767 , n358768 );
buf ( n358770 , n38686 );
nand ( n358771 , n358761 , n358770 );
nand ( n358772 , n38677 , n358771 );
buf ( n358773 , n358772 );
buf ( n358774 , n358751 );
buf ( n358775 , n358759 );
nand ( n38693 , n358774 , n358775 );
buf ( n38694 , n38693 );
buf ( n38695 , n38694 );
nand ( n38696 , n358773 , n38695 );
buf ( n358780 , n38696 );
and ( n38698 , n358727 , n358780 );
not ( n358782 , n358727 );
not ( n358783 , n358780 );
and ( n38701 , n358782 , n358783 );
nor ( n38702 , n38698 , n38701 );
buf ( n358786 , n36450 );
not ( n358787 , n358786 );
buf ( n358788 , n344014 );
not ( n38706 , n358788 );
and ( n38707 , n358787 , n38706 );
buf ( n358791 , n358744 );
buf ( n358792 , n344018 );
and ( n358793 , n358791 , n358792 );
nor ( n38711 , n38707 , n358793 );
buf ( n358795 , n38711 );
buf ( n358796 , n358795 );
xnor ( n358797 , n356405 , n356756 );
not ( n38715 , n358797 );
and ( n38716 , n356753 , n38715 );
not ( n358800 , n356753 );
and ( n358801 , n358800 , n358797 );
nor ( n38719 , n38716 , n358801 );
buf ( n358803 , n38719 );
xor ( n358804 , n358796 , n358803 );
not ( n358805 , n23911 );
not ( n38723 , n356640 );
or ( n38724 , n358805 , n38723 );
nand ( n358808 , n38724 , n358661 );
not ( n38726 , n358808 );
nand ( n38727 , n38726 , n358683 );
and ( n358811 , n38727 , n358670 );
and ( n38729 , n358679 , n358808 );
nor ( n38730 , n358811 , n38729 );
buf ( n358814 , n38730 );
xor ( n38732 , n358804 , n358814 );
buf ( n358816 , n38732 );
xor ( n38734 , n38702 , n358816 );
buf ( n358818 , n38734 );
xor ( n38736 , n358717 , n358818 );
xor ( n358820 , n38351 , n358463 );
and ( n358821 , n358820 , n358489 );
and ( n38739 , n38351 , n358463 );
or ( n38740 , n358821 , n38739 );
buf ( n358824 , n38740 );
buf ( n358825 , n358824 );
not ( n38743 , n358825 );
xor ( n38744 , n358759 , n358771 );
xnor ( n38745 , n38744 , n358751 );
buf ( n358829 , n38745 );
nand ( n38747 , n38743 , n358829 );
buf ( n358831 , n38747 );
buf ( n358832 , n358831 );
not ( n358833 , n358832 );
or ( n38751 , n358397 , n358344 );
nand ( n358835 , n38751 , n358325 );
buf ( n358836 , n358397 );
buf ( n358837 , n358344 );
nand ( n358838 , n358836 , n358837 );
buf ( n358839 , n358838 );
nand ( n38757 , n358835 , n358839 );
buf ( n358841 , n38757 );
not ( n358842 , n358841 );
or ( n38760 , n358833 , n358842 );
buf ( n358844 , n38745 );
not ( n38762 , n358844 );
buf ( n358846 , n358824 );
nand ( n358847 , n38762 , n358846 );
buf ( n358848 , n358847 );
buf ( n358849 , n358848 );
nand ( n38767 , n38760 , n358849 );
buf ( n358851 , n38767 );
buf ( n358852 , n358851 );
xor ( n38770 , n38736 , n358852 );
buf ( n358854 , n38770 );
not ( n358855 , n358854 );
buf ( n38773 , n358855 );
buf ( n358857 , n38615 );
buf ( n358858 , n358705 );
xor ( n358859 , n358857 , n358858 );
buf ( n358860 , n38608 );
xnor ( n358861 , n358859 , n358860 );
buf ( n358862 , n358861 );
buf ( n358863 , n358862 );
not ( n358864 , n358406 );
buf ( n358865 , n358491 );
buf ( n38783 , n358865 );
buf ( n358867 , n38783 );
buf ( n358868 , n358867 );
not ( n358869 , n358868 );
buf ( n358870 , n358869 );
buf ( n358871 , n358870 );
buf ( n358872 , n358511 );
nand ( n358873 , n358871 , n358872 );
buf ( n358874 , n358873 );
not ( n38792 , n358874 );
or ( n38793 , n358864 , n38792 );
buf ( n358877 , n358511 );
not ( n38795 , n358877 );
buf ( n358879 , n358867 );
nand ( n358880 , n38795 , n358879 );
buf ( n358881 , n358880 );
nand ( n358882 , n38793 , n358881 );
buf ( n358883 , n358882 );
xor ( n358884 , n358863 , n358883 );
buf ( n358885 , n358824 );
not ( n358886 , n358885 );
buf ( n358887 , n38745 );
not ( n38800 , n358887 );
or ( n38801 , n358886 , n38800 );
buf ( n358890 , n358824 );
buf ( n358891 , n38745 );
or ( n38804 , n358890 , n358891 );
nand ( n358893 , n38801 , n38804 );
buf ( n358894 , n358893 );
buf ( n358895 , n358894 );
buf ( n358896 , n38757 );
and ( n358897 , n358895 , n358896 );
not ( n358898 , n358895 );
buf ( n358899 , n38757 );
not ( n358900 , n358899 );
buf ( n358901 , n358900 );
buf ( n358902 , n358901 );
and ( n38815 , n358898 , n358902 );
nor ( n38816 , n358897 , n38815 );
buf ( n358905 , n38816 );
buf ( n358906 , n358905 );
and ( n38819 , n358884 , n358906 );
and ( n38820 , n358863 , n358883 );
or ( n38821 , n38819 , n38820 );
buf ( n358910 , n38821 );
buf ( n358911 , n358910 );
not ( n358912 , n358911 );
buf ( n358913 , n358912 );
buf ( n358914 , n358913 );
nand ( n38827 , n38773 , n358914 );
buf ( n358916 , n38827 );
buf ( n358917 , n358916 );
xor ( n358918 , n358863 , n358883 );
xor ( n358919 , n358918 , n358906 );
buf ( n358920 , n358919 );
not ( n38833 , n358920 );
buf ( n358922 , n38833 );
buf ( n358923 , n358531 );
not ( n38836 , n358923 );
buf ( n358925 , n38440 );
buf ( n358926 , n358925 );
not ( n38839 , n358926 );
or ( n358928 , n38836 , n38839 );
buf ( n358929 , n358925 );
buf ( n358930 , n358531 );
or ( n358931 , n358929 , n358930 );
buf ( n358932 , n38318 );
nand ( n358933 , n358931 , n358932 );
buf ( n38844 , n358933 );
buf ( n358935 , n38844 );
nand ( n358936 , n358928 , n358935 );
buf ( n358937 , n358936 );
buf ( n358938 , n358937 );
not ( n358939 , n358938 );
buf ( n358940 , n358939 );
buf ( n358941 , n358940 );
nand ( n358942 , n358922 , n358941 );
buf ( n358943 , n358942 );
buf ( n358944 , n358943 );
and ( n358945 , n358917 , n358944 );
buf ( n358946 , n358945 );
xor ( n358947 , n358796 , n358803 );
and ( n38858 , n358947 , n358814 );
and ( n38859 , n358796 , n358803 );
or ( n358950 , n38858 , n38859 );
buf ( n358951 , n358950 );
not ( n358952 , n358951 );
buf ( n358953 , n358727 );
and ( n38864 , n358783 , n358953 );
nor ( n358955 , n38864 , n358816 );
buf ( n358956 , n358780 );
not ( n358957 , n358956 );
buf ( n358958 , n358953 );
nor ( n38869 , n358957 , n358958 );
buf ( n38870 , n38869 );
nor ( n358961 , n358955 , n38870 );
and ( n358962 , n358952 , n358961 );
not ( n358963 , n358952 );
not ( n358964 , n358961 );
and ( n358965 , n358963 , n358964 );
nor ( n358966 , n358962 , n358965 );
not ( n358967 , n36659 );
not ( n358968 , n36527 );
or ( n38873 , n358967 , n358968 );
nand ( n358970 , n356780 , n356716 );
nand ( n38875 , n38873 , n358970 );
not ( n38876 , n38875 );
not ( n38877 , n356777 );
or ( n38878 , n38876 , n38877 );
or ( n38879 , n356777 , n38875 );
nand ( n358976 , n38878 , n38879 );
not ( n358977 , n358976 );
and ( n38882 , n358966 , n358977 );
not ( n358979 , n358966 );
and ( n38884 , n358979 , n358976 );
nor ( n38885 , n38882 , n38884 );
not ( n358982 , n38885 );
xor ( n358983 , n358717 , n358818 );
and ( n38888 , n358983 , n358852 );
and ( n358985 , n358717 , n358818 );
or ( n358986 , n38888 , n358985 );
buf ( n358987 , n358986 );
or ( n358988 , n358982 , n358987 );
nand ( n358989 , n358946 , n358988 );
xor ( n38894 , n356797 , n356809 );
xnor ( n358991 , n38894 , n36720 );
buf ( n358992 , n358991 );
nand ( n38897 , n358964 , n358952 );
not ( n38898 , n38897 );
not ( n38899 , n358976 );
or ( n38900 , n38898 , n38899 );
nand ( n38901 , n358961 , n358951 );
nand ( n38902 , n38900 , n38901 );
buf ( n358999 , n38902 );
and ( n38904 , n358992 , n358999 );
buf ( n359001 , n38904 );
nor ( n38906 , n358989 , n359001 );
nand ( n38907 , n358654 , n38906 );
buf ( n38908 , n358608 );
buf ( n38909 , n358594 );
nand ( n38910 , n38908 , n38909 );
buf ( n38911 , n38910 );
buf ( n359008 , n38911 );
buf ( n359009 , n38464 );
nor ( n359010 , n359008 , n359009 );
buf ( n359011 , n359010 );
not ( n359012 , n357557 );
not ( n38917 , n357535 );
or ( n359014 , n359012 , n38917 );
nand ( n38919 , n359014 , n351742 );
buf ( n359016 , n38919 );
buf ( n359017 , n357240 );
buf ( n359018 , n359017 );
buf ( n359019 , n359018 );
nand ( n359020 , n352110 , n359019 );
buf ( n359021 , n359020 );
nor ( n38926 , n359016 , n359021 );
buf ( n359023 , n38926 );
and ( n359024 , n359023 , n351407 );
nand ( n38929 , n38906 , n359011 , n359024 );
buf ( n359026 , n359001 );
not ( n359027 , n359026 );
buf ( n359028 , n359027 );
buf ( n359029 , n358855 );
buf ( n359030 , n358913 );
nand ( n38935 , n359029 , n359030 );
buf ( n359032 , n38935 );
buf ( n359033 , n359032 );
buf ( n359034 , n358854 );
buf ( n359035 , n358910 );
nand ( n38940 , n359034 , n359035 );
buf ( n359037 , n38940 );
buf ( n359038 , n359037 );
buf ( n359039 , n358920 );
buf ( n359040 , n358937 );
nand ( n38945 , n359039 , n359040 );
buf ( n359042 , n38945 );
buf ( n359043 , n359042 );
nand ( n359044 , n359038 , n359043 );
buf ( n359045 , n359044 );
buf ( n359046 , n359045 );
nand ( n38951 , n359033 , n359046 );
buf ( n359048 , n38951 );
buf ( n359049 , n359048 );
buf ( n359050 , n38885 );
not ( n38955 , n359050 );
buf ( n359052 , n358987 );
nor ( n359053 , n38955 , n359052 );
buf ( n359054 , n359053 );
buf ( n359055 , n359054 );
nor ( n38960 , n359049 , n359055 );
buf ( n359057 , n38960 );
and ( n359058 , n359028 , n359057 );
not ( n38963 , n38885 );
nand ( n38964 , n38963 , n358987 );
buf ( n359061 , n38964 );
not ( n38966 , n358991 );
not ( n38967 , n38902 );
nor ( n38968 , n38966 , n38967 );
buf ( n359065 , n38968 );
or ( n38970 , n359061 , n359065 );
buf ( n359067 , n38966 );
buf ( n359068 , n38967 );
nand ( n38973 , n359067 , n359068 );
buf ( n359070 , n38973 );
buf ( n359071 , n359070 );
nand ( n38976 , n38970 , n359071 );
buf ( n359073 , n38976 );
nor ( n38978 , n359058 , n359073 );
nand ( n359075 , n38907 , n38929 , n38978 );
not ( n38980 , n359075 );
or ( n38981 , n356858 , n38980 );
not ( n38982 , n356299 );
buf ( n38983 , n36516 );
buf ( n359080 , n356814 );
nand ( n359081 , n38983 , n359080 );
buf ( n359082 , n359081 );
buf ( n359083 , n359082 );
buf ( n359084 , n356853 );
or ( n359085 , n359083 , n359084 );
buf ( n359086 , n356833 );
buf ( n359087 , n356850 );
nand ( n359088 , n359086 , n359087 );
buf ( n359089 , n359088 );
buf ( n359090 , n359089 );
nand ( n359091 , n359085 , n359090 );
buf ( n359092 , n359091 );
not ( n359093 , n359092 );
or ( n359094 , n38982 , n359093 );
buf ( n359095 , n356147 );
buf ( n359096 , n356296 );
or ( n359097 , n359095 , n359096 );
buf ( n359098 , n359097 );
nand ( n359099 , n359094 , n359098 );
and ( n39004 , n359099 , n356320 );
not ( n359101 , n36283 );
nand ( n359102 , n359101 , n356309 );
not ( n39007 , n359102 );
nor ( n359104 , n39004 , n39007 );
nand ( n359105 , n38981 , n359104 );
not ( n39010 , n359105 );
or ( n39011 , n35954 , n39010 );
buf ( n359108 , n355983 );
not ( n359109 , n359108 );
buf ( n359110 , n355962 );
nand ( n359111 , n355876 , n355928 );
buf ( n359112 , n359111 );
or ( n39017 , n359110 , n359112 );
buf ( n359114 , n355935 );
buf ( n359115 , n355959 );
nand ( n39020 , n359114 , n359115 );
buf ( n39021 , n39020 );
buf ( n359118 , n39021 );
nand ( n39023 , n39017 , n359118 );
buf ( n359120 , n39023 );
buf ( n359121 , n359120 );
not ( n39026 , n359121 );
or ( n359123 , n359109 , n39026 );
buf ( n359124 , n355980 );
not ( n39029 , n359124 );
buf ( n359126 , n355972 );
nand ( n359127 , n39029 , n359126 );
buf ( n359128 , n359127 );
buf ( n359129 , n359128 );
nand ( n359130 , n359123 , n359129 );
buf ( n359131 , n359130 );
buf ( n359132 , n359131 );
not ( n359133 , n359132 );
buf ( n359134 , n359133 );
nand ( n39039 , n39011 , n359134 );
nand ( n359136 , n35622 , n39039 );
buf ( n359137 , n355652 );
not ( n39042 , n359137 );
buf ( n359139 , n355589 );
nor ( n39044 , n39042 , n359139 );
buf ( n359141 , n39044 );
not ( n39046 , n359141 );
nand ( n39047 , n359136 , n39046 );
not ( n359144 , n39047 );
buf ( n359145 , n359144 );
not ( n39050 , n359145 );
buf ( n359147 , n39050 );
xnor ( n359148 , n355582 , n359147 );
buf ( n359149 , n359148 );
buf ( n359150 , n355561 );
not ( n359151 , n359150 );
buf ( n359152 , n35531 );
nand ( n359153 , n359151 , n359152 );
buf ( n359154 , n359153 );
not ( n359155 , n355559 );
nor ( n359156 , n359154 , n359155 );
not ( n39061 , n359156 );
and ( n359158 , n35505 , n355530 );
nor ( n39063 , n359158 , n35513 );
nand ( n39064 , n35440 , n39063 );
buf ( n359161 , n39064 );
not ( n359162 , n359161 );
buf ( n359163 , n359162 );
buf ( n359164 , n359163 );
buf ( n359165 , n35397 );
not ( n39070 , n359165 );
buf ( n359167 , n34586 );
not ( n359168 , n359167 );
buf ( n359169 , n34684 );
not ( n359170 , n359169 );
or ( n39075 , n359168 , n359170 );
buf ( n359172 , n354737 );
nand ( n39077 , n39075 , n359172 );
buf ( n359174 , n39077 );
buf ( n359175 , n359174 );
nand ( n359176 , n39070 , n359175 );
buf ( n359177 , n359176 );
buf ( n359178 , n359177 );
nand ( n39083 , n359164 , n359178 );
buf ( n359180 , n39083 );
nand ( n39085 , n355519 , n35489 );
buf ( n359182 , n39085 );
not ( n39087 , n359182 );
buf ( n359184 , n355484 );
nand ( n359185 , n39087 , n359184 );
buf ( n359186 , n359185 );
buf ( n359187 , n359186 );
not ( n39092 , n359187 );
buf ( n359189 , n39092 );
or ( n359190 , n359180 , n359189 );
buf ( n359191 , n355093 );
buf ( n39096 , n359191 );
buf ( n359193 , n39096 );
nand ( n359194 , n359190 , n359193 );
not ( n359195 , n359194 );
or ( n39100 , n39061 , n359195 );
and ( n39101 , n359189 , n359193 );
nor ( n39102 , n39101 , n359155 );
not ( n359199 , n39102 );
nand ( n359200 , n359180 , n359193 );
not ( n39105 , n359200 );
or ( n359202 , n359199 , n39105 );
nand ( n359203 , n359202 , n359154 );
nand ( n39108 , n39100 , n359203 );
buf ( n359205 , n39108 );
not ( n359206 , n359205 );
buf ( n359207 , n359206 );
not ( n39112 , n359207 );
not ( n359209 , n355536 );
buf ( n359210 , n354643 );
not ( n39115 , n359210 );
buf ( n359212 , n354726 );
buf ( n359213 , n34699 );
and ( n39118 , n359212 , n359213 );
buf ( n359215 , n39118 );
buf ( n359216 , n359215 );
nand ( n359217 , n39115 , n359216 );
buf ( n359218 , n359217 );
buf ( n359219 , n359218 );
buf ( n359220 , n359215 );
not ( n359221 , n354615 );
buf ( n359222 , n359221 );
nand ( n39127 , n359220 , n359222 );
buf ( n359224 , n39127 );
buf ( n359225 , n359224 );
buf ( n359226 , n359215 );
not ( n39131 , n34680 );
buf ( n359228 , n39131 );
nand ( n359229 , n359226 , n359228 );
buf ( n359230 , n359229 );
buf ( n359231 , n359230 );
and ( n359232 , n355340 , n355427 , n354456 , n355412 );
buf ( n359233 , n359232 );
nand ( n39138 , n359219 , n359225 , n359231 , n359233 );
buf ( n39139 , n39138 );
or ( n359236 , n355411 , n35335 );
and ( n39141 , n359236 , n35494 );
nor ( n359238 , n39141 , n35502 );
buf ( n359239 , n359238 );
nand ( n39144 , n35510 , n35509 );
nand ( n359241 , n39144 , n355541 );
buf ( n359242 , n359241 );
nor ( n359243 , n359239 , n359242 );
buf ( n359244 , n359243 );
nand ( n359245 , n39139 , n359244 );
not ( n359246 , n359245 );
or ( n39151 , n359209 , n359246 );
buf ( n359248 , n342675 );
not ( n359249 , n359248 );
buf ( n359250 , n341897 );
buf ( n359251 , n359250 );
not ( n359252 , n359251 );
or ( n39157 , n359249 , n359252 );
buf ( n359254 , n355521 );
nand ( n359255 , n39157 , n359254 );
buf ( n359256 , n359255 );
not ( n39161 , n359256 );
buf ( n359258 , n355500 );
buf ( n359259 , n359258 );
buf ( n359260 , n359259 );
not ( n39165 , n359260 );
or ( n359262 , n39161 , n39165 );
not ( n359263 , n355515 );
not ( n359264 , n35478 );
or ( n39169 , n359263 , n359264 );
buf ( n359266 , n355461 );
not ( n359267 , n359266 );
buf ( n359268 , n359267 );
nand ( n359269 , n39169 , n359268 );
buf ( n359270 , n359269 );
not ( n39175 , n359270 );
buf ( n359272 , n39175 );
buf ( n359273 , n359272 );
buf ( n359274 , n359273 );
buf ( n359275 , n359274 );
nand ( n39180 , n359262 , n359275 );
nand ( n39181 , n355484 , n39180 );
nand ( n359278 , n39151 , n39181 );
buf ( n39183 , n359193 );
buf ( n359280 , n355559 );
nand ( n39185 , n39183 , n359280 );
buf ( n359282 , n39185 );
xnor ( n359283 , n359278 , n359282 );
not ( n39188 , n359283 );
or ( n39189 , n39112 , n39188 );
buf ( n359286 , n359283 );
not ( n359287 , n359286 );
buf ( n359288 , n39108 );
nand ( n39193 , n359287 , n359288 );
buf ( n359290 , n39193 );
nand ( n359291 , n39189 , n359290 );
not ( n359292 , n359291 );
not ( n39197 , n359156 );
not ( n359294 , n359194 );
or ( n39199 , n39197 , n359294 );
nand ( n359296 , n39199 , n359203 );
not ( n359297 , n355578 );
or ( n359298 , n359296 , n359297 );
not ( n39203 , n355578 );
nand ( n39204 , n359296 , n39203 );
nand ( n39205 , n359298 , n39204 );
nand ( n359302 , n359292 , n39205 );
buf ( n39207 , n359302 );
not ( n39208 , n39207 );
buf ( n359305 , n39208 );
buf ( n359306 , n359305 );
buf ( n359307 , n359306 );
buf ( n359308 , n359307 );
not ( n359309 , n359308 );
buf ( n359310 , n359309 );
buf ( n359311 , n359310 );
buf ( n359312 , n359291 );
buf ( n39217 , n359312 );
not ( n39218 , n39217 );
buf ( n359315 , n39218 );
nand ( n359316 , n359311 , n359315 );
buf ( n359317 , n359316 );
buf ( n359318 , n359317 );
and ( n359319 , n359149 , n359318 );
buf ( n359320 , n359319 );
buf ( n359321 , n359320 );
not ( n359322 , n32847 );
nand ( n39227 , n359322 , n576 );
buf ( n359324 , n353109 );
buf ( n359325 , n576 );
nand ( n359326 , n359324 , n359325 );
buf ( n359327 , n359326 );
or ( n39232 , n39227 , n359327 );
buf ( n359329 , n359327 );
not ( n39234 , n359329 );
buf ( n359331 , n39227 );
not ( n359332 , n359331 );
or ( n39237 , n39234 , n359332 );
buf ( n359334 , n14890 );
not ( n39239 , n359334 );
buf ( n359336 , n15711 );
not ( n359337 , n359336 );
or ( n39242 , n39239 , n359337 );
buf ( n359339 , n576 );
not ( n359340 , n359339 );
buf ( n359341 , n352857 );
not ( n359342 , n359341 );
or ( n359343 , n359340 , n359342 );
buf ( n359344 , n32830 );
buf ( n359345 , n332672 );
nand ( n359346 , n359344 , n359345 );
buf ( n359347 , n359346 );
buf ( n359348 , n359347 );
nand ( n359349 , n359343 , n359348 );
buf ( n359350 , n359349 );
buf ( n359351 , n359350 );
nand ( n39256 , n39242 , n359351 );
buf ( n39257 , n39256 );
buf ( n359354 , n39257 );
nand ( n39259 , n39237 , n359354 );
buf ( n39260 , n39259 );
nand ( n359357 , n39232 , n39260 );
buf ( n359358 , n359357 );
buf ( n359359 , n32830 );
buf ( n359360 , n576 );
nand ( n39265 , n359359 , n359360 );
buf ( n359362 , n39265 );
buf ( n359363 , n359362 );
nor ( n359364 , n359358 , n359363 );
buf ( n359365 , n359364 );
buf ( n359366 , n359365 );
buf ( n359367 , n359357 );
buf ( n359368 , n359362 );
and ( n39273 , n359367 , n359368 );
buf ( n359370 , n39273 );
buf ( n359371 , n359370 );
or ( n39276 , n359366 , n359371 );
buf ( n359373 , n39276 );
not ( n359374 , n359373 );
and ( n39279 , n33331 , n354977 );
xor ( n359376 , n32841 , n353065 );
and ( n359377 , n359376 , n33137 );
and ( n39282 , n32841 , n353065 );
or ( n39283 , n359377 , n39282 );
xor ( n359380 , n352835 , n352843 );
and ( n359381 , n359380 , n352873 );
and ( n39286 , n352835 , n352843 );
or ( n359383 , n359381 , n39286 );
not ( n359384 , n359383 );
nand ( n39289 , n353077 , n576 );
not ( n359386 , n39289 );
not ( n359387 , n353009 );
not ( n359388 , n353140 );
or ( n39293 , n359387 , n359388 );
buf ( n359390 , n578 );
not ( n359391 , n359390 );
buf ( n359392 , n352857 );
not ( n359393 , n359392 );
or ( n359394 , n359391 , n359393 );
buf ( n359395 , n32830 );
buf ( n359396 , n334748 );
nand ( n39301 , n359395 , n359396 );
buf ( n359398 , n39301 );
buf ( n359399 , n359398 );
nand ( n359400 , n359394 , n359399 );
buf ( n359401 , n359400 );
buf ( n359402 , n359401 );
buf ( n359403 , n334850 );
nand ( n359404 , n359402 , n359403 );
buf ( n359405 , n359404 );
nand ( n359406 , n39293 , n359405 );
xor ( n359407 , n359386 , n359406 );
not ( n39312 , n334786 );
not ( n359409 , n353162 );
or ( n359410 , n39312 , n359409 );
and ( n39315 , n353109 , n332672 );
not ( n39316 , n353109 );
and ( n359413 , n39316 , n576 );
or ( n359414 , n39315 , n359413 );
buf ( n359415 , n359414 );
buf ( n359416 , n14891 );
nand ( n359417 , n359415 , n359416 );
buf ( n359418 , n359417 );
nand ( n359419 , n359410 , n359418 );
xnor ( n359420 , n359407 , n359419 );
xor ( n39325 , n359384 , n359420 );
buf ( n359422 , n353164 );
not ( n39327 , n359422 );
buf ( n359424 , n353147 );
nand ( n359425 , n39327 , n359424 );
buf ( n359426 , n359425 );
not ( n39331 , n359426 );
not ( n39332 , n353128 );
or ( n359429 , n39331 , n39332 );
buf ( n359430 , n353147 );
not ( n359431 , n359430 );
buf ( n359432 , n353164 );
nand ( n39337 , n359431 , n359432 );
buf ( n359434 , n39337 );
nand ( n39339 , n359429 , n359434 );
xnor ( n359436 , n39325 , n39339 );
nand ( n359437 , n39283 , n359436 );
buf ( n359438 , n359437 );
buf ( n359439 , n39227 );
not ( n359440 , n359439 );
buf ( n359441 , n39257 );
not ( n39346 , n359441 );
or ( n359443 , n359440 , n39346 );
buf ( n359444 , n39257 );
buf ( n359445 , n39227 );
or ( n39350 , n359444 , n359445 );
nand ( n359447 , n359443 , n39350 );
buf ( n359448 , n359447 );
buf ( n359449 , n359448 );
not ( n359450 , n359449 );
buf ( n359451 , n359327 );
not ( n359452 , n359451 );
and ( n39357 , n359450 , n359452 );
buf ( n359454 , n359448 );
buf ( n359455 , n359327 );
and ( n39360 , n359454 , n359455 );
nor ( n39361 , n39357 , n39360 );
buf ( n359458 , n39361 );
buf ( n359459 , n359458 );
not ( n39364 , n359459 );
buf ( n359461 , n359327 );
buf ( n359462 , n334786 );
not ( n359463 , n359462 );
buf ( n359464 , n576 );
not ( n359465 , n359464 );
buf ( n359466 , n32847 );
not ( n39371 , n359466 );
or ( n359468 , n359465 , n39371 );
buf ( n39373 , n32846 );
buf ( n359470 , n332672 );
nand ( n359471 , n39373 , n359470 );
buf ( n359472 , n359471 );
buf ( n359473 , n359472 );
nand ( n39378 , n359468 , n359473 );
buf ( n359475 , n39378 );
buf ( n359476 , n359475 );
not ( n39381 , n359476 );
or ( n359478 , n359463 , n39381 );
buf ( n359479 , n359350 );
buf ( n359480 , n14891 );
nand ( n359481 , n359479 , n359480 );
buf ( n359482 , n359481 );
buf ( n359483 , n359482 );
nand ( n359484 , n359478 , n359483 );
buf ( n359485 , n359484 );
buf ( n359486 , n359485 );
xor ( n359487 , n359461 , n359486 );
buf ( n359488 , n338094 );
not ( n359489 , n359488 );
buf ( n359490 , n353145 );
not ( n359491 , n359490 );
or ( n359492 , n359489 , n359491 );
buf ( n359493 , n359401 );
nand ( n359494 , n359492 , n359493 );
buf ( n359495 , n359494 );
buf ( n359496 , n359495 );
not ( n359497 , n359496 );
buf ( n359498 , n32951 );
buf ( n359499 , n576 );
nand ( n359500 , n359498 , n359499 );
buf ( n359501 , n359500 );
buf ( n359502 , n359501 );
nand ( n39407 , n359497 , n359502 );
buf ( n359504 , n39407 );
buf ( n359505 , n359504 );
not ( n39410 , n359505 );
buf ( n359507 , n334786 );
not ( n359508 , n359507 );
buf ( n359509 , n359414 );
not ( n39414 , n359509 );
or ( n359511 , n359508 , n39414 );
buf ( n359512 , n359475 );
buf ( n359513 , n14891 );
nand ( n359514 , n359512 , n359513 );
buf ( n359515 , n359514 );
buf ( n359516 , n359515 );
nand ( n359517 , n359511 , n359516 );
buf ( n359518 , n359517 );
buf ( n359519 , n359518 );
not ( n39424 , n359519 );
or ( n39425 , n39410 , n39424 );
buf ( n359522 , n359501 );
not ( n359523 , n359522 );
buf ( n359524 , n359495 );
nand ( n39429 , n359523 , n359524 );
buf ( n359526 , n39429 );
buf ( n359527 , n359526 );
nand ( n39432 , n39425 , n359527 );
buf ( n359529 , n39432 );
buf ( n359530 , n359529 );
and ( n359531 , n359487 , n359530 );
and ( n359532 , n359461 , n359486 );
or ( n39437 , n359531 , n359532 );
buf ( n359534 , n39437 );
buf ( n359535 , n359534 );
nand ( n359536 , n39364 , n359535 );
buf ( n359537 , n359536 );
buf ( n359538 , n359537 );
nand ( n39443 , n359438 , n359538 );
buf ( n359540 , n39443 );
buf ( n359541 , n359540 );
not ( n359542 , n359541 );
buf ( n359543 , n359542 );
nand ( n39448 , n359543 , n353365 );
nor ( n39449 , n39279 , n39448 );
not ( n359546 , n359458 );
nor ( n359547 , n359546 , n359534 );
not ( n39452 , n359547 );
buf ( n359549 , n359386 );
xnor ( n39454 , n359501 , n359495 );
xor ( n39455 , n39454 , n359518 );
buf ( n359552 , n39455 );
xor ( n359553 , n359549 , n359552 );
not ( n39458 , n39289 );
not ( n359555 , n359419 );
or ( n39460 , n39458 , n359555 );
or ( n359557 , n359419 , n39289 );
nand ( n39462 , n359557 , n359406 );
nand ( n359559 , n39460 , n39462 );
buf ( n359560 , n359559 );
xor ( n39465 , n359553 , n359560 );
buf ( n359562 , n39465 );
not ( n39467 , n359420 );
nand ( n359564 , n39467 , n359384 );
not ( n359565 , n359564 );
not ( n359566 , n39339 );
or ( n39471 , n359565 , n359566 );
nand ( n359568 , n359420 , n359383 );
nand ( n39473 , n39471 , n359568 );
nand ( n39474 , n359562 , n39473 );
buf ( n359571 , n39474 );
xor ( n359572 , n359549 , n359552 );
and ( n39477 , n359572 , n359560 );
and ( n359574 , n359549 , n359552 );
or ( n359575 , n39477 , n359574 );
buf ( n359576 , n359575 );
buf ( n359577 , n359576 );
xor ( n359578 , n359461 , n359486 );
xor ( n39483 , n359578 , n359530 );
buf ( n359580 , n39483 );
buf ( n359581 , n359580 );
nor ( n39486 , n359577 , n359581 );
buf ( n359583 , n39486 );
buf ( n359584 , n359583 );
or ( n359585 , n359571 , n359584 );
buf ( n39490 , n359576 );
buf ( n359587 , n359580 );
nand ( n39492 , n39490 , n359587 );
buf ( n39493 , n39492 );
buf ( n359590 , n39493 );
nand ( n39495 , n359585 , n359590 );
buf ( n39496 , n39495 );
nand ( n359593 , n39452 , n39496 );
and ( n39498 , n39449 , n359593 );
not ( n359595 , n359593 );
or ( n359596 , n359562 , n39473 );
not ( n359597 , n359583 );
nand ( n39502 , n359596 , n359597 );
nor ( n359599 , n39502 , n359547 );
not ( n359600 , n359537 );
or ( n39505 , n359599 , n359600 );
or ( n359602 , n39283 , n359436 );
or ( n359603 , n359540 , n359602 );
nand ( n359604 , n39505 , n359603 );
not ( n39509 , n359604 );
or ( n359606 , n359595 , n39509 );
and ( n39511 , n353365 , n35531 );
nand ( n39512 , n359593 , n359543 , n39511 , n355559 );
nand ( n359609 , n359606 , n39512 );
nor ( n359610 , n39498 , n359609 );
not ( n39515 , n359610 );
buf ( n359612 , n359186 );
not ( n39517 , n359612 );
buf ( n359614 , n359163 );
not ( n359615 , n359614 );
or ( n39520 , n39517 , n359615 );
not ( n39521 , n33138 );
nand ( n39522 , n39521 , n353363 );
nand ( n359619 , n35062 , n39522 , n359602 );
not ( n359620 , n359619 );
and ( n39525 , n359620 , n359599 );
buf ( n359622 , n39525 );
nand ( n359623 , n39520 , n359622 );
buf ( n359624 , n359623 );
not ( n359625 , n359177 );
nand ( n359626 , n359625 , n39525 );
nand ( n39531 , n39515 , n359624 , n359626 );
not ( n359628 , n39531 );
or ( n359629 , n359374 , n359628 );
not ( n39534 , n359610 );
not ( n359631 , n359373 );
nand ( n359632 , n39534 , n359631 , n359624 , n359626 );
nand ( n39537 , n359629 , n359632 );
not ( n359634 , n39537 );
nor ( n39539 , n359600 , n359547 );
not ( n359636 , n39539 );
not ( n39541 , n359636 );
buf ( n39542 , n359245 );
buf ( n359639 , n39542 );
buf ( n359640 , n355536 );
not ( n359641 , n359640 );
not ( n39546 , n39502 );
nand ( n39547 , n359620 , n39546 );
buf ( n359644 , n39547 );
nor ( n359645 , n359641 , n359644 );
buf ( n359646 , n359645 );
buf ( n359647 , n359646 );
nand ( n359648 , n359639 , n359647 );
buf ( n359649 , n359648 );
not ( n39554 , n39547 );
not ( n359651 , n359260 );
not ( n359652 , n359256 );
or ( n39557 , n359651 , n359652 );
nand ( n359654 , n39557 , n359275 );
nand ( n359655 , n39554 , n359654 , n355484 );
not ( n39560 , n39546 );
not ( n39561 , n359602 );
not ( n39562 , n355567 );
not ( n359659 , n33331 );
or ( n359660 , n39562 , n359659 );
nand ( n39565 , n359660 , n353365 );
not ( n39566 , n39565 );
or ( n39567 , n39561 , n39566 );
buf ( n359664 , n359437 );
nand ( n359665 , n39567 , n359664 );
not ( n39570 , n359665 );
or ( n39571 , n39560 , n39570 );
not ( n359668 , n39496 );
nand ( n359669 , n39571 , n359668 );
not ( n39574 , n359669 );
nand ( n359671 , n359649 , n359655 , n39574 );
not ( n39576 , n359671 );
or ( n359673 , n39541 , n39576 );
not ( n39578 , n39539 );
nor ( n39579 , n39578 , n359669 );
nand ( n359676 , n39579 , n359649 , n359655 );
nand ( n39581 , n359673 , n359676 );
and ( n39582 , n359634 , n39581 );
not ( n359679 , n359634 );
buf ( n359680 , n39581 );
not ( n39585 , n359680 );
buf ( n359682 , n39585 );
and ( n359683 , n359679 , n359682 );
nor ( n39588 , n39582 , n359683 );
not ( n359685 , n39588 );
buf ( n359686 , n359685 );
buf ( n39591 , n359686 );
buf ( n39592 , n39591 );
buf ( n359689 , n39592 );
not ( n359690 , n359689 );
buf ( n359691 , n359620 );
buf ( n359692 , n359691 );
buf ( n359693 , n359692 );
buf ( n359694 , n359365 );
not ( n359695 , n359694 );
buf ( n359696 , n359695 );
and ( n39601 , n359599 , n359696 );
and ( n359698 , n359693 , n39601 );
not ( n39603 , n359698 );
not ( n359700 , n359278 );
or ( n39605 , n39603 , n359700 );
not ( n39606 , n359665 );
not ( n359703 , n39606 );
and ( n359704 , n359703 , n39601 );
not ( n39609 , n359600 );
nand ( n359706 , n39609 , n359593 );
buf ( n359707 , n359706 );
buf ( n359708 , n359696 );
and ( n359709 , n359707 , n359708 );
buf ( n359710 , n359370 );
nor ( n359711 , n359709 , n359710 );
buf ( n359712 , n359711 );
not ( n359713 , n359712 );
nor ( n39618 , n359704 , n359713 );
nand ( n359715 , n39605 , n39618 );
buf ( n39620 , n359715 );
not ( n39621 , n39620 );
buf ( n39622 , n39621 );
buf ( n359719 , n39622 );
buf ( n359720 , n359719 );
buf ( n359721 , n36285 );
not ( n359722 , n359721 );
buf ( n359723 , n359102 );
nand ( n359724 , n359722 , n359723 );
buf ( n359725 , n359724 );
not ( n39630 , n359725 );
not ( n359727 , n39630 );
buf ( n359728 , n356299 );
not ( n359729 , n359728 );
and ( n359730 , n356817 , n356856 );
buf ( n359731 , n359730 );
not ( n359732 , n359731 );
buf ( n359733 , n359075 );
not ( n39638 , n359733 );
or ( n359735 , n359732 , n39638 );
buf ( n39640 , n359092 );
not ( n39641 , n39640 );
buf ( n39642 , n39641 );
buf ( n359739 , n39642 );
nand ( n39644 , n359735 , n359739 );
buf ( n359741 , n39644 );
buf ( n359742 , n359741 );
not ( n359743 , n359742 );
or ( n39648 , n359729 , n359743 );
buf ( n359745 , n359098 );
nand ( n359746 , n39648 , n359745 );
buf ( n359747 , n359746 );
not ( n359748 , n359747 );
not ( n359749 , n359748 );
or ( n359750 , n359727 , n359749 );
buf ( n359751 , n359747 );
buf ( n359752 , n359725 );
nand ( n359753 , n359751 , n359752 );
buf ( n359754 , n359753 );
nand ( n359755 , n359750 , n359754 );
buf ( n359756 , n359755 );
not ( n39655 , n359756 );
and ( n359758 , n359720 , n39655 );
not ( n359759 , n359720 );
not ( n39658 , n39655 );
and ( n39659 , n359759 , n39658 );
or ( n359762 , n359758 , n39659 );
buf ( n359763 , n359762 );
not ( n39662 , n359763 );
or ( n39663 , n359690 , n39662 );
buf ( n359766 , n359741 );
buf ( n359767 , n359766 );
buf ( n359768 , n359767 );
buf ( n359769 , n359098 );
buf ( n359770 , n356299 );
nand ( n39666 , n359769 , n359770 );
buf ( n39667 , n39666 );
not ( n359773 , n39667 );
and ( n359774 , n359768 , n359773 );
not ( n39670 , n359768 );
and ( n39671 , n39670 , n39667 );
nor ( n39672 , n359774 , n39671 );
buf ( n359778 , n39672 );
buf ( n359779 , n359778 );
buf ( n39675 , n359779 );
buf ( n359781 , n39675 );
buf ( n359782 , n359781 );
not ( n359783 , n359782 );
buf ( n359784 , n359783 );
and ( n359785 , n359784 , n359720 );
not ( n39681 , n359784 );
buf ( n359787 , n359720 );
not ( n359788 , n359787 );
buf ( n359789 , n359788 );
and ( n359790 , n39681 , n359789 );
or ( n359791 , n359785 , n359790 );
buf ( n359792 , n359791 );
not ( n359793 , n359715 );
buf ( n359794 , n359793 );
not ( n39690 , n359794 );
buf ( n359796 , n359634 );
not ( n359797 , n359796 );
or ( n359798 , n39690 , n359797 );
not ( n39694 , n359634 );
not ( n359800 , n359793 );
nand ( n359801 , n39694 , n359800 );
buf ( n359802 , n359801 );
nand ( n359803 , n359798 , n359802 );
buf ( n359804 , n359803 );
nand ( n39700 , n359804 , n39588 );
not ( n39701 , n39700 );
buf ( n359807 , n39701 );
buf ( n39703 , n359807 );
buf ( n359809 , n39703 );
buf ( n359810 , n359809 );
not ( n39706 , n359810 );
buf ( n39707 , n39706 );
buf ( n359813 , n39707 );
not ( n39709 , n359813 );
buf ( n359815 , n39709 );
buf ( n359816 , n359815 );
nand ( n359817 , n359792 , n359816 );
buf ( n359818 , n359817 );
buf ( n359819 , n359818 );
nand ( n359820 , n39663 , n359819 );
buf ( n359821 , n359820 );
buf ( n359822 , n359821 );
xor ( n359823 , n359321 , n359822 );
and ( n359824 , n39493 , n359597 );
buf ( n359825 , n359596 );
buf ( n359826 , n359825 );
buf ( n359827 , n359826 );
not ( n359828 , n359827 );
nand ( n39724 , n35062 , n39522 );
not ( n359830 , n39724 );
and ( n39726 , n359830 , n355536 , n359602 );
not ( n359832 , n39726 );
not ( n39728 , n39542 );
or ( n359834 , n359832 , n39728 );
nand ( n359835 , n359834 , n39606 );
not ( n359836 , n359835 );
or ( n39732 , n359828 , n359836 );
buf ( n359838 , n359693 );
buf ( n359839 , n359827 );
and ( n39735 , n359838 , n359839 );
buf ( n359841 , n39735 );
not ( n359842 , n39181 );
and ( n359843 , n359841 , n359842 );
buf ( n359844 , n39474 );
not ( n359845 , n359844 );
buf ( n359846 , n359845 );
nor ( n359847 , n359843 , n359846 );
nand ( n359848 , n39732 , n359847 );
xor ( n359849 , n359824 , n359848 );
not ( n39745 , n359620 );
not ( n359851 , n39064 );
or ( n359852 , n39745 , n359851 );
not ( n39748 , n359665 );
nand ( n39749 , n359852 , n39748 );
not ( n359855 , n39749 );
not ( n359856 , n359855 );
buf ( n359857 , n359177 );
not ( n39753 , n359857 );
not ( n39754 , n39085 );
nand ( n359860 , n355484 , n39754 );
buf ( n359861 , n359860 );
not ( n39757 , n359861 );
or ( n39758 , n39753 , n39757 );
buf ( n359864 , n359693 );
nand ( n359865 , n39758 , n359864 );
buf ( n359866 , n359865 );
not ( n39762 , n359866 );
or ( n359868 , n359856 , n39762 );
buf ( n359869 , n359827 );
buf ( n359870 , n39474 );
nand ( n359871 , n359869 , n359870 );
buf ( n359872 , n359871 );
nand ( n39768 , n359868 , n359872 );
nor ( n359874 , n39749 , n359872 );
nand ( n359875 , n359874 , n359866 );
nand ( n39771 , n39768 , n359875 );
buf ( n359877 , n39771 );
buf ( n359878 , n359877 );
buf ( n359879 , n359878 );
xnor ( n39775 , n359849 , n359879 );
buf ( n359881 , n39775 );
not ( n359882 , n359827 );
not ( n359883 , n359835 );
or ( n39779 , n359882 , n359883 );
nand ( n359885 , n39779 , n359847 );
not ( n359886 , n359824 );
and ( n39782 , n359885 , n359886 );
not ( n39783 , n359885 );
and ( n39784 , n39783 , n359824 );
nor ( n359890 , n39782 , n39784 );
buf ( n359891 , n359890 );
not ( n359892 , n359891 );
not ( n359893 , n359636 );
not ( n359894 , n359671 );
or ( n359895 , n359893 , n359894 );
nand ( n359896 , n359895 , n359676 );
buf ( n359897 , n359896 );
not ( n39790 , n359897 );
or ( n359899 , n359892 , n39790 );
buf ( n39792 , n359890 );
not ( n359901 , n39792 );
buf ( n359902 , n359901 );
buf ( n359903 , n359902 );
not ( n359904 , n359896 );
buf ( n359905 , n359904 );
nand ( n359906 , n359903 , n359905 );
buf ( n359907 , n359906 );
buf ( n359908 , n359907 );
nand ( n359909 , n359899 , n359908 );
buf ( n359910 , n359909 );
buf ( n359911 , n359910 );
nand ( n359912 , n359881 , n359911 );
buf ( n359913 , n359912 );
buf ( n359914 , n359913 );
not ( n359915 , n359914 );
buf ( n359916 , n359915 );
buf ( n359917 , n359916 );
buf ( n359918 , n359917 );
buf ( n359919 , n359918 );
buf ( n359920 , n359919 );
not ( n359921 , n359920 );
buf ( n39814 , n359105 );
buf ( n39815 , n39814 );
buf ( n39816 , n39815 );
not ( n359925 , n35893 );
buf ( n359926 , n359925 );
buf ( n359927 , n359111 );
buf ( n359928 , n359927 );
nand ( n39821 , n359926 , n359928 );
buf ( n39822 , n39821 );
buf ( n359931 , n39822 );
not ( n39824 , n359931 );
buf ( n359933 , n39824 );
and ( n39826 , n39816 , n359933 );
not ( n359935 , n39816 );
and ( n359936 , n359935 , n39822 );
nor ( n359937 , n39826 , n359936 );
buf ( n39830 , n359937 );
not ( n359939 , n39830 );
not ( n39832 , n359939 );
not ( n39833 , n39832 );
buf ( n39834 , n359896 );
buf ( n359943 , n39834 );
buf ( n359944 , n359943 );
buf ( n359945 , n359944 );
not ( n359946 , n359945 );
buf ( n359947 , n359946 );
buf ( n359948 , n359947 );
not ( n359949 , n359948 );
buf ( n359950 , n359949 );
and ( n39843 , n39833 , n359950 );
not ( n39844 , n39833 );
buf ( n359953 , n359950 );
not ( n359954 , n359953 );
buf ( n359955 , n359954 );
and ( n39848 , n39844 , n359955 );
or ( n39849 , n39843 , n39848 );
buf ( n359958 , n39849 );
not ( n359959 , n359958 );
or ( n39852 , n359921 , n359959 );
buf ( n39853 , n359950 );
not ( n39854 , n39853 );
not ( n359963 , n359925 );
not ( n39856 , n359105 );
or ( n39857 , n359963 , n39856 );
nand ( n359966 , n39857 , n359927 );
not ( n39859 , n355962 );
and ( n39860 , n39859 , n39021 );
and ( n39861 , n359966 , n39860 );
not ( n359970 , n359966 );
not ( n39863 , n39860 );
and ( n39864 , n359970 , n39863 );
nor ( n359973 , n39861 , n39864 );
buf ( n359974 , n359973 );
buf ( n39867 , n359974 );
not ( n359976 , n39867 );
not ( n359977 , n359976 );
buf ( n39870 , n359977 );
not ( n359979 , n39870 );
buf ( n359980 , n359979 );
not ( n359981 , n359980 );
or ( n39874 , n39854 , n359981 );
buf ( n359983 , n39870 );
buf ( n359984 , n359955 );
nand ( n39877 , n359983 , n359984 );
buf ( n39878 , n39877 );
buf ( n359987 , n39878 );
nand ( n39880 , n39874 , n359987 );
buf ( n39881 , n39880 );
buf ( n359990 , n39881 );
buf ( n359991 , n39775 );
not ( n359992 , n359991 );
buf ( n359993 , n359992 );
buf ( n359994 , n359993 );
not ( n359995 , n359994 );
buf ( n359996 , n359995 );
buf ( n39889 , n359996 );
not ( n39890 , n39889 );
buf ( n39891 , n39890 );
buf ( n360000 , n39891 );
nand ( n39893 , n359990 , n360000 );
buf ( n360002 , n39893 );
buf ( n360003 , n360002 );
nand ( n39896 , n39852 , n360003 );
buf ( n39897 , n39896 );
buf ( n360006 , n39897 );
xor ( n39899 , n359823 , n360006 );
buf ( n360008 , n39899 );
buf ( n360009 , n360008 );
buf ( n360010 , n355497 );
not ( n360011 , n360010 );
buf ( n360012 , n360011 );
buf ( n360013 , n360012 );
not ( n360014 , n360013 );
buf ( n360015 , n342010 );
not ( n360016 , n360015 );
or ( n39909 , n360014 , n360016 );
buf ( n360018 , n35478 );
not ( n360019 , n360018 );
buf ( n360020 , n360019 );
buf ( n360021 , n360020 );
nand ( n360022 , n39909 , n360021 );
buf ( n360023 , n360022 );
buf ( n360024 , n355514 );
not ( n360025 , n360024 );
buf ( n360026 , n360025 );
and ( n360027 , n360026 , n39522 , n354977 , n355093 );
and ( n39920 , n355480 , n35449 , n360027 );
nand ( n39921 , n360023 , n39920 );
nor ( n360030 , n35397 , n39724 );
nand ( n39923 , n360030 , n354740 );
nand ( n360032 , n359830 , n35515 );
and ( n360033 , n355474 , n359830 );
buf ( n39926 , n39565 );
nor ( n360035 , n360033 , n39926 );
nand ( n360036 , n39921 , n39923 , n360032 , n360035 );
nand ( n39929 , n359602 , n359437 );
xor ( n360038 , n360036 , n39929 );
not ( n360039 , n35544 );
or ( n39932 , n360038 , n360039 );
not ( n360041 , n39929 );
and ( n39934 , n360036 , n360041 );
not ( n360043 , n360036 );
and ( n360044 , n360043 , n39929 );
nor ( n39937 , n39934 , n360044 );
not ( n360046 , n39937 );
nand ( n360047 , n360039 , n360046 );
nand ( n360048 , n39932 , n360047 );
buf ( n360049 , n360048 );
buf ( n360050 , n360049 );
buf ( n360051 , n360050 );
buf ( n360052 , n360051 );
not ( n39945 , n360052 );
buf ( n39946 , n39945 );
buf ( n360055 , n39946 );
buf ( n39948 , n360055 );
buf ( n39949 , n39948 );
buf ( n39950 , n39949 );
buf ( n39951 , n39950 );
buf ( n39952 , n39951 );
buf ( n360061 , n39952 );
not ( n39954 , n360061 );
buf ( n360063 , n359879 );
buf ( n360064 , n360063 );
buf ( n360065 , n360064 );
buf ( n360066 , n360065 );
not ( n360067 , n360066 );
buf ( n360068 , n360067 );
buf ( n360069 , n360068 );
buf ( n39962 , n360069 );
buf ( n39963 , n39962 );
buf ( n360072 , n39963 );
not ( n39965 , n360072 );
buf ( n39966 , n39965 );
buf ( n360075 , n39966 );
not ( n39968 , n360075 );
not ( n360077 , n355965 );
and ( n360078 , n359075 , n36792 );
not ( n39971 , n360078 );
or ( n39972 , n360077 , n39971 );
buf ( n360081 , n356320 );
not ( n39974 , n360081 );
buf ( n360083 , n359099 );
not ( n39976 , n360083 );
or ( n39977 , n39974 , n39976 );
buf ( n360086 , n359102 );
nand ( n39979 , n39977 , n360086 );
buf ( n39980 , n39979 );
buf ( n39981 , n39980 );
buf ( n360090 , n355965 );
and ( n360091 , n39981 , n360090 );
buf ( n360092 , n360091 );
buf ( n360093 , n360092 );
buf ( n360094 , n359120 );
nor ( n360095 , n360093 , n360094 );
buf ( n360096 , n360095 );
nand ( n360097 , n39972 , n360096 );
buf ( n360098 , n355986 );
not ( n39991 , n360098 );
buf ( n360100 , n359128 );
nand ( n39993 , n39991 , n360100 );
buf ( n360102 , n39993 );
buf ( n360103 , n360102 );
not ( n39996 , n360103 );
buf ( n360105 , n39996 );
and ( n39998 , n360097 , n360105 );
not ( n39999 , n360097 );
buf ( n360108 , n360102 );
and ( n40001 , n39999 , n360108 );
nor ( n360110 , n39998 , n40001 );
buf ( n40003 , n360110 );
buf ( n40004 , n40003 );
buf ( n40005 , n40004 );
buf ( n360114 , n40005 );
not ( n40007 , n360114 );
buf ( n360116 , n40007 );
buf ( n360117 , n360116 );
not ( n40010 , n360117 );
or ( n360119 , n39968 , n40010 );
buf ( n360120 , n360116 );
not ( n360121 , n360120 );
buf ( n360122 , n360121 );
buf ( n360123 , n360122 );
buf ( n40016 , n39966 );
not ( n360125 , n40016 );
buf ( n360126 , n360125 );
buf ( n360127 , n360126 );
nand ( n360128 , n360123 , n360127 );
buf ( n360129 , n360128 );
buf ( n360130 , n360129 );
nand ( n360131 , n360119 , n360130 );
buf ( n360132 , n360131 );
buf ( n360133 , n360132 );
not ( n360134 , n360133 );
or ( n40027 , n39954 , n360134 );
buf ( n360136 , n39966 );
not ( n360137 , n360136 );
not ( n360138 , n39870 );
buf ( n360139 , n360138 );
not ( n360140 , n360139 );
or ( n40033 , n360137 , n360140 );
buf ( n360142 , n39870 );
buf ( n360143 , n360126 );
nand ( n40036 , n360142 , n360143 );
buf ( n360145 , n40036 );
buf ( n360146 , n360145 );
nand ( n40039 , n40033 , n360146 );
buf ( n360148 , n40039 );
buf ( n40041 , n360148 );
buf ( n360150 , n39937 );
not ( n40043 , n360150 );
buf ( n360152 , n359879 );
not ( n360153 , n360152 );
buf ( n360154 , n360153 );
buf ( n360155 , n360154 );
not ( n360156 , n360155 );
or ( n360157 , n40043 , n360156 );
buf ( n360158 , n359879 );
buf ( n360159 , n360046 );
nand ( n360160 , n360158 , n360159 );
buf ( n360161 , n360160 );
buf ( n360162 , n360161 );
nand ( n40055 , n360157 , n360162 );
buf ( n360164 , n40055 );
nand ( n360165 , n360164 , n360048 );
not ( n40058 , n360165 );
buf ( n40059 , n40058 );
buf ( n360168 , n40059 );
buf ( n40061 , n360168 );
nand ( n40062 , n40041 , n40061 );
buf ( n360171 , n40062 );
buf ( n360172 , n360171 );
nand ( n360173 , n40027 , n360172 );
buf ( n360174 , n360173 );
buf ( n360175 , n360174 );
not ( n40068 , n360175 );
buf ( n360177 , n359307 );
not ( n40070 , n360177 );
not ( n40071 , n355989 );
not ( n360180 , n360078 );
or ( n40073 , n40071 , n360180 );
buf ( n360182 , n360092 );
buf ( n360183 , n355983 );
and ( n360184 , n360182 , n360183 );
buf ( n360185 , n359131 );
nor ( n360186 , n360184 , n360185 );
buf ( n360187 , n360186 );
nand ( n40080 , n40073 , n360187 );
not ( n360189 , n359141 );
not ( n360190 , n355652 );
nand ( n40083 , n360190 , n355589 );
nand ( n360192 , n360189 , n40083 );
not ( n360193 , n360192 );
and ( n40086 , n40080 , n360193 );
not ( n40087 , n40080 );
and ( n40088 , n40087 , n360192 );
nor ( n40089 , n40086 , n40088 );
buf ( n40090 , n40089 );
not ( n40091 , n40090 );
buf ( n40092 , n40091 );
not ( n40093 , n40092 );
xor ( n40094 , n355582 , n40093 );
buf ( n360203 , n40094 );
not ( n40096 , n360203 );
or ( n40097 , n40070 , n40096 );
buf ( n360206 , n359148 );
buf ( n360207 , n39217 );
nand ( n40100 , n360206 , n360207 );
buf ( n360209 , n40100 );
buf ( n360210 , n360209 );
nand ( n40103 , n40097 , n360210 );
buf ( n360212 , n40103 );
buf ( n360213 , n360212 );
not ( n40106 , n360213 );
or ( n360215 , n40068 , n40106 );
buf ( n40108 , n360174 );
not ( n40109 , n40108 );
buf ( n360218 , n40109 );
buf ( n360219 , n360218 );
not ( n40112 , n360219 );
buf ( n360221 , n360212 );
not ( n360222 , n360221 );
buf ( n360223 , n360222 );
buf ( n360224 , n360223 );
not ( n360225 , n360224 );
or ( n40118 , n40112 , n360225 );
buf ( n360227 , n359919 );
not ( n40120 , n360227 );
buf ( n360229 , n359950 );
not ( n360230 , n360229 );
buf ( n360231 , n39655 );
not ( n360232 , n360231 );
or ( n360233 , n360230 , n360232 );
buf ( n360234 , n39658 );
buf ( n360235 , n359955 );
nand ( n360236 , n360234 , n360235 );
buf ( n360237 , n360236 );
buf ( n360238 , n360237 );
nand ( n360239 , n360233 , n360238 );
buf ( n360240 , n360239 );
buf ( n360241 , n360240 );
not ( n360242 , n360241 );
or ( n360243 , n40120 , n360242 );
buf ( n360244 , n39849 );
buf ( n360245 , n39891 );
nand ( n40138 , n360244 , n360245 );
buf ( n360247 , n40138 );
buf ( n360248 , n360247 );
nand ( n360249 , n360243 , n360248 );
buf ( n360250 , n360249 );
buf ( n360251 , n360250 );
nand ( n40144 , n40118 , n360251 );
buf ( n360253 , n40144 );
buf ( n360254 , n360253 );
nand ( n360255 , n360215 , n360254 );
buf ( n360256 , n360255 );
buf ( n360257 , n39952 );
not ( n40150 , n360257 );
buf ( n40151 , n39966 );
buf ( n360260 , n40151 );
not ( n360261 , n360260 );
buf ( n360262 , n40092 );
not ( n360263 , n360262 );
or ( n40156 , n360261 , n360263 );
buf ( n360265 , n40093 );
buf ( n360266 , n360126 );
nand ( n40159 , n360265 , n360266 );
buf ( n360268 , n40159 );
buf ( n360269 , n360268 );
nand ( n40162 , n40156 , n360269 );
buf ( n360271 , n40162 );
buf ( n360272 , n360271 );
not ( n40165 , n360272 );
or ( n360274 , n40150 , n40165 );
buf ( n360275 , n360132 );
buf ( n360276 , n360168 );
nand ( n360277 , n360275 , n360276 );
buf ( n360278 , n360277 );
buf ( n360279 , n360278 );
nand ( n40172 , n360274 , n360279 );
buf ( n360281 , n40172 );
buf ( n360282 , n39592 );
not ( n40175 , n360282 );
buf ( n360284 , n359791 );
not ( n40177 , n360284 );
or ( n40178 , n40175 , n40177 );
not ( n360287 , n356817 );
nand ( n40180 , n38907 , n38929 , n38978 );
not ( n40181 , n40180 );
or ( n40182 , n360287 , n40181 );
nand ( n360291 , n40182 , n359082 );
buf ( n360292 , n360291 );
buf ( n360293 , n359089 );
buf ( n360294 , n356856 );
nand ( n40187 , n360293 , n360294 );
buf ( n360296 , n40187 );
buf ( n360297 , n360296 );
not ( n40190 , n360297 );
buf ( n360299 , n40190 );
buf ( n360300 , n360299 );
and ( n360301 , n360292 , n360300 );
not ( n360302 , n360292 );
buf ( n360303 , n360296 );
and ( n40196 , n360302 , n360303 );
nor ( n360305 , n360301 , n40196 );
buf ( n360306 , n360305 );
buf ( n40199 , n360306 );
not ( n360308 , n40199 );
not ( n40201 , n360308 );
not ( n40202 , n40201 );
and ( n40203 , n40202 , n359720 );
not ( n360312 , n40202 );
and ( n40205 , n360312 , n359789 );
or ( n360314 , n40203 , n40205 );
buf ( n40207 , n360314 );
buf ( n360316 , n359815 );
nand ( n40209 , n40207 , n360316 );
buf ( n360318 , n40209 );
buf ( n360319 , n360318 );
nand ( n360320 , n40178 , n360319 );
buf ( n360321 , n360320 );
buf ( n360322 , n360321 );
not ( n360323 , n360322 );
buf ( n360324 , n360323 );
xor ( n40217 , n360281 , n360324 );
xor ( n360326 , n360256 , n40217 );
buf ( n40219 , n360326 );
xor ( n40220 , n360009 , n40219 );
buf ( n360329 , n360321 );
not ( n360330 , n360329 );
buf ( n360331 , n359815 );
not ( n360332 , n360331 );
buf ( n360333 , n359720 );
not ( n40226 , n360333 );
buf ( n40227 , n358989 );
not ( n40228 , n40227 );
not ( n40229 , n40228 );
not ( n40230 , n359011 );
not ( n40231 , n351407 );
not ( n40232 , n359023 );
or ( n360341 , n40231 , n40232 );
not ( n360342 , n37499 );
nand ( n360343 , n360341 , n360342 );
not ( n360344 , n360343 );
or ( n360345 , n40230 , n360344 );
buf ( n360346 , n38540 );
not ( n360347 , n360346 );
buf ( n360348 , n38556 );
not ( n360349 , n360348 );
or ( n360350 , n360347 , n360349 );
buf ( n360351 , n358652 );
nand ( n360352 , n360350 , n360351 );
buf ( n360353 , n360352 );
nand ( n360354 , n360345 , n360353 );
buf ( n360355 , n360354 );
buf ( n360356 , n360355 );
buf ( n360357 , n360356 );
not ( n40235 , n360357 );
or ( n360359 , n40229 , n40235 );
buf ( n360360 , n359057 );
buf ( n360361 , n38964 );
not ( n40239 , n360361 );
buf ( n360363 , n40239 );
buf ( n360364 , n360363 );
nor ( n40242 , n360360 , n360364 );
buf ( n360366 , n40242 );
nand ( n360367 , n360359 , n360366 );
nand ( n40245 , n359028 , n359070 );
not ( n360369 , n40245 );
and ( n360370 , n360367 , n360369 );
not ( n40248 , n360367 );
and ( n360372 , n40248 , n40245 );
nor ( n360373 , n360370 , n360372 );
buf ( n40251 , n360373 );
not ( n40252 , n40251 );
buf ( n360376 , n40252 );
not ( n360377 , n360376 );
or ( n40255 , n40226 , n360377 );
not ( n360379 , n40252 );
buf ( n360380 , n360379 );
buf ( n360381 , n359789 );
nand ( n360382 , n360380 , n360381 );
buf ( n360383 , n360382 );
buf ( n360384 , n360383 );
nand ( n40262 , n40255 , n360384 );
buf ( n360386 , n40262 );
buf ( n360387 , n360386 );
not ( n360388 , n360387 );
or ( n360389 , n360332 , n360388 );
buf ( n40267 , n40180 );
and ( n40268 , n356817 , n359082 );
and ( n40269 , n40267 , n40268 );
not ( n40270 , n40267 );
not ( n40271 , n40268 );
and ( n360395 , n40270 , n40271 );
nor ( n40273 , n40269 , n360395 );
not ( n360397 , n40273 );
not ( n40275 , n360397 );
buf ( n360399 , n40275 );
not ( n360400 , n360399 );
buf ( n360401 , n360400 );
buf ( n360402 , n360401 );
not ( n360403 , n360402 );
buf ( n360404 , n360403 );
buf ( n360405 , n360404 );
not ( n360406 , n360405 );
buf ( n360407 , n360406 );
and ( n360408 , n360407 , n359720 );
not ( n40286 , n360407 );
and ( n40287 , n40286 , n359789 );
or ( n40288 , n360408 , n40287 );
buf ( n360412 , n40288 );
buf ( n360413 , n39592 );
nand ( n40291 , n360412 , n360413 );
buf ( n360415 , n40291 );
buf ( n360416 , n360415 );
nand ( n360417 , n360389 , n360416 );
buf ( n360418 , n360417 );
buf ( n360419 , n360418 );
buf ( n360420 , n39891 );
not ( n360421 , n360420 );
buf ( n360422 , n360240 );
not ( n360423 , n360422 );
or ( n360424 , n360421 , n360423 );
buf ( n360425 , n359950 );
not ( n360426 , n360425 );
buf ( n40304 , n359784 );
not ( n40305 , n40304 );
or ( n40306 , n360426 , n40305 );
buf ( n360430 , n359781 );
buf ( n360431 , n360430 );
buf ( n360432 , n359955 );
nand ( n360433 , n360431 , n360432 );
buf ( n360434 , n360433 );
buf ( n360435 , n360434 );
nand ( n360436 , n40306 , n360435 );
buf ( n360437 , n360436 );
buf ( n360438 , n360437 );
buf ( n360439 , n359919 );
nand ( n40317 , n360438 , n360439 );
buf ( n360441 , n40317 );
buf ( n360442 , n360441 );
nand ( n360443 , n360424 , n360442 );
buf ( n360444 , n360443 );
buf ( n360445 , n360444 );
xor ( n40323 , n360419 , n360445 );
buf ( n40324 , n360168 );
not ( n40325 , n40324 );
and ( n360449 , n39833 , n39966 );
not ( n40327 , n39833 );
and ( n40328 , n40327 , n360126 );
or ( n360452 , n360449 , n40328 );
buf ( n360453 , n360452 );
not ( n40331 , n360453 );
or ( n360455 , n40325 , n40331 );
buf ( n360456 , n360148 );
buf ( n360457 , n39952 );
nand ( n360458 , n360456 , n360457 );
buf ( n360459 , n360458 );
buf ( n360460 , n360459 );
nand ( n40338 , n360455 , n360460 );
buf ( n40339 , n40338 );
buf ( n360463 , n40339 );
and ( n40341 , n40323 , n360463 );
and ( n360465 , n360419 , n360445 );
or ( n360466 , n40341 , n360465 );
buf ( n360467 , n360466 );
buf ( n360468 , n360467 );
not ( n360469 , n360468 );
buf ( n360470 , n360469 );
buf ( n360471 , n360470 );
not ( n360472 , n360471 );
or ( n40350 , n360330 , n360472 );
or ( n360474 , n355337 , n355313 );
buf ( n40352 , n360474 );
buf ( n360476 , n355340 );
buf ( n40354 , n360476 );
buf ( n40355 , n40354 );
buf ( n360479 , n40355 );
nand ( n40357 , n40352 , n360479 );
buf ( n40358 , n40357 );
buf ( n40359 , n40358 );
not ( n360483 , n40359 );
buf ( n360484 , n360483 );
not ( n360485 , n360484 );
not ( n40363 , n355429 );
nand ( n40364 , n354615 , n355439 );
nand ( n40365 , n354456 , n354643 );
nor ( n40366 , n40364 , n40365 );
not ( n40367 , n40366 );
buf ( n360491 , n355500 );
not ( n360492 , n360491 );
buf ( n360493 , n342007 );
not ( n360494 , n360493 );
or ( n40372 , n360492 , n360494 );
buf ( n360496 , n359272 );
nand ( n360497 , n40372 , n360496 );
buf ( n360498 , n360497 );
not ( n360499 , n360498 );
or ( n360500 , n40367 , n360499 );
and ( n40378 , n34684 , n34586 );
nor ( n360502 , n40378 , n354734 );
nand ( n360503 , n360500 , n360502 );
not ( n40381 , n360503 );
or ( n360505 , n40363 , n40381 );
buf ( n360506 , n355427 );
buf ( n360507 , n360506 );
buf ( n360508 , n360507 );
buf ( n360509 , n360508 );
buf ( n360510 , n35496 );
buf ( n360511 , n360510 );
not ( n360512 , n360511 );
buf ( n360513 , n360512 );
buf ( n360514 , n360513 );
and ( n360515 , n360509 , n360514 );
buf ( n360516 , n35494 );
not ( n360517 , n360516 );
buf ( n360518 , n360517 );
buf ( n360519 , n360518 );
nor ( n360520 , n360515 , n360519 );
buf ( n360521 , n360520 );
nand ( n360522 , n360505 , n360521 );
buf ( n360523 , n360522 );
not ( n360524 , n360523 );
buf ( n360525 , n360524 );
not ( n40403 , n360525 );
or ( n40404 , n360485 , n40403 );
buf ( n40405 , n360522 );
buf ( n360529 , n40358 );
nand ( n40407 , n40405 , n360529 );
buf ( n40408 , n40407 );
nand ( n360532 , n40404 , n40408 );
not ( n360533 , n360532 );
not ( n40411 , n360533 );
buf ( n360535 , n39144 );
buf ( n360536 , n355536 );
nand ( n40414 , n360535 , n360536 );
buf ( n360538 , n40414 );
not ( n40416 , n360538 );
buf ( n360540 , n359654 );
and ( n360541 , n40366 , n355429 , n40355 );
buf ( n360542 , n360541 );
nand ( n360543 , n360540 , n360542 );
buf ( n360544 , n360543 );
buf ( n360545 , n39139 );
buf ( n40423 , n360545 );
buf ( n360547 , n40423 );
buf ( n360548 , n360474 );
not ( n40426 , n360548 );
buf ( n360550 , n359238 );
nor ( n360551 , n40426 , n360550 );
buf ( n360552 , n360551 );
nand ( n40430 , n360544 , n360547 , n360552 );
not ( n360554 , n40430 );
or ( n40432 , n40416 , n360554 );
not ( n360556 , n360552 );
nor ( n40434 , n360556 , n360538 );
nand ( n40435 , n360544 , n40434 , n360547 );
nand ( n360559 , n40432 , n40435 );
not ( n360560 , n360559 );
or ( n40438 , n40411 , n360560 );
not ( n360562 , n360559 );
not ( n360563 , n360484 );
not ( n40441 , n360525 );
or ( n360565 , n360563 , n40441 );
nand ( n360566 , n360565 , n40408 );
nand ( n40444 , n360562 , n360566 );
nand ( n40445 , n40438 , n40444 );
buf ( n40446 , n40445 );
not ( n360570 , n40446 );
buf ( n360571 , n360570 );
buf ( n360572 , n360571 );
not ( n360573 , n360572 );
buf ( n360574 , n360573 );
buf ( n360575 , n360574 );
buf ( n360576 , n360575 );
buf ( n360577 , n360576 );
buf ( n360578 , n360577 );
not ( n40456 , n360578 );
buf ( n360580 , n40456 );
buf ( n360581 , n360580 );
not ( n360582 , n360581 );
not ( n360583 , n40445 );
not ( n40461 , n360562 );
not ( n360585 , n40461 );
xnor ( n40463 , n359278 , n359282 );
buf ( n360587 , n40463 );
not ( n40465 , n360587 );
buf ( n360589 , n40465 );
not ( n40467 , n360589 );
or ( n360591 , n360585 , n40467 );
buf ( n360592 , n40463 );
buf ( n360593 , n360562 );
nand ( n40471 , n360592 , n360593 );
buf ( n360595 , n40471 );
nand ( n40473 , n360591 , n360595 );
nand ( n40474 , n360583 , n40473 );
not ( n40475 , n40474 );
buf ( n360599 , n40475 );
buf ( n360600 , n360599 );
buf ( n360601 , n360600 );
buf ( n360602 , n360601 );
not ( n360603 , n360602 );
buf ( n360604 , n360603 );
buf ( n360605 , n360604 );
not ( n360606 , n360605 );
or ( n40484 , n360582 , n360606 );
buf ( n360608 , n360589 );
not ( n360609 , n360608 );
buf ( n360610 , n360609 );
buf ( n360611 , n360610 );
not ( n40489 , n360611 );
buf ( n360613 , n40489 );
buf ( n360614 , n360613 );
not ( n360615 , n360614 );
buf ( n360616 , n360615 );
buf ( n360617 , n360616 );
not ( n360618 , n360617 );
buf ( n360619 , n359147 );
not ( n40497 , n360619 );
or ( n360621 , n360618 , n40497 );
buf ( n40499 , n359147 );
not ( n360623 , n40499 );
buf ( n360624 , n360623 );
buf ( n360625 , n360624 );
buf ( n360626 , n360613 );
nand ( n360627 , n360625 , n360626 );
buf ( n360628 , n360627 );
buf ( n360629 , n360628 );
nand ( n360630 , n360621 , n360629 );
buf ( n360631 , n360630 );
buf ( n360632 , n360631 );
nand ( n360633 , n40484 , n360632 );
buf ( n360634 , n360633 );
not ( n40512 , n359815 );
not ( n360636 , n40288 );
or ( n360637 , n40512 , n360636 );
nand ( n40515 , n360314 , n39592 );
nand ( n40516 , n360637 , n40515 );
xor ( n360640 , n360634 , n40516 );
buf ( n360641 , n39217 );
not ( n360642 , n360641 );
buf ( n360643 , n40094 );
not ( n40521 , n360643 );
or ( n360645 , n360642 , n40521 );
buf ( n360646 , n355582 );
buf ( n360647 , n360122 );
and ( n360648 , n360646 , n360647 );
not ( n360649 , n360646 );
buf ( n360650 , n360116 );
and ( n360651 , n360649 , n360650 );
nor ( n360652 , n360648 , n360651 );
buf ( n360653 , n360652 );
buf ( n360654 , n360653 );
buf ( n360655 , n359307 );
nand ( n360656 , n360654 , n360655 );
buf ( n360657 , n360656 );
buf ( n360658 , n360657 );
nand ( n360659 , n360645 , n360658 );
buf ( n360660 , n360659 );
and ( n40538 , n360640 , n360660 );
and ( n360662 , n360634 , n40516 );
or ( n40540 , n40538 , n360662 );
buf ( n360664 , n40540 );
nand ( n360665 , n40350 , n360664 );
buf ( n360666 , n360665 );
buf ( n360667 , n360666 );
buf ( n360668 , n360467 );
buf ( n360669 , n360324 );
nand ( n360670 , n360668 , n360669 );
buf ( n360671 , n360670 );
buf ( n360672 , n360671 );
and ( n360673 , n360667 , n360672 );
buf ( n360674 , n360673 );
buf ( n360675 , n360674 );
and ( n360676 , n40220 , n360675 );
and ( n360677 , n360009 , n40219 );
or ( n40555 , n360676 , n360677 );
buf ( n360679 , n40555 );
buf ( n360680 , n360679 );
not ( n40558 , n360680 );
buf ( n360682 , n359320 );
not ( n360683 , n360682 );
buf ( n360684 , n360683 );
buf ( n360685 , n360684 );
not ( n360686 , n360685 );
buf ( n360687 , n39897 );
not ( n360688 , n360687 );
or ( n40566 , n360686 , n360688 );
buf ( n360690 , n359320 );
not ( n360691 , n360690 );
buf ( n360692 , n39897 );
not ( n40570 , n360692 );
buf ( n40571 , n40570 );
buf ( n360695 , n40571 );
not ( n40573 , n360695 );
or ( n360697 , n360691 , n40573 );
buf ( n360698 , n359821 );
nand ( n40576 , n360697 , n360698 );
buf ( n360700 , n40576 );
buf ( n360701 , n360700 );
nand ( n40579 , n40566 , n360701 );
buf ( n360703 , n40579 );
buf ( n360704 , n360703 );
buf ( n360705 , n359950 );
not ( n360706 , n360705 );
buf ( n360707 , n360116 );
not ( n360708 , n360707 );
or ( n360709 , n360706 , n360708 );
buf ( n360710 , n360122 );
buf ( n360711 , n359955 );
nand ( n360712 , n360710 , n360711 );
buf ( n360713 , n360712 );
buf ( n360714 , n360713 );
nand ( n40589 , n360709 , n360714 );
buf ( n360716 , n40589 );
and ( n40591 , n360716 , n39891 );
and ( n360718 , n39881 , n359919 );
nor ( n40593 , n40591 , n360718 );
buf ( n360720 , n40593 );
buf ( n360721 , n360168 );
not ( n360722 , n360721 );
buf ( n360723 , n360271 );
not ( n360724 , n360723 );
or ( n360725 , n360722 , n360724 );
and ( n40600 , n39966 , n359147 );
not ( n360727 , n39966 );
and ( n360728 , n360727 , n360624 );
or ( n40603 , n40600 , n360728 );
buf ( n360730 , n40603 );
buf ( n360731 , n39952 );
nand ( n40606 , n360730 , n360731 );
buf ( n360733 , n40606 );
buf ( n360734 , n360733 );
nand ( n40609 , n360725 , n360734 );
buf ( n360736 , n40609 );
buf ( n40611 , n360736 );
xor ( n40612 , n360720 , n40611 );
buf ( n360739 , n359815 );
not ( n360740 , n360739 );
buf ( n360741 , n359762 );
not ( n360742 , n360741 );
or ( n360743 , n360740 , n360742 );
and ( n360744 , n39833 , n359720 );
not ( n40619 , n39833 );
and ( n360746 , n40619 , n359789 );
or ( n360747 , n360744 , n360746 );
buf ( n360748 , n360747 );
buf ( n360749 , n39592 );
nand ( n360750 , n360748 , n360749 );
buf ( n360751 , n360750 );
buf ( n360752 , n360751 );
nand ( n360753 , n360743 , n360752 );
buf ( n360754 , n360753 );
buf ( n360755 , n360754 );
xor ( n40630 , n40612 , n360755 );
buf ( n360757 , n40630 );
buf ( n360758 , n360757 );
xor ( n360759 , n360704 , n360758 );
buf ( n360760 , n360281 );
not ( n40635 , n360760 );
buf ( n360762 , n360324 );
nand ( n360763 , n40635 , n360762 );
buf ( n360764 , n360763 );
buf ( n360765 , n360764 );
not ( n360766 , n360765 );
buf ( n360767 , n360256 );
not ( n360768 , n360767 );
or ( n360769 , n360766 , n360768 );
buf ( n360770 , n360281 );
buf ( n360771 , n360321 );
nand ( n360772 , n360770 , n360771 );
buf ( n360773 , n360772 );
buf ( n360774 , n360773 );
nand ( n360775 , n360769 , n360774 );
buf ( n360776 , n360775 );
buf ( n360777 , n360776 );
xor ( n360778 , n360759 , n360777 );
buf ( n360779 , n360778 );
buf ( n360780 , n360779 );
nand ( n40653 , n40558 , n360780 );
buf ( n360782 , n40653 );
buf ( n360783 , n360782 );
buf ( n360784 , n360779 );
not ( n360785 , n360784 );
buf ( n360786 , n360679 );
nand ( n360787 , n360785 , n360786 );
buf ( n360788 , n360787 );
buf ( n40658 , n360788 );
nand ( n40659 , n360783 , n40658 );
buf ( n40660 , n40659 );
buf ( n360792 , n40660 );
buf ( n360793 , n40660 );
not ( n360794 , n360793 );
buf ( n360795 , n360794 );
buf ( n360796 , n360795 );
buf ( n360797 , n360418 );
not ( n360798 , n360797 );
buf ( n360799 , n360798 );
buf ( n360800 , n360799 );
buf ( n360801 , n360601 );
not ( n360802 , n360801 );
buf ( n360803 , n360616 );
not ( n360804 , n360803 );
buf ( n360805 , n40092 );
not ( n40675 , n360805 );
or ( n360807 , n360804 , n40675 );
buf ( n40677 , n40093 );
buf ( n40678 , n360613 );
nand ( n40679 , n40677 , n40678 );
buf ( n40680 , n40679 );
buf ( n360812 , n40680 );
nand ( n40682 , n360807 , n360812 );
buf ( n360814 , n40682 );
buf ( n360815 , n360814 );
not ( n40685 , n360815 );
or ( n360817 , n360802 , n40685 );
buf ( n360818 , n360631 );
buf ( n360819 , n360577 );
nand ( n360820 , n360818 , n360819 );
buf ( n360821 , n360820 );
buf ( n360822 , n360821 );
nand ( n40692 , n360817 , n360822 );
buf ( n360824 , n40692 );
buf ( n360825 , n360824 );
xor ( n40695 , n360800 , n360825 );
buf ( n40696 , n39592 );
not ( n40697 , n40696 );
buf ( n360829 , n359720 );
not ( n40699 , n360829 );
buf ( n40700 , n358946 );
not ( n360832 , n40700 );
not ( n360833 , n360354 );
or ( n40703 , n360832 , n360833 );
nand ( n360835 , n40703 , n359048 );
buf ( n360836 , n360363 );
buf ( n360837 , n359054 );
or ( n360838 , n360836 , n360837 );
buf ( n360839 , n360838 );
and ( n40709 , n360835 , n360839 );
not ( n40710 , n360835 );
not ( n360842 , n360839 );
and ( n360843 , n40710 , n360842 );
nor ( n40713 , n40709 , n360843 );
not ( n360845 , n40713 );
buf ( n360846 , n360845 );
not ( n360847 , n360846 );
buf ( n360848 , n360847 );
buf ( n360849 , n360848 );
buf ( n360850 , n360849 );
buf ( n360851 , n360850 );
buf ( n360852 , n360851 );
not ( n360853 , n360852 );
or ( n40723 , n40699 , n360853 );
buf ( n360855 , n360851 );
not ( n40725 , n360855 );
buf ( n360857 , n40725 );
buf ( n360858 , n360857 );
buf ( n360859 , n359789 );
nand ( n360860 , n360858 , n360859 );
buf ( n360861 , n360860 );
buf ( n360862 , n360861 );
nand ( n360863 , n40723 , n360862 );
buf ( n360864 , n360863 );
buf ( n360865 , n360864 );
not ( n360866 , n360865 );
or ( n40736 , n40697 , n360866 );
buf ( n360868 , n359720 );
not ( n40738 , n360868 );
buf ( n40739 , n358943 );
not ( n40740 , n40739 );
not ( n40741 , n360354 );
or ( n40742 , n40740 , n40741 );
buf ( n360874 , n359042 );
buf ( n360875 , n360874 );
buf ( n360876 , n360875 );
buf ( n40746 , n360876 );
nand ( n360878 , n40742 , n40746 );
nand ( n360879 , n359032 , n359037 );
not ( n40749 , n360879 );
and ( n40750 , n360878 , n40749 );
not ( n360882 , n360878 );
and ( n40752 , n360882 , n360879 );
nor ( n40753 , n40750 , n40752 );
buf ( n360885 , n40753 );
not ( n360886 , n360885 );
buf ( n40756 , n360886 );
buf ( n360888 , n40756 );
not ( n360889 , n360888 );
or ( n40759 , n40738 , n360889 );
buf ( n360891 , n360885 );
buf ( n360892 , n360891 );
buf ( n360893 , n360892 );
buf ( n360894 , n360893 );
buf ( n360895 , n359789 );
nand ( n360896 , n360894 , n360895 );
buf ( n360897 , n360896 );
buf ( n360898 , n360897 );
nand ( n360899 , n40759 , n360898 );
buf ( n360900 , n360899 );
buf ( n360901 , n360900 );
buf ( n360902 , n359815 );
nand ( n360903 , n360901 , n360902 );
buf ( n360904 , n360903 );
buf ( n360905 , n360904 );
nand ( n360906 , n40736 , n360905 );
buf ( n360907 , n360906 );
buf ( n360908 , n360907 );
buf ( n360909 , n39592 );
not ( n360910 , n360909 );
buf ( n360911 , n360386 );
not ( n360912 , n360911 );
or ( n360913 , n360910 , n360912 );
buf ( n360914 , n360864 );
buf ( n360915 , n359815 );
nand ( n40782 , n360914 , n360915 );
buf ( n360917 , n40782 );
buf ( n360918 , n360917 );
nand ( n40785 , n360913 , n360918 );
buf ( n360920 , n40785 );
buf ( n360921 , n360920 );
xor ( n40788 , n360908 , n360921 );
buf ( n360923 , n39891 );
not ( n360924 , n360923 );
buf ( n360925 , n359950 );
not ( n360926 , n360925 );
buf ( n360927 , n40202 );
not ( n40794 , n360927 );
or ( n40795 , n360926 , n40794 );
buf ( n360930 , n40199 );
not ( n40797 , n360930 );
not ( n40798 , n40797 );
buf ( n360933 , n40798 );
buf ( n360934 , n359955 );
nand ( n40801 , n360933 , n360934 );
buf ( n360936 , n40801 );
buf ( n360937 , n360936 );
nand ( n360938 , n40795 , n360937 );
buf ( n360939 , n360938 );
buf ( n360940 , n360939 );
not ( n40807 , n360940 );
or ( n40808 , n360924 , n40807 );
buf ( n360943 , n359950 );
not ( n40810 , n360943 );
buf ( n360945 , n360407 );
not ( n360946 , n360945 );
or ( n360947 , n40810 , n360946 );
buf ( n360948 , n360404 );
buf ( n360949 , n359955 );
nand ( n360950 , n360948 , n360949 );
buf ( n360951 , n360950 );
buf ( n360952 , n360951 );
nand ( n360953 , n360947 , n360952 );
buf ( n360954 , n360953 );
buf ( n360955 , n360954 );
buf ( n360956 , n359919 );
nand ( n40823 , n360955 , n360956 );
buf ( n360958 , n40823 );
buf ( n360959 , n360958 );
nand ( n360960 , n40808 , n360959 );
buf ( n360961 , n360960 );
buf ( n360962 , n360961 );
and ( n40829 , n40788 , n360962 );
and ( n40830 , n360908 , n360921 );
or ( n40831 , n40829 , n40830 );
buf ( n360966 , n40831 );
buf ( n360967 , n360966 );
xor ( n40834 , n40695 , n360967 );
buf ( n360969 , n40834 );
buf ( n360970 , n360969 );
buf ( n360971 , n360907 );
not ( n40838 , n360971 );
buf ( n360973 , n40838 );
buf ( n360974 , n360973 );
buf ( n40841 , n355412 );
not ( n360976 , n40841 );
not ( n360977 , n360503 );
or ( n40844 , n360976 , n360977 );
nand ( n360979 , n40844 , n360510 );
nand ( n40846 , n360508 , n35494 );
not ( n40847 , n40846 );
and ( n40848 , n360979 , n40847 );
not ( n40849 , n360979 );
and ( n40850 , n40849 , n40846 );
nor ( n360985 , n40848 , n40850 );
not ( n40852 , n360985 );
nand ( n360987 , n360532 , n40852 );
not ( n40854 , n360987 );
not ( n360989 , n360566 );
buf ( n40856 , n360985 );
nand ( n40857 , n360989 , n40856 );
not ( n360992 , n40857 );
or ( n360993 , n40854 , n360992 );
nand ( n40860 , n40841 , n360510 );
not ( n360995 , n40860 );
not ( n360996 , n360995 );
not ( n40863 , n40366 );
not ( n360998 , n360498 );
or ( n360999 , n40863 , n360998 );
nand ( n40866 , n360999 , n360502 );
not ( n40867 , n40866 );
not ( n361002 , n40867 );
or ( n40869 , n360996 , n361002 );
nand ( n361004 , n360503 , n40860 );
nand ( n40871 , n40869 , n361004 );
not ( n361006 , n40871 );
not ( n361007 , n360985 );
or ( n40874 , n361006 , n361007 );
not ( n361009 , n40871 );
nand ( n40876 , n361009 , n40852 );
nand ( n361011 , n40874 , n40876 );
nand ( n40878 , n360993 , n361011 );
not ( n361013 , n40878 );
buf ( n361014 , n361013 );
not ( n40881 , n361014 );
buf ( n361016 , n40881 );
buf ( n361017 , n361016 );
not ( n40884 , n361017 );
buf ( n361019 , n40884 );
buf ( n40886 , n361019 );
buf ( n361021 , n40886 );
buf ( n361022 , n361021 );
buf ( n361023 , n361022 );
not ( n361024 , n361023 );
buf ( n40891 , n360989 );
buf ( n361026 , n40891 );
not ( n40893 , n361026 );
buf ( n361028 , n40893 );
not ( n40895 , n361028 );
buf ( n361030 , n40092 );
not ( n40897 , n361030 );
or ( n361032 , n40895 , n40897 );
buf ( n40899 , n40090 );
buf ( n361034 , n40899 );
buf ( n361035 , n361026 );
nand ( n361036 , n361034 , n361035 );
buf ( n361037 , n361036 );
buf ( n361038 , n361037 );
nand ( n361039 , n361032 , n361038 );
buf ( n361040 , n361039 );
buf ( n361041 , n361040 );
not ( n361042 , n361041 );
or ( n40909 , n361024 , n361042 );
buf ( n361044 , n40893 );
not ( n40911 , n361044 );
buf ( n361046 , n359147 );
not ( n361047 , n361046 );
or ( n40914 , n40911 , n361047 );
buf ( n361049 , n360624 );
buf ( n361050 , n361026 );
nand ( n361051 , n361049 , n361050 );
buf ( n361052 , n361051 );
buf ( n361053 , n361052 );
nand ( n40920 , n40914 , n361053 );
buf ( n40921 , n40920 );
buf ( n361056 , n40921 );
not ( n40923 , n361011 );
buf ( n361058 , n40923 );
buf ( n40925 , n361058 );
buf ( n361060 , n40925 );
buf ( n361061 , n361060 );
nand ( n40928 , n361056 , n361061 );
buf ( n361063 , n40928 );
buf ( n361064 , n361063 );
nand ( n361065 , n40909 , n361064 );
buf ( n361066 , n361065 );
buf ( n361067 , n361066 );
xor ( n40934 , n360974 , n361067 );
buf ( n361069 , n39217 );
not ( n361070 , n361069 );
buf ( n361071 , n355582 );
not ( n40938 , n361071 );
not ( n361073 , n39830 );
buf ( n361074 , n361073 );
not ( n361075 , n361074 );
or ( n361076 , n40938 , n361075 );
buf ( n40943 , n39830 );
buf ( n361078 , n40943 );
not ( n40945 , n355582 );
buf ( n361080 , n40945 );
nand ( n361081 , n361078 , n361080 );
buf ( n361082 , n361081 );
buf ( n361083 , n361082 );
nand ( n40950 , n361076 , n361083 );
buf ( n40951 , n40950 );
buf ( n361086 , n40951 );
not ( n40953 , n361086 );
or ( n361088 , n361070 , n40953 );
buf ( n361089 , n355582 );
not ( n361090 , n361089 );
buf ( n361091 , n39655 );
not ( n40958 , n361091 );
or ( n361093 , n361090 , n40958 );
buf ( n361094 , n359756 );
buf ( n361095 , n40945 );
nand ( n361096 , n361094 , n361095 );
buf ( n361097 , n361096 );
buf ( n361098 , n361097 );
nand ( n361099 , n361093 , n361098 );
buf ( n361100 , n361099 );
buf ( n361101 , n361100 );
buf ( n361102 , n359307 );
nand ( n361103 , n361101 , n361102 );
buf ( n361104 , n361103 );
buf ( n361105 , n361104 );
nand ( n361106 , n361088 , n361105 );
buf ( n361107 , n361106 );
buf ( n361108 , n361107 );
and ( n361109 , n40934 , n361108 );
and ( n40976 , n360974 , n361067 );
or ( n40977 , n361109 , n40976 );
buf ( n361112 , n40977 );
buf ( n361113 , n361112 );
buf ( n361114 , n361060 );
not ( n361115 , n361114 );
buf ( n361116 , n361115 );
buf ( n361117 , n361116 );
not ( n361118 , n361117 );
buf ( n361119 , n361022 );
not ( n361120 , n361119 );
buf ( n361121 , n361120 );
buf ( n361122 , n361121 );
not ( n40989 , n361122 );
or ( n40990 , n361118 , n40989 );
buf ( n361125 , n40921 );
nand ( n40992 , n40990 , n361125 );
buf ( n361127 , n40992 );
buf ( n361128 , n361127 );
buf ( n361129 , n39952 );
not ( n361130 , n361129 );
buf ( n361131 , n39966 );
not ( n361132 , n361131 );
not ( n40999 , n359756 );
buf ( n361134 , n40999 );
not ( n41001 , n361134 );
or ( n41002 , n361132 , n41001 );
buf ( n361137 , n39658 );
buf ( n361138 , n360126 );
nand ( n41005 , n361137 , n361138 );
buf ( n361140 , n41005 );
buf ( n361141 , n361140 );
nand ( n41008 , n41002 , n361141 );
buf ( n361143 , n41008 );
buf ( n361144 , n361143 );
not ( n41011 , n361144 );
or ( n41012 , n361130 , n41011 );
buf ( n361147 , n39966 );
not ( n41014 , n361147 );
buf ( n361149 , n359784 );
not ( n41016 , n361149 );
or ( n361151 , n41014 , n41016 );
buf ( n361152 , n359781 );
buf ( n361153 , n360126 );
nand ( n361154 , n361152 , n361153 );
buf ( n361155 , n361154 );
buf ( n361156 , n361155 );
nand ( n361157 , n361151 , n361156 );
buf ( n361158 , n361157 );
buf ( n361159 , n361158 );
buf ( n361160 , n360168 );
nand ( n361161 , n361159 , n361160 );
buf ( n361162 , n361161 );
buf ( n361163 , n361162 );
nand ( n361164 , n41012 , n361163 );
buf ( n361165 , n361164 );
buf ( n361166 , n361165 );
xor ( n41033 , n361128 , n361166 );
buf ( n361168 , n359307 );
not ( n361169 , n361168 );
buf ( n361170 , n40951 );
not ( n41037 , n361170 );
or ( n41038 , n361169 , n41037 );
buf ( n361173 , n355582 );
not ( n361174 , n361173 );
buf ( n361175 , n360138 );
not ( n361176 , n361175 );
or ( n41043 , n361174 , n361176 );
buf ( n361178 , n39870 );
buf ( n361179 , n40945 );
nand ( n361180 , n361178 , n361179 );
buf ( n361181 , n361180 );
buf ( n361182 , n361181 );
nand ( n41049 , n41043 , n361182 );
buf ( n361184 , n41049 );
buf ( n361185 , n361184 );
buf ( n361186 , n39217 );
nand ( n361187 , n361185 , n361186 );
buf ( n361188 , n361187 );
buf ( n361189 , n361188 );
nand ( n361190 , n41038 , n361189 );
buf ( n361191 , n361190 );
buf ( n361192 , n361191 );
xor ( n41059 , n41033 , n361192 );
buf ( n361194 , n41059 );
buf ( n361195 , n361194 );
xor ( n41062 , n361113 , n361195 );
buf ( n361197 , n360577 );
not ( n41064 , n361197 );
buf ( n361199 , n360814 );
not ( n361200 , n361199 );
or ( n41067 , n41064 , n361200 );
buf ( n361202 , n360601 );
buf ( n361203 , n360616 );
not ( n361204 , n361203 );
buf ( n361205 , n360116 );
not ( n361206 , n361205 );
or ( n41073 , n361204 , n361206 );
buf ( n361208 , n360122 );
buf ( n361209 , n360613 );
nand ( n361210 , n361208 , n361209 );
buf ( n361211 , n361210 );
buf ( n41078 , n361211 );
nand ( n41079 , n41073 , n41078 );
buf ( n41080 , n41079 );
buf ( n361215 , n41080 );
nand ( n41082 , n361202 , n361215 );
buf ( n41083 , n41082 );
buf ( n361218 , n41083 );
nand ( n41085 , n41067 , n361218 );
buf ( n361220 , n41085 );
buf ( n361221 , n361220 );
xor ( n361222 , n360908 , n360921 );
xor ( n41089 , n361222 , n360962 );
buf ( n361224 , n41089 );
buf ( n361225 , n361224 );
xor ( n41092 , n361221 , n361225 );
buf ( n361227 , n359919 );
not ( n361228 , n361227 );
buf ( n361229 , n359950 );
not ( n361230 , n361229 );
buf ( n361231 , n40252 );
not ( n361232 , n361231 );
or ( n41099 , n361230 , n361232 );
buf ( n361234 , n360379 );
buf ( n361235 , n359955 );
nand ( n361236 , n361234 , n361235 );
buf ( n361237 , n361236 );
buf ( n361238 , n361237 );
nand ( n361239 , n41099 , n361238 );
buf ( n361240 , n361239 );
buf ( n361241 , n361240 );
not ( n41108 , n361241 );
or ( n361243 , n361228 , n41108 );
buf ( n361244 , n360954 );
buf ( n361245 , n39891 );
nand ( n361246 , n361244 , n361245 );
buf ( n361247 , n361246 );
buf ( n361248 , n361247 );
nand ( n41115 , n361243 , n361248 );
buf ( n361250 , n41115 );
buf ( n361251 , n361250 );
not ( n361252 , n361251 );
not ( n41119 , n360601 );
buf ( n361254 , n360616 );
not ( n361255 , n361254 );
buf ( n361256 , n359979 );
not ( n361257 , n361256 );
or ( n361258 , n361255 , n361257 );
buf ( n361259 , n39870 );
buf ( n361260 , n360613 );
nand ( n361261 , n361259 , n361260 );
buf ( n361262 , n361261 );
buf ( n361263 , n361262 );
nand ( n361264 , n361258 , n361263 );
buf ( n361265 , n361264 );
not ( n361266 , n361265 );
or ( n361267 , n41119 , n361266 );
nand ( n361268 , n360577 , n41080 );
nand ( n361269 , n361267 , n361268 );
buf ( n361270 , n361269 );
not ( n41132 , n361270 );
or ( n41133 , n361252 , n41132 );
buf ( n361273 , n361269 );
buf ( n361274 , n361250 );
or ( n361275 , n361273 , n361274 );
buf ( n361276 , n39952 );
not ( n41138 , n361276 );
buf ( n361278 , n361158 );
not ( n361279 , n361278 );
or ( n41141 , n41138 , n361279 );
buf ( n361281 , n39966 );
not ( n361282 , n361281 );
buf ( n361283 , n40202 );
not ( n361284 , n361283 );
or ( n361285 , n361282 , n361284 );
buf ( n361286 , n40798 );
buf ( n361287 , n360126 );
nand ( n41149 , n361286 , n361287 );
buf ( n361289 , n41149 );
buf ( n361290 , n361289 );
nand ( n41152 , n361285 , n361290 );
buf ( n361292 , n41152 );
buf ( n361293 , n361292 );
buf ( n361294 , n360168 );
nand ( n41156 , n361293 , n361294 );
buf ( n361296 , n41156 );
buf ( n361297 , n361296 );
nand ( n361298 , n41141 , n361297 );
buf ( n361299 , n361298 );
buf ( n361300 , n361299 );
nand ( n361301 , n361275 , n361300 );
buf ( n361302 , n361301 );
buf ( n361303 , n361302 );
nand ( n361304 , n41133 , n361303 );
buf ( n361305 , n361304 );
buf ( n361306 , n361305 );
xor ( n361307 , n41092 , n361306 );
buf ( n361308 , n361307 );
buf ( n361309 , n361308 );
and ( n361310 , n41062 , n361309 );
and ( n361311 , n361113 , n361195 );
or ( n41173 , n361310 , n361311 );
buf ( n361313 , n41173 );
buf ( n41175 , n361313 );
xor ( n41176 , n360970 , n41175 );
xor ( n361316 , n361128 , n361166 );
and ( n41178 , n361316 , n361192 );
and ( n361318 , n361128 , n361166 );
or ( n41180 , n41178 , n361318 );
buf ( n361320 , n41180 );
buf ( n361321 , n361320 );
buf ( n361322 , n39891 );
not ( n361323 , n361322 );
buf ( n361324 , n360437 );
not ( n41186 , n361324 );
or ( n361326 , n361323 , n41186 );
buf ( n361327 , n360939 );
buf ( n361328 , n359919 );
nand ( n361329 , n361327 , n361328 );
buf ( n361330 , n361329 );
buf ( n361331 , n361330 );
nand ( n41193 , n361326 , n361331 );
buf ( n361333 , n41193 );
buf ( n361334 , n361333 );
buf ( n361335 , n39217 );
not ( n361336 , n361335 );
buf ( n361337 , n360653 );
not ( n41199 , n361337 );
or ( n361339 , n361336 , n41199 );
buf ( n41201 , n361184 );
buf ( n361341 , n359307 );
nand ( n41203 , n41201 , n361341 );
buf ( n361343 , n41203 );
buf ( n361344 , n361343 );
nand ( n361345 , n361339 , n361344 );
buf ( n361346 , n361345 );
buf ( n361347 , n361346 );
xor ( n361348 , n361334 , n361347 );
buf ( n361349 , n39952 );
not ( n361350 , n361349 );
buf ( n361351 , n360452 );
not ( n41213 , n361351 );
or ( n41214 , n361350 , n41213 );
buf ( n361354 , n361143 );
buf ( n361355 , n360168 );
nand ( n41217 , n361354 , n361355 );
buf ( n361357 , n41217 );
buf ( n361358 , n361357 );
nand ( n41220 , n41214 , n361358 );
buf ( n41221 , n41220 );
buf ( n361361 , n41221 );
xor ( n41223 , n361348 , n361361 );
buf ( n361363 , n41223 );
buf ( n361364 , n361363 );
xor ( n41226 , n361321 , n361364 );
xor ( n361366 , n361221 , n361225 );
and ( n361367 , n361366 , n361306 );
and ( n41229 , n361221 , n361225 );
or ( n361369 , n361367 , n41229 );
buf ( n361370 , n361369 );
buf ( n361371 , n361370 );
xor ( n361372 , n41226 , n361371 );
buf ( n361373 , n361372 );
buf ( n361374 , n361373 );
and ( n41236 , n41176 , n361374 );
and ( n361376 , n360970 , n41175 );
or ( n361377 , n41236 , n361376 );
buf ( n361378 , n361377 );
buf ( n361379 , n361378 );
xor ( n361380 , n360800 , n360825 );
and ( n41242 , n361380 , n360967 );
and ( n361382 , n360800 , n360825 );
or ( n361383 , n41242 , n361382 );
buf ( n361384 , n361383 );
buf ( n361385 , n361384 );
xor ( n361386 , n360634 , n40516 );
xor ( n41248 , n361386 , n360660 );
buf ( n361388 , n41248 );
xor ( n361389 , n361334 , n361347 );
and ( n361390 , n361389 , n361361 );
and ( n41252 , n361334 , n361347 );
or ( n41253 , n361390 , n41252 );
buf ( n361393 , n41253 );
buf ( n361394 , n361393 );
xor ( n361395 , n361388 , n361394 );
xor ( n361396 , n360419 , n360445 );
xor ( n41258 , n361396 , n360463 );
buf ( n361398 , n41258 );
buf ( n361399 , n361398 );
xor ( n41261 , n361395 , n361399 );
buf ( n361401 , n41261 );
buf ( n361402 , n361401 );
xor ( n41264 , n361385 , n361402 );
xor ( n41265 , n361321 , n361364 );
and ( n361405 , n41265 , n361371 );
and ( n41267 , n361321 , n361364 );
or ( n41268 , n361405 , n41267 );
buf ( n361408 , n41268 );
buf ( n361409 , n361408 );
xor ( n41271 , n41264 , n361409 );
buf ( n361411 , n41271 );
buf ( n361412 , n361411 );
or ( n41274 , n361379 , n361412 );
buf ( n361414 , n41274 );
buf ( n361415 , n361414 );
xor ( n41277 , n361388 , n361394 );
and ( n361417 , n41277 , n361399 );
and ( n361418 , n361388 , n361394 );
or ( n41280 , n361417 , n361418 );
buf ( n361420 , n41280 );
buf ( n361421 , n360467 );
buf ( n361422 , n360321 );
and ( n361423 , n361421 , n361422 );
not ( n41285 , n361421 );
buf ( n361425 , n360324 );
and ( n361426 , n41285 , n361425 );
nor ( n361427 , n361423 , n361426 );
buf ( n361428 , n361427 );
xnor ( n361429 , n361428 , n40540 );
xor ( n361430 , n361420 , n361429 );
buf ( n361431 , n360212 );
buf ( n361432 , n360174 );
and ( n361433 , n361431 , n361432 );
not ( n41295 , n361431 );
buf ( n361435 , n360218 );
and ( n41297 , n41295 , n361435 );
nor ( n361437 , n361433 , n41297 );
buf ( n361438 , n361437 );
buf ( n361439 , n361438 );
buf ( n361440 , n360250 );
xnor ( n41302 , n361439 , n361440 );
buf ( n361442 , n41302 );
xnor ( n41304 , n361430 , n361442 );
buf ( n361444 , n41304 );
xor ( n361445 , n361385 , n361402 );
and ( n41307 , n361445 , n361409 );
and ( n361447 , n361385 , n361402 );
or ( n41309 , n41307 , n361447 );
buf ( n361449 , n41309 );
buf ( n361450 , n361449 );
nor ( n41312 , n361444 , n361450 );
buf ( n41313 , n41312 );
buf ( n361453 , n41313 );
not ( n41315 , n361453 );
buf ( n361455 , n41315 );
buf ( n361456 , n361455 );
nand ( n41318 , n361415 , n361456 );
buf ( n361458 , n41318 );
buf ( n361459 , n361458 );
buf ( n361460 , n361442 );
not ( n361461 , n361460 );
buf ( n361462 , n361429 );
not ( n41324 , n361462 );
buf ( n41325 , n41324 );
buf ( n361465 , n41325 );
not ( n41327 , n361465 );
or ( n361467 , n361461 , n41327 );
buf ( n361468 , n361420 );
nand ( n41330 , n361467 , n361468 );
buf ( n361470 , n41330 );
buf ( n361471 , n361470 );
buf ( n361472 , n361442 );
not ( n361473 , n361472 );
buf ( n361474 , n361429 );
nand ( n361475 , n361473 , n361474 );
buf ( n361476 , n361475 );
buf ( n361477 , n361476 );
and ( n361478 , n361471 , n361477 );
buf ( n361479 , n361478 );
buf ( n361480 , n361479 );
xor ( n361481 , n360009 , n40219 );
xor ( n361482 , n361481 , n360675 );
buf ( n361483 , n361482 );
buf ( n361484 , n361483 );
nand ( n41346 , n361480 , n361484 );
buf ( n361486 , n41346 );
buf ( n361487 , n361486 );
not ( n361488 , n361487 );
buf ( n361489 , n361488 );
buf ( n361490 , n361489 );
nor ( n361491 , n361459 , n361490 );
buf ( n361492 , n361491 );
buf ( n361493 , n361492 );
not ( n361494 , n361493 );
not ( n361495 , n40364 );
not ( n41354 , n361495 );
not ( n361497 , n39754 );
or ( n41356 , n41354 , n361497 );
buf ( n361499 , n359268 );
not ( n361500 , n361499 );
buf ( n361501 , n361500 );
not ( n41360 , n361501 );
not ( n361503 , n361495 );
or ( n361504 , n41360 , n361503 );
buf ( n41363 , n354651 );
not ( n361506 , n41363 );
not ( n361507 , n34679 );
or ( n41366 , n361506 , n361507 );
not ( n361509 , n359221 );
nand ( n41368 , n41366 , n361509 );
nand ( n361511 , n361504 , n41368 );
not ( n41370 , n361511 );
nand ( n41371 , n41356 , n41370 );
buf ( n361514 , n34694 );
buf ( n361515 , n361514 );
not ( n41374 , n361515 );
buf ( n361517 , n354643 );
buf ( n361518 , n361517 );
buf ( n361519 , n361518 );
buf ( n361520 , n361519 );
nand ( n361521 , n41374 , n361520 );
buf ( n361522 , n361521 );
and ( n361523 , n41371 , n361522 );
not ( n361524 , n41371 );
not ( n41383 , n361522 );
and ( n41384 , n361524 , n41383 );
nor ( n41385 , n361523 , n41384 );
buf ( n41386 , n41385 );
buf ( n361529 , n41386 );
not ( n361530 , n361529 );
buf ( n361531 , n361530 );
buf ( n361532 , n361531 );
not ( n361533 , n361532 );
buf ( n361534 , n361533 );
buf ( n361535 , n361534 );
buf ( n361536 , n361535 );
buf ( n361537 , n361536 );
buf ( n361538 , n361537 );
not ( n361539 , n361538 );
buf ( n361540 , n361539 );
buf ( n361541 , n361540 );
not ( n361542 , n361541 );
buf ( n361543 , n360116 );
not ( n41402 , n361543 );
or ( n361545 , n361542 , n41402 );
buf ( n361546 , n40005 );
buf ( n41405 , n361546 );
buf ( n41406 , n41405 );
buf ( n361549 , n41406 );
buf ( n361550 , n361537 );
nand ( n361551 , n361549 , n361550 );
buf ( n361552 , n361551 );
buf ( n361553 , n361552 );
nand ( n361554 , n361545 , n361553 );
buf ( n361555 , n361554 );
buf ( n361556 , n361555 );
not ( n361557 , n35448 );
not ( n41416 , n361557 );
not ( n41417 , n39180 );
or ( n41418 , n41416 , n41417 );
buf ( n41419 , n34679 );
buf ( n41420 , n41419 );
nand ( n361563 , n41418 , n41420 );
not ( n361564 , n41363 );
not ( n41423 , n361564 );
nand ( n361566 , n41423 , n361509 );
and ( n361567 , n361563 , n361566 );
not ( n41426 , n361563 );
not ( n41427 , n361566 );
and ( n41428 , n41426 , n41427 );
nor ( n41429 , n361567 , n41428 );
not ( n41430 , n41429 );
not ( n361573 , n41430 );
not ( n361574 , n41385 );
not ( n41433 , n361574 );
not ( n361576 , n41433 );
or ( n361577 , n361573 , n361576 );
not ( n41436 , n41385 );
nand ( n361579 , n41436 , n41429 );
nand ( n361580 , n361577 , n361579 );
buf ( n361581 , n41419 );
buf ( n361582 , n361557 );
nand ( n41441 , n361581 , n361582 );
buf ( n361584 , n41441 );
and ( n361585 , n359654 , n361584 );
not ( n361586 , n359654 );
not ( n41445 , n361584 );
and ( n41446 , n361586 , n41445 );
nor ( n41447 , n361585 , n41446 );
buf ( n41448 , n41447 );
not ( n361591 , n41448 );
and ( n361592 , n41429 , n361591 );
not ( n41451 , n41429 );
not ( n41452 , n41447 );
buf ( n361595 , n41452 );
not ( n41454 , n361595 );
buf ( n361597 , n41454 );
and ( n361598 , n41451 , n361597 );
nor ( n41457 , n361592 , n361598 );
nand ( n361600 , n361580 , n41457 );
buf ( n361601 , n361600 );
buf ( n361602 , n361601 );
buf ( n361603 , n361602 );
buf ( n361604 , n361603 );
not ( n361605 , n361604 );
buf ( n361606 , n361605 );
buf ( n361607 , n361606 );
buf ( n361608 , n361607 );
buf ( n361609 , n361608 );
buf ( n361610 , n361609 );
nand ( n361611 , n361556 , n361610 );
buf ( n361612 , n361611 );
not ( n361613 , n361540 );
not ( n41472 , n40089 );
not ( n361615 , n41472 );
or ( n41474 , n361613 , n361615 );
not ( n361617 , n40091 );
buf ( n361618 , n361617 );
buf ( n361619 , n361537 );
nand ( n361620 , n361618 , n361619 );
buf ( n361621 , n361620 );
nand ( n41480 , n41474 , n361621 );
buf ( n41481 , n41457 );
buf ( n41482 , n41481 );
not ( n361625 , n41482 );
not ( n361626 , n361625 );
not ( n41485 , n361626 );
nand ( n361628 , n41480 , n41485 );
nand ( n361629 , n361612 , n361628 );
buf ( n361630 , n361629 );
buf ( n361631 , n39620 );
buf ( n361632 , n361631 );
buf ( n41491 , n358594 );
buf ( n361634 , n41491 );
buf ( n361635 , n38539 );
not ( n41494 , n361635 );
buf ( n361637 , n41494 );
buf ( n361638 , n361637 );
nand ( n361639 , n361634 , n361638 );
buf ( n361640 , n361639 );
buf ( n361641 , n361640 );
not ( n361642 , n361641 );
buf ( n361643 , n361642 );
buf ( n361644 , n361643 );
not ( n41503 , n361644 );
buf ( n361646 , n360343 );
not ( n361647 , n361646 );
buf ( n361648 , n361647 );
buf ( n361649 , n361648 );
not ( n41508 , n361649 );
or ( n361651 , n41503 , n41508 );
buf ( n361652 , n361648 );
not ( n361653 , n361652 );
buf ( n361654 , n361653 );
buf ( n361655 , n361654 );
buf ( n361656 , n361640 );
nand ( n41515 , n361655 , n361656 );
buf ( n361658 , n41515 );
buf ( n41517 , n361658 );
nand ( n361660 , n361651 , n41517 );
buf ( n361661 , n361660 );
buf ( n361662 , n361661 );
not ( n361663 , n361662 );
buf ( n361664 , n361663 );
buf ( n361665 , n361664 );
not ( n41524 , n361665 );
buf ( n361667 , n41524 );
buf ( n361668 , n361667 );
buf ( n41527 , n361668 );
buf ( n41528 , n41527 );
buf ( n361671 , n41528 );
buf ( n361672 , n361671 );
buf ( n361673 , n361672 );
buf ( n361674 , n361673 );
and ( n361675 , n361632 , n361674 );
not ( n41534 , n361632 );
buf ( n361677 , n361673 );
not ( n361678 , n361677 );
buf ( n361679 , n361678 );
buf ( n361680 , n361679 );
and ( n361681 , n41534 , n361680 );
nor ( n41540 , n361675 , n361681 );
buf ( n361683 , n41540 );
not ( n361684 , n361683 );
buf ( n361685 , n39592 );
not ( n361686 , n361685 );
buf ( n361687 , n361686 );
not ( n41546 , n361687 );
and ( n41547 , n361684 , n41546 );
buf ( n361690 , n39621 );
not ( n361691 , n361690 );
buf ( n361692 , n359020 );
not ( n41551 , n361692 );
buf ( n361694 , n41551 );
not ( n41553 , n361694 );
not ( n41554 , n31757 );
or ( n361697 , n41553 , n41554 );
not ( n361698 , n37181 );
nand ( n41557 , n361697 , n361698 );
buf ( n361700 , n37465 );
not ( n361701 , n361700 );
buf ( n361702 , n357557 );
nand ( n361703 , n361701 , n361702 );
buf ( n361704 , n361703 );
and ( n41563 , n361704 , n357567 );
and ( n361706 , n41557 , n41563 );
not ( n41565 , n41557 );
not ( n361708 , n41563 );
and ( n41567 , n41565 , n361708 );
nor ( n361710 , n361706 , n41567 );
buf ( n41569 , n361710 );
not ( n361712 , n41569 );
buf ( n361713 , n361712 );
not ( n361714 , n361713 );
or ( n41573 , n361691 , n361714 );
buf ( n361716 , n361710 );
buf ( n361717 , n361716 );
buf ( n361718 , n361717 );
buf ( n361719 , n361631 );
nand ( n361720 , n361718 , n361719 );
buf ( n361721 , n361720 );
buf ( n361722 , n361721 );
nand ( n41581 , n41573 , n361722 );
buf ( n41582 , n41581 );
not ( n361725 , n41582 );
nor ( n361726 , n361725 , n39707 );
nor ( n41585 , n41547 , n361726 );
buf ( n361728 , n41585 );
not ( n361729 , n41491 );
not ( n41588 , n360343 );
or ( n41589 , n361729 , n41588 );
buf ( n361732 , n361637 );
nand ( n41591 , n41589 , n361732 );
buf ( n361734 , n358608 );
not ( n361735 , n361734 );
buf ( n361736 , n358631 );
not ( n41595 , n361736 );
buf ( n361738 , n41595 );
buf ( n361739 , n361738 );
nor ( n41598 , n361735 , n361739 );
buf ( n41599 , n41598 );
and ( n361742 , n41591 , n41599 );
not ( n41601 , n41591 );
buf ( n361744 , n41599 );
not ( n41603 , n361744 );
buf ( n361746 , n41603 );
and ( n41605 , n41601 , n361746 );
nor ( n361748 , n361742 , n41605 );
buf ( n41607 , n361748 );
buf ( n361750 , n41607 );
not ( n361751 , n361750 );
buf ( n361752 , n361751 );
not ( n361753 , n361752 );
buf ( n361754 , n359950 );
not ( n41613 , n361754 );
or ( n361756 , n361753 , n41613 );
not ( n41615 , n41607 );
not ( n41616 , n41615 );
buf ( n41617 , n41616 );
buf ( n361760 , n359944 );
buf ( n361761 , n361760 );
buf ( n361762 , n361761 );
buf ( n361763 , n361762 );
not ( n41622 , n361763 );
buf ( n41623 , n41622 );
buf ( n361766 , n41623 );
nand ( n41625 , n41617 , n361766 );
buf ( n41626 , n41625 );
buf ( n41627 , n41626 );
nand ( n41628 , n361756 , n41627 );
buf ( n41629 , n41628 );
buf ( n361772 , n41629 );
not ( n41631 , n361772 );
buf ( n361774 , n359919 );
not ( n41633 , n361774 );
or ( n361776 , n41631 , n41633 );
buf ( n361777 , n359950 );
not ( n41636 , n361777 );
buf ( n361779 , n38911 );
not ( n41638 , n361779 );
buf ( n361781 , n41638 );
not ( n41640 , n361781 );
not ( n41641 , n360343 );
or ( n41642 , n41640 , n41641 );
buf ( n361785 , n38540 );
not ( n41644 , n361785 );
buf ( n361787 , n361738 );
nor ( n41646 , n41644 , n361787 );
buf ( n41647 , n41646 );
nand ( n361790 , n41642 , n41647 );
buf ( n361791 , n358643 );
buf ( n41650 , n361791 );
buf ( n361793 , n41650 );
buf ( n41652 , n38552 );
nand ( n41653 , n361793 , n41652 );
not ( n41654 , n41653 );
and ( n41655 , n361790 , n41654 );
not ( n41656 , n361790 );
and ( n41657 , n41656 , n41653 );
nor ( n361800 , n41655 , n41657 );
not ( n41659 , n361800 );
not ( n361802 , n41659 );
buf ( n41661 , n361802 );
buf ( n41662 , n41661 );
buf ( n41663 , n41662 );
buf ( n41664 , n41663 );
not ( n41665 , n41664 );
buf ( n41666 , n41665 );
buf ( n361809 , n41666 );
not ( n41668 , n361809 );
or ( n361811 , n41636 , n41668 );
buf ( n361812 , n41663 );
buf ( n361813 , n359955 );
nand ( n361814 , n361812 , n361813 );
buf ( n361815 , n361814 );
buf ( n361816 , n361815 );
nand ( n361817 , n361811 , n361816 );
buf ( n361818 , n361817 );
buf ( n361819 , n361818 );
buf ( n361820 , n39891 );
nand ( n361821 , n361819 , n361820 );
buf ( n361822 , n361821 );
buf ( n361823 , n361822 );
nand ( n361824 , n361776 , n361823 );
buf ( n361825 , n361824 );
buf ( n361826 , n361825 );
xor ( n41685 , n361728 , n361826 );
buf ( n361828 , n39217 );
not ( n361829 , n361828 );
buf ( n361830 , n355582 );
not ( n41689 , n361830 );
buf ( n361832 , n360851 );
not ( n361833 , n361832 );
or ( n41692 , n41689 , n361833 );
buf ( n361835 , n360857 );
buf ( n361836 , n40945 );
nand ( n41695 , n361835 , n361836 );
buf ( n361838 , n41695 );
buf ( n361839 , n361838 );
nand ( n361840 , n41692 , n361839 );
buf ( n361841 , n361840 );
buf ( n361842 , n361841 );
not ( n41701 , n361842 );
or ( n41702 , n361829 , n41701 );
buf ( n361845 , n355582 );
not ( n41704 , n361845 );
buf ( n361847 , n40756 );
not ( n361848 , n361847 );
or ( n41707 , n41704 , n361848 );
buf ( n361850 , n360893 );
buf ( n361851 , n35547 );
buf ( n361852 , n361851 );
nand ( n361853 , n361850 , n361852 );
buf ( n361854 , n361853 );
buf ( n361855 , n361854 );
nand ( n41714 , n41707 , n361855 );
buf ( n361857 , n41714 );
buf ( n361858 , n361857 );
buf ( n361859 , n359307 );
nand ( n41718 , n361858 , n361859 );
buf ( n361861 , n41718 );
buf ( n361862 , n361861 );
nand ( n361863 , n41702 , n361862 );
buf ( n361864 , n361863 );
buf ( n361865 , n361864 );
and ( n41724 , n41685 , n361865 );
and ( n361867 , n361728 , n361826 );
or ( n41726 , n41724 , n361867 );
buf ( n361869 , n41726 );
buf ( n361870 , n361869 );
xor ( n41729 , n361630 , n361870 );
buf ( n361872 , n361060 );
not ( n361873 , n361872 );
buf ( n361874 , n40893 );
not ( n361875 , n361874 );
buf ( n361876 , n39655 );
not ( n41735 , n361876 );
or ( n361878 , n361875 , n41735 );
buf ( n361879 , n39658 );
buf ( n361880 , n361026 );
nand ( n361881 , n361879 , n361880 );
buf ( n361882 , n361881 );
buf ( n361883 , n361882 );
nand ( n361884 , n361878 , n361883 );
buf ( n361885 , n361884 );
buf ( n361886 , n361885 );
not ( n361887 , n361886 );
or ( n361888 , n361873 , n361887 );
buf ( n361889 , n361022 );
buf ( n361890 , n40893 );
not ( n361891 , n361890 );
buf ( n361892 , n359784 );
not ( n361893 , n361892 );
or ( n361894 , n361891 , n361893 );
buf ( n361895 , n359781 );
buf ( n361896 , n361026 );
nand ( n361897 , n361895 , n361896 );
buf ( n361898 , n361897 );
buf ( n361899 , n361898 );
nand ( n361900 , n361894 , n361899 );
buf ( n361901 , n361900 );
buf ( n361902 , n361901 );
nand ( n361903 , n361889 , n361902 );
buf ( n361904 , n361903 );
buf ( n361905 , n361904 );
nand ( n41764 , n361888 , n361905 );
buf ( n361907 , n41764 );
buf ( n361908 , n361907 );
xor ( n361909 , n41729 , n361908 );
buf ( n361910 , n361909 );
not ( n361911 , n41448 );
buf ( n41770 , n361911 );
not ( n41771 , n41770 );
buf ( n41772 , n41771 );
buf ( n361915 , n41772 );
buf ( n41774 , n361915 );
buf ( n361917 , n41774 );
buf ( n41776 , n361917 );
not ( n41777 , n41776 );
buf ( n41778 , n41777 );
buf ( n361921 , n41778 );
not ( n361922 , n361921 );
buf ( n361923 , n359147 );
not ( n41782 , n361923 );
or ( n41783 , n361922 , n41782 );
buf ( n361926 , n360624 );
buf ( n361927 , n361917 );
nand ( n361928 , n361926 , n361927 );
buf ( n361929 , n361928 );
buf ( n361930 , n361929 );
nand ( n361931 , n41783 , n361930 );
buf ( n361932 , n361931 );
buf ( n361933 , n360023 );
buf ( n361934 , n361501 );
not ( n41793 , n361934 );
buf ( n361936 , n360026 );
nand ( n41795 , n41793 , n361936 );
buf ( n361938 , n41795 );
buf ( n41797 , n361938 );
not ( n41798 , n41797 );
buf ( n41799 , n41798 );
buf ( n361942 , n41799 );
and ( n41801 , n361933 , n361942 );
not ( n361944 , n361933 );
buf ( n41803 , n361938 );
and ( n41804 , n361944 , n41803 );
nor ( n361947 , n41801 , n41804 );
buf ( n361948 , n361947 );
or ( n41807 , n41452 , n361948 );
buf ( n361950 , n41807 );
buf ( n361951 , n342334 );
not ( n41810 , n361951 );
buf ( n361953 , n41810 );
buf ( n361954 , n361953 );
not ( n361955 , n361948 );
buf ( n361956 , n361955 );
and ( n361957 , n361954 , n361956 );
not ( n41816 , n361954 );
buf ( n361959 , n361948 );
and ( n41818 , n41816 , n361959 );
nor ( n41819 , n361957 , n41818 );
buf ( n361962 , n41819 );
buf ( n361963 , n361962 );
buf ( n361964 , n41452 );
buf ( n361965 , n361948 );
nand ( n361966 , n361964 , n361965 );
buf ( n361967 , n361966 );
buf ( n361968 , n361967 );
nand ( n41827 , n361950 , n361963 , n361968 );
buf ( n361970 , n41827 );
buf ( n361971 , n361970 );
not ( n41830 , n361971 );
not ( n41831 , n41830 );
buf ( n361974 , n41831 );
buf ( n361975 , n361962 );
not ( n41834 , n361975 );
buf ( n41835 , n41834 );
not ( n41836 , n41835 );
buf ( n361979 , n41836 );
nand ( n361980 , n361974 , n361979 );
buf ( n361981 , n361980 );
and ( n361982 , n361932 , n361981 );
not ( n41841 , n361982 );
buf ( n361984 , n41371 );
buf ( n361985 , n41383 );
and ( n41844 , n361984 , n361985 );
not ( n361987 , n361984 );
buf ( n361988 , n361522 );
and ( n41847 , n361987 , n361988 );
nor ( n361990 , n41844 , n41847 );
buf ( n361991 , n361990 );
not ( n361992 , n361991 );
and ( n41851 , n361519 , n361495 );
not ( n361994 , n41851 );
not ( n361995 , n39754 );
or ( n41854 , n361994 , n361995 );
and ( n361997 , n361511 , n361519 );
nor ( n361998 , n361997 , n361514 );
nand ( n41857 , n41854 , n361998 );
nand ( n41858 , n354733 , n354456 );
not ( n362001 , n41858 );
and ( n362002 , n41857 , n362001 );
not ( n41861 , n41857 );
and ( n41862 , n41861 , n41858 );
nor ( n362005 , n362002 , n41862 );
not ( n41864 , n362005 );
or ( n362007 , n361992 , n41864 );
not ( n362008 , n362005 );
not ( n41867 , n361991 );
nand ( n41868 , n362008 , n41867 );
nand ( n41869 , n362007 , n41868 );
buf ( n362012 , n361009 );
not ( n362013 , n362012 );
buf ( n362014 , n362005 );
not ( n362015 , n362014 );
or ( n362016 , n362013 , n362015 );
nand ( n41875 , n362008 , n40871 );
buf ( n362018 , n41875 );
nand ( n362019 , n362016 , n362018 );
buf ( n362020 , n362019 );
nand ( n362021 , n41869 , n362020 );
buf ( n41880 , n362021 );
buf ( n41881 , n41880 );
buf ( n41882 , n41881 );
buf ( n362025 , n41882 );
not ( n41884 , n362025 );
buf ( n362027 , n41884 );
buf ( n362028 , n362027 );
buf ( n41887 , n362028 );
buf ( n362030 , n41887 );
buf ( n362031 , n362030 );
not ( n41890 , n362031 );
buf ( n362033 , n40871 );
buf ( n41892 , n362033 );
buf ( n362035 , n41892 );
not ( n41894 , n362035 );
buf ( n362037 , n41894 );
buf ( n362038 , n362037 );
buf ( n362039 , n361073 );
and ( n41898 , n362038 , n362039 );
not ( n362041 , n362038 );
buf ( n41900 , n39832 );
and ( n41901 , n362041 , n41900 );
nor ( n362044 , n41898 , n41901 );
buf ( n362045 , n362044 );
buf ( n362046 , n362045 );
not ( n41905 , n362046 );
or ( n362048 , n41890 , n41905 );
not ( n41907 , n359974 );
and ( n362050 , n41907 , n41892 );
not ( n362051 , n41907 );
and ( n362052 , n362051 , n362037 );
or ( n41911 , n362050 , n362052 );
buf ( n362054 , n41911 );
buf ( n41913 , n41869 );
not ( n41914 , n41913 );
buf ( n41915 , n41914 );
buf ( n41916 , n41915 );
buf ( n41917 , n41916 );
buf ( n41918 , n41917 );
buf ( n362061 , n41918 );
not ( n362062 , n362061 );
buf ( n362063 , n362062 );
buf ( n362064 , n362063 );
not ( n362065 , n362064 );
buf ( n362066 , n362065 );
buf ( n362067 , n362066 );
nand ( n362068 , n362054 , n362067 );
buf ( n362069 , n362068 );
buf ( n362070 , n362069 );
nand ( n362071 , n362048 , n362070 );
buf ( n362072 , n362071 );
nor ( n41931 , n41841 , n362072 );
not ( n41932 , n41931 );
not ( n362075 , n361982 );
nand ( n362076 , n362075 , n362072 );
nand ( n41935 , n41932 , n362076 );
buf ( n362078 , n41585 );
not ( n41937 , n362078 );
buf ( n362080 , n41937 );
buf ( n362081 , n362080 );
buf ( n362082 , n39592 );
not ( n41941 , n362082 );
buf ( n362084 , n39621 );
buf ( n362085 , n361751 );
and ( n362086 , n362084 , n362085 );
not ( n41945 , n362084 );
not ( n41946 , n41615 );
buf ( n362089 , n41946 );
and ( n362090 , n41945 , n362089 );
nor ( n362091 , n362086 , n362090 );
buf ( n362092 , n362091 );
buf ( n362093 , n362092 );
not ( n362094 , n362093 );
buf ( n362095 , n362094 );
buf ( n362096 , n362095 );
not ( n362097 , n362096 );
or ( n41956 , n41941 , n362097 );
buf ( n362099 , n39707 );
buf ( n362100 , n361683 );
or ( n41959 , n362099 , n362100 );
buf ( n362102 , n41959 );
buf ( n362103 , n362102 );
nand ( n41962 , n41956 , n362103 );
buf ( n362105 , n41962 );
buf ( n362106 , n362105 );
xor ( n41965 , n362081 , n362106 );
buf ( n362108 , n39891 );
not ( n362109 , n362108 );
buf ( n362110 , n359950 );
not ( n362111 , n362110 );
nand ( n362112 , n358649 , n38463 );
buf ( n362113 , n362112 );
and ( n41972 , n362113 , n361793 );
not ( n41973 , n41972 );
not ( n362116 , n361790 );
not ( n41975 , n362116 );
not ( n41976 , n41975 );
or ( n41977 , n41973 , n41976 );
not ( n41978 , n41652 );
nor ( n41979 , n362113 , n41978 );
and ( n41980 , n362116 , n41979 );
and ( n41981 , n362113 , n41978 );
not ( n41982 , n362113 );
not ( n41983 , n41652 );
nor ( n41984 , n41983 , n361793 );
and ( n362127 , n41982 , n41984 );
or ( n41986 , n41981 , n362127 );
nor ( n41987 , n41980 , n41986 );
nand ( n362130 , n41977 , n41987 );
buf ( n362131 , n362130 );
buf ( n41990 , n362131 );
buf ( n362133 , n41990 );
buf ( n41992 , n362133 );
buf ( n362135 , n41992 );
buf ( n362136 , n362135 );
buf ( n362137 , n362136 );
not ( n362138 , n362137 );
buf ( n362139 , n362138 );
buf ( n362140 , n362139 );
not ( n362141 , n362140 );
or ( n41999 , n362111 , n362141 );
buf ( n362143 , n362133 );
not ( n362144 , n362143 );
buf ( n362145 , n362144 );
buf ( n362146 , n362145 );
not ( n362147 , n362146 );
buf ( n362148 , n362147 );
buf ( n362149 , n362148 );
buf ( n362150 , n359955 );
nand ( n362151 , n362149 , n362150 );
buf ( n362152 , n362151 );
buf ( n362153 , n362152 );
nand ( n362154 , n41999 , n362153 );
buf ( n362155 , n362154 );
buf ( n42011 , n362155 );
not ( n42012 , n42011 );
or ( n42013 , n362109 , n42012 );
buf ( n42014 , n359919 );
buf ( n362160 , n361818 );
nand ( n42016 , n42014 , n362160 );
buf ( n42017 , n42016 );
buf ( n362163 , n42017 );
nand ( n42019 , n42013 , n362163 );
buf ( n42020 , n42019 );
buf ( n362166 , n42020 );
xor ( n42022 , n41965 , n362166 );
buf ( n362168 , n42022 );
xor ( n362169 , n41935 , n362168 );
buf ( n362170 , n362169 );
not ( n362171 , n362170 );
buf ( n362172 , n362171 );
buf ( n362173 , n362172 );
not ( n42029 , n362173 );
buf ( n362175 , n41830 );
not ( n362176 , n362175 );
buf ( n362177 , n41778 );
not ( n362178 , n362177 );
not ( n362179 , n40899 );
buf ( n362180 , n362179 );
not ( n42036 , n362180 );
or ( n42037 , n362178 , n42036 );
buf ( n362183 , n361617 );
buf ( n362184 , n361917 );
nand ( n42040 , n362183 , n362184 );
buf ( n362186 , n42040 );
buf ( n362187 , n362186 );
nand ( n362188 , n42037 , n362187 );
buf ( n362189 , n362188 );
buf ( n362190 , n362189 );
not ( n362191 , n362190 );
or ( n362192 , n362176 , n362191 );
buf ( n362193 , n361932 );
buf ( n362194 , n41835 );
nand ( n362195 , n362193 , n362194 );
buf ( n362196 , n362195 );
buf ( n362197 , n362196 );
nand ( n362198 , n362192 , n362197 );
buf ( n362199 , n362198 );
buf ( n362200 , n362199 );
buf ( n362201 , n362066 );
not ( n362202 , n362201 );
buf ( n362203 , n362045 );
not ( n42059 , n362203 );
or ( n362205 , n362202 , n42059 );
buf ( n362206 , n41892 );
not ( n362207 , n362206 );
not ( n362208 , n359756 );
buf ( n362209 , n362208 );
not ( n42065 , n362209 );
or ( n362211 , n362207 , n42065 );
not ( n362212 , n359756 );
not ( n42068 , n362212 );
buf ( n362214 , n42068 );
buf ( n362215 , n362037 );
nand ( n42071 , n362214 , n362215 );
buf ( n42072 , n42071 );
buf ( n362218 , n42072 );
nand ( n42074 , n362211 , n362218 );
buf ( n42075 , n42074 );
buf ( n362221 , n42075 );
buf ( n42077 , n362030 );
nand ( n42078 , n362221 , n42077 );
buf ( n362224 , n42078 );
buf ( n362225 , n362224 );
nand ( n42081 , n362205 , n362225 );
buf ( n42082 , n42081 );
buf ( n362228 , n42082 );
xor ( n42084 , n362200 , n362228 );
buf ( n362230 , n39952 );
not ( n362231 , n362230 );
buf ( n362232 , n39966 );
not ( n42088 , n362232 );
buf ( n362234 , n362139 );
not ( n362235 , n362234 );
or ( n42091 , n42088 , n362235 );
buf ( n42092 , n362148 );
buf ( n362238 , n39963 );
nand ( n362239 , n42092 , n362238 );
buf ( n362240 , n362239 );
buf ( n362241 , n362240 );
nand ( n362242 , n42091 , n362241 );
buf ( n362243 , n362242 );
buf ( n362244 , n362243 );
not ( n362245 , n362244 );
or ( n362246 , n362231 , n362245 );
buf ( n362247 , n40059 );
buf ( n362248 , n39966 );
not ( n362249 , n362248 );
buf ( n362250 , n41666 );
not ( n42106 , n362250 );
or ( n42107 , n362249 , n42106 );
buf ( n362253 , n361802 );
buf ( n362254 , n39963 );
nand ( n42110 , n362253 , n362254 );
buf ( n362256 , n42110 );
buf ( n362257 , n362256 );
nand ( n42113 , n42107 , n362257 );
buf ( n42114 , n42113 );
buf ( n362260 , n42114 );
nand ( n362261 , n362247 , n362260 );
buf ( n362262 , n362261 );
buf ( n362263 , n362262 );
nand ( n42119 , n362246 , n362263 );
buf ( n362265 , n42119 );
buf ( n362266 , n362265 );
buf ( n362267 , n359307 );
not ( n362268 , n362267 );
buf ( n42124 , n355582 );
not ( n42125 , n42124 );
buf ( n362271 , n360357 );
not ( n42127 , n362271 );
buf ( n362273 , n42127 );
buf ( n42129 , n360876 );
buf ( n362275 , n40739 );
nand ( n42131 , n42129 , n362275 );
buf ( n42132 , n42131 );
and ( n362278 , n362273 , n42132 );
not ( n42134 , n362273 );
not ( n362280 , n42132 );
and ( n362281 , n42134 , n362280 );
nor ( n42137 , n362278 , n362281 );
buf ( n362283 , n42137 );
buf ( n362284 , n362283 );
buf ( n362285 , n362284 );
buf ( n362286 , n362285 );
not ( n362287 , n362286 );
buf ( n362288 , n362287 );
buf ( n362289 , n362288 );
not ( n42145 , n362289 );
or ( n42146 , n42125 , n42145 );
buf ( n42147 , n362285 );
buf ( n42148 , n42147 );
buf ( n42149 , n42148 );
buf ( n42150 , n42149 );
buf ( n362296 , n40945 );
nand ( n362297 , n42150 , n362296 );
buf ( n362298 , n362297 );
buf ( n362299 , n362298 );
nand ( n362300 , n42146 , n362299 );
buf ( n362301 , n362300 );
buf ( n362302 , n362301 );
not ( n362303 , n362302 );
or ( n42159 , n362268 , n362303 );
buf ( n362305 , n361857 );
buf ( n362306 , n39217 );
nand ( n362307 , n362305 , n362306 );
buf ( n362308 , n362307 );
buf ( n362309 , n362308 );
nand ( n362310 , n42159 , n362309 );
buf ( n362311 , n362310 );
buf ( n362312 , n362311 );
xor ( n362313 , n362266 , n362312 );
buf ( n362314 , n361022 );
not ( n362315 , n362314 );
not ( n42171 , n361026 );
buf ( n362317 , n42171 );
not ( n362318 , n362317 );
buf ( n362319 , n360401 );
not ( n362320 , n362319 );
or ( n362321 , n362318 , n362320 );
buf ( n362322 , n40275 );
buf ( n362323 , n361026 );
nand ( n362324 , n362322 , n362323 );
buf ( n362325 , n362324 );
buf ( n362326 , n362325 );
nand ( n362327 , n362321 , n362326 );
buf ( n362328 , n362327 );
buf ( n362329 , n362328 );
not ( n362330 , n362329 );
or ( n362331 , n362315 , n362330 );
buf ( n362332 , n40893 );
not ( n362333 , n362332 );
buf ( n362334 , n40202 );
not ( n42190 , n362334 );
or ( n362336 , n362333 , n42190 );
buf ( n362337 , n360930 );
buf ( n362338 , n361026 );
nand ( n362339 , n362337 , n362338 );
buf ( n362340 , n362339 );
buf ( n362341 , n362340 );
nand ( n362342 , n362336 , n362341 );
buf ( n362343 , n362342 );
buf ( n362344 , n362343 );
buf ( n362345 , n361060 );
nand ( n42201 , n362344 , n362345 );
buf ( n42202 , n42201 );
buf ( n362348 , n42202 );
nand ( n42204 , n362331 , n362348 );
buf ( n42205 , n42204 );
buf ( n362351 , n42205 );
and ( n42207 , n362313 , n362351 );
and ( n362353 , n362266 , n362312 );
or ( n42209 , n42207 , n362353 );
buf ( n362355 , n42209 );
buf ( n362356 , n362355 );
and ( n362357 , n42084 , n362356 );
and ( n42213 , n362200 , n362228 );
or ( n42214 , n362357 , n42213 );
buf ( n362360 , n42214 );
buf ( n362361 , n362360 );
not ( n42217 , n362361 );
buf ( n362363 , n42217 );
buf ( n362364 , n362363 );
not ( n362365 , n362364 );
or ( n42221 , n42029 , n362365 );
buf ( n362367 , n362169 );
buf ( n362368 , n362360 );
nand ( n42224 , n362367 , n362368 );
buf ( n362370 , n42224 );
buf ( n362371 , n362370 );
nand ( n42227 , n42221 , n362371 );
buf ( n42228 , n42227 );
xor ( n42229 , n361910 , n42228 );
buf ( n42230 , n42229 );
buf ( n362376 , n342714 );
not ( n362377 , n362376 );
not ( n42233 , n362377 );
not ( n362379 , n42233 );
not ( n362380 , n342018 );
not ( n362381 , n362380 );
or ( n42237 , n362379 , n362381 );
nand ( n362383 , n362377 , n342018 );
nand ( n42239 , n42237 , n362383 );
buf ( n362385 , n42239 );
not ( n362386 , n362385 );
buf ( n42242 , n362386 );
not ( n362388 , n42242 );
buf ( n362389 , n362388 );
not ( n42245 , n362389 );
not ( n362391 , n362383 );
nand ( n362392 , n362380 , n42233 );
not ( n42248 , n362392 );
or ( n362394 , n362391 , n42248 );
not ( n362395 , n336227 );
not ( n42251 , n342014 );
or ( n362397 , n362395 , n42251 );
nand ( n362398 , n342013 , n336228 );
nand ( n42254 , n362397 , n362398 );
and ( n362400 , n42254 , n342334 );
not ( n42256 , n42254 );
and ( n362402 , n42256 , n361953 );
nor ( n362403 , n362400 , n362402 );
nand ( n42259 , n362394 , n362403 );
not ( n362405 , n42259 );
buf ( n42261 , n362405 );
buf ( n42262 , n42261 );
buf ( n42263 , n42262 );
buf ( n42264 , n42263 );
not ( n42265 , n42264 );
buf ( n42266 , n42265 );
buf ( n362412 , n42266 );
not ( n42268 , n362412 );
or ( n362414 , n42245 , n42268 );
buf ( n362415 , n342334 );
not ( n362416 , n362415 );
buf ( n362417 , n362416 );
buf ( n362418 , n362417 );
not ( n42274 , n362418 );
buf ( n362420 , n42274 );
buf ( n362421 , n362420 );
not ( n362422 , n362421 );
buf ( n362423 , n362422 );
buf ( n362424 , n362423 );
buf ( n362425 , n362424 );
buf ( n362426 , n362425 );
buf ( n362427 , n362426 );
not ( n42283 , n362427 );
buf ( n362429 , n359147 );
not ( n362430 , n362429 );
or ( n42286 , n42283 , n362430 );
buf ( n362432 , n360624 );
buf ( n362433 , n362426 );
not ( n42289 , n362433 );
buf ( n362435 , n42289 );
buf ( n362436 , n362435 );
buf ( n42292 , n362436 );
buf ( n362438 , n42292 );
buf ( n362439 , n362438 );
nand ( n42295 , n362432 , n362439 );
buf ( n362441 , n42295 );
buf ( n362442 , n362441 );
nand ( n42298 , n42286 , n362442 );
buf ( n42299 , n42298 );
buf ( n42300 , n42299 );
nand ( n42301 , n362414 , n42300 );
buf ( n42302 , n42301 );
buf ( n42303 , n42302 );
not ( n362449 , n360601 );
buf ( n362450 , n359283 );
buf ( n362451 , n362450 );
buf ( n362452 , n362451 );
buf ( n362453 , n362452 );
not ( n362454 , n362453 );
not ( n362455 , n40713 );
buf ( n362456 , n362455 );
buf ( n362457 , n362456 );
buf ( n362458 , n362457 );
buf ( n362459 , n362458 );
not ( n362460 , n362459 );
buf ( n362461 , n362460 );
buf ( n362462 , n362461 );
not ( n362463 , n362462 );
or ( n362464 , n362454 , n362463 );
buf ( n362465 , n362461 );
not ( n362466 , n362465 );
buf ( n362467 , n362466 );
buf ( n362468 , n362467 );
buf ( n362469 , n362452 );
not ( n42325 , n362469 );
buf ( n362471 , n42325 );
buf ( n362472 , n362471 );
nand ( n42328 , n362468 , n362472 );
buf ( n362474 , n42328 );
buf ( n362475 , n362474 );
nand ( n42331 , n362464 , n362475 );
buf ( n362477 , n42331 );
not ( n42333 , n362477 );
or ( n362479 , n362449 , n42333 );
buf ( n362480 , n360616 );
not ( n362481 , n362480 );
buf ( n362482 , n40252 );
not ( n42338 , n362482 );
or ( n362484 , n362481 , n42338 );
buf ( n362485 , n40251 );
buf ( n362486 , n362485 );
buf ( n362487 , n360616 );
not ( n42343 , n362487 );
buf ( n362489 , n42343 );
buf ( n362490 , n362489 );
nand ( n362491 , n362486 , n362490 );
buf ( n362492 , n362491 );
buf ( n362493 , n362492 );
nand ( n362494 , n362484 , n362493 );
buf ( n362495 , n362494 );
nand ( n362496 , n362495 , n360577 );
nand ( n42352 , n362479 , n362496 );
buf ( n362498 , n42352 );
xor ( n362499 , n42303 , n362498 );
buf ( n42355 , n32084 );
buf ( n362501 , n42355 );
not ( n362502 , n362501 );
buf ( n362503 , n361631 );
not ( n42359 , n362503 );
or ( n42360 , n362502 , n42359 );
buf ( n362506 , n352119 );
buf ( n362507 , n39621 );
nand ( n42363 , n362506 , n362507 );
buf ( n362509 , n42363 );
buf ( n362510 , n362509 );
nand ( n42366 , n42360 , n362510 );
buf ( n362512 , n42366 );
buf ( n362513 , n362512 );
not ( n362514 , n362513 );
buf ( n362515 , n359809 );
not ( n362516 , n362515 );
or ( n42372 , n362514 , n362516 );
not ( n42373 , n359685 );
buf ( n362519 , n42373 );
not ( n42375 , n362519 );
buf ( n362521 , n42375 );
buf ( n362522 , n362521 );
not ( n362523 , n352110 );
not ( n362524 , n31757 );
or ( n42380 , n362523 , n362524 );
buf ( n362526 , n32075 );
nand ( n362527 , n42380 , n362526 );
nand ( n42383 , n359019 , n357249 );
not ( n362529 , n42383 );
and ( n362530 , n362527 , n362529 );
not ( n42386 , n362527 );
and ( n42387 , n42386 , n42383 );
nor ( n42388 , n362530 , n42387 );
buf ( n362534 , n42388 );
buf ( n362535 , n362534 );
not ( n42391 , n362535 );
buf ( n362537 , n42391 );
buf ( n362538 , n362537 );
not ( n362539 , n362538 );
buf ( n362540 , n362539 );
buf ( n362541 , n362540 );
not ( n42397 , n362541 );
buf ( n362543 , n361631 );
not ( n362544 , n362543 );
or ( n42400 , n42397 , n362544 );
buf ( n42401 , n39621 );
buf ( n362547 , n362534 );
buf ( n362548 , n362547 );
buf ( n362549 , n362548 );
buf ( n362550 , n362549 );
not ( n42406 , n362550 );
buf ( n362552 , n42406 );
buf ( n362553 , n362552 );
nand ( n362554 , n42401 , n362553 );
buf ( n362555 , n362554 );
buf ( n362556 , n362555 );
nand ( n362557 , n42400 , n362556 );
buf ( n362558 , n362557 );
buf ( n362559 , n362558 );
nand ( n362560 , n362522 , n362559 );
buf ( n362561 , n362560 );
buf ( n362562 , n362561 );
nand ( n362563 , n42372 , n362562 );
buf ( n362564 , n362563 );
buf ( n362565 , n362564 );
not ( n42421 , n362565 );
buf ( n362567 , n42421 );
buf ( n42423 , n362567 );
buf ( n362569 , n40059 );
not ( n362570 , n362569 );
buf ( n362571 , n39966 );
not ( n42427 , n362571 );
buf ( n362573 , n41615 );
not ( n362574 , n362573 );
or ( n42430 , n42427 , n362574 );
not ( n42431 , n361751 );
nand ( n362577 , n42431 , n39963 );
buf ( n362578 , n362577 );
nand ( n362579 , n42430 , n362578 );
buf ( n362580 , n362579 );
buf ( n362581 , n362580 );
not ( n362582 , n362581 );
or ( n362583 , n362570 , n362582 );
buf ( n362584 , n42114 );
buf ( n362585 , n39949 );
nand ( n362586 , n362584 , n362585 );
buf ( n362587 , n362586 );
buf ( n362588 , n362587 );
nand ( n42444 , n362583 , n362588 );
buf ( n42445 , n42444 );
buf ( n362591 , n42445 );
xor ( n362592 , n42423 , n362591 );
not ( n42448 , n361717 );
buf ( n362594 , n42448 );
buf ( n362595 , n361762 );
and ( n362596 , n362594 , n362595 );
buf ( n362597 , n361717 );
buf ( n42453 , n359904 );
buf ( n42454 , n42453 );
buf ( n42455 , n42454 );
buf ( n362601 , n42455 );
and ( n42457 , n362597 , n362601 );
nor ( n362603 , n362596 , n42457 );
buf ( n362604 , n362603 );
buf ( n362605 , n362604 );
not ( n362606 , n362605 );
buf ( n362607 , n362606 );
buf ( n362608 , n362607 );
not ( n42464 , n362608 );
buf ( n362610 , n359919 );
not ( n362611 , n362610 );
or ( n42467 , n42464 , n362611 );
buf ( n362613 , n39891 );
buf ( n362614 , n359950 );
not ( n42470 , n362614 );
buf ( n362616 , n361679 );
not ( n362617 , n362616 );
or ( n42473 , n42470 , n362617 );
buf ( n362619 , n361673 );
buf ( n362620 , n41623 );
nand ( n42476 , n362619 , n362620 );
buf ( n42477 , n42476 );
buf ( n362623 , n42477 );
nand ( n42479 , n42473 , n362623 );
buf ( n362625 , n42479 );
buf ( n362626 , n362625 );
nand ( n42482 , n362613 , n362626 );
buf ( n362628 , n42482 );
buf ( n362629 , n362628 );
nand ( n362630 , n42467 , n362629 );
buf ( n362631 , n362630 );
buf ( n362632 , n362631 );
and ( n42488 , n362592 , n362632 );
and ( n42489 , n42423 , n362591 );
or ( n362635 , n42488 , n42489 );
buf ( n362636 , n362635 );
buf ( n362637 , n362636 );
and ( n362638 , n362499 , n362637 );
and ( n362639 , n42303 , n362498 );
or ( n42495 , n362638 , n362639 );
buf ( n362641 , n42495 );
buf ( n362642 , n362641 );
not ( n42498 , n362243 );
not ( n362644 , n40059 );
or ( n362645 , n42498 , n362644 );
buf ( n362646 , n39966 );
not ( n362647 , n362646 );
buf ( n362648 , n362288 );
not ( n362649 , n362648 );
or ( n362650 , n362647 , n362649 );
buf ( n362651 , n42149 );
buf ( n362652 , n39963 );
nand ( n42508 , n362651 , n362652 );
buf ( n362654 , n42508 );
buf ( n362655 , n362654 );
nand ( n362656 , n362650 , n362655 );
buf ( n362657 , n362656 );
buf ( n362658 , n362657 );
not ( n362659 , n362658 );
buf ( n362660 , n362659 );
buf ( n362661 , n39952 );
not ( n362662 , n362661 );
buf ( n362663 , n362662 );
or ( n362664 , n362660 , n362663 );
nand ( n42520 , n362645 , n362664 );
buf ( n362666 , n42520 );
buf ( n362667 , n360601 );
not ( n42523 , n362667 );
buf ( n362669 , n362495 );
not ( n362670 , n362669 );
or ( n42526 , n42523 , n362670 );
buf ( n362672 , n360616 );
not ( n362673 , n362672 );
buf ( n362674 , n360401 );
not ( n362675 , n362674 );
or ( n362676 , n362673 , n362675 );
buf ( n362677 , n362489 );
buf ( n362678 , n40275 );
nand ( n362679 , n362677 , n362678 );
buf ( n362680 , n362679 );
buf ( n362681 , n362680 );
nand ( n362682 , n362676 , n362681 );
buf ( n362683 , n362682 );
buf ( n362684 , n362683 );
buf ( n362685 , n360577 );
nand ( n362686 , n362684 , n362685 );
buf ( n362687 , n362686 );
buf ( n362688 , n362687 );
nand ( n362689 , n42526 , n362688 );
buf ( n362690 , n362689 );
buf ( n362691 , n362690 );
xor ( n362692 , n362666 , n362691 );
buf ( n362693 , n361060 );
not ( n362694 , n362693 );
buf ( n362695 , n361901 );
not ( n42551 , n362695 );
or ( n42552 , n362694 , n42551 );
buf ( n362698 , n362343 );
buf ( n362699 , n361022 );
nand ( n362700 , n362698 , n362699 );
buf ( n362701 , n362700 );
buf ( n362702 , n362701 );
nand ( n42558 , n42552 , n362702 );
buf ( n362704 , n42558 );
buf ( n362705 , n362704 );
xor ( n42561 , n362692 , n362705 );
buf ( n362707 , n42561 );
buf ( n362708 , n362707 );
xor ( n42564 , n362642 , n362708 );
buf ( n362710 , n362564 );
buf ( n362711 , n362558 );
not ( n362712 , n362711 );
buf ( n362713 , n359809 );
not ( n362714 , n362713 );
or ( n42570 , n362712 , n362714 );
buf ( n42571 , n41582 );
buf ( n362717 , n39592 );
nand ( n362718 , n42571 , n362717 );
buf ( n362719 , n362718 );
buf ( n362720 , n362719 );
nand ( n42576 , n42570 , n362720 );
buf ( n362722 , n42576 );
buf ( n362723 , n362722 );
xor ( n362724 , n362710 , n362723 );
buf ( n362725 , n362625 );
not ( n362726 , n362725 );
buf ( n362727 , n359919 );
not ( n42583 , n362727 );
or ( n362729 , n362726 , n42583 );
buf ( n362730 , n41629 );
buf ( n362731 , n39891 );
nand ( n362732 , n362730 , n362731 );
buf ( n362733 , n362732 );
buf ( n362734 , n362733 );
nand ( n42590 , n362729 , n362734 );
buf ( n362736 , n42590 );
buf ( n362737 , n362736 );
and ( n42593 , n362724 , n362737 );
and ( n42594 , n362710 , n362723 );
or ( n42595 , n42593 , n42594 );
buf ( n362741 , n42595 );
buf ( n362742 , n362741 );
buf ( n362743 , n41485 );
not ( n42599 , n362743 );
buf ( n362745 , n361555 );
not ( n362746 , n362745 );
or ( n362747 , n42599 , n362746 );
not ( n42603 , n361537 );
not ( n362749 , n359977 );
or ( n362750 , n42603 , n362749 );
not ( n42606 , n41907 );
not ( n362752 , n42606 );
nand ( n362753 , n362752 , n361540 );
nand ( n362754 , n362750 , n362753 );
buf ( n362755 , n362754 );
buf ( n362756 , n361609 );
nand ( n42612 , n362755 , n362756 );
buf ( n42613 , n42612 );
buf ( n362759 , n42613 );
nand ( n42615 , n362747 , n362759 );
buf ( n42616 , n42615 );
buf ( n362762 , n42616 );
xor ( n362763 , n362742 , n362762 );
xor ( n42619 , n361728 , n361826 );
xor ( n362765 , n42619 , n361865 );
buf ( n362766 , n362765 );
buf ( n362767 , n362766 );
xor ( n362768 , n362763 , n362767 );
buf ( n362769 , n362768 );
buf ( n362770 , n362769 );
and ( n362771 , n42564 , n362770 );
and ( n42627 , n362642 , n362708 );
or ( n362773 , n362771 , n42627 );
buf ( n362774 , n362773 );
buf ( n362775 , n362774 );
buf ( n362776 , n40059 );
not ( n362777 , n362776 );
buf ( n362778 , n362657 );
not ( n362779 , n362778 );
or ( n362780 , n362777 , n362779 );
buf ( n362781 , n39966 );
not ( n362782 , n362781 );
buf ( n362783 , n40756 );
not ( n42639 , n362783 );
or ( n42640 , n362782 , n42639 );
buf ( n362786 , n360893 );
buf ( n362787 , n39963 );
nand ( n362788 , n362786 , n362787 );
buf ( n362789 , n362788 );
buf ( n362790 , n362789 );
nand ( n42646 , n42640 , n362790 );
buf ( n362792 , n42646 );
buf ( n362793 , n362792 );
buf ( n362794 , n39952 );
nand ( n42650 , n362793 , n362794 );
buf ( n362796 , n42650 );
buf ( n362797 , n362796 );
nand ( n42653 , n362780 , n362797 );
buf ( n362799 , n42653 );
buf ( n42655 , n362799 );
buf ( n362801 , n39217 );
not ( n42657 , n362801 );
not ( n362803 , n40251 );
not ( n42659 , n362803 );
buf ( n42660 , n361851 );
and ( n42661 , n42659 , n42660 );
not ( n42662 , n42659 );
and ( n42663 , n42662 , n355582 );
or ( n42664 , n42661 , n42663 );
buf ( n362810 , n42664 );
not ( n362811 , n362810 );
or ( n42667 , n42657 , n362811 );
buf ( n362813 , n361841 );
buf ( n362814 , n359307 );
nand ( n42670 , n362813 , n362814 );
buf ( n362816 , n42670 );
buf ( n362817 , n362816 );
nand ( n362818 , n42667 , n362817 );
buf ( n362819 , n362818 );
buf ( n362820 , n362819 );
xor ( n42676 , n42655 , n362820 );
buf ( n362822 , n360601 );
not ( n362823 , n362822 );
buf ( n362824 , n362683 );
not ( n362825 , n362824 );
or ( n42681 , n362823 , n362825 );
buf ( n362827 , n360616 );
not ( n362828 , n362827 );
not ( n42684 , n360930 );
buf ( n362830 , n42684 );
not ( n362831 , n362830 );
or ( n42687 , n362828 , n362831 );
buf ( n362833 , n40201 );
buf ( n362834 , n362489 );
nand ( n42690 , n362833 , n362834 );
buf ( n362836 , n42690 );
buf ( n362837 , n362836 );
nand ( n42693 , n42687 , n362837 );
buf ( n362839 , n42693 );
buf ( n362840 , n362839 );
buf ( n362841 , n360577 );
nand ( n362842 , n362840 , n362841 );
buf ( n362843 , n362842 );
buf ( n362844 , n362843 );
nand ( n362845 , n42681 , n362844 );
buf ( n362846 , n362845 );
buf ( n362847 , n362846 );
xor ( n362848 , n42676 , n362847 );
buf ( n362849 , n362848 );
buf ( n362850 , n362849 );
xor ( n42706 , n362666 , n362691 );
and ( n42707 , n42706 , n362705 );
and ( n42708 , n362666 , n362691 );
or ( n42709 , n42707 , n42708 );
buf ( n362855 , n42709 );
buf ( n362856 , n362855 );
xor ( n42712 , n362850 , n362856 );
buf ( n362858 , n42712 );
buf ( n362859 , n362858 );
xor ( n362860 , n362742 , n362762 );
and ( n362861 , n362860 , n362767 );
and ( n42717 , n362742 , n362762 );
or ( n362863 , n362861 , n42717 );
buf ( n362864 , n362863 );
buf ( n362865 , n362864 );
xor ( n42721 , n362859 , n362865 );
buf ( n362867 , n42721 );
buf ( n362868 , n362867 );
xor ( n362869 , n362775 , n362868 );
xor ( n42725 , n362710 , n362723 );
xor ( n362871 , n42725 , n362737 );
buf ( n362872 , n362871 );
buf ( n362873 , n362872 );
buf ( n362874 , n362066 );
not ( n42730 , n362874 );
buf ( n362876 , n42075 );
not ( n362877 , n362876 );
or ( n42733 , n42730 , n362877 );
buf ( n362879 , n41892 );
not ( n42735 , n362879 );
buf ( n362881 , n359784 );
not ( n362882 , n362881 );
or ( n42738 , n42735 , n362882 );
buf ( n362884 , n359781 );
buf ( n362885 , n362037 );
nand ( n362886 , n362884 , n362885 );
buf ( n362887 , n362886 );
buf ( n362888 , n362887 );
nand ( n42744 , n42738 , n362888 );
buf ( n362890 , n42744 );
buf ( n362891 , n362890 );
buf ( n362892 , n362030 );
nand ( n362893 , n362891 , n362892 );
buf ( n362894 , n362893 );
buf ( n362895 , n362894 );
nand ( n362896 , n42733 , n362895 );
buf ( n362897 , n362896 );
buf ( n362898 , n362897 );
xor ( n362899 , n362873 , n362898 );
buf ( n362900 , n361609 );
not ( n362901 , n362900 );
buf ( n362902 , n361540 );
buf ( n362903 , n39832 );
and ( n42759 , n362902 , n362903 );
not ( n42760 , n362902 );
buf ( n362906 , n361073 );
and ( n42762 , n42760 , n362906 );
nor ( n362908 , n42759 , n42762 );
buf ( n362909 , n362908 );
buf ( n362910 , n362909 );
not ( n362911 , n362910 );
or ( n362912 , n362901 , n362911 );
buf ( n362913 , n362754 );
buf ( n362914 , n41485 );
nand ( n362915 , n362913 , n362914 );
buf ( n362916 , n362915 );
buf ( n362917 , n362916 );
nand ( n362918 , n362912 , n362917 );
buf ( n362919 , n362918 );
buf ( n362920 , n362919 );
and ( n362921 , n362899 , n362920 );
and ( n362922 , n362873 , n362898 );
or ( n42778 , n362921 , n362922 );
buf ( n362924 , n42778 );
buf ( n362925 , n362924 );
buf ( n362926 , n41835 );
not ( n42782 , n362926 );
buf ( n362928 , n362189 );
not ( n362929 , n362928 );
or ( n42785 , n42782 , n362929 );
buf ( n362931 , n41778 );
buf ( n362932 , n41406 );
and ( n362933 , n362931 , n362932 );
not ( n42789 , n362931 );
buf ( n362935 , n360116 );
and ( n362936 , n42789 , n362935 );
nor ( n42792 , n362933 , n362936 );
buf ( n362938 , n42792 );
buf ( n362939 , n362938 );
buf ( n362940 , n41830 );
nand ( n362941 , n362939 , n362940 );
buf ( n362942 , n362941 );
buf ( n362943 , n362942 );
nand ( n362944 , n42785 , n362943 );
buf ( n362945 , n362944 );
buf ( n362946 , n362945 );
buf ( n362947 , n360577 );
not ( n362948 , n362947 );
buf ( n362949 , n362477 );
not ( n362950 , n362949 );
or ( n362951 , n362948 , n362950 );
buf ( n362952 , n360893 );
buf ( n362953 , n362471 );
nand ( n362954 , n362952 , n362953 );
buf ( n362955 , n362954 );
nand ( n42811 , n362452 , n360886 );
nand ( n362957 , n362955 , n42811 );
buf ( n42813 , n362957 );
buf ( n362959 , n360601 );
nand ( n42815 , n42813 , n362959 );
buf ( n362961 , n42815 );
buf ( n362962 , n362961 );
nand ( n42818 , n362951 , n362962 );
buf ( n362964 , n42818 );
buf ( n362965 , n362964 );
not ( n42821 , n362965 );
buf ( n362967 , n42171 );
buf ( n362968 , n40251 );
xor ( n42824 , n362967 , n362968 );
buf ( n42825 , n42824 );
buf ( n362971 , n42825 );
not ( n42827 , n362971 );
buf ( n362973 , n42827 );
buf ( n362974 , n362973 );
not ( n42830 , n362974 );
buf ( n362976 , n361121 );
not ( n362977 , n362976 );
and ( n42833 , n42830 , n362977 );
buf ( n362979 , n362328 );
buf ( n362980 , n361060 );
and ( n42836 , n362979 , n362980 );
nor ( n362982 , n42833 , n42836 );
buf ( n362983 , n362982 );
buf ( n362984 , n362983 );
not ( n362985 , n362984 );
buf ( n362986 , n362985 );
buf ( n362987 , n362986 );
not ( n42843 , n362987 );
or ( n362989 , n42821 , n42843 );
buf ( n42845 , n362964 );
not ( n42846 , n42845 );
buf ( n42847 , n42846 );
not ( n42848 , n42847 );
not ( n42849 , n362983 );
or ( n42850 , n42848 , n42849 );
not ( n42851 , n362301 );
not ( n362997 , n39217 );
or ( n362998 , n42851 , n362997 );
and ( n362999 , n355582 , n362145 );
not ( n363000 , n355582 );
and ( n363001 , n363000 , n362148 );
or ( n363002 , n362999 , n363001 );
buf ( n42852 , n363002 );
buf ( n363004 , n359307 );
nand ( n363005 , n42852 , n363004 );
buf ( n363006 , n363005 );
nand ( n42856 , n362998 , n363006 );
nand ( n363008 , n42850 , n42856 );
buf ( n363009 , n363008 );
nand ( n363010 , n362989 , n363009 );
buf ( n363011 , n363010 );
buf ( n363012 , n363011 );
xor ( n363013 , n362946 , n363012 );
xor ( n363014 , n362266 , n362312 );
xor ( n42864 , n363014 , n362351 );
buf ( n363016 , n42864 );
buf ( n363017 , n363016 );
and ( n42867 , n363013 , n363017 );
and ( n363019 , n362946 , n363012 );
or ( n42869 , n42867 , n363019 );
buf ( n363021 , n42869 );
buf ( n363022 , n363021 );
xor ( n363023 , n362925 , n363022 );
xor ( n42873 , n362200 , n362228 );
xor ( n363025 , n42873 , n362356 );
buf ( n363026 , n363025 );
buf ( n363027 , n363026 );
and ( n363028 , n363023 , n363027 );
and ( n42878 , n362925 , n363022 );
or ( n363030 , n363028 , n42878 );
buf ( n363031 , n363030 );
buf ( n363032 , n363031 );
xor ( n363033 , n362869 , n363032 );
buf ( n363034 , n363033 );
buf ( n363035 , n363034 );
xor ( n363036 , n42230 , n363035 );
buf ( n42886 , n39700 );
not ( n363038 , n42886 );
buf ( n363039 , n363038 );
not ( n42889 , n363039 );
not ( n363041 , n30911 );
not ( n42891 , n363041 );
buf ( n363043 , n42891 );
not ( n42893 , n363043 );
buf ( n42894 , n361631 );
not ( n42895 , n42894 );
or ( n42896 , n42893 , n42895 );
buf ( n363048 , n39621 );
not ( n42898 , n42891 );
buf ( n363050 , n42898 );
nand ( n363051 , n363048 , n363050 );
buf ( n363052 , n363051 );
buf ( n363053 , n363052 );
nand ( n42903 , n42896 , n363053 );
buf ( n363055 , n42903 );
buf ( n363056 , n363055 );
not ( n42906 , n363056 );
or ( n363058 , n42889 , n42906 );
buf ( n42908 , n362521 );
buf ( n363060 , n351762 );
buf ( n42910 , n363060 );
buf ( n42911 , n42910 );
buf ( n363063 , n42911 );
not ( n42913 , n363063 );
buf ( n363065 , n361631 );
not ( n363066 , n363065 );
or ( n42916 , n42913 , n363066 );
buf ( n363068 , n39621 );
buf ( n363069 , n42911 );
not ( n363070 , n363069 );
buf ( n363071 , n363070 );
buf ( n363072 , n363071 );
nand ( n363073 , n363068 , n363072 );
buf ( n363074 , n363073 );
buf ( n363075 , n363074 );
nand ( n42925 , n42916 , n363075 );
buf ( n42926 , n42925 );
buf ( n363078 , n42926 );
nand ( n42928 , n42908 , n363078 );
buf ( n42929 , n42928 );
buf ( n363081 , n42929 );
nand ( n363082 , n363058 , n363081 );
buf ( n363083 , n363082 );
buf ( n363084 , n363083 );
buf ( n42934 , n42926 );
not ( n42935 , n42934 );
buf ( n42936 , n359809 );
not ( n42937 , n42936 );
or ( n42938 , n42935 , n42937 );
buf ( n42939 , n39592 );
buf ( n363091 , n362512 );
nand ( n363092 , n42939 , n363091 );
buf ( n363093 , n363092 );
buf ( n363094 , n363093 );
nand ( n42944 , n42938 , n363094 );
buf ( n42945 , n42944 );
buf ( n363097 , n42945 );
xor ( n42947 , n363084 , n363097 );
buf ( n363099 , n39949 );
not ( n363100 , n363099 );
buf ( n363101 , n362580 );
not ( n42951 , n363101 );
or ( n363103 , n363100 , n42951 );
buf ( n363104 , n40059 );
buf ( n363105 , n39963 );
not ( n363106 , n363105 );
buf ( n363107 , n363106 );
buf ( n363108 , n363107 );
not ( n42958 , n363108 );
buf ( n363110 , n361679 );
not ( n363111 , n363110 );
or ( n363112 , n42958 , n363111 );
buf ( n363113 , n361673 );
buf ( n363114 , n359879 );
not ( n363115 , n363114 );
buf ( n363116 , n363115 );
buf ( n363117 , n363116 );
not ( n363118 , n363117 );
buf ( n363119 , n363118 );
buf ( n363120 , n363119 );
not ( n42970 , n363120 );
buf ( n363122 , n42970 );
buf ( n363123 , n363122 );
nand ( n363124 , n363113 , n363123 );
buf ( n363125 , n363124 );
buf ( n363126 , n363125 );
nand ( n42976 , n363112 , n363126 );
buf ( n363128 , n42976 );
buf ( n42978 , n363128 );
nand ( n42979 , n363104 , n42978 );
buf ( n42980 , n42979 );
buf ( n42981 , n42980 );
nand ( n42982 , n363103 , n42981 );
buf ( n42983 , n42982 );
buf ( n363135 , n42983 );
and ( n42985 , n42947 , n363135 );
and ( n42986 , n363084 , n363097 );
or ( n363138 , n42985 , n42986 );
buf ( n363139 , n363138 );
buf ( n42989 , n363139 );
buf ( n363141 , n362066 );
not ( n363142 , n363141 );
buf ( n42992 , n362890 );
not ( n42993 , n42992 );
or ( n42994 , n363142 , n42993 );
buf ( n363146 , n41892 );
not ( n363147 , n363146 );
buf ( n363148 , n360308 );
not ( n363149 , n363148 );
or ( n363150 , n363147 , n363149 );
buf ( n363151 , n360930 );
buf ( n363152 , n362037 );
nand ( n363153 , n363151 , n363152 );
buf ( n363154 , n363153 );
buf ( n363155 , n363154 );
nand ( n363156 , n363150 , n363155 );
buf ( n363157 , n363156 );
buf ( n363158 , n363157 );
buf ( n363159 , n362030 );
nand ( n363160 , n363158 , n363159 );
buf ( n363161 , n363160 );
buf ( n363162 , n363161 );
nand ( n363163 , n42994 , n363162 );
buf ( n363164 , n363163 );
buf ( n363165 , n363164 );
xor ( n43015 , n42989 , n363165 );
buf ( n363167 , n41830 );
not ( n363168 , n363167 );
buf ( n363169 , n41778 );
not ( n43019 , n363169 );
buf ( n363171 , n359974 );
not ( n363172 , n363171 );
buf ( n363173 , n363172 );
not ( n363174 , n363173 );
or ( n363175 , n43019 , n363174 );
buf ( n363176 , n42606 );
buf ( n363177 , n361917 );
nand ( n363178 , n363176 , n363177 );
buf ( n363179 , n363178 );
buf ( n363180 , n363179 );
nand ( n43030 , n363175 , n363180 );
buf ( n43031 , n43030 );
buf ( n43032 , n43031 );
not ( n43033 , n43032 );
or ( n43034 , n363168 , n43033 );
buf ( n43035 , n362938 );
buf ( n43036 , n41835 );
nand ( n43037 , n43035 , n43036 );
buf ( n43038 , n43037 );
buf ( n43039 , n43038 );
nand ( n43040 , n43034 , n43039 );
buf ( n43041 , n43040 );
buf ( n363193 , n43041 );
and ( n363194 , n43015 , n363193 );
and ( n43044 , n42989 , n363165 );
or ( n363196 , n363194 , n43044 );
buf ( n363197 , n363196 );
buf ( n363198 , n363197 );
xor ( n363199 , n42303 , n362498 );
xor ( n363200 , n363199 , n362637 );
buf ( n363201 , n363200 );
buf ( n363202 , n363201 );
xor ( n363203 , n363198 , n363202 );
xor ( n363204 , n42423 , n362591 );
xor ( n363205 , n363204 , n362632 );
buf ( n363206 , n363205 );
buf ( n43051 , n363206 );
buf ( n363208 , n42266 );
not ( n363209 , n363208 );
buf ( n363210 , n363209 );
buf ( n363211 , n363210 );
not ( n43056 , n363211 );
not ( n363213 , n362438 );
not ( n43058 , n361617 );
or ( n363215 , n363213 , n43058 );
buf ( n363216 , n362438 );
not ( n43061 , n363216 );
buf ( n363218 , n43061 );
nand ( n43063 , n40091 , n363218 );
nand ( n43064 , n363215 , n43063 );
buf ( n363221 , n43064 );
not ( n43066 , n363221 );
or ( n363223 , n43056 , n43066 );
buf ( n363224 , n42299 );
buf ( n363225 , n42242 );
nand ( n363226 , n363224 , n363225 );
buf ( n363227 , n363226 );
buf ( n363228 , n363227 );
nand ( n363229 , n363223 , n363228 );
buf ( n363230 , n363229 );
buf ( n363231 , n363230 );
xor ( n363232 , n43051 , n363231 );
buf ( n363233 , n41485 );
not ( n363234 , n363233 );
buf ( n363235 , n362909 );
not ( n363236 , n363235 );
or ( n43081 , n363234 , n363236 );
buf ( n363238 , n361540 );
not ( n43083 , n363238 );
buf ( n363240 , n362208 );
not ( n43085 , n363240 );
or ( n43086 , n43083 , n43085 );
buf ( n363243 , n42068 );
buf ( n363244 , n361537 );
nand ( n363245 , n363243 , n363244 );
buf ( n363246 , n363245 );
buf ( n363247 , n363246 );
nand ( n363248 , n43086 , n363247 );
buf ( n363249 , n363248 );
buf ( n363250 , n363249 );
buf ( n363251 , n361609 );
nand ( n363252 , n363250 , n363251 );
buf ( n363253 , n363252 );
buf ( n363254 , n363253 );
nand ( n363255 , n43081 , n363254 );
buf ( n363256 , n363255 );
buf ( n363257 , n363256 );
and ( n363258 , n363232 , n363257 );
and ( n43103 , n43051 , n363231 );
or ( n363260 , n363258 , n43103 );
buf ( n363261 , n363260 );
buf ( n363262 , n363261 );
and ( n43107 , n363203 , n363262 );
and ( n363264 , n363198 , n363202 );
or ( n363265 , n43107 , n363264 );
buf ( n363266 , n363265 );
buf ( n363267 , n363266 );
xor ( n363268 , n362642 , n362708 );
xor ( n363269 , n363268 , n362770 );
buf ( n363270 , n363269 );
buf ( n363271 , n363270 );
xor ( n363272 , n363267 , n363271 );
xor ( n43117 , n362925 , n363022 );
xor ( n43118 , n43117 , n363027 );
buf ( n363275 , n43118 );
buf ( n43120 , n363275 );
and ( n43121 , n363272 , n43120 );
and ( n43122 , n363267 , n363271 );
or ( n43123 , n43121 , n43122 );
buf ( n43124 , n43123 );
buf ( n43125 , n43124 );
xor ( n43126 , n363036 , n43125 );
buf ( n43127 , n43126 );
buf ( n363284 , n43127 );
xor ( n43129 , n362873 , n362898 );
xor ( n43130 , n43129 , n362920 );
buf ( n43131 , n43130 );
buf ( n363288 , n43131 );
buf ( n363289 , n359913 );
buf ( n43134 , n363289 );
buf ( n363291 , n43134 );
buf ( n363292 , n363291 );
buf ( n363293 , n362540 );
buf ( n363294 , n42455 );
and ( n363295 , n363293 , n363294 );
not ( n43140 , n363293 );
buf ( n363297 , n361762 );
and ( n43142 , n43140 , n363297 );
nor ( n43143 , n363295 , n43142 );
buf ( n363300 , n43143 );
buf ( n363301 , n363300 );
or ( n363302 , n363292 , n363301 );
buf ( n363303 , n359996 );
buf ( n363304 , n362604 );
or ( n363305 , n363303 , n363304 );
nand ( n43150 , n363302 , n363305 );
buf ( n363307 , n43150 );
buf ( n363308 , n363307 );
buf ( n363309 , n39217 );
not ( n363310 , n363309 );
buf ( n363311 , n363002 );
not ( n43156 , n363311 );
or ( n363313 , n363310 , n43156 );
buf ( n363314 , n359307 );
buf ( n363315 , n355582 );
not ( n363316 , n363315 );
buf ( n363317 , n41659 );
buf ( n363318 , n363317 );
not ( n43163 , n363318 );
or ( n43164 , n363316 , n43163 );
buf ( n363321 , n41663 );
buf ( n363322 , n361851 );
nand ( n43167 , n363321 , n363322 );
buf ( n43168 , n43167 );
buf ( n363325 , n43168 );
nand ( n363326 , n43164 , n363325 );
buf ( n363327 , n363326 );
buf ( n363328 , n363327 );
nand ( n363329 , n363314 , n363328 );
buf ( n363330 , n363329 );
buf ( n363331 , n363330 );
nand ( n363332 , n363313 , n363331 );
buf ( n363333 , n363332 );
buf ( n363334 , n363333 );
xor ( n43179 , n363308 , n363334 );
buf ( n363336 , n361060 );
not ( n43181 , n363336 );
buf ( n363338 , n42825 );
not ( n43183 , n363338 );
or ( n363340 , n43181 , n43183 );
and ( n363341 , n42171 , n360851 );
not ( n363342 , n42171 );
and ( n43187 , n363342 , n362467 );
or ( n363344 , n363341 , n43187 );
buf ( n363345 , n363344 );
buf ( n363346 , n361022 );
nand ( n363347 , n363345 , n363346 );
buf ( n363348 , n363347 );
buf ( n363349 , n363348 );
nand ( n43194 , n363340 , n363349 );
buf ( n363351 , n43194 );
buf ( n363352 , n363351 );
and ( n43197 , n43179 , n363352 );
and ( n363354 , n363308 , n363334 );
or ( n363355 , n43197 , n363354 );
buf ( n363356 , n363355 );
buf ( n363357 , n363356 );
buf ( n363358 , n360616 );
not ( n363359 , n363358 );
buf ( n363360 , n42149 );
not ( n363361 , n363360 );
buf ( n363362 , n363361 );
buf ( n363363 , n363362 );
not ( n43208 , n363363 );
or ( n363365 , n363359 , n43208 );
buf ( n363366 , n42149 );
buf ( n363367 , n362489 );
nand ( n363368 , n363366 , n363367 );
buf ( n363369 , n363368 );
buf ( n363370 , n363369 );
nand ( n43215 , n363365 , n363370 );
buf ( n363372 , n43215 );
buf ( n363373 , n363372 );
buf ( n363374 , n360601 );
and ( n363375 , n363373 , n363374 );
not ( n43220 , n362957 );
nor ( n363377 , n43220 , n360580 );
buf ( n363378 , n363377 );
nor ( n43223 , n363375 , n363378 );
buf ( n363380 , n43223 );
buf ( n363381 , n363380 );
not ( n43226 , n363381 );
buf ( n363383 , n363157 );
not ( n43228 , n363383 );
buf ( n363385 , n362066 );
not ( n363386 , n363385 );
or ( n43231 , n43228 , n363386 );
not ( n363388 , n360397 );
buf ( n43233 , n363388 );
not ( n363390 , n43233 );
buf ( n363391 , n363390 );
and ( n363392 , n363391 , n41892 );
not ( n363393 , n363391 );
and ( n43238 , n363393 , n362037 );
or ( n363395 , n363392 , n43238 );
buf ( n363396 , n363395 );
buf ( n363397 , n362030 );
nand ( n363398 , n363396 , n363397 );
buf ( n363399 , n363398 );
buf ( n363400 , n363399 );
nand ( n363401 , n43231 , n363400 );
buf ( n363402 , n363401 );
buf ( n363403 , n363402 );
not ( n363404 , n363403 );
buf ( n363405 , n363404 );
buf ( n363406 , n363405 );
not ( n363407 , n363406 );
or ( n43252 , n43226 , n363407 );
and ( n43253 , n342654 , n342687 );
not ( n363410 , n342654 );
not ( n363411 , n342687 );
and ( n43256 , n363410 , n363411 );
nor ( n363413 , n43253 , n43256 );
not ( n43258 , n363413 );
not ( n363415 , n43258 );
not ( n363416 , n363415 );
not ( n43261 , n363416 );
buf ( n363418 , n43261 );
not ( n363419 , n363418 );
buf ( n363420 , n363419 );
buf ( n363421 , n363420 );
not ( n363422 , n363421 );
and ( n363423 , n342715 , n342687 );
not ( n43268 , n342715 );
and ( n363425 , n43268 , n363411 );
nor ( n363426 , n363423 , n363425 );
nand ( n43271 , n363426 , n43258 );
not ( n363428 , n43271 );
buf ( n363429 , n363428 );
not ( n43274 , n363429 );
buf ( n363431 , n43274 );
not ( n363432 , n363431 );
or ( n43277 , n363422 , n363432 );
buf ( n363434 , n359147 );
buf ( n363435 , n22772 );
and ( n43280 , n363434 , n363435 );
buf ( n363437 , n359144 );
not ( n363438 , n363437 );
buf ( n363439 , n363438 );
buf ( n363440 , n363439 );
not ( n363441 , n363440 );
buf ( n363442 , n363441 );
buf ( n363443 , n363442 );
not ( n363444 , n22772 );
buf ( n363445 , n363444 );
and ( n363446 , n363443 , n363445 );
nor ( n43282 , n43280 , n363446 );
buf ( n43283 , n43282 );
buf ( n363449 , n43283 );
not ( n363450 , n363449 );
buf ( n363451 , n363450 );
buf ( n363452 , n363451 );
nand ( n363453 , n43277 , n363452 );
buf ( n363454 , n363453 );
buf ( n363455 , n363454 );
nand ( n43291 , n43252 , n363455 );
buf ( n363457 , n43291 );
buf ( n363458 , n363457 );
buf ( n363459 , n363380 );
not ( n43295 , n363459 );
buf ( n363461 , n363402 );
nand ( n363462 , n43295 , n363461 );
buf ( n363463 , n363462 );
buf ( n363464 , n363463 );
nand ( n43300 , n363458 , n363464 );
buf ( n363466 , n43300 );
buf ( n363467 , n363466 );
xor ( n363468 , n363357 , n363467 );
xor ( n43304 , n42856 , n362964 );
xor ( n43305 , n43304 , n362986 );
buf ( n363471 , n43305 );
and ( n43307 , n363468 , n363471 );
and ( n363473 , n363357 , n363467 );
or ( n363474 , n43307 , n363473 );
buf ( n363475 , n363474 );
buf ( n363476 , n363475 );
xor ( n363477 , n363288 , n363476 );
xor ( n43313 , n362946 , n363012 );
xor ( n363479 , n43313 , n363017 );
buf ( n363480 , n363479 );
buf ( n363481 , n363480 );
and ( n43317 , n363477 , n363481 );
and ( n363483 , n363288 , n363476 );
or ( n363484 , n43317 , n363483 );
buf ( n363485 , n363484 );
buf ( n363486 , n363485 );
xor ( n363487 , n42989 , n363165 );
xor ( n43323 , n363487 , n363193 );
buf ( n363489 , n43323 );
buf ( n363490 , n363489 );
not ( n43326 , n42242 );
not ( n363492 , n43064 );
or ( n43328 , n43326 , n363492 );
buf ( n363494 , n363218 );
not ( n363495 , n363494 );
buf ( n363496 , n360116 );
not ( n363497 , n363496 );
or ( n363498 , n363495 , n363497 );
buf ( n363499 , n41406 );
buf ( n363500 , n362438 );
nand ( n363501 , n363499 , n363500 );
buf ( n363502 , n363501 );
buf ( n363503 , n363502 );
nand ( n43339 , n363498 , n363503 );
buf ( n363505 , n43339 );
buf ( n43341 , n363505 );
buf ( n43342 , n363210 );
nand ( n43343 , n43341 , n43342 );
buf ( n43344 , n43343 );
nand ( n363510 , n43328 , n43344 );
buf ( n363511 , n363510 );
not ( n363512 , n41835 );
not ( n363513 , n43031 );
or ( n43349 , n363512 , n363513 );
and ( n43350 , n359939 , n361917 );
and ( n363516 , n40943 , n41778 );
nor ( n363517 , n43350 , n363516 );
nand ( n43353 , n363517 , n41830 );
nand ( n363519 , n43349 , n43353 );
buf ( n363520 , n363519 );
xor ( n43356 , n363511 , n363520 );
xor ( n363522 , n363308 , n363334 );
xor ( n363523 , n363522 , n363352 );
buf ( n363524 , n363523 );
buf ( n363525 , n363524 );
and ( n43361 , n43356 , n363525 );
and ( n363527 , n363511 , n363520 );
or ( n363528 , n43361 , n363527 );
buf ( n363529 , n363528 );
buf ( n363530 , n363529 );
xor ( n363531 , n363490 , n363530 );
xor ( n43367 , n363084 , n363097 );
xor ( n363533 , n43367 , n363135 );
buf ( n363534 , n363533 );
buf ( n363535 , n363534 );
buf ( n363536 , n363083 );
not ( n363537 , n363536 );
buf ( n363538 , n363537 );
buf ( n363539 , n363538 );
buf ( n363540 , n363107 );
not ( n363541 , n363540 );
not ( n43377 , n361716 );
buf ( n363543 , n43377 );
not ( n363544 , n363543 );
or ( n43380 , n363541 , n363544 );
not ( n363546 , n361716 );
not ( n363547 , n363546 );
buf ( n363548 , n363547 );
buf ( n363549 , n363122 );
nand ( n43385 , n363548 , n363549 );
buf ( n43386 , n43385 );
buf ( n363552 , n43386 );
nand ( n43388 , n43380 , n363552 );
buf ( n43389 , n43388 );
buf ( n363555 , n43389 );
not ( n43391 , n363555 );
buf ( n363557 , n40059 );
not ( n363558 , n363557 );
or ( n43394 , n43391 , n363558 );
buf ( n363560 , n39949 );
buf ( n363561 , n363128 );
nand ( n43397 , n363560 , n363561 );
buf ( n363563 , n43397 );
buf ( n363564 , n363563 );
nand ( n363565 , n43394 , n363564 );
buf ( n363566 , n363565 );
buf ( n363567 , n363566 );
xor ( n363568 , n363539 , n363567 );
buf ( n363569 , n363291 );
buf ( n363570 , n32087 );
not ( n43406 , n363570 );
buf ( n363572 , n41623 );
not ( n363573 , n363572 );
or ( n43409 , n43406 , n363573 );
buf ( n363575 , n352119 );
buf ( n363576 , n359950 );
nand ( n363577 , n363575 , n363576 );
buf ( n363578 , n363577 );
buf ( n363579 , n363578 );
nand ( n363580 , n43409 , n363579 );
buf ( n363581 , n363580 );
buf ( n363582 , n363581 );
not ( n363583 , n363582 );
buf ( n363584 , n363583 );
buf ( n363585 , n363584 );
or ( n363586 , n363569 , n363585 );
buf ( n363587 , n359996 );
buf ( n363588 , n363300 );
or ( n43424 , n363587 , n363588 );
nand ( n363590 , n363586 , n43424 );
buf ( n363591 , n363590 );
buf ( n363592 , n363591 );
and ( n43428 , n363568 , n363592 );
and ( n363594 , n363539 , n363567 );
or ( n43430 , n43428 , n363594 );
buf ( n363596 , n43430 );
buf ( n363597 , n363596 );
xor ( n43433 , n363535 , n363597 );
buf ( n363599 , n361609 );
not ( n363600 , n363599 );
buf ( n363601 , n361531 );
buf ( n363602 , n363601 );
buf ( n363603 , n363602 );
and ( n43439 , n363603 , n359784 );
not ( n363605 , n363603 );
and ( n43441 , n363605 , n359781 );
or ( n363607 , n43439 , n43441 );
buf ( n363608 , n363607 );
not ( n363609 , n363608 );
or ( n43445 , n363600 , n363609 );
buf ( n363611 , n363249 );
buf ( n43447 , n41485 );
nand ( n43448 , n363611 , n43447 );
buf ( n43449 , n43448 );
buf ( n43450 , n43449 );
nand ( n43451 , n43445 , n43450 );
buf ( n43452 , n43451 );
buf ( n363618 , n43452 );
and ( n363619 , n43433 , n363618 );
and ( n43455 , n363535 , n363597 );
or ( n363621 , n363619 , n43455 );
buf ( n363622 , n363621 );
buf ( n363623 , n363622 );
and ( n363624 , n363531 , n363623 );
and ( n363625 , n363490 , n363530 );
or ( n43461 , n363624 , n363625 );
buf ( n363627 , n43461 );
buf ( n43463 , n363627 );
xor ( n363629 , n363198 , n363202 );
xor ( n363630 , n363629 , n363262 );
buf ( n363631 , n363630 );
buf ( n363632 , n363631 );
xor ( n363633 , n43463 , n363632 );
xor ( n43469 , n363288 , n363476 );
xor ( n363635 , n43469 , n363481 );
buf ( n363636 , n363635 );
buf ( n363637 , n363636 );
and ( n43473 , n363633 , n363637 );
and ( n363639 , n43463 , n363632 );
or ( n363640 , n43473 , n363639 );
buf ( n363641 , n363640 );
buf ( n363642 , n363641 );
xor ( n43478 , n363486 , n363642 );
xor ( n43479 , n363267 , n363271 );
xor ( n363645 , n43479 , n43120 );
buf ( n363646 , n363645 );
buf ( n363647 , n363646 );
and ( n43483 , n43478 , n363647 );
and ( n363649 , n363486 , n363642 );
or ( n363650 , n43483 , n363649 );
buf ( n363651 , n363650 );
buf ( n363652 , n363651 );
or ( n363653 , n363284 , n363652 );
buf ( n363654 , n363653 );
xor ( n363655 , n361630 , n361870 );
and ( n43491 , n363655 , n361908 );
and ( n363657 , n361630 , n361870 );
or ( n43493 , n43491 , n363657 );
buf ( n363659 , n43493 );
buf ( n43495 , n363659 );
buf ( n363661 , n362076 );
not ( n43497 , n361982 );
buf ( n363663 , n362072 );
not ( n43499 , n363663 );
buf ( n363665 , n43499 );
not ( n363666 , n363665 );
or ( n43502 , n43497 , n363666 );
nand ( n363668 , n43502 , n362168 );
buf ( n363669 , n363668 );
nand ( n363670 , n363661 , n363669 );
buf ( n363671 , n363670 );
buf ( n363672 , n363671 );
xor ( n363673 , n43495 , n363672 );
xor ( n43509 , n362081 , n362106 );
and ( n363675 , n43509 , n362166 );
and ( n363676 , n362081 , n362106 );
or ( n43512 , n363675 , n363676 );
buf ( n363678 , n43512 );
buf ( n363679 , n363678 );
buf ( n363680 , n361540 );
not ( n363681 , n363680 );
buf ( n363682 , n359147 );
not ( n43518 , n363682 );
or ( n363684 , n363681 , n43518 );
buf ( n363685 , n360624 );
buf ( n363686 , n361537 );
nand ( n363687 , n363685 , n363686 );
buf ( n363688 , n363687 );
buf ( n363689 , n363688 );
nand ( n43525 , n363684 , n363689 );
buf ( n363691 , n43525 );
and ( n363692 , n363691 , n41485 );
and ( n363693 , n41480 , n361609 );
nor ( n43529 , n363692 , n363693 );
buf ( n363695 , n43529 );
not ( n363696 , n363695 );
buf ( n363697 , n363696 );
buf ( n363698 , n363697 );
and ( n363699 , n363679 , n363698 );
not ( n43535 , n363679 );
buf ( n363701 , n43529 );
and ( n363702 , n43535 , n363701 );
nor ( n43538 , n363699 , n363702 );
buf ( n363704 , n43538 );
buf ( n363705 , n363704 );
buf ( n363706 , n361060 );
not ( n43542 , n363706 );
and ( n43543 , n40893 , n361073 );
not ( n363709 , n40893 );
and ( n43545 , n363709 , n39832 );
or ( n363711 , n43543 , n43545 );
buf ( n363712 , n363711 );
not ( n43548 , n363712 );
or ( n43549 , n43542 , n43548 );
buf ( n363715 , n361885 );
buf ( n363716 , n361022 );
nand ( n43552 , n363715 , n363716 );
buf ( n43553 , n43552 );
buf ( n363719 , n43553 );
nand ( n43555 , n43549 , n363719 );
buf ( n363721 , n43555 );
buf ( n363722 , n363721 );
xor ( n43558 , n363705 , n363722 );
buf ( n363724 , n43558 );
buf ( n363725 , n363724 );
xor ( n363726 , n363673 , n363725 );
buf ( n363727 , n363726 );
buf ( n363728 , n363727 );
xor ( n43564 , n362775 , n362868 );
and ( n43565 , n43564 , n363032 );
and ( n363731 , n362775 , n362868 );
or ( n43567 , n43565 , n363731 );
buf ( n363733 , n43567 );
buf ( n363734 , n363733 );
xor ( n43570 , n363728 , n363734 );
buf ( n43571 , n362855 );
buf ( n43572 , n362849 );
or ( n43573 , n43571 , n43572 );
buf ( n43574 , n43573 );
buf ( n363740 , n43574 );
buf ( n363741 , n362864 );
and ( n363742 , n363740 , n363741 );
and ( n363743 , n362850 , n362856 );
buf ( n363744 , n363743 );
buf ( n363745 , n363744 );
nor ( n363746 , n363742 , n363745 );
buf ( n363747 , n363746 );
xor ( n43583 , n42655 , n362820 );
and ( n363749 , n43583 , n362847 );
and ( n363750 , n42655 , n362820 );
or ( n43586 , n363749 , n363750 );
buf ( n363752 , n43586 );
buf ( n363753 , n363752 );
buf ( n363754 , n361631 );
buf ( n363755 , n41666 );
and ( n363756 , n363754 , n363755 );
not ( n363757 , n363754 );
buf ( n363758 , n41663 );
and ( n363759 , n363757 , n363758 );
or ( n363760 , n363756 , n363759 );
buf ( n363761 , n363760 );
or ( n43597 , n363761 , n361687 );
or ( n43598 , n362092 , n39707 );
nand ( n363764 , n43597 , n43598 );
not ( n363765 , n363764 );
buf ( n363766 , n39952 );
not ( n363767 , n363766 );
buf ( n363768 , n39966 );
not ( n363769 , n363768 );
buf ( n363770 , n360851 );
not ( n363771 , n363770 );
or ( n363772 , n363769 , n363771 );
buf ( n363773 , n360857 );
buf ( n363774 , n39963 );
nand ( n43610 , n363773 , n363774 );
buf ( n363776 , n43610 );
buf ( n363777 , n363776 );
nand ( n363778 , n363772 , n363777 );
buf ( n363779 , n363778 );
buf ( n363780 , n363779 );
not ( n363781 , n363780 );
or ( n43617 , n363767 , n363781 );
buf ( n363783 , n362792 );
buf ( n363784 , n40059 );
nand ( n363785 , n363783 , n363784 );
buf ( n363786 , n363785 );
buf ( n363787 , n363786 );
nand ( n363788 , n43617 , n363787 );
buf ( n363789 , n363788 );
xor ( n363790 , n363765 , n363789 );
buf ( n363791 , n39217 );
not ( n363792 , n363791 );
and ( n43628 , n361851 , n40275 );
not ( n363794 , n361851 );
and ( n363795 , n363794 , n360401 );
or ( n43631 , n43628 , n363795 );
buf ( n363797 , n43631 );
not ( n363798 , n363797 );
or ( n363799 , n363792 , n363798 );
buf ( n363800 , n42664 );
buf ( n363801 , n359307 );
nand ( n43637 , n363800 , n363801 );
buf ( n363803 , n43637 );
buf ( n363804 , n363803 );
nand ( n363805 , n363799 , n363804 );
buf ( n363806 , n363805 );
xor ( n43642 , n363790 , n363806 );
buf ( n363808 , n43642 );
xor ( n363809 , n363753 , n363808 );
buf ( n43645 , n39891 );
not ( n43646 , n43645 );
buf ( n363812 , n359950 );
not ( n43648 , n363812 );
buf ( n363814 , n362288 );
not ( n363815 , n363814 );
or ( n43651 , n43648 , n363815 );
buf ( n363817 , n362285 );
buf ( n363818 , n359955 );
nand ( n363819 , n363817 , n363818 );
buf ( n363820 , n363819 );
buf ( n363821 , n363820 );
nand ( n43657 , n43651 , n363821 );
buf ( n43658 , n43657 );
buf ( n363824 , n43658 );
not ( n43660 , n363824 );
or ( n363826 , n43646 , n43660 );
buf ( n363827 , n362155 );
buf ( n363828 , n359919 );
nand ( n363829 , n363827 , n363828 );
buf ( n363830 , n363829 );
buf ( n363831 , n363830 );
nand ( n43667 , n363826 , n363831 );
buf ( n363833 , n43667 );
buf ( n363834 , n363833 );
buf ( n363835 , n360577 );
not ( n43671 , n363835 );
buf ( n363837 , n360616 );
not ( n43673 , n363837 );
buf ( n363839 , n359784 );
not ( n43675 , n363839 );
or ( n363841 , n43673 , n43675 );
buf ( n363842 , n359781 );
buf ( n363843 , n362489 );
nand ( n363844 , n363842 , n363843 );
buf ( n363845 , n363844 );
buf ( n363846 , n363845 );
nand ( n363847 , n363841 , n363846 );
buf ( n363848 , n363847 );
buf ( n363849 , n363848 );
not ( n363850 , n363849 );
or ( n363851 , n43671 , n363850 );
buf ( n363852 , n362839 );
buf ( n363853 , n360601 );
nand ( n363854 , n363852 , n363853 );
buf ( n363855 , n363854 );
buf ( n363856 , n363855 );
nand ( n363857 , n363851 , n363856 );
buf ( n363858 , n363857 );
buf ( n363859 , n363858 );
xor ( n363860 , n363834 , n363859 );
buf ( n363861 , n362066 );
not ( n363862 , n363861 );
buf ( n363863 , n41892 );
buf ( n363864 , n40005 );
not ( n363865 , n363864 );
buf ( n363866 , n363865 );
buf ( n363867 , n363866 );
not ( n363868 , n363867 );
buf ( n363869 , n363868 );
buf ( n363870 , n363869 );
and ( n363871 , n363863 , n363870 );
not ( n363872 , n363863 );
buf ( n363873 , n363866 );
and ( n363874 , n363872 , n363873 );
nor ( n43710 , n363871 , n363874 );
buf ( n43711 , n43710 );
buf ( n363877 , n43711 );
not ( n43713 , n363877 );
or ( n363879 , n363862 , n43713 );
buf ( n363880 , n41911 );
buf ( n363881 , n362030 );
nand ( n363882 , n363880 , n363881 );
buf ( n363883 , n363882 );
buf ( n363884 , n363883 );
nand ( n363885 , n363879 , n363884 );
buf ( n363886 , n363885 );
buf ( n363887 , n363886 );
xor ( n43723 , n363860 , n363887 );
buf ( n363889 , n43723 );
buf ( n363890 , n363889 );
xor ( n43726 , n363809 , n363890 );
buf ( n363892 , n43726 );
xor ( n363893 , n363747 , n363892 );
not ( n363894 , n362172 );
not ( n363895 , n362360 );
or ( n43731 , n363894 , n363895 );
not ( n43732 , n362169 );
not ( n363898 , n362363 );
or ( n43734 , n43732 , n363898 );
nand ( n43735 , n43734 , n361910 );
nand ( n363901 , n43731 , n43735 );
xnor ( n363902 , n363893 , n363901 );
buf ( n363903 , n363902 );
xor ( n363904 , n43570 , n363903 );
buf ( n363905 , n363904 );
buf ( n363906 , n363905 );
xor ( n363907 , n42230 , n363035 );
and ( n363908 , n363907 , n43125 );
and ( n43744 , n42230 , n363035 );
or ( n363910 , n363908 , n43744 );
buf ( n363911 , n363910 );
buf ( n363912 , n363911 );
nor ( n43748 , n363906 , n363912 );
buf ( n363914 , n43748 );
buf ( n363915 , n363914 );
not ( n363916 , n363915 );
buf ( n363917 , n363916 );
nand ( n363918 , n363654 , n363917 );
not ( n43754 , n363761 );
not ( n363920 , n39707 );
and ( n363921 , n43754 , n363920 );
and ( n43757 , n359789 , n362136 );
not ( n363923 , n359789 );
and ( n363924 , n363923 , n362139 );
or ( n363925 , n43757 , n363924 );
and ( n43761 , n363925 , n39592 );
nor ( n363927 , n363921 , n43761 );
xor ( n43763 , n363764 , n363927 );
buf ( n363929 , n355582 );
not ( n43765 , n363929 );
buf ( n363931 , n40797 );
not ( n363932 , n363931 );
or ( n43768 , n43765 , n363932 );
buf ( n363934 , n40201 );
buf ( n363935 , n40945 );
nand ( n43771 , n363934 , n363935 );
buf ( n363937 , n43771 );
buf ( n363938 , n363937 );
nand ( n43774 , n43768 , n363938 );
buf ( n363940 , n43774 );
buf ( n363941 , n363940 );
not ( n363942 , n363941 );
buf ( n363943 , n39218 );
nor ( n43779 , n363942 , n363943 );
buf ( n363945 , n43779 );
buf ( n363946 , n363945 );
buf ( n363947 , n43631 );
not ( n363948 , n363947 );
buf ( n363949 , n359310 );
nor ( n43785 , n363948 , n363949 );
buf ( n43786 , n43785 );
buf ( n363952 , n43786 );
nor ( n363953 , n363946 , n363952 );
buf ( n363954 , n363953 );
buf ( n363955 , n363954 );
xnor ( n363956 , n43763 , n363955 );
buf ( n363957 , n363956 );
buf ( n363958 , n363721 );
buf ( n363959 , n363697 );
or ( n43795 , n363958 , n363959 );
buf ( n363961 , n363678 );
nand ( n43797 , n43795 , n363961 );
buf ( n43798 , n43797 );
buf ( n363964 , n43798 );
buf ( n43800 , n363721 );
buf ( n363966 , n363697 );
nand ( n363967 , n43800 , n363966 );
buf ( n363968 , n363967 );
buf ( n363969 , n363968 );
and ( n363970 , n363964 , n363969 );
buf ( n363971 , n363970 );
buf ( n363972 , n363971 );
xor ( n363973 , n363957 , n363972 );
buf ( n363974 , n41892 );
not ( n43810 , n363974 );
buf ( n363976 , n40092 );
not ( n43812 , n363976 );
or ( n363978 , n43810 , n43812 );
buf ( n363979 , n40899 );
buf ( n363980 , n363979 );
buf ( n363981 , n362037 );
nand ( n363982 , n363980 , n363981 );
buf ( n363983 , n363982 );
buf ( n363984 , n363983 );
nand ( n43820 , n363978 , n363984 );
buf ( n43821 , n43820 );
buf ( n363987 , n43821 );
buf ( n43823 , n362066 );
buf ( n363989 , n43823 );
and ( n363990 , n363987 , n363989 );
buf ( n363991 , n43711 );
not ( n363992 , n363991 );
buf ( n363993 , n362030 );
not ( n363994 , n363993 );
buf ( n363995 , n363994 );
buf ( n363996 , n363995 );
nor ( n43832 , n363992 , n363996 );
buf ( n363998 , n43832 );
buf ( n363999 , n363998 );
nor ( n364000 , n363990 , n363999 );
buf ( n364001 , n364000 );
buf ( n364002 , n364001 );
buf ( n364003 , n360616 );
not ( n43839 , n364003 );
buf ( n364005 , n39655 );
not ( n364006 , n364005 );
or ( n364007 , n43839 , n364006 );
buf ( n364008 , n359756 );
buf ( n364009 , n360613 );
nand ( n43845 , n364008 , n364009 );
buf ( n364011 , n43845 );
buf ( n364012 , n364011 );
nand ( n43848 , n364007 , n364012 );
buf ( n364014 , n43848 );
buf ( n364015 , n364014 );
buf ( n364016 , n360577 );
and ( n364017 , n364015 , n364016 );
buf ( n364018 , n363848 );
buf ( n364019 , n360601 );
and ( n364020 , n364018 , n364019 );
buf ( n364021 , n364020 );
buf ( n364022 , n364021 );
nor ( n364023 , n364017 , n364022 );
buf ( n364024 , n364023 );
buf ( n364025 , n364024 );
xor ( n364026 , n364002 , n364025 );
xor ( n364027 , n361026 , n39870 );
buf ( n364028 , n364027 );
not ( n364029 , n364028 );
buf ( n364030 , n361116 );
not ( n364031 , n364030 );
and ( n43867 , n364029 , n364031 );
buf ( n364033 , n363711 );
buf ( n43869 , n361022 );
and ( n43870 , n364033 , n43869 );
nor ( n43871 , n43867 , n43870 );
buf ( n43872 , n43871 );
buf ( n364038 , n43872 );
xor ( n43874 , n364026 , n364038 );
buf ( n364040 , n43874 );
buf ( n364041 , n364040 );
xor ( n364042 , n363973 , n364041 );
buf ( n364043 , n364042 );
buf ( n364044 , n364043 );
buf ( n364045 , n363901 );
buf ( n364046 , n363892 );
not ( n43882 , n364046 );
buf ( n364048 , n363747 );
nand ( n43884 , n43882 , n364048 );
buf ( n43885 , n43884 );
buf ( n364051 , n43885 );
nand ( n364052 , n364045 , n364051 );
buf ( n364053 , n364052 );
buf ( n364054 , n364053 );
buf ( n364055 , n363747 );
not ( n43891 , n364055 );
buf ( n364057 , n363892 );
nand ( n364058 , n43891 , n364057 );
buf ( n364059 , n364058 );
buf ( n364060 , n364059 );
and ( n43896 , n364054 , n364060 );
buf ( n364062 , n43896 );
buf ( n364063 , n364062 );
xor ( n364064 , n364044 , n364063 );
xor ( n43900 , n363765 , n363789 );
and ( n364066 , n43900 , n363806 );
and ( n43902 , n363765 , n363789 );
or ( n43903 , n364066 , n43902 );
buf ( n364069 , n43903 );
not ( n43905 , n40059 );
not ( n43906 , n363779 );
or ( n364072 , n43905 , n43906 );
buf ( n43908 , n40251 );
xnor ( n364074 , n39963 , n43908 );
nand ( n43910 , n364074 , n39952 );
nand ( n364076 , n364072 , n43910 );
buf ( n364077 , n359919 );
not ( n364078 , n364077 );
buf ( n364079 , n43658 );
not ( n43915 , n364079 );
or ( n364081 , n364078 , n43915 );
and ( n364082 , n359950 , n40756 );
not ( n43918 , n359950 );
and ( n364084 , n43918 , n360893 );
or ( n364085 , n364082 , n364084 );
buf ( n364086 , n364085 );
buf ( n364087 , n39891 );
nand ( n43923 , n364086 , n364087 );
buf ( n364089 , n43923 );
buf ( n364090 , n364089 );
nand ( n364091 , n364081 , n364090 );
buf ( n364092 , n364091 );
not ( n364093 , n364092 );
xor ( n43929 , n364076 , n364093 );
buf ( n364095 , n363691 );
buf ( n364096 , n361609 );
not ( n43932 , n364096 );
not ( n364098 , n41485 );
buf ( n364099 , n364098 );
nand ( n364100 , n43932 , n364099 );
buf ( n364101 , n364100 );
buf ( n364102 , n364101 );
and ( n364103 , n364095 , n364102 );
buf ( n364104 , n364103 );
xor ( n43940 , n43929 , n364104 );
buf ( n364106 , n43940 );
xor ( n43942 , n364069 , n364106 );
xor ( n43943 , n363834 , n363859 );
and ( n364109 , n43943 , n363887 );
and ( n43945 , n363834 , n363859 );
or ( n364111 , n364109 , n43945 );
buf ( n364112 , n364111 );
buf ( n364113 , n364112 );
xor ( n43949 , n43942 , n364113 );
buf ( n364115 , n43949 );
buf ( n364116 , n364115 );
xor ( n43952 , n363753 , n363808 );
and ( n43953 , n43952 , n363890 );
and ( n364119 , n363753 , n363808 );
or ( n364120 , n43953 , n364119 );
buf ( n364121 , n364120 );
buf ( n364122 , n364121 );
and ( n43958 , n364116 , n364122 );
not ( n364124 , n364116 );
buf ( n364125 , n364121 );
not ( n43961 , n364125 );
buf ( n364127 , n43961 );
buf ( n43963 , n364127 );
and ( n364129 , n364124 , n43963 );
nor ( n43965 , n43958 , n364129 );
buf ( n43966 , n43965 );
xor ( n364132 , n43495 , n363672 );
and ( n43968 , n364132 , n363725 );
and ( n364134 , n43495 , n363672 );
or ( n364135 , n43968 , n364134 );
buf ( n364136 , n364135 );
xnor ( n364137 , n43966 , n364136 );
buf ( n364138 , n364137 );
xor ( n43974 , n364064 , n364138 );
buf ( n364140 , n43974 );
xor ( n43976 , n363728 , n363734 );
and ( n43977 , n43976 , n363903 );
and ( n364143 , n363728 , n363734 );
or ( n43979 , n43977 , n364143 );
buf ( n364145 , n43979 );
not ( n43981 , n364145 );
nand ( n364147 , n364140 , n43981 );
not ( n364148 , n364147 );
nor ( n43984 , n363918 , n364148 );
xor ( n364150 , n364044 , n364063 );
and ( n364151 , n364150 , n364138 );
and ( n43987 , n364044 , n364063 );
or ( n364153 , n364151 , n43987 );
buf ( n364154 , n364153 );
buf ( n364155 , n364154 );
buf ( n364156 , n40059 );
not ( n364157 , n364156 );
buf ( n364158 , n364074 );
not ( n364159 , n364158 );
or ( n43995 , n364157 , n364159 );
buf ( n364161 , n39966 );
not ( n364162 , n364161 );
buf ( n364163 , n360401 );
not ( n364164 , n364163 );
or ( n44000 , n364162 , n364164 );
buf ( n364166 , n40275 );
buf ( n364167 , n39963 );
nand ( n44003 , n364166 , n364167 );
buf ( n44004 , n44003 );
buf ( n364170 , n44004 );
nand ( n364171 , n44000 , n364170 );
buf ( n364172 , n364171 );
buf ( n364173 , n364172 );
buf ( n364174 , n39952 );
nand ( n44010 , n364173 , n364174 );
buf ( n44011 , n44010 );
buf ( n364177 , n44011 );
nand ( n44013 , n43995 , n364177 );
buf ( n364179 , n44013 );
not ( n364180 , n359815 );
not ( n364181 , n363925 );
or ( n44017 , n364180 , n364181 );
and ( n364183 , n362285 , n359789 );
not ( n364184 , n362285 );
and ( n44020 , n364184 , n359720 );
or ( n364186 , n364183 , n44020 );
nand ( n44022 , n364186 , n39592 );
nand ( n364188 , n44017 , n44022 );
xor ( n44024 , n364179 , n364188 );
buf ( n364190 , n39217 );
not ( n364191 , n364190 );
buf ( n364192 , n355582 );
not ( n44028 , n364192 );
buf ( n364194 , n359784 );
not ( n44030 , n364194 );
or ( n364196 , n44028 , n44030 );
buf ( n364197 , n359781 );
buf ( n364198 , n40945 );
nand ( n364199 , n364197 , n364198 );
buf ( n364200 , n364199 );
buf ( n364201 , n364200 );
nand ( n364202 , n364196 , n364201 );
buf ( n364203 , n364202 );
buf ( n364204 , n364203 );
not ( n364205 , n364204 );
or ( n44041 , n364191 , n364205 );
buf ( n364207 , n363940 );
buf ( n364208 , n359307 );
nand ( n44044 , n364207 , n364208 );
buf ( n364210 , n44044 );
buf ( n364211 , n364210 );
nand ( n44047 , n44041 , n364211 );
buf ( n364213 , n44047 );
xnor ( n44049 , n44024 , n364213 );
buf ( n364215 , n44049 );
buf ( n364216 , n39891 );
not ( n364217 , n364216 );
buf ( n364218 , n359950 );
not ( n364219 , n364218 );
buf ( n364220 , n360851 );
not ( n44056 , n364220 );
or ( n364222 , n364219 , n44056 );
buf ( n364223 , n360857 );
buf ( n364224 , n359955 );
nand ( n364225 , n364223 , n364224 );
buf ( n364226 , n364225 );
buf ( n364227 , n364226 );
nand ( n44063 , n364222 , n364227 );
buf ( n44064 , n44063 );
buf ( n364230 , n44064 );
not ( n44066 , n364230 );
or ( n364232 , n364217 , n44066 );
buf ( n44068 , n364085 );
buf ( n364234 , n359919 );
nand ( n44070 , n44068 , n364234 );
buf ( n364236 , n44070 );
buf ( n364237 , n364236 );
nand ( n364238 , n364232 , n364237 );
buf ( n364239 , n364238 );
buf ( n364240 , n364239 );
buf ( n364241 , n364027 );
not ( n364242 , n364241 );
buf ( n364243 , n361121 );
not ( n364244 , n364243 );
and ( n44080 , n364242 , n364244 );
buf ( n364246 , n40893 );
not ( n364247 , n364246 );
buf ( n364248 , n360116 );
not ( n364249 , n364248 );
or ( n364250 , n364247 , n364249 );
buf ( n364251 , n360122 );
buf ( n364252 , n361026 );
nand ( n44088 , n364251 , n364252 );
buf ( n364254 , n44088 );
buf ( n364255 , n364254 );
nand ( n44091 , n364250 , n364255 );
buf ( n364257 , n44091 );
buf ( n364258 , n364257 );
buf ( n364259 , n361060 );
and ( n364260 , n364258 , n364259 );
nor ( n364261 , n44080 , n364260 );
buf ( n364262 , n364261 );
buf ( n364263 , n364262 );
xor ( n364264 , n364240 , n364263 );
buf ( n364265 , n41892 );
buf ( n364266 , n359147 );
and ( n44102 , n364265 , n364266 );
not ( n44103 , n364265 );
buf ( n44104 , n360624 );
and ( n364270 , n44103 , n44104 );
nor ( n44106 , n44102 , n364270 );
buf ( n44107 , n44106 );
buf ( n364273 , n44107 );
not ( n44109 , n364273 );
buf ( n364275 , n362063 );
not ( n364276 , n364275 );
and ( n44112 , n44109 , n364276 );
buf ( n364278 , n43821 );
buf ( n364279 , n362030 );
and ( n364280 , n364278 , n364279 );
nor ( n44116 , n44112 , n364280 );
buf ( n364282 , n44116 );
buf ( n364283 , n364282 );
xor ( n44119 , n364264 , n364283 );
buf ( n364285 , n44119 );
buf ( n364286 , n364285 );
xor ( n44122 , n364215 , n364286 );
xor ( n44123 , n364002 , n364025 );
and ( n364289 , n44123 , n364038 );
and ( n44125 , n364002 , n364025 );
or ( n364291 , n364289 , n44125 );
buf ( n364292 , n364291 );
buf ( n364293 , n364292 );
xor ( n44129 , n44122 , n364293 );
buf ( n364295 , n44129 );
buf ( n364296 , n364295 );
buf ( n364297 , n364121 );
not ( n364298 , n364297 );
not ( n44134 , n364115 );
not ( n364300 , n44134 );
buf ( n44136 , n364300 );
not ( n44137 , n44136 );
or ( n44138 , n364298 , n44137 );
buf ( n364304 , n44134 );
not ( n44140 , n364304 );
buf ( n364306 , n364127 );
not ( n364307 , n364306 );
or ( n364308 , n44140 , n364307 );
buf ( n364309 , n364136 );
nand ( n364310 , n364308 , n364309 );
buf ( n364311 , n364310 );
buf ( n364312 , n364311 );
nand ( n364313 , n44138 , n364312 );
buf ( n364314 , n364313 );
buf ( n364315 , n364314 );
not ( n44151 , n364315 );
buf ( n364317 , n44151 );
buf ( n364318 , n364317 );
xor ( n44154 , n364296 , n364318 );
buf ( n364320 , n360613 );
buf ( n364321 , n361073 );
and ( n364322 , n364320 , n364321 );
not ( n364323 , n364320 );
buf ( n364324 , n39832 );
and ( n44160 , n364323 , n364324 );
or ( n364326 , n364322 , n44160 );
buf ( n364327 , n364326 );
not ( n364328 , n364327 );
not ( n364329 , n360580 );
and ( n364330 , n364328 , n364329 );
buf ( n364331 , n364014 );
not ( n364332 , n364331 );
buf ( n364333 , n360604 );
nor ( n44169 , n364332 , n364333 );
buf ( n44170 , n44169 );
nor ( n44171 , n364330 , n44170 );
buf ( n364337 , n44171 );
not ( n364338 , n364076 );
not ( n44174 , n364092 );
and ( n44175 , n364338 , n44174 );
nor ( n44176 , n44175 , n364104 );
not ( n364342 , n364076 );
nor ( n44178 , n364342 , n364093 );
nor ( n364344 , n44176 , n44178 );
buf ( n364345 , n364344 );
xor ( n44181 , n364337 , n364345 );
or ( n44182 , n363927 , n363955 );
nand ( n44183 , n44182 , n363765 );
nand ( n44184 , n363955 , n363927 );
nand ( n44185 , n44183 , n44184 );
buf ( n364351 , n44185 );
xor ( n364352 , n44181 , n364351 );
buf ( n364353 , n364352 );
buf ( n364354 , n364353 );
buf ( n364355 , n43903 );
not ( n44191 , n364355 );
buf ( n364357 , n43940 );
not ( n44193 , n364357 );
buf ( n364359 , n44193 );
buf ( n364360 , n364359 );
nand ( n44196 , n44191 , n364360 );
buf ( n364362 , n44196 );
buf ( n364363 , n364362 );
buf ( n364364 , n364112 );
and ( n364365 , n364363 , n364364 );
buf ( n364366 , n43903 );
not ( n44202 , n364366 );
buf ( n364368 , n364359 );
nor ( n44204 , n44202 , n364368 );
buf ( n364370 , n44204 );
buf ( n364371 , n364370 );
nor ( n44207 , n364365 , n364371 );
buf ( n364373 , n44207 );
buf ( n364374 , n364373 );
xor ( n364375 , n364354 , n364374 );
xor ( n364376 , n363957 , n363972 );
and ( n44212 , n364376 , n364041 );
and ( n44213 , n363957 , n363972 );
or ( n364379 , n44212 , n44213 );
buf ( n364380 , n364379 );
buf ( n364381 , n364380 );
xor ( n364382 , n364375 , n364381 );
buf ( n364383 , n364382 );
buf ( n364384 , n364383 );
xor ( n364385 , n44154 , n364384 );
buf ( n364386 , n364385 );
buf ( n364387 , n364386 );
nand ( n44223 , n364155 , n364387 );
buf ( n364389 , n44223 );
and ( n364390 , n43984 , n364389 );
buf ( n364391 , n359815 );
not ( n364392 , n364391 );
buf ( n364393 , n364186 );
not ( n44229 , n364393 );
or ( n364395 , n364392 , n44229 );
buf ( n364396 , n360900 );
buf ( n364397 , n39592 );
nand ( n364398 , n364396 , n364397 );
buf ( n364399 , n364398 );
buf ( n364400 , n364399 );
nand ( n364401 , n364395 , n364400 );
buf ( n364402 , n364401 );
buf ( n364403 , n364402 );
buf ( n364404 , n39952 );
not ( n364405 , n364404 );
buf ( n364406 , n361292 );
not ( n364407 , n364406 );
or ( n44243 , n364405 , n364407 );
buf ( n364409 , n364172 );
buf ( n364410 , n40059 );
nand ( n364411 , n364409 , n364410 );
buf ( n364412 , n364411 );
buf ( n364413 , n364412 );
nand ( n364414 , n44243 , n364413 );
buf ( n364415 , n364414 );
buf ( n364416 , n364415 );
xor ( n364417 , n364403 , n364416 );
buf ( n364418 , n39891 );
not ( n364419 , n364418 );
buf ( n364420 , n361240 );
not ( n364421 , n364420 );
or ( n44257 , n364419 , n364421 );
buf ( n364423 , n44064 );
buf ( n364424 , n359919 );
nand ( n44260 , n364423 , n364424 );
buf ( n364426 , n44260 );
buf ( n364427 , n364426 );
nand ( n44263 , n44257 , n364427 );
buf ( n364429 , n44263 );
buf ( n364430 , n364429 );
xor ( n44266 , n364417 , n364430 );
buf ( n364432 , n44266 );
xor ( n364433 , n364240 , n364263 );
and ( n44269 , n364433 , n364283 );
and ( n364435 , n364240 , n364263 );
or ( n44271 , n44269 , n364435 );
buf ( n364437 , n44271 );
not ( n44273 , n364437 );
and ( n44274 , n364432 , n44273 );
not ( n364440 , n364432 );
and ( n364441 , n364440 , n364437 );
nor ( n44277 , n44274 , n364441 );
buf ( n364443 , n364239 );
not ( n364444 , n364443 );
buf ( n364445 , n364444 );
buf ( n364446 , n364445 );
and ( n364447 , n363995 , n362063 );
nor ( n44283 , n364447 , n44107 );
buf ( n364449 , n44283 );
xor ( n364450 , n364446 , n364449 );
buf ( n364451 , n361040 );
buf ( n364452 , n361060 );
buf ( n364453 , n364452 );
and ( n364454 , n364451 , n364453 );
buf ( n364455 , n364257 );
not ( n44291 , n364455 );
buf ( n364457 , n361121 );
nor ( n44293 , n44291 , n364457 );
buf ( n364459 , n44293 );
buf ( n364460 , n364459 );
nor ( n364461 , n364454 , n364460 );
buf ( n364462 , n364461 );
buf ( n364463 , n364462 );
xor ( n44299 , n364450 , n364463 );
buf ( n364465 , n44299 );
and ( n364466 , n44277 , n364465 );
not ( n44302 , n44277 );
buf ( n364468 , n364465 );
not ( n364469 , n364468 );
buf ( n364470 , n364469 );
and ( n44306 , n44302 , n364470 );
nor ( n364472 , n364466 , n44306 );
xor ( n364473 , n364337 , n364345 );
and ( n44309 , n364473 , n364351 );
and ( n364475 , n364337 , n364345 );
or ( n44311 , n44309 , n364475 );
buf ( n364477 , n44311 );
buf ( n364478 , n364477 );
and ( n364479 , n361100 , n39217 );
and ( n44315 , n364203 , n359307 );
nor ( n364481 , n364479 , n44315 );
buf ( n364482 , n364481 );
not ( n44318 , n364482 );
buf ( n364484 , n44318 );
buf ( n44320 , n361265 );
not ( n364486 , n44320 );
buf ( n364487 , n364486 );
buf ( n364488 , n364487 );
not ( n364489 , n364488 );
buf ( n364490 , n360580 );
not ( n364491 , n364490 );
and ( n44327 , n364489 , n364491 );
buf ( n364493 , n364327 );
not ( n44329 , n364493 );
buf ( n364495 , n44329 );
buf ( n364496 , n364495 );
buf ( n364497 , n360601 );
and ( n44333 , n364496 , n364497 );
nor ( n364499 , n44327 , n44333 );
buf ( n364500 , n364499 );
xor ( n364501 , n364484 , n364500 );
buf ( n364502 , n364179 );
not ( n364503 , n364502 );
buf ( n44339 , n364213 );
not ( n44340 , n44339 );
or ( n44341 , n364503 , n44340 );
buf ( n364507 , n364213 );
buf ( n364508 , n364179 );
or ( n44344 , n364507 , n364508 );
buf ( n364510 , n364188 );
nand ( n364511 , n44344 , n364510 );
buf ( n364512 , n364511 );
buf ( n364513 , n364512 );
nand ( n364514 , n44341 , n364513 );
buf ( n364515 , n364514 );
xor ( n44351 , n364501 , n364515 );
buf ( n364517 , n44351 );
xor ( n44353 , n364478 , n364517 );
xor ( n44354 , n364215 , n364286 );
and ( n364520 , n44354 , n364293 );
and ( n364521 , n364215 , n364286 );
or ( n44357 , n364520 , n364521 );
buf ( n364523 , n44357 );
buf ( n364524 , n364523 );
xor ( n44360 , n44353 , n364524 );
buf ( n364526 , n44360 );
xor ( n44362 , n364472 , n364526 );
xor ( n44363 , n364354 , n364374 );
and ( n364529 , n44363 , n364381 );
and ( n44365 , n364354 , n364374 );
or ( n364531 , n364529 , n44365 );
buf ( n364532 , n364531 );
xor ( n44368 , n44362 , n364532 );
buf ( n364534 , n44368 );
xor ( n44370 , n364296 , n364318 );
and ( n364536 , n44370 , n364384 );
and ( n364537 , n364296 , n364318 );
or ( n44373 , n364536 , n364537 );
buf ( n364539 , n44373 );
buf ( n364540 , n364539 );
nand ( n364541 , n364534 , n364540 );
buf ( n364542 , n364541 );
xor ( n44378 , n364446 , n364449 );
and ( n364544 , n44378 , n364463 );
and ( n44380 , n364446 , n364449 );
or ( n364546 , n364544 , n44380 );
buf ( n364547 , n364546 );
buf ( n364548 , n364547 );
xor ( n44384 , n364403 , n364416 );
and ( n364550 , n44384 , n364430 );
and ( n364551 , n364403 , n364416 );
or ( n44387 , n364550 , n364551 );
buf ( n364553 , n44387 );
buf ( n364554 , n364553 );
xnor ( n44390 , n364548 , n364554 );
buf ( n44391 , n44390 );
buf ( n364557 , n44391 );
xor ( n44393 , n361269 , n361250 );
xnor ( n364559 , n44393 , n361299 );
buf ( n364560 , n364559 );
and ( n44396 , n364557 , n364560 );
not ( n364562 , n364557 );
buf ( n364563 , n364559 );
not ( n44399 , n364563 );
buf ( n44400 , n44399 );
buf ( n364566 , n44400 );
and ( n44402 , n364562 , n364566 );
nor ( n364568 , n44396 , n44402 );
buf ( n364569 , n364568 );
buf ( n364570 , n364569 );
buf ( n364571 , n364500 );
not ( n364572 , n364571 );
buf ( n364573 , n364572 );
buf ( n364574 , n364573 );
not ( n364575 , n364574 );
buf ( n364576 , n364484 );
not ( n44412 , n364576 );
or ( n364578 , n364575 , n44412 );
buf ( n44414 , n364515 );
buf ( n364580 , n364481 );
buf ( n364581 , n364500 );
nand ( n44417 , n364580 , n364581 );
buf ( n364583 , n44417 );
buf ( n364584 , n364583 );
nand ( n44420 , n44414 , n364584 );
buf ( n364586 , n44420 );
buf ( n364587 , n364586 );
nand ( n44423 , n364578 , n364587 );
buf ( n364589 , n44423 );
buf ( n364590 , n364589 );
xor ( n364591 , n360974 , n361067 );
xor ( n364592 , n364591 , n361108 );
buf ( n364593 , n364592 );
buf ( n364594 , n364593 );
and ( n364595 , n364590 , n364594 );
not ( n44431 , n364590 );
buf ( n364597 , n364593 );
not ( n364598 , n364597 );
buf ( n364599 , n364598 );
buf ( n364600 , n364599 );
and ( n364601 , n44431 , n364600 );
nor ( n364602 , n364595 , n364601 );
buf ( n364603 , n364602 );
buf ( n364604 , n364603 );
buf ( n364605 , n364465 );
not ( n44441 , n364605 );
buf ( n364607 , n364437 );
not ( n364608 , n364607 );
or ( n44444 , n44441 , n364608 );
buf ( n364610 , n364432 );
nand ( n44446 , n44444 , n364610 );
buf ( n364612 , n44446 );
buf ( n44448 , n364612 );
buf ( n364614 , n364437 );
not ( n44450 , n364614 );
buf ( n364616 , n364470 );
nand ( n364617 , n44450 , n364616 );
buf ( n364618 , n364617 );
buf ( n364619 , n364618 );
nand ( n364620 , n44448 , n364619 );
buf ( n364621 , n364620 );
buf ( n364622 , n364621 );
xnor ( n44458 , n364604 , n364622 );
buf ( n364624 , n44458 );
buf ( n364625 , n364624 );
xor ( n364626 , n364570 , n364625 );
xor ( n44462 , n364478 , n364517 );
and ( n364628 , n44462 , n364524 );
and ( n44464 , n364478 , n364517 );
or ( n44465 , n364628 , n44464 );
buf ( n364631 , n44465 );
buf ( n364632 , n364631 );
xor ( n44468 , n364626 , n364632 );
buf ( n364634 , n44468 );
buf ( n364635 , n364634 );
xor ( n44471 , n364472 , n364526 );
and ( n364637 , n44471 , n364532 );
and ( n364638 , n364472 , n364526 );
or ( n44474 , n364637 , n364638 );
buf ( n364640 , n44474 );
nand ( n44476 , n364635 , n364640 );
buf ( n364642 , n44476 );
nand ( n364643 , n364542 , n364642 );
not ( n44479 , n364643 );
xor ( n364645 , n364570 , n364625 );
and ( n44481 , n364645 , n364632 );
and ( n44482 , n364570 , n364625 );
or ( n44483 , n44481 , n44482 );
buf ( n364649 , n44483 );
buf ( n364650 , n364559 );
not ( n44486 , n364650 );
buf ( n364652 , n364547 );
not ( n44488 , n364652 );
or ( n364654 , n44486 , n44488 );
buf ( n364655 , n364553 );
nand ( n364656 , n364654 , n364655 );
buf ( n364657 , n364656 );
buf ( n364658 , n364657 );
buf ( n364659 , n364547 );
not ( n44495 , n364659 );
buf ( n364661 , n44400 );
nand ( n44497 , n44495 , n364661 );
buf ( n364663 , n44497 );
buf ( n364664 , n364663 );
nand ( n44500 , n364658 , n364664 );
buf ( n364666 , n44500 );
buf ( n364667 , n364666 );
not ( n364668 , n364667 );
xor ( n44504 , n361113 , n361195 );
xor ( n44505 , n44504 , n361309 );
buf ( n364671 , n44505 );
buf ( n364672 , n364671 );
not ( n44508 , n364672 );
buf ( n364674 , n44508 );
buf ( n364675 , n364674 );
not ( n44511 , n364675 );
or ( n44512 , n364668 , n44511 );
buf ( n364678 , n364671 );
buf ( n364679 , n364666 );
not ( n44515 , n364679 );
buf ( n364681 , n44515 );
buf ( n364682 , n364681 );
nand ( n44518 , n364678 , n364682 );
buf ( n364684 , n44518 );
buf ( n364685 , n364684 );
nand ( n44521 , n44512 , n364685 );
buf ( n364687 , n44521 );
buf ( n364688 , n364589 );
not ( n364689 , n364688 );
buf ( n364690 , n364599 );
nand ( n44526 , n364689 , n364690 );
buf ( n44527 , n44526 );
buf ( n364693 , n44527 );
not ( n44529 , n364693 );
buf ( n364695 , n364621 );
not ( n364696 , n364695 );
or ( n44532 , n44529 , n364696 );
buf ( n364698 , n364589 );
buf ( n364699 , n364593 );
nand ( n44535 , n364698 , n364699 );
buf ( n364701 , n44535 );
buf ( n364702 , n364701 );
nand ( n364703 , n44532 , n364702 );
buf ( n364704 , n364703 );
xnor ( n44540 , n364687 , n364704 );
nand ( n44541 , n364649 , n44540 );
buf ( n364707 , n364681 );
not ( n364708 , n364707 );
buf ( n364709 , n364674 );
not ( n364710 , n364709 );
or ( n364711 , n364708 , n364710 );
buf ( n364712 , n364704 );
nand ( n364713 , n364711 , n364712 );
buf ( n364714 , n364713 );
buf ( n364715 , n364714 );
buf ( n364716 , n364671 );
buf ( n364717 , n364666 );
nand ( n44553 , n364716 , n364717 );
buf ( n364719 , n44553 );
buf ( n364720 , n364719 );
nand ( n364721 , n364715 , n364720 );
buf ( n364722 , n364721 );
xor ( n44558 , n360970 , n41175 );
xor ( n44559 , n44558 , n361374 );
buf ( n44560 , n44559 );
or ( n364726 , n364722 , n44560 );
and ( n44562 , n44479 , n44541 , n364726 );
nand ( n364728 , n364390 , n44562 );
not ( n44564 , n364728 );
buf ( n364730 , n44564 );
not ( n364731 , n364730 );
not ( n44567 , n41835 );
buf ( n44568 , n41772 );
not ( n44569 , n44568 );
buf ( n44570 , n44569 );
buf ( n364736 , n44570 );
not ( n44572 , n364736 );
not ( n44573 , n42355 );
buf ( n364739 , n44573 );
not ( n44575 , n364739 );
or ( n44576 , n44572 , n44575 );
buf ( n364742 , n361911 );
buf ( n44578 , n364742 );
buf ( n364744 , n44578 );
buf ( n364745 , n364744 );
not ( n44581 , n364745 );
not ( n364747 , n32085 );
buf ( n364748 , n364747 );
nand ( n364749 , n44581 , n364748 );
buf ( n364750 , n364749 );
buf ( n364751 , n364750 );
nand ( n364752 , n44576 , n364751 );
buf ( n364753 , n364752 );
not ( n364754 , n364753 );
or ( n44590 , n44567 , n364754 );
not ( n44591 , n361971 );
buf ( n364757 , n44591 );
buf ( n364758 , n41452 );
buf ( n364759 , n364758 );
buf ( n364760 , n364759 );
buf ( n364761 , n364760 );
not ( n364762 , n364761 );
buf ( n364763 , n364762 );
buf ( n364764 , n364763 );
not ( n364765 , n364764 );
buf ( n364766 , n364765 );
buf ( n364767 , n364766 );
not ( n364768 , n364767 );
buf ( n44604 , n351762 );
not ( n364770 , n44604 );
buf ( n364771 , n364770 );
buf ( n364772 , n364771 );
not ( n364773 , n364772 );
buf ( n364774 , n364773 );
buf ( n364775 , n364774 );
not ( n364776 , n364775 );
buf ( n364777 , n364776 );
buf ( n364778 , n364777 );
not ( n364779 , n364778 );
or ( n44615 , n364768 , n364779 );
buf ( n364781 , n361911 );
not ( n364782 , n364781 );
buf ( n364783 , n364782 );
buf ( n364784 , n364783 );
buf ( n364785 , n31730 );
nand ( n364786 , n364784 , n364785 );
buf ( n364787 , n364786 );
buf ( n364788 , n364787 );
nand ( n364789 , n44615 , n364788 );
buf ( n364790 , n364789 );
buf ( n364791 , n364790 );
nand ( n44627 , n364757 , n364791 );
buf ( n364793 , n44627 );
nand ( n44629 , n44590 , n364793 );
buf ( n364795 , n41882 );
not ( n364796 , n364795 );
buf ( n364797 , n364796 );
not ( n364798 , n364797 );
not ( n44634 , n362033 );
buf ( n364800 , n44634 );
not ( n364801 , n364800 );
nand ( n44637 , n351310 , n351315 );
buf ( n44638 , n44637 );
not ( n364804 , n44638 );
buf ( n364805 , n364804 );
not ( n44641 , n364805 );
or ( n364807 , n364801 , n44641 );
not ( n364808 , n44637 );
buf ( n364809 , n364808 );
not ( n364810 , n364809 );
buf ( n364811 , n41892 );
nand ( n364812 , n364810 , n364811 );
buf ( n364813 , n364812 );
buf ( n364814 , n364813 );
nand ( n364815 , n364807 , n364814 );
buf ( n364816 , n364815 );
not ( n364817 , n364816 );
or ( n364818 , n364798 , n364817 );
buf ( n364819 , n41915 );
not ( n44655 , n364819 );
buf ( n364821 , n44655 );
buf ( n364822 , n364821 );
not ( n44658 , n364822 );
buf ( n364824 , n44658 );
buf ( n364825 , n364824 );
not ( n44661 , n31072 );
not ( n364827 , n44661 );
buf ( n364828 , n364827 );
not ( n44664 , n364828 );
buf ( n364830 , n362033 );
not ( n364831 , n364830 );
buf ( n364832 , n364831 );
buf ( n364833 , n364832 );
not ( n44669 , n364833 );
or ( n364835 , n44664 , n44669 );
buf ( n364836 , n41892 );
buf ( n364837 , n44661 );
nand ( n44673 , n364836 , n364837 );
buf ( n364839 , n44673 );
buf ( n364840 , n364839 );
nand ( n364841 , n364835 , n364840 );
buf ( n364842 , n364841 );
buf ( n364843 , n364842 );
nand ( n364844 , n364825 , n364843 );
buf ( n364845 , n364844 );
nand ( n44681 , n364818 , n364845 );
xor ( n364847 , n44629 , n44681 );
buf ( n364848 , n361600 );
not ( n364849 , n364848 );
buf ( n364850 , n364849 );
not ( n44686 , n364850 );
buf ( n364852 , n44686 );
buf ( n364853 , n351364 );
not ( n364854 , n364853 );
buf ( n364855 , n364854 );
buf ( n364856 , n364855 );
not ( n44692 , n364856 );
buf ( n364858 , n44692 );
buf ( n364859 , n364858 );
not ( n364860 , n364859 );
buf ( n364861 , n361534 );
not ( n44697 , n364861 );
or ( n364863 , n364860 , n44697 );
buf ( n364864 , n361531 );
buf ( n364865 , n351364 );
not ( n364866 , n364865 );
buf ( n364867 , n364866 );
buf ( n364868 , n364867 );
buf ( n364869 , n364868 );
buf ( n364870 , n364869 );
buf ( n44706 , n364870 );
nand ( n44707 , n364864 , n44706 );
buf ( n364873 , n44707 );
buf ( n364874 , n364873 );
nand ( n44710 , n364863 , n364874 );
buf ( n364876 , n44710 );
buf ( n364877 , n364876 );
not ( n364878 , n364877 );
buf ( n364879 , n364878 );
or ( n44715 , n364852 , n364879 );
buf ( n364881 , n30912 );
not ( n44717 , n361574 );
buf ( n364883 , n44717 );
and ( n364884 , n364881 , n364883 );
not ( n364885 , n364881 );
buf ( n364886 , n361531 );
and ( n364887 , n364885 , n364886 );
nor ( n364888 , n364884 , n364887 );
buf ( n364889 , n364888 );
not ( n364890 , n364889 );
nand ( n364891 , n364890 , n361625 );
nand ( n44727 , n44715 , n364891 );
and ( n44728 , n364847 , n44727 );
and ( n364894 , n44629 , n44681 );
or ( n364895 , n44728 , n364894 );
not ( n44731 , n364895 );
buf ( n364897 , n359916 );
not ( n364898 , n364897 );
buf ( n364899 , n364898 );
not ( n364900 , n352268 );
not ( n364901 , n364900 );
not ( n44737 , n364901 );
buf ( n364903 , n42455 );
not ( n44739 , n364903 );
buf ( n364905 , n44739 );
and ( n364906 , n44737 , n364905 );
not ( n364907 , n44737 );
buf ( n44743 , n359896 );
not ( n364909 , n44743 );
and ( n364910 , n364907 , n364909 );
nor ( n44746 , n364906 , n364910 );
or ( n364912 , n364899 , n44746 );
buf ( n364913 , n351160 );
not ( n44749 , n364913 );
buf ( n364915 , n44749 );
buf ( n364916 , n364915 );
buf ( n364917 , n359944 );
not ( n364918 , n364917 );
buf ( n364919 , n364918 );
buf ( n364920 , n364919 );
not ( n364921 , n364920 );
buf ( n364922 , n364921 );
buf ( n364923 , n364922 );
and ( n364924 , n364916 , n364923 );
not ( n364925 , n364916 );
buf ( n364926 , n41623 );
and ( n364927 , n364925 , n364926 );
nor ( n44763 , n364924 , n364927 );
buf ( n364929 , n44763 );
or ( n364930 , n364929 , n359996 );
nand ( n44766 , n364912 , n364930 );
not ( n44767 , n44766 );
buf ( n364933 , n43261 );
not ( n364934 , n364933 );
not ( n44770 , n22772 );
not ( n364936 , n363317 );
or ( n364937 , n44770 , n364936 );
buf ( n364938 , n361802 );
buf ( n364939 , n363444 );
nand ( n44775 , n364938 , n364939 );
buf ( n44776 , n44775 );
nand ( n364942 , n364937 , n44776 );
buf ( n364943 , n364942 );
not ( n44779 , n364943 );
or ( n364945 , n364934 , n44779 );
buf ( n364946 , n342719 );
not ( n364947 , n364946 );
not ( n44783 , n41607 );
buf ( n364949 , n44783 );
not ( n364950 , n364949 );
or ( n44786 , n364947 , n364950 );
buf ( n364952 , n41607 );
not ( n364953 , n342719 );
buf ( n364954 , n364953 );
nand ( n44790 , n364952 , n364954 );
buf ( n364956 , n44790 );
buf ( n364957 , n364956 );
nand ( n364958 , n44786 , n364957 );
buf ( n364959 , n364958 );
buf ( n364960 , n364959 );
not ( n44796 , n43274 );
buf ( n364962 , n44796 );
nand ( n44798 , n364960 , n364962 );
buf ( n364964 , n44798 );
buf ( n364965 , n364964 );
nand ( n364966 , n364945 , n364965 );
buf ( n364967 , n364966 );
not ( n364968 , n364967 );
nand ( n44804 , n44767 , n364968 );
not ( n44805 , n44804 );
or ( n364971 , n44731 , n44805 );
nand ( n364972 , n44766 , n364967 );
nand ( n44808 , n364971 , n364972 );
not ( n364974 , n44808 );
buf ( n364975 , n22556 );
buf ( n364976 , n364975 );
not ( n364977 , n364976 );
buf ( n364978 , n364977 );
buf ( n364979 , n364978 );
not ( n44815 , n364979 );
buf ( n364981 , n44815 );
buf ( n364982 , n364981 );
buf ( n44818 , n364982 );
buf ( n44819 , n44818 );
buf ( n364985 , n44819 );
not ( n44821 , n364985 );
not ( n364987 , n359778 );
buf ( n364988 , n364987 );
not ( n44824 , n364988 );
or ( n44825 , n44821 , n44824 );
buf ( n44826 , n359778 );
buf ( n364992 , n44819 );
not ( n44828 , n364992 );
buf ( n364994 , n44828 );
buf ( n364995 , n364994 );
buf ( n364996 , n364995 );
buf ( n364997 , n364996 );
buf ( n364998 , n364997 );
nand ( n44834 , n44826 , n364998 );
buf ( n365000 , n44834 );
buf ( n365001 , n365000 );
nand ( n44837 , n44825 , n365001 );
buf ( n365003 , n44837 );
buf ( n365004 , n365003 );
not ( n365005 , n365004 );
not ( n44841 , n342879 );
not ( n365007 , n22899 );
or ( n44843 , n44841 , n365007 );
nand ( n44844 , n342846 , n342878 );
nand ( n365010 , n44843 , n44844 );
not ( n365011 , n365010 );
buf ( n365012 , n22556 );
not ( n365013 , n365012 );
buf ( n365014 , n22899 );
nand ( n44850 , n365013 , n365014 );
buf ( n44851 , n44850 );
nand ( n365017 , n22556 , n342846 );
nand ( n44853 , n365011 , n44851 , n365017 );
buf ( n365019 , n44853 );
not ( n365020 , n365019 );
buf ( n365021 , n365020 );
buf ( n365022 , n365021 );
buf ( n365023 , n365022 );
buf ( n365024 , n365023 );
buf ( n365025 , n365024 );
not ( n44861 , n365025 );
buf ( n44862 , n44861 );
buf ( n365028 , n44862 );
not ( n44864 , n365028 );
buf ( n365030 , n44864 );
buf ( n44866 , n365030 );
buf ( n365032 , n44866 );
buf ( n365033 , n365032 );
buf ( n365034 , n365033 );
not ( n365035 , n365034 );
buf ( n365036 , n365035 );
buf ( n365037 , n365036 );
nor ( n365038 , n365005 , n365037 );
buf ( n365039 , n365038 );
not ( n365040 , n365039 );
buf ( n365041 , n342965 );
buf ( n365042 , n365041 );
not ( n365043 , n365042 );
buf ( n365044 , n359147 );
not ( n44880 , n365044 );
or ( n44881 , n365043 , n44880 );
nand ( n365047 , n359136 , n39046 );
buf ( n365048 , n365047 );
not ( n44884 , n365048 );
buf ( n365050 , n365041 );
not ( n365051 , n365050 );
buf ( n365052 , n365051 );
buf ( n365053 , n365052 );
nand ( n44889 , n44884 , n365053 );
buf ( n365055 , n44889 );
buf ( n365056 , n365055 );
nand ( n44892 , n44881 , n365056 );
buf ( n365058 , n44892 );
buf ( n365059 , n365058 );
buf ( n365060 , n22499 );
not ( n365061 , n365060 );
buf ( n365062 , n365061 );
and ( n44898 , n342965 , n365062 );
not ( n44899 , n342965 );
and ( n365065 , n44899 , n342445 );
or ( n365066 , n44898 , n365065 );
not ( n44902 , n365062 );
not ( n365068 , n23037 );
or ( n44904 , n44902 , n365068 );
buf ( n365070 , n22499 );
not ( n44906 , n23034 );
buf ( n365072 , n44906 );
nand ( n44908 , n365070 , n365072 );
buf ( n365074 , n44908 );
nand ( n365075 , n44904 , n365074 );
not ( n365076 , n365075 );
nand ( n44912 , n365066 , n365076 );
buf ( n44913 , n44912 );
buf ( n44914 , n44913 );
buf ( n44915 , n365075 );
buf ( n365081 , n44915 );
not ( n365082 , n365081 );
buf ( n365083 , n365082 );
buf ( n365084 , n365083 );
nand ( n365085 , n44914 , n365084 );
buf ( n365086 , n365085 );
buf ( n365087 , n365086 );
and ( n44923 , n365059 , n365087 );
buf ( n365089 , n44923 );
not ( n44925 , n359755 );
not ( n44926 , n44925 );
buf ( n365092 , n44926 );
not ( n365093 , n365092 );
buf ( n365094 , n364994 );
not ( n44930 , n365094 );
and ( n365096 , n365093 , n44930 );
buf ( n365097 , n44926 );
buf ( n365098 , n364997 );
and ( n365099 , n365097 , n365098 );
nor ( n365100 , n365096 , n365099 );
buf ( n365101 , n365100 );
not ( n44937 , n365101 );
buf ( n365103 , n365010 );
buf ( n365104 , n365103 );
buf ( n365105 , n365104 );
buf ( n365106 , n365105 );
buf ( n365107 , n365106 );
buf ( n365108 , n365107 );
buf ( n44944 , n365108 );
not ( n44945 , n44944 );
buf ( n44946 , n44945 );
buf ( n365112 , n44946 );
buf ( n365113 , n365112 );
not ( n365114 , n365113 );
buf ( n365115 , n365114 );
buf ( n365116 , n365115 );
buf ( n365117 , n365116 );
buf ( n365118 , n365117 );
nand ( n44954 , n44937 , n365118 );
nand ( n365120 , n365040 , n365089 , n44954 );
not ( n44956 , n365120 );
or ( n44957 , n364974 , n44956 );
not ( n365123 , n365089 );
not ( n365124 , n365039 );
nand ( n44960 , n365124 , n44954 );
nand ( n365126 , n365123 , n44960 );
nand ( n365127 , n44957 , n365126 );
and ( n44963 , n22961 , n362179 );
not ( n365129 , n22961 );
and ( n365130 , n365129 , n40899 );
or ( n44966 , n44963 , n365130 );
not ( n365132 , n44966 );
not ( n365133 , n365132 );
buf ( n365134 , n342965 );
not ( n365135 , n365134 );
buf ( n365136 , n365135 );
and ( n365137 , n342931 , n365136 );
not ( n365138 , n342931 );
and ( n365139 , n365138 , n342965 );
or ( n44970 , n365137 , n365139 );
buf ( n365141 , n44970 );
not ( n365142 , n365141 );
buf ( n365143 , n365142 );
buf ( n365144 , n365143 );
buf ( n365145 , n365144 );
buf ( n365146 , n365145 );
buf ( n365147 , n365146 );
not ( n365148 , n365147 );
buf ( n365149 , n365148 );
buf ( n365150 , n365149 );
buf ( n365151 , n365150 );
buf ( n365152 , n365151 );
buf ( n365153 , n365152 );
not ( n365154 , n365153 );
buf ( n365155 , n365154 );
not ( n44986 , n365155 );
and ( n365157 , n365133 , n44986 );
not ( n44988 , n22959 );
not ( n365159 , n363866 );
or ( n365160 , n44988 , n365159 );
and ( n44991 , n360097 , n360105 );
not ( n365162 , n360097 );
and ( n365163 , n365162 , n360108 );
or ( n365164 , n44991 , n365163 );
buf ( n365165 , n365164 );
not ( n365166 , n365165 );
buf ( n365167 , n365166 );
buf ( n365168 , n365167 );
buf ( n365169 , n365168 );
buf ( n365170 , n365169 );
buf ( n365171 , n365170 );
buf ( n365172 , n342909 );
nand ( n365173 , n365171 , n365172 );
buf ( n365174 , n365173 );
nand ( n45005 , n365160 , n365174 );
buf ( n365176 , n45005 );
not ( n365177 , n365176 );
xor ( n45008 , n342934 , n22954 );
and ( n365179 , n45008 , n365143 );
not ( n45010 , n365179 );
not ( n365181 , n45010 );
buf ( n45012 , n365181 );
buf ( n365183 , n45012 );
buf ( n45014 , n365183 );
buf ( n45015 , n45014 );
buf ( n365186 , n45015 );
buf ( n365187 , n365186 );
buf ( n45018 , n365187 );
buf ( n365189 , n45018 );
not ( n365190 , n365189 );
buf ( n45021 , n365190 );
buf ( n365192 , n45021 );
buf ( n365193 , n365192 );
nor ( n45024 , n365177 , n365193 );
buf ( n365195 , n45024 );
nor ( n365196 , n365157 , n365195 );
buf ( n365197 , n365196 );
not ( n45028 , n365197 );
buf ( n45029 , n45028 );
buf ( n365200 , n45029 );
not ( n45031 , n365200 );
not ( n365202 , n342881 );
not ( n365203 , n365202 );
not ( n45034 , n40943 );
or ( n365205 , n365203 , n45034 );
not ( n365206 , n39830 );
nand ( n365207 , n365206 , n342881 );
nand ( n365208 , n365205 , n365207 );
not ( n45039 , n342475 );
not ( n365210 , n342879 );
or ( n365211 , n45039 , n365210 );
not ( n45042 , n342475 );
xor ( n365213 , n342829 , n342867 );
not ( n365214 , n365213 );
and ( n45045 , n45042 , n365214 );
or ( n45046 , n342475 , n22956 );
not ( n365217 , n22525 );
not ( n365218 , n22529 );
or ( n45049 , n365217 , n365218 );
not ( n45050 , n22954 );
nand ( n45051 , n45049 , n45050 );
nand ( n45052 , n45046 , n45051 );
nor ( n45053 , n45045 , n45052 );
nand ( n365224 , n365211 , n45053 );
not ( n45055 , n365224 );
buf ( n365226 , n45055 );
not ( n365227 , n365226 );
not ( n45058 , n365227 );
and ( n365229 , n365208 , n45058 );
not ( n45060 , n365202 );
not ( n45061 , n45060 );
not ( n45062 , n41907 );
or ( n45063 , n45061 , n45062 );
buf ( n365234 , n39867 );
not ( n45065 , n342881 );
buf ( n365236 , n45065 );
nand ( n365237 , n365234 , n365236 );
buf ( n365238 , n365237 );
nand ( n365239 , n45063 , n365238 );
buf ( n365240 , n45052 );
buf ( n45071 , n365240 );
buf ( n365242 , n45071 );
buf ( n45073 , n365242 );
buf ( n45074 , n45073 );
buf ( n45075 , n45074 );
and ( n45076 , n365239 , n45075 );
nor ( n45077 , n365229 , n45076 );
buf ( n365248 , n45077 );
not ( n45079 , n365248 );
buf ( n365250 , n45079 );
buf ( n365251 , n365250 );
not ( n365252 , n365251 );
or ( n45083 , n45031 , n365252 );
not ( n365254 , n45077 );
not ( n45085 , n365196 );
or ( n365256 , n365254 , n45085 );
buf ( n365257 , n352212 );
not ( n365258 , n365257 );
buf ( n365259 , n365258 );
buf ( n365260 , n365259 );
not ( n45091 , n360989 );
buf ( n45092 , n45091 );
buf ( n365263 , n45092 );
and ( n365264 , n365260 , n365263 );
not ( n45095 , n365260 );
not ( n365266 , n360989 );
not ( n365267 , n365266 );
buf ( n365268 , n365267 );
and ( n365269 , n45095 , n365268 );
nor ( n365270 , n365264 , n365269 );
buf ( n365271 , n365270 );
buf ( n365272 , n365271 );
not ( n45103 , n365272 );
buf ( n365274 , n45103 );
buf ( n365275 , n365274 );
not ( n365276 , n365275 );
buf ( n365277 , n361013 );
buf ( n365278 , n365277 );
buf ( n365279 , n365278 );
buf ( n365280 , n365279 );
not ( n365281 , n365280 );
or ( n365282 , n365276 , n365281 );
buf ( n45113 , n352192 );
buf ( n365284 , n45113 );
not ( n365285 , n365284 );
buf ( n45116 , n40891 );
buf ( n365287 , n45116 );
not ( n45118 , n365287 );
or ( n365289 , n365285 , n45118 );
not ( n365290 , n360532 );
buf ( n365291 , n365290 );
not ( n45122 , n365291 );
buf ( n365293 , n45122 );
buf ( n365294 , n365293 );
not ( n45125 , n352192 );
buf ( n365296 , n45125 );
nand ( n365297 , n365294 , n365296 );
buf ( n365298 , n365297 );
buf ( n365299 , n365298 );
nand ( n365300 , n365289 , n365299 );
buf ( n365301 , n365300 );
buf ( n365302 , n365301 );
not ( n365303 , n361011 );
buf ( n365304 , n365303 );
nand ( n365305 , n365302 , n365304 );
buf ( n365306 , n365305 );
buf ( n365307 , n365306 );
nand ( n365308 , n365282 , n365307 );
buf ( n365309 , n365308 );
buf ( n365310 , n365309 );
not ( n365311 , n361975 );
not ( n365312 , n365311 );
not ( n45143 , n365312 );
not ( n365314 , n45143 );
not ( n365315 , n364790 );
or ( n45146 , n365314 , n365315 );
buf ( n365317 , n364760 );
buf ( n365318 , n365317 );
buf ( n365319 , n365318 );
buf ( n365320 , n365319 );
not ( n365321 , n365320 );
not ( n45152 , n30911 );
buf ( n365323 , n45152 );
not ( n45154 , n365323 );
or ( n365325 , n365321 , n45154 );
buf ( n365326 , n361911 );
not ( n45157 , n365326 );
not ( n365328 , n30911 );
not ( n365329 , n365328 );
buf ( n365330 , n365329 );
nand ( n365331 , n45157 , n365330 );
buf ( n365332 , n365331 );
buf ( n365333 , n365332 );
nand ( n365334 , n365325 , n365333 );
buf ( n365335 , n365334 );
nand ( n45166 , n365335 , n44591 );
nand ( n365337 , n45146 , n45166 );
buf ( n365338 , n365337 );
buf ( n45169 , n365338 );
buf ( n45170 , n45169 );
buf ( n365341 , n45170 );
xor ( n45172 , n365310 , n365341 );
not ( n365343 , n39217 );
not ( n365344 , n31231 );
buf ( n365345 , n365344 );
not ( n45176 , n365345 );
buf ( n45177 , n45176 );
buf ( n365348 , n45177 );
not ( n45179 , n365348 );
buf ( n365350 , n361851 );
not ( n45181 , n365350 );
or ( n365352 , n45179 , n45181 );
not ( n365353 , n355579 );
buf ( n365354 , n365353 );
buf ( n365355 , n45177 );
not ( n45186 , n365355 );
buf ( n365357 , n45186 );
buf ( n365358 , n365357 );
nand ( n45189 , n365354 , n365358 );
buf ( n365360 , n45189 );
buf ( n365361 , n365360 );
nand ( n365362 , n365352 , n365361 );
buf ( n365363 , n365362 );
not ( n45194 , n365363 );
or ( n45195 , n365343 , n45194 );
not ( n45196 , n351229 );
buf ( n365367 , n355578 );
not ( n365368 , n365367 );
not ( n45199 , n365368 );
or ( n45200 , n45196 , n45199 );
or ( n45201 , n365368 , n351229 );
nand ( n365372 , n45200 , n45201 );
not ( n365373 , n365372 );
not ( n45204 , n39207 );
nand ( n365375 , n365373 , n45204 );
nand ( n365376 , n45195 , n365375 );
buf ( n365377 , n365376 );
and ( n45208 , n45172 , n365377 );
and ( n45209 , n365310 , n365341 );
or ( n45210 , n45208 , n45209 );
buf ( n365381 , n45210 );
buf ( n365382 , n351062 );
not ( n45213 , n365382 );
buf ( n365384 , n45213 );
buf ( n365385 , n365384 );
buf ( n365386 , n365385 );
buf ( n365387 , n365386 );
buf ( n365388 , n365387 );
not ( n45219 , n365388 );
buf ( n365390 , n45219 );
buf ( n365391 , n365390 );
buf ( n365392 , n365391 );
buf ( n365393 , n365392 );
buf ( n365394 , n365393 );
not ( n365395 , n365394 );
buf ( n365396 , n361631 );
not ( n365397 , n365396 );
or ( n365398 , n365395 , n365397 );
buf ( n365399 , n359800 );
buf ( n45230 , n365399 );
buf ( n45231 , n45230 );
buf ( n365402 , n45231 );
not ( n45233 , n365402 );
buf ( n45234 , n45233 );
buf ( n365405 , n45234 );
buf ( n365406 , n365393 );
not ( n45237 , n365406 );
buf ( n365408 , n45237 );
buf ( n45239 , n365408 );
nand ( n45240 , n365405 , n45239 );
buf ( n45241 , n45240 );
buf ( n45242 , n45241 );
nand ( n45243 , n365398 , n45242 );
buf ( n45244 , n45243 );
buf ( n365415 , n45244 );
not ( n365416 , n365415 );
buf ( n365417 , n363038 );
not ( n365418 , n365417 );
or ( n365419 , n365416 , n365418 );
buf ( n365420 , n362521 );
buf ( n365421 , n39621 );
not ( n365422 , n351345 );
buf ( n365423 , n365422 );
and ( n365424 , n365421 , n365423 );
not ( n45250 , n365421 );
buf ( n365426 , n365422 );
not ( n365427 , n365426 );
buf ( n365428 , n365427 );
buf ( n365429 , n365428 );
and ( n365430 , n45250 , n365429 );
or ( n365431 , n365424 , n365430 );
buf ( n365432 , n365431 );
buf ( n365433 , n365432 );
nand ( n365434 , n365420 , n365433 );
buf ( n365435 , n365434 );
buf ( n365436 , n365435 );
nand ( n365437 , n365419 , n365436 );
buf ( n365438 , n365437 );
not ( n365439 , n365438 );
buf ( n365440 , n32202 );
buf ( n45266 , n365440 );
not ( n45267 , n45266 );
buf ( n45268 , n362452 );
not ( n45269 , n45268 );
buf ( n45270 , n45269 );
buf ( n365446 , n45270 );
not ( n365447 , n365446 );
or ( n45273 , n45267 , n365447 );
buf ( n365449 , n362452 );
buf ( n45275 , n365440 );
not ( n365451 , n45275 );
buf ( n365452 , n365451 );
buf ( n365453 , n365452 );
nand ( n365454 , n365449 , n365453 );
buf ( n365455 , n365454 );
buf ( n365456 , n365455 );
nand ( n365457 , n45273 , n365456 );
buf ( n365458 , n365457 );
buf ( n45284 , n365458 );
not ( n45285 , n45284 );
buf ( n365461 , n40475 );
not ( n45287 , n365461 );
or ( n365463 , n45285 , n45287 );
not ( n365464 , n351294 );
not ( n45290 , n365464 );
buf ( n365466 , n360589 );
buf ( n365467 , n365466 );
buf ( n365468 , n365467 );
buf ( n365469 , n365468 );
not ( n365470 , n365469 );
buf ( n365471 , n365470 );
not ( n45297 , n365471 );
or ( n365473 , n45290 , n45297 );
not ( n365474 , n31260 );
not ( n45300 , n365474 );
nand ( n365476 , n45270 , n45300 );
nand ( n365477 , n365473 , n365476 );
nand ( n45303 , n365477 , n360574 );
buf ( n365479 , n45303 );
nand ( n365480 , n365463 , n365479 );
buf ( n365481 , n365480 );
buf ( n365482 , n365481 );
not ( n365483 , n365482 );
buf ( n365484 , n360051 );
not ( n365485 , n365484 );
buf ( n365486 , n365485 );
not ( n45312 , n365486 );
buf ( n365488 , n351195 );
buf ( n365489 , n365488 );
buf ( n365490 , n365489 );
buf ( n365491 , n365490 );
not ( n45317 , n365491 );
buf ( n365493 , n360065 );
buf ( n45319 , n365493 );
buf ( n365495 , n45319 );
buf ( n365496 , n365495 );
not ( n45322 , n365496 );
buf ( n365498 , n45322 );
buf ( n365499 , n365498 );
not ( n45325 , n365499 );
or ( n365501 , n45317 , n45325 );
buf ( n365502 , n360154 );
buf ( n365503 , n365502 );
buf ( n365504 , n365503 );
buf ( n365505 , n365504 );
not ( n45331 , n365505 );
buf ( n365507 , n45331 );
buf ( n45333 , n365507 );
buf ( n365509 , n365490 );
not ( n45335 , n365509 );
buf ( n45336 , n45335 );
buf ( n365512 , n45336 );
nand ( n45338 , n45333 , n365512 );
buf ( n45339 , n45338 );
buf ( n365515 , n45339 );
nand ( n45341 , n365501 , n365515 );
buf ( n365517 , n45341 );
not ( n365518 , n365517 );
or ( n365519 , n45312 , n365518 );
not ( n45345 , n360165 );
buf ( n365521 , n351160 );
not ( n365522 , n365521 );
buf ( n365523 , n363122 );
not ( n365524 , n365523 );
or ( n365525 , n365522 , n365524 );
buf ( n365526 , n363116 );
not ( n45352 , n365526 );
buf ( n365528 , n45352 );
buf ( n365529 , n365528 );
buf ( n365530 , n364915 );
nand ( n45356 , n365529 , n365530 );
buf ( n365532 , n45356 );
buf ( n365533 , n365532 );
nand ( n365534 , n365525 , n365533 );
buf ( n365535 , n365534 );
nand ( n365536 , n45345 , n365535 );
nand ( n45362 , n365519 , n365536 );
buf ( n365538 , n45362 );
not ( n45364 , n365538 );
buf ( n365540 , n45364 );
buf ( n365541 , n365540 );
nand ( n365542 , n365483 , n365541 );
buf ( n365543 , n365542 );
not ( n45369 , n365543 );
or ( n45370 , n365439 , n45369 );
nand ( n45371 , n365481 , n45362 );
nand ( n45372 , n45370 , n45371 );
or ( n45373 , n365381 , n45372 );
buf ( n45374 , n365279 );
not ( n45375 , n45374 );
buf ( n45376 , n45375 );
buf ( n365552 , n45376 );
buf ( n365553 , n365301 );
not ( n45379 , n365553 );
buf ( n45380 , n45379 );
buf ( n365556 , n45380 );
or ( n365557 , n365552 , n365556 );
not ( n365558 , n361011 );
not ( n45384 , n365558 );
buf ( n365560 , n45384 );
not ( n365561 , n351318 );
buf ( n365562 , n365561 );
not ( n365563 , n365562 );
buf ( n365564 , n365267 );
not ( n365565 , n365564 );
or ( n45391 , n365563 , n365565 );
buf ( n365567 , n365290 );
not ( n45393 , n365567 );
buf ( n365569 , n45393 );
buf ( n365570 , n365569 );
buf ( n365571 , n351318 );
nand ( n45397 , n365570 , n365571 );
buf ( n365573 , n45397 );
buf ( n365574 , n365573 );
nand ( n45400 , n45391 , n365574 );
buf ( n45401 , n45400 );
buf ( n365577 , n45401 );
not ( n45403 , n365577 );
buf ( n45404 , n45403 );
buf ( n365580 , n45404 );
or ( n45406 , n365560 , n365580 );
nand ( n365582 , n365557 , n45406 );
buf ( n365583 , n365582 );
buf ( n365584 , n361603 );
not ( n45410 , n365584 );
buf ( n365586 , n364889 );
not ( n45412 , n365586 );
and ( n365588 , n45410 , n45412 );
not ( n45414 , n44717 );
and ( n365590 , n364777 , n45414 );
not ( n365591 , n364777 );
and ( n45417 , n365591 , n361534 );
nor ( n365593 , n365590 , n45417 );
buf ( n365594 , n365593 );
buf ( n365595 , n41482 );
nor ( n365596 , n365594 , n365595 );
buf ( n365597 , n365596 );
buf ( n365598 , n365597 );
nor ( n365599 , n365588 , n365598 );
buf ( n365600 , n365599 );
and ( n365601 , n365583 , n365600 );
not ( n365602 , n365583 );
buf ( n365603 , n365600 );
not ( n45429 , n365603 );
buf ( n365605 , n45429 );
and ( n365606 , n365602 , n365605 );
or ( n365607 , n365601 , n365606 );
buf ( n365608 , n365607 );
buf ( n365609 , n364842 );
not ( n365610 , n365609 );
buf ( n365611 , n362021 );
not ( n45437 , n365611 );
buf ( n45438 , n45437 );
buf ( n365614 , n45438 );
not ( n45440 , n365614 );
or ( n45441 , n365610 , n45440 );
buf ( n365617 , n41869 );
buf ( n365618 , n365617 );
buf ( n365619 , n365618 );
buf ( n365620 , n365619 );
not ( n365621 , n365620 );
buf ( n365622 , n365621 );
buf ( n365623 , n365622 );
buf ( n365624 , n364858 );
not ( n45450 , n365624 );
buf ( n365626 , n361009 );
buf ( n365627 , n365626 );
not ( n45453 , n365627 );
or ( n45454 , n45450 , n45453 );
not ( n45455 , n361009 );
buf ( n365631 , n45455 );
buf ( n45457 , n364858 );
not ( n45458 , n45457 );
buf ( n45459 , n45458 );
buf ( n365635 , n45459 );
nand ( n365636 , n365631 , n365635 );
buf ( n365637 , n365636 );
buf ( n365638 , n365637 );
nand ( n365639 , n45454 , n365638 );
buf ( n365640 , n365639 );
buf ( n365641 , n365640 );
nand ( n365642 , n365623 , n365641 );
buf ( n365643 , n365642 );
buf ( n365644 , n365643 );
nand ( n365645 , n45441 , n365644 );
buf ( n365646 , n365645 );
buf ( n365647 , n365646 );
xor ( n45473 , n365608 , n365647 );
buf ( n365649 , n45473 );
nand ( n365650 , n45373 , n365649 );
nand ( n365651 , n45372 , n365381 );
nand ( n45477 , n365650 , n365651 );
nand ( n45478 , n365256 , n45477 );
buf ( n365654 , n45478 );
nand ( n365655 , n45083 , n365654 );
buf ( n365656 , n365655 );
xor ( n365657 , n365127 , n365656 );
not ( n45483 , n22556 );
and ( n45484 , n45483 , n342528 );
not ( n45485 , n45483 );
buf ( n365661 , n342528 );
not ( n45487 , n365661 );
buf ( n365663 , n45487 );
and ( n45489 , n45485 , n365663 );
nor ( n365665 , n45484 , n45489 );
not ( n45491 , n365665 );
buf ( n45492 , n45491 );
buf ( n45493 , n45492 );
not ( n45494 , n45493 );
not ( n365670 , n342564 );
buf ( n365671 , n365670 );
buf ( n45497 , n365671 );
buf ( n365673 , n45497 );
buf ( n365674 , n365673 );
not ( n365675 , n365674 );
buf ( n365676 , n365675 );
buf ( n365677 , n365676 );
not ( n45503 , n365677 );
buf ( n45504 , n359778 );
not ( n365680 , n45504 );
buf ( n365681 , n365680 );
buf ( n365682 , n365681 );
not ( n45508 , n365682 );
or ( n365684 , n45503 , n45508 );
buf ( n45510 , n359778 );
buf ( n365686 , n365673 );
nand ( n45512 , n45510 , n365686 );
buf ( n365688 , n45512 );
buf ( n365689 , n365688 );
nand ( n45515 , n365684 , n365689 );
buf ( n365691 , n45515 );
buf ( n365692 , n365691 );
not ( n365693 , n365692 );
or ( n45519 , n45494 , n365693 );
not ( n45520 , n365676 );
not ( n45521 , n360308 );
or ( n45522 , n45520 , n45521 );
not ( n45523 , n40199 );
buf ( n365699 , n45523 );
not ( n365700 , n365699 );
buf ( n45526 , n365673 );
nand ( n45527 , n365700 , n45526 );
buf ( n45528 , n45527 );
nand ( n365704 , n45522 , n45528 );
buf ( n365705 , n365704 );
buf ( n365706 , n342564 );
not ( n365707 , n365706 );
buf ( n365708 , n365663 );
nand ( n45534 , n365707 , n365708 );
buf ( n365710 , n45534 );
buf ( n365711 , n365710 );
buf ( n365712 , n342564 );
buf ( n365713 , n342528 );
nand ( n365714 , n365712 , n365713 );
buf ( n365715 , n365714 );
buf ( n365716 , n365715 );
buf ( n365717 , n365665 );
nand ( n45543 , n365711 , n365716 , n365717 );
buf ( n45544 , n45543 );
buf ( n365720 , n45544 );
buf ( n45546 , n365720 );
buf ( n365722 , n45546 );
buf ( n365723 , n365722 );
not ( n45549 , n365723 );
buf ( n365725 , n45549 );
buf ( n365726 , n365725 );
buf ( n45552 , n365726 );
buf ( n45553 , n45552 );
buf ( n365729 , n45553 );
nand ( n45555 , n365705 , n365729 );
buf ( n45556 , n45555 );
buf ( n365732 , n45556 );
nand ( n45558 , n45519 , n365732 );
buf ( n365734 , n45558 );
buf ( n365735 , n365734 );
not ( n365736 , n365735 );
buf ( n365737 , n41607 );
not ( n45563 , n365737 );
buf ( n365739 , n362435 );
not ( n45565 , n365739 );
and ( n45566 , n45563 , n45565 );
buf ( n365742 , n362435 );
buf ( n365743 , n41607 );
and ( n45569 , n365742 , n365743 );
nor ( n45570 , n45566 , n45569 );
buf ( n365746 , n45570 );
buf ( n365747 , n365746 );
not ( n45573 , n365747 );
buf ( n365749 , n45573 );
buf ( n365750 , n365749 );
buf ( n365751 , n42242 );
and ( n365752 , n365750 , n365751 );
buf ( n365753 , n362426 );
not ( n45579 , n365753 );
buf ( n365755 , n361661 );
buf ( n365756 , n365755 );
buf ( n365757 , n365756 );
buf ( n365758 , n365757 );
not ( n365759 , n365758 );
buf ( n365760 , n365759 );
buf ( n45586 , n365760 );
not ( n45587 , n45586 );
or ( n45588 , n45579 , n45587 );
buf ( n45589 , n361667 );
buf ( n365765 , n342335 );
not ( n45591 , n365765 );
buf ( n45592 , n45591 );
buf ( n365768 , n45592 );
buf ( n45594 , n365768 );
buf ( n45595 , n45594 );
buf ( n365771 , n45595 );
not ( n45597 , n365771 );
buf ( n365773 , n45597 );
buf ( n365774 , n365773 );
nand ( n365775 , n45589 , n365774 );
buf ( n365776 , n365775 );
buf ( n365777 , n365776 );
nand ( n365778 , n45588 , n365777 );
buf ( n365779 , n365778 );
buf ( n365780 , n365779 );
not ( n365781 , n365780 );
buf ( n365782 , n42266 );
nor ( n45608 , n365781 , n365782 );
buf ( n45609 , n45608 );
buf ( n365785 , n45609 );
nor ( n45611 , n365752 , n365785 );
buf ( n365787 , n45611 );
buf ( n365788 , n365787 );
not ( n45614 , n365788 );
buf ( n45615 , n39775 );
buf ( n365791 , n359910 );
nand ( n365792 , n45615 , n365791 );
buf ( n365793 , n365792 );
buf ( n365794 , n365793 );
not ( n45620 , n365794 );
buf ( n365796 , n364929 );
not ( n365797 , n365796 );
and ( n45623 , n45620 , n365797 );
buf ( n365799 , n39775 );
buf ( n365800 , n365799 );
buf ( n365801 , n365800 );
buf ( n365802 , n365801 );
buf ( n365803 , n45336 );
buf ( n365804 , n364922 );
and ( n365805 , n365803 , n365804 );
not ( n45631 , n365803 );
buf ( n365807 , n41623 );
and ( n45633 , n45631 , n365807 );
nor ( n365809 , n365805 , n45633 );
buf ( n365810 , n365809 );
buf ( n365811 , n365810 );
nor ( n45637 , n365802 , n365811 );
buf ( n365813 , n45637 );
buf ( n365814 , n365813 );
nor ( n45640 , n45623 , n365814 );
buf ( n365816 , n45640 );
buf ( n365817 , n365816 );
not ( n365818 , n365817 );
or ( n45644 , n45614 , n365818 );
not ( n45645 , n365646 );
nand ( n365821 , n45645 , n365600 );
not ( n45647 , n365821 );
not ( n365823 , n365583 );
or ( n45649 , n45647 , n365823 );
buf ( n365825 , n365605 );
buf ( n365826 , n365646 );
nand ( n45652 , n365825 , n365826 );
buf ( n365828 , n45652 );
nand ( n365829 , n45649 , n365828 );
buf ( n365830 , n365829 );
nand ( n45656 , n45644 , n365830 );
buf ( n45657 , n45656 );
buf ( n365833 , n45657 );
buf ( n365834 , n365816 );
not ( n365835 , n365834 );
buf ( n365836 , n365835 );
buf ( n365837 , n365836 );
buf ( n365838 , n365787 );
not ( n365839 , n365838 );
buf ( n365840 , n365839 );
buf ( n365841 , n365840 );
nand ( n365842 , n365837 , n365841 );
buf ( n365843 , n365842 );
buf ( n365844 , n365843 );
and ( n45670 , n365833 , n365844 );
buf ( n365846 , n45670 );
buf ( n365847 , n365846 );
not ( n365848 , n365847 );
or ( n45674 , n365736 , n365848 );
buf ( n365850 , n365734 );
buf ( n365851 , n365846 );
or ( n365852 , n365850 , n365851 );
nand ( n365853 , n45674 , n365852 );
buf ( n365854 , n365853 );
buf ( n365855 , n365854 );
buf ( n365856 , n45075 );
not ( n365857 , n365856 );
buf ( n365858 , n342881 );
not ( n365859 , n365858 );
buf ( n365860 , n363866 );
not ( n365861 , n365860 );
or ( n45687 , n365859 , n365861 );
buf ( n365863 , n365170 );
buf ( n45689 , n365202 );
nand ( n45690 , n365863 , n45689 );
buf ( n45691 , n45690 );
buf ( n365867 , n45691 );
nand ( n45693 , n45687 , n365867 );
buf ( n45694 , n45693 );
buf ( n365870 , n45694 );
not ( n45696 , n365870 );
or ( n365872 , n365857 , n45696 );
nand ( n45698 , n365239 , n45058 );
buf ( n365874 , n45698 );
nand ( n45700 , n365872 , n365874 );
buf ( n365876 , n45700 );
buf ( n45702 , n365876 );
buf ( n365878 , n45702 );
and ( n45704 , n365855 , n365878 );
not ( n45705 , n365855 );
not ( n45706 , n45702 );
buf ( n365882 , n45706 );
and ( n45708 , n45705 , n365882 );
nor ( n45709 , n45704 , n45708 );
buf ( n365885 , n45709 );
xor ( n45711 , n365657 , n365885 );
buf ( n365887 , n45711 );
not ( n45713 , n43261 );
buf ( n365889 , n22772 );
not ( n45715 , n365889 );
buf ( n365891 , n362130 );
not ( n45717 , n365891 );
buf ( n45718 , n45717 );
buf ( n365894 , n45718 );
not ( n365895 , n365894 );
or ( n365896 , n45715 , n365895 );
buf ( n365897 , n362133 );
buf ( n365898 , n363444 );
nand ( n365899 , n365897 , n365898 );
buf ( n365900 , n365899 );
buf ( n365901 , n365900 );
nand ( n365902 , n365896 , n365901 );
buf ( n365903 , n365902 );
not ( n45729 , n365903 );
or ( n365905 , n45713 , n45729 );
not ( n365906 , n43274 );
nand ( n45732 , n365906 , n364942 );
nand ( n45733 , n365905 , n45732 );
not ( n45734 , n45733 );
not ( n365910 , n45734 );
buf ( n365911 , n42263 );
not ( n365912 , n365911 );
buf ( n365913 , n362417 );
buf ( n45739 , n365913 );
buf ( n365915 , n45739 );
buf ( n365916 , n365915 );
not ( n45742 , n365916 );
buf ( n365918 , n45742 );
and ( n45744 , n361716 , n365918 );
not ( n45745 , n361716 );
and ( n45746 , n45745 , n362426 );
or ( n45747 , n45744 , n45746 );
buf ( n365923 , n45747 );
not ( n45749 , n365923 );
or ( n365925 , n365912 , n45749 );
buf ( n45751 , n365779 );
buf ( n365927 , n42242 );
nand ( n365928 , n45751 , n365927 );
buf ( n365929 , n365928 );
buf ( n365930 , n365929 );
nand ( n365931 , n365925 , n365930 );
buf ( n365932 , n365931 );
buf ( n365933 , n365932 );
not ( n365934 , n365933 );
buf ( n365935 , n365517 );
not ( n45761 , n365935 );
buf ( n365937 , n45345 );
not ( n365938 , n365937 );
or ( n45764 , n45761 , n365938 );
not ( n365940 , n31197 );
not ( n365941 , n365498 );
or ( n45767 , n365940 , n365941 );
buf ( n365943 , n360065 );
not ( n365944 , n365943 );
buf ( n365945 , n365944 );
buf ( n365946 , n365945 );
not ( n365947 , n365946 );
buf ( n365948 , n365947 );
nand ( n365949 , n365948 , n351229 );
nand ( n365950 , n45767 , n365949 );
buf ( n365951 , n365950 );
buf ( n365952 , n360051 );
not ( n45778 , n365952 );
buf ( n365954 , n45778 );
buf ( n365955 , n365954 );
nand ( n45781 , n365951 , n365955 );
buf ( n365957 , n45781 );
buf ( n365958 , n365957 );
nand ( n365959 , n45764 , n365958 );
buf ( n365960 , n365959 );
buf ( n365961 , n365960 );
not ( n45787 , n365961 );
buf ( n365963 , n45787 );
buf ( n45789 , n365963 );
nand ( n45790 , n365934 , n45789 );
buf ( n365966 , n45790 );
buf ( n365967 , n365966 );
buf ( n365968 , n365432 );
not ( n45794 , n365968 );
not ( n45795 , n42886 );
buf ( n365971 , n45795 );
not ( n45797 , n365971 );
or ( n45798 , n45794 , n45797 );
buf ( n365974 , n39592 );
buf ( n45800 , n31093 );
buf ( n45801 , n45800 );
buf ( n45802 , n45801 );
buf ( n365978 , n45802 );
buf ( n45804 , n365978 );
buf ( n365980 , n45804 );
buf ( n365981 , n365980 );
not ( n365982 , n365981 );
buf ( n365983 , n361631 );
not ( n45809 , n365983 );
or ( n365985 , n365982 , n45809 );
buf ( n365986 , n39621 );
buf ( n365987 , n365980 );
not ( n365988 , n365987 );
buf ( n365989 , n365988 );
buf ( n365990 , n365989 );
nand ( n365991 , n365986 , n365990 );
buf ( n365992 , n365991 );
buf ( n365993 , n365992 );
nand ( n45819 , n365985 , n365993 );
buf ( n365995 , n45819 );
buf ( n365996 , n365995 );
nand ( n365997 , n365974 , n365996 );
buf ( n365998 , n365997 );
buf ( n365999 , n365998 );
nand ( n366000 , n45798 , n365999 );
buf ( n366001 , n366000 );
buf ( n366002 , n366001 );
and ( n366003 , n365967 , n366002 );
buf ( n366004 , n365932 );
buf ( n366005 , n365960 );
and ( n45831 , n366004 , n366005 );
buf ( n366007 , n45831 );
buf ( n366008 , n366007 );
nor ( n45834 , n366003 , n366008 );
buf ( n366010 , n45834 );
not ( n45836 , n366010 );
and ( n366012 , n365910 , n45836 );
buf ( n366013 , n45734 );
buf ( n366014 , n366010 );
nand ( n366015 , n366013 , n366014 );
buf ( n366016 , n366015 );
buf ( n366017 , n45401 );
not ( n366018 , n366017 );
not ( n366019 , n360987 );
not ( n45845 , n40857 );
or ( n366021 , n366019 , n45845 );
nand ( n366022 , n366021 , n361011 );
buf ( n366023 , n366022 );
not ( n366024 , n366023 );
buf ( n366025 , n366024 );
buf ( n366026 , n366025 );
not ( n45852 , n366026 );
or ( n366028 , n366018 , n45852 );
buf ( n366029 , n40923 );
not ( n45855 , n360533 );
and ( n366031 , n45855 , n31073 );
not ( n366032 , n45855 );
and ( n45858 , n366032 , n351107 );
or ( n45859 , n366031 , n45858 );
buf ( n366035 , n45859 );
nand ( n366036 , n366029 , n366035 );
buf ( n366037 , n366036 );
buf ( n366038 , n366037 );
nand ( n45864 , n366028 , n366038 );
buf ( n366040 , n45864 );
buf ( n366041 , n366040 );
buf ( n366042 , n365640 );
not ( n366043 , n366042 );
buf ( n366044 , n41882 );
not ( n366045 , n366044 );
buf ( n366046 , n366045 );
buf ( n366047 , n366046 );
not ( n45873 , n366047 );
or ( n45874 , n366043 , n45873 );
buf ( n366050 , n41918 );
buf ( n366051 , n30912 );
not ( n45877 , n366051 );
buf ( n366053 , n44634 );
not ( n366054 , n366053 );
or ( n45880 , n45877 , n366054 );
buf ( n366056 , n41892 );
buf ( n366057 , n363041 );
nand ( n366058 , n366056 , n366057 );
buf ( n366059 , n366058 );
buf ( n366060 , n366059 );
nand ( n45886 , n45880 , n366060 );
buf ( n366062 , n45886 );
buf ( n366063 , n366062 );
nand ( n366064 , n366050 , n366063 );
buf ( n366065 , n366064 );
buf ( n366066 , n366065 );
nand ( n366067 , n45874 , n366066 );
buf ( n366068 , n366067 );
buf ( n366069 , n366068 );
not ( n366070 , n366069 );
buf ( n366071 , n366070 );
buf ( n366072 , n366071 );
xor ( n366073 , n366041 , n366072 );
not ( n366074 , n361603 );
not ( n45900 , n365593 );
and ( n45901 , n366074 , n45900 );
not ( n366077 , n32084 );
not ( n366078 , n366077 );
buf ( n366079 , n366078 );
not ( n366080 , n366079 );
buf ( n366081 , n41386 );
not ( n45907 , n366081 );
buf ( n45908 , n45907 );
buf ( n366084 , n45908 );
not ( n45910 , n366084 );
buf ( n366086 , n45910 );
buf ( n366087 , n366086 );
not ( n366088 , n366087 );
or ( n45914 , n366080 , n366088 );
not ( n45915 , n32084 );
not ( n45916 , n45915 );
buf ( n366092 , n45916 );
not ( n366093 , n366092 );
buf ( n366094 , n44717 );
not ( n366095 , n366094 );
buf ( n366096 , n366095 );
buf ( n366097 , n366096 );
nand ( n366098 , n366093 , n366097 );
buf ( n366099 , n366098 );
buf ( n366100 , n366099 );
nand ( n45926 , n45914 , n366100 );
buf ( n366102 , n45926 );
not ( n366103 , n41481 );
and ( n45929 , n366102 , n366103 );
nor ( n366105 , n45901 , n45929 );
buf ( n366106 , n366105 );
xor ( n45932 , n366073 , n366106 );
buf ( n366108 , n45932 );
and ( n45934 , n366016 , n366108 );
nor ( n45935 , n366012 , n45934 );
buf ( n366111 , n45935 );
not ( n45937 , n366111 );
buf ( n366113 , n45937 );
not ( n366114 , n366113 );
buf ( n366115 , n45859 );
not ( n366116 , n366115 );
buf ( n366117 , n366116 );
buf ( n366118 , n366117 );
not ( n45944 , n366118 );
buf ( n366120 , n366022 );
not ( n366121 , n366120 );
and ( n45947 , n45944 , n366121 );
buf ( n366123 , n364858 );
not ( n45949 , n366123 );
buf ( n366125 , n365290 );
not ( n366126 , n366125 );
or ( n366127 , n45949 , n366126 );
buf ( n366128 , n365266 );
buf ( n366129 , n351367 );
not ( n366130 , n366129 );
buf ( n366131 , n366130 );
buf ( n366132 , n366131 );
nand ( n366133 , n366128 , n366132 );
buf ( n366134 , n366133 );
buf ( n366135 , n366134 );
nand ( n366136 , n366127 , n366135 );
buf ( n366137 , n366136 );
buf ( n366138 , n366137 );
not ( n366139 , n366138 );
buf ( n366140 , n45384 );
nor ( n45966 , n366139 , n366140 );
buf ( n366142 , n45966 );
buf ( n366143 , n366142 );
nor ( n366144 , n45947 , n366143 );
buf ( n366145 , n366144 );
not ( n45971 , n360613 );
not ( n366147 , n45113 );
or ( n366148 , n45971 , n366147 );
buf ( n366149 , n365468 );
not ( n366150 , n366149 );
buf ( n366151 , n366150 );
nand ( n45977 , n366151 , n352194 );
nand ( n45978 , n366148 , n45977 );
not ( n366154 , n45978 );
buf ( n366155 , n40445 );
not ( n366156 , n366155 );
buf ( n366157 , n366156 );
nand ( n45983 , n366157 , n40473 );
buf ( n366159 , n45983 );
not ( n45985 , n366159 );
buf ( n366161 , n45985 );
not ( n45987 , n366161 );
or ( n45988 , n366154 , n45987 );
not ( n366164 , n351318 );
not ( n45990 , n365471 );
or ( n366166 , n366164 , n45990 );
nand ( n366167 , n360613 , n351320 );
nand ( n45993 , n366166 , n366167 );
nand ( n366169 , n45993 , n360574 );
nand ( n366170 , n45988 , n366169 );
buf ( n45996 , n366170 );
xor ( n45997 , n366145 , n45996 );
buf ( n366173 , n366062 );
not ( n366174 , n366173 );
buf ( n366175 , n364797 );
not ( n46001 , n366175 );
or ( n366177 , n366174 , n46001 );
buf ( n366178 , n41918 );
buf ( n366179 , n351762 );
not ( n366180 , n366179 );
buf ( n366181 , n365626 );
not ( n46007 , n366181 );
or ( n46008 , n366180 , n46007 );
buf ( n366184 , n362033 );
buf ( n366185 , n351762 );
not ( n46011 , n366185 );
buf ( n366187 , n46011 );
buf ( n46013 , n366187 );
nand ( n46014 , n366184 , n46013 );
buf ( n366190 , n46014 );
buf ( n366191 , n366190 );
nand ( n366192 , n46008 , n366191 );
buf ( n366193 , n366192 );
buf ( n366194 , n366193 );
nand ( n366195 , n366178 , n366194 );
buf ( n366196 , n366195 );
buf ( n366197 , n366196 );
nand ( n46023 , n366177 , n366197 );
buf ( n366199 , n46023 );
xor ( n46025 , n45997 , n366199 );
not ( n366201 , n46025 );
not ( n366202 , n366201 );
buf ( n366203 , n42266 );
buf ( n366204 , n365746 );
or ( n46030 , n366203 , n366204 );
buf ( n46031 , n361800 );
buf ( n366207 , n365915 );
buf ( n46033 , n366207 );
buf ( n366209 , n46033 );
buf ( n46035 , n366209 );
not ( n46036 , n46035 );
buf ( n366212 , n46036 );
and ( n46038 , n46031 , n366212 );
not ( n46039 , n46031 );
and ( n46040 , n46039 , n366209 );
nor ( n46041 , n46038 , n46040 );
buf ( n366217 , n46041 );
buf ( n366218 , n362388 );
or ( n46044 , n366217 , n366218 );
nand ( n366220 , n46030 , n46044 );
buf ( n366221 , n366220 );
buf ( n366222 , n366221 );
not ( n46048 , n366222 );
buf ( n366224 , n365793 );
not ( n46050 , n366224 );
buf ( n366226 , n46050 );
buf ( n366227 , n366226 );
not ( n46053 , n366227 );
buf ( n366229 , n46053 );
buf ( n366230 , n366229 );
not ( n366231 , n366230 );
buf ( n366232 , n365810 );
not ( n46058 , n366232 );
and ( n366234 , n366231 , n46058 );
buf ( n366235 , n359993 );
not ( n46061 , n366235 );
buf ( n366237 , n46061 );
buf ( n46063 , n366237 );
and ( n46064 , n31197 , n359947 );
not ( n366240 , n31197 );
buf ( n366241 , n359947 );
not ( n46067 , n366241 );
buf ( n366243 , n46067 );
and ( n46069 , n366240 , n366243 );
nor ( n366245 , n46064 , n46069 );
buf ( n366246 , n366245 );
nor ( n46072 , n46063 , n366246 );
buf ( n366248 , n46072 );
buf ( n366249 , n366248 );
nor ( n46075 , n366234 , n366249 );
buf ( n366251 , n46075 );
buf ( n366252 , n366251 );
not ( n366253 , n366252 );
or ( n366254 , n46048 , n366253 );
buf ( n366255 , n366251 );
buf ( n366256 , n366221 );
or ( n366257 , n366255 , n366256 );
nand ( n46083 , n366254 , n366257 );
buf ( n46084 , n46083 );
not ( n366260 , n46084 );
not ( n366261 , n366260 );
or ( n46087 , n366202 , n366261 );
nand ( n366263 , n46025 , n46084 );
nand ( n46089 , n46087 , n366263 );
not ( n46090 , n46089 );
not ( n366266 , n46090 );
or ( n366267 , n366114 , n366266 );
buf ( n366268 , n46089 );
buf ( n366269 , n45935 );
nand ( n366270 , n366268 , n366269 );
buf ( n366271 , n366270 );
nand ( n366272 , n366267 , n366271 );
buf ( n46098 , n352212 );
not ( n46099 , n46098 );
buf ( n366275 , n360610 );
not ( n46101 , n366275 );
buf ( n366277 , n46101 );
buf ( n366278 , n366277 );
not ( n366279 , n366278 );
or ( n46105 , n46099 , n366279 );
buf ( n366281 , n362452 );
buf ( n366282 , n365259 );
nand ( n46108 , n366281 , n366282 );
buf ( n46109 , n46108 );
buf ( n366285 , n46109 );
nand ( n46111 , n46105 , n366285 );
buf ( n366287 , n46111 );
not ( n366288 , n366287 );
and ( n46113 , n40473 , n360583 );
not ( n366290 , n46113 );
or ( n366291 , n366288 , n366290 );
buf ( n366292 , n45978 );
buf ( n366293 , n360574 );
nand ( n366294 , n366292 , n366293 );
buf ( n366295 , n366294 );
nand ( n366296 , n366291 , n366295 );
not ( n46121 , n366296 );
buf ( n366298 , n364766 );
not ( n366299 , n366298 );
buf ( n46124 , n362534 );
not ( n46125 , n46124 );
buf ( n46126 , n46125 );
buf ( n366303 , n46126 );
not ( n46128 , n366303 );
or ( n366305 , n366299 , n46128 );
buf ( n366306 , n362534 );
buf ( n366307 , n364783 );
nand ( n366308 , n366306 , n366307 );
buf ( n366309 , n366308 );
buf ( n366310 , n366309 );
nand ( n366311 , n366305 , n366310 );
buf ( n366312 , n366311 );
not ( n366313 , n366312 );
not ( n366314 , n366313 );
not ( n366315 , n361970 );
buf ( n46135 , n366315 );
not ( n366317 , n46135 );
not ( n366318 , n366317 );
and ( n46138 , n366314 , n366318 );
buf ( n366320 , n44570 );
not ( n366321 , n366320 );
not ( n366322 , n41569 );
buf ( n366323 , n366322 );
not ( n46143 , n366323 );
or ( n46144 , n366321 , n46143 );
buf ( n366326 , n41569 );
buf ( n366327 , n361597 );
not ( n46147 , n366327 );
buf ( n366329 , n46147 );
buf ( n366330 , n366329 );
not ( n46150 , n366330 );
buf ( n366332 , n46150 );
buf ( n366333 , n366332 );
nand ( n46153 , n366326 , n366333 );
buf ( n366335 , n46153 );
buf ( n366336 , n366335 );
nand ( n46156 , n46144 , n366336 );
buf ( n46157 , n46156 );
buf ( n366339 , n361975 );
not ( n46159 , n366339 );
and ( n366341 , n46157 , n46159 );
nor ( n366342 , n46138 , n366341 );
and ( n46162 , n46121 , n366342 );
not ( n366344 , n46121 );
buf ( n366345 , n366342 );
not ( n366346 , n366345 );
buf ( n366347 , n366346 );
and ( n46167 , n366344 , n366347 );
nor ( n46168 , n46162 , n46167 );
not ( n366350 , n39207 );
xor ( n366351 , n365367 , n365452 );
not ( n46171 , n366351 );
and ( n366353 , n366350 , n46171 );
buf ( n366354 , n45300 );
not ( n46174 , n366354 );
not ( n366356 , n355578 );
buf ( n366357 , n366356 );
not ( n46177 , n366357 );
or ( n366359 , n46174 , n46177 );
not ( n366360 , n359297 );
buf ( n366361 , n366360 );
buf ( n366362 , n365464 );
nand ( n366363 , n366361 , n366362 );
buf ( n366364 , n366363 );
buf ( n366365 , n366364 );
nand ( n46185 , n366359 , n366365 );
buf ( n366367 , n46185 );
not ( n46187 , n366367 );
not ( n46188 , n359312 );
nor ( n46189 , n46187 , n46188 );
nor ( n46190 , n366353 , n46189 );
and ( n366372 , n46168 , n46190 );
not ( n46192 , n46168 );
not ( n46193 , n46190 );
and ( n366375 , n46192 , n46193 );
nor ( n366376 , n366372 , n366375 );
not ( n366377 , n366376 );
buf ( n366378 , n342653 );
not ( n46198 , n366378 );
not ( n366380 , n342759 );
buf ( n366381 , n366380 );
nand ( n46201 , n46198 , n366381 );
buf ( n46202 , n46201 );
buf ( n366384 , n46202 );
nand ( n46204 , n342653 , n22810 );
buf ( n366386 , n46204 );
not ( n366387 , n342614 );
not ( n46207 , n22810 );
or ( n46208 , n366387 , n46207 );
not ( n366390 , n22810 );
not ( n366391 , n342614 );
nand ( n46211 , n366390 , n366391 );
nand ( n366393 , n46208 , n46211 );
buf ( n366394 , n366393 );
and ( n366395 , n366384 , n366386 , n366394 );
buf ( n366396 , n366395 );
buf ( n366397 , n366396 );
buf ( n366398 , n366397 );
buf ( n366399 , n366398 );
buf ( n366400 , n366399 );
buf ( n366401 , n366400 );
buf ( n366402 , n366401 );
buf ( n366403 , n366402 );
not ( n366404 , n366403 );
buf ( n46224 , n362285 );
not ( n46225 , n46224 );
buf ( n366407 , n46225 );
and ( n46227 , n22710 , n366407 );
not ( n366409 , n22710 );
and ( n46229 , n366409 , n42149 );
or ( n366411 , n46227 , n46229 );
buf ( n366412 , n366411 );
not ( n46232 , n366412 );
or ( n366414 , n366404 , n46232 );
buf ( n366415 , n360885 );
not ( n46235 , n366415 );
buf ( n46236 , n46235 );
and ( n366418 , n46236 , n342656 );
not ( n46238 , n46236 );
and ( n366420 , n46238 , n342657 );
or ( n366421 , n366418 , n366420 );
buf ( n366422 , n366421 );
buf ( n366423 , n366393 );
not ( n366424 , n366423 );
buf ( n366425 , n366424 );
buf ( n366426 , n366425 );
buf ( n366427 , n366426 );
buf ( n366428 , n366427 );
buf ( n366429 , n366428 );
not ( n366430 , n366429 );
buf ( n366431 , n366430 );
buf ( n366432 , n366431 );
not ( n366433 , n366432 );
buf ( n366434 , n366433 );
buf ( n366435 , n366434 );
nand ( n46255 , n366422 , n366435 );
buf ( n366437 , n46255 );
buf ( n366438 , n366437 );
nand ( n366439 , n366414 , n366438 );
buf ( n366440 , n366439 );
buf ( n366441 , n366440 );
not ( n46261 , n366441 );
buf ( n366443 , n46261 );
not ( n366444 , n366443 );
and ( n46264 , n366377 , n366444 );
buf ( n366446 , n366443 );
buf ( n366447 , n366376 );
nand ( n366448 , n366446 , n366447 );
buf ( n366449 , n366448 );
not ( n46269 , n44591 );
not ( n46270 , n364753 );
or ( n46271 , n46269 , n46270 );
buf ( n366453 , n366312 );
buf ( n46273 , n46159 );
nand ( n46274 , n366453 , n46273 );
buf ( n366456 , n46274 );
nand ( n46276 , n46271 , n366456 );
buf ( n366458 , n365950 );
not ( n46278 , n366458 );
buf ( n366460 , n45345 );
not ( n46280 , n366460 );
or ( n366462 , n46278 , n46280 );
buf ( n366463 , n45177 );
not ( n46283 , n366463 );
buf ( n366465 , n365498 );
not ( n366466 , n366465 );
or ( n46286 , n46283 , n366466 );
buf ( n366468 , n365495 );
buf ( n366469 , n365357 );
nand ( n46289 , n366468 , n366469 );
buf ( n46290 , n46289 );
buf ( n366472 , n46290 );
nand ( n366473 , n46286 , n366472 );
buf ( n366474 , n366473 );
buf ( n366475 , n366474 );
buf ( n366476 , n365954 );
nand ( n46296 , n366475 , n366476 );
buf ( n366478 , n46296 );
buf ( n366479 , n366478 );
nand ( n46299 , n366462 , n366479 );
buf ( n366481 , n46299 );
xor ( n46301 , n46276 , n366481 );
not ( n366483 , n362521 );
not ( n46303 , n44737 );
buf ( n366485 , n46303 );
not ( n366486 , n366485 );
buf ( n366487 , n45231 );
not ( n46307 , n366487 );
or ( n366489 , n366486 , n46307 );
buf ( n366490 , n45234 );
buf ( n366491 , n44737 );
nand ( n366492 , n366490 , n366491 );
buf ( n366493 , n366492 );
buf ( n366494 , n366493 );
nand ( n46314 , n366489 , n366494 );
buf ( n46315 , n46314 );
not ( n366497 , n46315 );
or ( n46317 , n366483 , n366497 );
nand ( n366499 , n365995 , n45795 );
nand ( n366500 , n46317 , n366499 );
xor ( n46320 , n46301 , n366500 );
and ( n366502 , n366449 , n46320 );
nor ( n46322 , n46264 , n366502 );
and ( n366504 , n366272 , n46322 );
not ( n46324 , n366272 );
buf ( n366506 , n46322 );
not ( n46326 , n366506 );
buf ( n366508 , n46326 );
and ( n366509 , n46324 , n366508 );
nor ( n366510 , n366504 , n366509 );
buf ( n46330 , n366510 );
not ( n366512 , n361606 );
not ( n366513 , n366102 );
or ( n46333 , n366512 , n366513 );
xor ( n366515 , n362549 , n366096 );
buf ( n366516 , n366515 );
not ( n46336 , n41481 );
buf ( n366518 , n46336 );
buf ( n46338 , n366518 );
nand ( n46339 , n366516 , n46338 );
buf ( n46340 , n46339 );
nand ( n366522 , n46333 , n46340 );
not ( n46342 , n366522 );
buf ( n366524 , n46315 );
not ( n366525 , n366524 );
buf ( n366526 , n45795 );
not ( n366527 , n366526 );
or ( n46347 , n366525 , n366527 );
buf ( n366529 , n362521 );
buf ( n366530 , n351160 );
not ( n46350 , n366530 );
buf ( n366532 , n359793 );
buf ( n366533 , n366532 );
buf ( n366534 , n366533 );
buf ( n366535 , n366534 );
not ( n46355 , n366535 );
buf ( n366537 , n46355 );
buf ( n366538 , n366537 );
not ( n366539 , n366538 );
or ( n46359 , n46350 , n366539 );
buf ( n366541 , n39621 );
buf ( n366542 , n364915 );
nand ( n46362 , n366541 , n366542 );
buf ( n366544 , n46362 );
buf ( n366545 , n366544 );
nand ( n366546 , n46359 , n366545 );
buf ( n366547 , n366546 );
buf ( n366548 , n366547 );
nand ( n366549 , n366529 , n366548 );
buf ( n366550 , n366549 );
buf ( n366551 , n366550 );
nand ( n366552 , n46347 , n366551 );
buf ( n366553 , n366552 );
buf ( n366554 , n366553 );
not ( n366555 , n366554 );
buf ( n366556 , n366555 );
xor ( n46376 , n46342 , n366556 );
buf ( n366558 , n366105 );
not ( n366559 , n366558 );
buf ( n366560 , n366071 );
not ( n366561 , n366560 );
or ( n366562 , n366559 , n366561 );
buf ( n366563 , n366040 );
nand ( n46383 , n366562 , n366563 );
buf ( n46384 , n46383 );
buf ( n46385 , n46384 );
buf ( n366567 , n366105 );
not ( n366568 , n366567 );
buf ( n366569 , n366068 );
nand ( n46389 , n366568 , n366569 );
buf ( n46390 , n46389 );
buf ( n366572 , n46390 );
nand ( n46392 , n46385 , n366572 );
buf ( n46393 , n46392 );
xor ( n366575 , n46376 , n46393 );
not ( n366576 , n365192 );
and ( n46396 , n366576 , n44966 );
not ( n46397 , n342909 );
not ( n366579 , n46397 );
not ( n46399 , n365047 );
or ( n46400 , n366579 , n46399 );
buf ( n366582 , n359144 );
buf ( n366583 , n342909 );
nand ( n366584 , n366582 , n366583 );
buf ( n366585 , n366584 );
nand ( n366586 , n46400 , n366585 );
not ( n366587 , n366586 );
nor ( n366588 , n366587 , n365155 );
nor ( n366589 , n46396 , n366588 );
xor ( n366590 , n366575 , n366589 );
not ( n366591 , n365101 );
not ( n46404 , n365036 );
and ( n366593 , n366591 , n46404 );
buf ( n366594 , n364997 );
not ( n46407 , n366594 );
buf ( n46408 , n46407 );
buf ( n366597 , n46408 );
not ( n46410 , n366597 );
not ( n366599 , n359937 );
buf ( n366600 , n366599 );
buf ( n366601 , n366600 );
not ( n366602 , n366601 );
or ( n366603 , n46410 , n366602 );
buf ( n366604 , n39830 );
buf ( n366605 , n364994 );
nand ( n46418 , n366604 , n366605 );
buf ( n366607 , n46418 );
buf ( n366608 , n366607 );
nand ( n46421 , n366603 , n366608 );
buf ( n366610 , n46421 );
buf ( n366611 , n366610 );
not ( n366612 , n366611 );
buf ( n366613 , n365118 );
not ( n46426 , n366613 );
buf ( n366615 , n46426 );
buf ( n46428 , n366615 );
nor ( n46429 , n366612 , n46428 );
buf ( n46430 , n46429 );
nor ( n366619 , n366593 , n46430 );
xor ( n46432 , n366590 , n366619 );
buf ( n366621 , n46432 );
buf ( n366622 , n365787 );
not ( n46435 , n366622 );
buf ( n366624 , n365836 );
not ( n46437 , n366624 );
or ( n46438 , n46435 , n46437 );
buf ( n46439 , n365816 );
buf ( n366628 , n365840 );
nand ( n366629 , n46439 , n366628 );
buf ( n366630 , n366629 );
buf ( n366631 , n366630 );
nand ( n46444 , n46438 , n366631 );
buf ( n366633 , n46444 );
buf ( n366634 , n366633 );
buf ( n366635 , n365829 );
xor ( n366636 , n366634 , n366635 );
buf ( n366637 , n366636 );
buf ( n366638 , n366637 );
not ( n366639 , n342564 );
and ( n366640 , n366639 , n342590 );
not ( n46453 , n366639 );
and ( n46454 , n22640 , n22633 );
not ( n366643 , n22640 );
not ( n366644 , n22633 );
and ( n46457 , n366643 , n366644 );
nor ( n366646 , n46454 , n46457 );
and ( n46459 , n46453 , n366646 );
nor ( n366648 , n366640 , n46459 );
buf ( n366649 , n366648 );
buf ( n366650 , n366649 );
not ( n46463 , n366650 );
buf ( n366652 , n46463 );
buf ( n366653 , n366652 );
buf ( n366654 , n366653 );
buf ( n366655 , n366654 );
not ( n366656 , n366655 );
buf ( n46469 , n342617 );
not ( n366658 , n46469 );
buf ( n366659 , n366658 );
buf ( n366660 , n366659 );
buf ( n46473 , n366660 );
buf ( n46474 , n46473 );
buf ( n366663 , n46474 );
not ( n46476 , n366663 );
buf ( n46477 , n46476 );
buf ( n366666 , n46477 );
not ( n46479 , n366666 );
buf ( n366668 , n362461 );
not ( n366669 , n366668 );
or ( n366670 , n46479 , n366669 );
buf ( n366671 , n360845 );
not ( n366672 , n366671 );
buf ( n366673 , n366672 );
buf ( n366674 , n366673 );
buf ( n366675 , n366674 );
buf ( n366676 , n366675 );
buf ( n366677 , n366676 );
not ( n46490 , n366677 );
buf ( n46491 , n46490 );
buf ( n366680 , n46491 );
buf ( n366681 , n46477 );
not ( n46494 , n366681 );
buf ( n366683 , n46494 );
buf ( n366684 , n366683 );
nand ( n366685 , n366680 , n366684 );
buf ( n366686 , n366685 );
buf ( n366687 , n366686 );
nand ( n46500 , n366670 , n366687 );
buf ( n366689 , n46500 );
buf ( n366690 , n366689 );
not ( n366691 , n366690 );
or ( n366692 , n366656 , n366691 );
not ( n46505 , n366683 );
not ( n366694 , n360893 );
or ( n46507 , n46505 , n366694 );
nand ( n366696 , n46477 , n360886 );
nand ( n46509 , n46507 , n366696 );
buf ( n366698 , n342614 );
not ( n46511 , n366698 );
buf ( n366700 , n366646 );
nand ( n46513 , n46511 , n366700 );
buf ( n366702 , n46513 );
buf ( n366703 , n342614 );
buf ( n366704 , n342590 );
nand ( n46517 , n366703 , n366704 );
buf ( n366706 , n46517 );
and ( n366707 , n366702 , n366648 , n366706 );
not ( n366708 , n366707 );
not ( n46521 , n366708 );
nand ( n46522 , n46509 , n46521 );
buf ( n366711 , n46522 );
nand ( n366712 , n366692 , n366711 );
buf ( n366713 , n366712 );
not ( n46526 , n366713 );
not ( n366715 , n45492 );
not ( n366716 , n365673 );
buf ( n366717 , n363391 );
not ( n366718 , n366717 );
buf ( n366719 , n366718 );
not ( n46532 , n366719 );
or ( n366721 , n366716 , n46532 );
buf ( n366722 , n40273 );
buf ( n366723 , n366722 );
not ( n366724 , n366723 );
buf ( n366725 , n366724 );
nand ( n46538 , n366725 , n365676 );
nand ( n366727 , n366721 , n46538 );
not ( n366728 , n366727 );
or ( n366729 , n366715 , n366728 );
buf ( n366730 , n45553 );
not ( n366731 , n366730 );
buf ( n366732 , n366731 );
not ( n46545 , n366732 );
xnor ( n46546 , n365673 , n40251 );
nand ( n46547 , n46545 , n46546 );
nand ( n46548 , n366729 , n46547 );
not ( n46549 , n46548 );
nand ( n366738 , n46526 , n46549 );
not ( n366739 , n366738 );
buf ( n366740 , n46276 );
not ( n46553 , n366740 );
buf ( n366742 , n46553 );
buf ( n46555 , n366742 );
not ( n46556 , n365477 );
not ( n46557 , n40474 );
not ( n366746 , n46557 );
or ( n366747 , n46556 , n366746 );
buf ( n366748 , n366287 );
buf ( n366749 , n366157 );
not ( n46562 , n366749 );
buf ( n366751 , n46562 );
buf ( n366752 , n366751 );
not ( n46565 , n366752 );
buf ( n366754 , n46565 );
buf ( n366755 , n366754 );
not ( n366756 , n366755 );
buf ( n366757 , n366756 );
buf ( n366758 , n366757 );
nand ( n366759 , n366748 , n366758 );
buf ( n366760 , n366759 );
nand ( n366761 , n366747 , n366760 );
buf ( n366762 , n366761 );
xor ( n366763 , n46555 , n366762 );
buf ( n366764 , n39207 );
buf ( n366765 , n365363 );
not ( n366766 , n366765 );
buf ( n366767 , n366766 );
buf ( n366768 , n366767 );
or ( n46581 , n366764 , n366768 );
buf ( n46582 , n359312 );
not ( n46583 , n46582 );
buf ( n366772 , n46583 );
buf ( n366773 , n366351 );
or ( n46586 , n366772 , n366773 );
nand ( n46587 , n46581 , n46586 );
buf ( n366776 , n46587 );
buf ( n366777 , n366776 );
xor ( n46590 , n366763 , n366777 );
buf ( n366779 , n46590 );
not ( n366780 , n366779 );
or ( n46593 , n366739 , n366780 );
nand ( n366782 , n366713 , n46548 );
nand ( n366783 , n46593 , n366782 );
buf ( n366784 , n366783 );
xor ( n366785 , n366638 , n366784 );
buf ( n46598 , n366010 );
buf ( n366787 , n366108 );
buf ( n366788 , n45734 );
and ( n46601 , n366787 , n366788 );
not ( n46602 , n366787 );
buf ( n366791 , n45733 );
and ( n366792 , n46602 , n366791 );
nor ( n46605 , n46601 , n366792 );
buf ( n46606 , n46605 );
xor ( n46607 , n46598 , n46606 );
buf ( n366796 , n46607 );
and ( n46609 , n366785 , n366796 );
and ( n46610 , n366638 , n366784 );
or ( n46611 , n46609 , n46610 );
buf ( n366800 , n46611 );
buf ( n366801 , n366800 );
xor ( n46614 , n366621 , n366801 );
buf ( n366803 , n46614 );
xor ( n366804 , n46330 , n366803 );
buf ( n366805 , n366804 );
xor ( n366806 , n365887 , n366805 );
xor ( n46619 , n366638 , n366784 );
xor ( n46620 , n46619 , n366796 );
buf ( n366809 , n46620 );
buf ( n366810 , n366809 );
not ( n366811 , n45492 );
not ( n46624 , n46546 );
or ( n46625 , n366811 , n46624 );
buf ( n366814 , n365676 );
not ( n46627 , n366814 );
buf ( n366816 , n362461 );
not ( n46629 , n366816 );
or ( n46630 , n46627 , n46629 );
buf ( n46631 , n362458 );
buf ( n366820 , n365673 );
nand ( n366821 , n46631 , n366820 );
buf ( n366822 , n366821 );
buf ( n366823 , n366822 );
nand ( n46636 , n46630 , n366823 );
buf ( n366825 , n46636 );
buf ( n366826 , n366825 );
buf ( n366827 , n45553 );
nand ( n46640 , n366826 , n366827 );
buf ( n46641 , n46640 );
nand ( n366830 , n46625 , n46641 );
buf ( n366831 , n366830 );
xor ( n46644 , n365310 , n365341 );
xor ( n366833 , n46644 , n365377 );
buf ( n366834 , n366833 );
buf ( n366835 , n366834 );
xor ( n366836 , n366831 , n366835 );
xor ( n366837 , n365481 , n365540 );
xnor ( n46650 , n366837 , n365438 );
buf ( n366839 , n46650 );
and ( n46652 , n366836 , n366839 );
and ( n46653 , n366831 , n366835 );
or ( n46654 , n46652 , n46653 );
buf ( n366843 , n46654 );
buf ( n366844 , n366843 );
not ( n46657 , n366844 );
buf ( n366846 , n46657 );
buf ( n366847 , n366846 );
not ( n366848 , n366847 );
buf ( n366849 , n365381 );
xor ( n46662 , n45372 , n366849 );
xnor ( n366851 , n46662 , n365649 );
buf ( n366852 , n366851 );
not ( n46665 , n366852 );
or ( n46666 , n366848 , n46665 );
buf ( n366855 , n45113 );
not ( n366856 , n366855 );
buf ( n366857 , n364832 );
not ( n366858 , n366857 );
or ( n46671 , n366856 , n366858 );
buf ( n366860 , n45455 );
buf ( n366861 , n45125 );
nand ( n366862 , n366860 , n366861 );
buf ( n366863 , n366862 );
buf ( n366864 , n366863 );
nand ( n46677 , n46671 , n366864 );
buf ( n46678 , n46677 );
buf ( n366867 , n46678 );
not ( n46680 , n366867 );
buf ( n366869 , n362027 );
not ( n46682 , n366869 );
or ( n366871 , n46680 , n46682 );
buf ( n366872 , n365622 );
buf ( n366873 , n364816 );
nand ( n46686 , n366872 , n366873 );
buf ( n366875 , n46686 );
buf ( n366876 , n366875 );
nand ( n366877 , n366871 , n366876 );
buf ( n366878 , n366877 );
buf ( n366879 , n366878 );
not ( n366880 , n44796 );
not ( n46693 , n22768 );
not ( n366882 , n46693 );
not ( n366883 , n361712 );
or ( n46696 , n366882 , n366883 );
buf ( n366885 , n361716 );
buf ( n366886 , n364953 );
nand ( n46699 , n366885 , n366886 );
buf ( n366888 , n46699 );
nand ( n46701 , n46696 , n366888 );
not ( n46702 , n46701 );
or ( n46703 , n366880 , n46702 );
buf ( n366892 , n342719 );
not ( n366893 , n366892 );
buf ( n366894 , n365760 );
not ( n366895 , n366894 );
or ( n366896 , n366893 , n366895 );
buf ( n366897 , n41528 );
buf ( n366898 , n364953 );
nand ( n366899 , n366897 , n366898 );
buf ( n366900 , n366899 );
buf ( n366901 , n366900 );
nand ( n46714 , n366896 , n366901 );
buf ( n366903 , n46714 );
buf ( n366904 , n366903 );
buf ( n366905 , n43261 );
nand ( n46718 , n366904 , n366905 );
buf ( n46719 , n46718 );
nand ( n46720 , n46703 , n46719 );
buf ( n46721 , n46720 );
xor ( n46722 , n366879 , n46721 );
buf ( n46723 , n45177 );
not ( n46724 , n46723 );
buf ( n366913 , n45270 );
not ( n46726 , n366913 );
or ( n366915 , n46724 , n46726 );
buf ( n366916 , n362452 );
buf ( n366917 , n365357 );
nand ( n366918 , n366916 , n366917 );
buf ( n366919 , n366918 );
buf ( n366920 , n366919 );
nand ( n366921 , n366915 , n366920 );
buf ( n366922 , n366921 );
buf ( n366923 , n366922 );
not ( n366924 , n366923 );
buf ( n46737 , n40475 );
not ( n46738 , n46737 );
or ( n46739 , n366924 , n46738 );
buf ( n46740 , n365458 );
buf ( n46741 , n366757 );
nand ( n46742 , n46740 , n46741 );
buf ( n46743 , n46742 );
buf ( n46744 , n46743 );
nand ( n46745 , n46739 , n46744 );
buf ( n46746 , n46745 );
buf ( n46747 , n46746 );
and ( n46748 , n46722 , n46747 );
and ( n46749 , n366879 , n46721 );
or ( n46750 , n46748 , n46749 );
buf ( n46751 , n46750 );
not ( n366940 , n46751 );
buf ( n366941 , n46521 );
not ( n46754 , n366941 );
buf ( n366943 , n46477 );
not ( n366944 , n366943 );
buf ( n366945 , n366407 );
not ( n46758 , n366945 );
or ( n46759 , n366944 , n46758 );
buf ( n366948 , n42149 );
buf ( n366949 , n366683 );
nand ( n366950 , n366948 , n366949 );
buf ( n366951 , n366950 );
buf ( n366952 , n366951 );
nand ( n46765 , n46759 , n366952 );
buf ( n366954 , n46765 );
buf ( n366955 , n366954 );
not ( n46768 , n366955 );
or ( n366957 , n46754 , n46768 );
buf ( n366958 , n46509 );
buf ( n366959 , n366654 );
nand ( n366960 , n366958 , n366959 );
buf ( n366961 , n366960 );
buf ( n366962 , n366961 );
nand ( n366963 , n366957 , n366962 );
buf ( n366964 , n366963 );
not ( n46777 , n366964 );
or ( n366966 , n366940 , n46777 );
nor ( n366967 , n366964 , n46751 );
buf ( n366968 , n45170 );
not ( n46781 , n366968 );
buf ( n366970 , n365490 );
not ( n366971 , n366970 );
buf ( n366972 , n35547 );
not ( n366973 , n366972 );
or ( n46786 , n366971 , n366973 );
buf ( n366975 , n365353 );
buf ( n366976 , n45336 );
nand ( n46789 , n366975 , n366976 );
buf ( n366978 , n46789 );
buf ( n366979 , n366978 );
nand ( n46792 , n46786 , n366979 );
buf ( n366981 , n46792 );
not ( n46794 , n366981 );
buf ( n366983 , n359292 );
buf ( n366984 , n39205 );
nand ( n46797 , n366983 , n366984 );
buf ( n366986 , n46797 );
buf ( n366987 , n366986 );
not ( n366988 , n366987 );
buf ( n366989 , n366988 );
not ( n366990 , n366989 );
or ( n46803 , n46794 , n366990 );
not ( n46804 , n365372 );
nand ( n366993 , n46804 , n359312 );
nand ( n366994 , n46803 , n366993 );
buf ( n366995 , n366994 );
not ( n366996 , n366995 );
buf ( n366997 , n366996 );
buf ( n366998 , n366997 );
not ( n366999 , n366998 );
or ( n46812 , n46781 , n366999 );
buf ( n367001 , n46303 );
not ( n367002 , n367001 );
buf ( n367003 , n365498 );
not ( n46816 , n367003 );
or ( n367005 , n367002 , n46816 );
buf ( n367006 , n46303 );
not ( n46819 , n367006 );
buf ( n367008 , n365528 );
nand ( n46821 , n46819 , n367008 );
buf ( n367010 , n46821 );
buf ( n367011 , n367010 );
nand ( n46824 , n367005 , n367011 );
buf ( n367013 , n46824 );
buf ( n367014 , n367013 );
not ( n367015 , n367014 );
buf ( n367016 , n45345 );
not ( n46829 , n367016 );
or ( n46830 , n367015 , n46829 );
buf ( n367019 , n365535 );
buf ( n367020 , n39949 );
nand ( n46833 , n367019 , n367020 );
buf ( n46834 , n46833 );
buf ( n367023 , n46834 );
nand ( n46836 , n46830 , n367023 );
buf ( n367025 , n46836 );
buf ( n367026 , n367025 );
nand ( n367027 , n46812 , n367026 );
buf ( n367028 , n367027 );
buf ( n367029 , n45170 );
not ( n46842 , n367029 );
buf ( n367031 , n366994 );
nand ( n367032 , n46842 , n367031 );
buf ( n367033 , n367032 );
and ( n367034 , n367028 , n367033 );
or ( n46847 , n366967 , n367034 );
nand ( n46848 , n366966 , n46847 );
buf ( n367037 , n46848 );
nand ( n46850 , n46666 , n367037 );
buf ( n367039 , n46850 );
buf ( n367040 , n367039 );
buf ( n367041 , n366843 );
buf ( n367042 , n366851 );
not ( n46855 , n367042 );
buf ( n367044 , n46855 );
buf ( n46857 , n367044 );
nand ( n46858 , n367041 , n46857 );
buf ( n46859 , n46858 );
buf ( n367048 , n46859 );
nand ( n46861 , n367040 , n367048 );
buf ( n46862 , n46861 );
buf ( n367051 , n46862 );
xor ( n367052 , n366810 , n367051 );
buf ( n367053 , n45029 );
not ( n367054 , n367053 );
buf ( n367055 , n45077 );
not ( n46868 , n367055 );
or ( n367057 , n367054 , n46868 );
buf ( n367058 , n365250 );
buf ( n367059 , n365196 );
nand ( n46872 , n367058 , n367059 );
buf ( n367061 , n46872 );
buf ( n367062 , n367061 );
nand ( n367063 , n367057 , n367062 );
buf ( n367064 , n367063 );
buf ( n367065 , n367064 );
buf ( n367066 , n45477 );
xor ( n46879 , n367065 , n367066 );
buf ( n46880 , n46879 );
buf ( n367069 , n46880 );
and ( n46882 , n367052 , n367069 );
and ( n46883 , n366810 , n367051 );
or ( n367072 , n46882 , n46883 );
buf ( n367073 , n367072 );
buf ( n367074 , n367073 );
and ( n367075 , n366806 , n367074 );
and ( n367076 , n365887 , n366805 );
or ( n46889 , n367075 , n367076 );
buf ( n367078 , n46889 );
buf ( n367079 , n367078 );
buf ( n367080 , n365118 );
not ( n367081 , n367080 );
buf ( n367082 , n365003 );
not ( n46895 , n367082 );
or ( n367084 , n367081 , n46895 );
buf ( n367085 , n44819 );
not ( n46898 , n367085 );
buf ( n367087 , n360308 );
not ( n46900 , n367087 );
or ( n367089 , n46898 , n46900 );
not ( n46902 , n40199 );
buf ( n367091 , n46902 );
not ( n46904 , n367091 );
buf ( n367093 , n364997 );
nand ( n46906 , n46904 , n367093 );
buf ( n367095 , n46906 );
buf ( n367096 , n367095 );
nand ( n46909 , n367089 , n367096 );
buf ( n46910 , n46909 );
buf ( n46911 , n46910 );
buf ( n367100 , n365033 );
nand ( n367101 , n46911 , n367100 );
buf ( n367102 , n367101 );
buf ( n367103 , n367102 );
nand ( n367104 , n367084 , n367103 );
buf ( n367105 , n367104 );
not ( n367106 , n367105 );
buf ( n367107 , n366434 );
not ( n46920 , n367107 );
buf ( n367109 , n366411 );
not ( n367110 , n367109 );
or ( n46923 , n46920 , n367110 );
buf ( n367112 , n22710 );
not ( n367113 , n367112 );
buf ( n367114 , n362136 );
not ( n46927 , n367114 );
buf ( n367116 , n46927 );
buf ( n367117 , n367116 );
not ( n367118 , n367117 );
or ( n46931 , n367113 , n367118 );
buf ( n367120 , n362136 );
buf ( n367121 , n342657 );
nand ( n46934 , n367120 , n367121 );
buf ( n367123 , n46934 );
buf ( n367124 , n367123 );
nand ( n46937 , n46931 , n367124 );
buf ( n367126 , n46937 );
buf ( n367127 , n367126 );
buf ( n367128 , n366402 );
nand ( n367129 , n367127 , n367128 );
buf ( n367130 , n367129 );
buf ( n367131 , n367130 );
nand ( n367132 , n46923 , n367131 );
buf ( n367133 , n367132 );
not ( n367134 , n367133 );
or ( n46947 , n367106 , n367134 );
nor ( n367136 , n367105 , n367133 );
xor ( n367137 , n365932 , n365963 );
xor ( n46950 , n367137 , n366001 );
or ( n367139 , n367136 , n46950 );
nand ( n367140 , n46947 , n367139 );
buf ( n367141 , n367140 );
and ( n367142 , n46320 , n366443 );
not ( n367143 , n46320 );
and ( n367144 , n367143 , n366440 );
nor ( n367145 , n367142 , n367144 );
buf ( n46958 , n366376 );
xor ( n367147 , n367145 , n46958 );
buf ( n46960 , n367147 );
xor ( n46961 , n367141 , n46960 );
xor ( n367150 , n46555 , n366762 );
and ( n367151 , n367150 , n366777 );
and ( n46964 , n46555 , n366762 );
or ( n367153 , n367151 , n46964 );
buf ( n367154 , n367153 );
not ( n46967 , n366654 );
buf ( n367156 , n46477 );
not ( n46969 , n367156 );
not ( n367158 , n40251 );
buf ( n367159 , n367158 );
not ( n46972 , n367159 );
or ( n367161 , n46969 , n46972 );
buf ( n367162 , n40251 );
buf ( n367163 , n366683 );
nand ( n46976 , n367162 , n367163 );
buf ( n367165 , n46976 );
buf ( n367166 , n367165 );
nand ( n367167 , n367161 , n367166 );
buf ( n367168 , n367167 );
not ( n46981 , n367168 );
or ( n46982 , n46967 , n46981 );
buf ( n367171 , n366689 );
buf ( n367172 , n46521 );
nand ( n46985 , n367171 , n367172 );
buf ( n367174 , n46985 );
nand ( n46987 , n46982 , n367174 );
buf ( n367176 , n45553 );
not ( n46989 , n367176 );
buf ( n367178 , n366727 );
not ( n367179 , n367178 );
or ( n46992 , n46989 , n367179 );
nand ( n367181 , n365704 , n45492 );
buf ( n367182 , n367181 );
nand ( n367183 , n46992 , n367182 );
buf ( n367184 , n367183 );
xor ( n46997 , n46987 , n367184 );
xor ( n46998 , n367154 , n46997 );
buf ( n367187 , n46998 );
and ( n47000 , n46961 , n367187 );
and ( n47001 , n367141 , n46960 );
or ( n367190 , n47000 , n47001 );
buf ( n367191 , n367190 );
buf ( n367192 , n367191 );
not ( n367193 , n367192 );
buf ( n367194 , n367193 );
buf ( n367195 , n367194 );
buf ( n367196 , n366434 );
not ( n367197 , n367196 );
buf ( n367198 , n22710 );
not ( n367199 , n367198 );
buf ( n367200 , n360848 );
not ( n47013 , n367200 );
or ( n47014 , n367199 , n47013 );
buf ( n367203 , n362458 );
buf ( n367204 , n342657 );
nand ( n47017 , n367203 , n367204 );
buf ( n367206 , n47017 );
buf ( n367207 , n367206 );
nand ( n47020 , n47014 , n367207 );
buf ( n367209 , n47020 );
buf ( n367210 , n367209 );
not ( n367211 , n367210 );
or ( n47024 , n367197 , n367211 );
buf ( n367213 , n366421 );
buf ( n367214 , n366402 );
nand ( n47027 , n367213 , n367214 );
buf ( n367216 , n47027 );
buf ( n367217 , n367216 );
nand ( n47030 , n47024 , n367217 );
buf ( n47031 , n47030 );
not ( n367220 , n47031 );
buf ( n367221 , n366347 );
not ( n367222 , n367221 );
buf ( n367223 , n366296 );
not ( n47036 , n367223 );
or ( n367225 , n367222 , n47036 );
buf ( n367226 , n366342 );
not ( n47039 , n367226 );
buf ( n367228 , n46121 );
not ( n367229 , n367228 );
or ( n47042 , n47039 , n367229 );
buf ( n367231 , n46193 );
nand ( n367232 , n47042 , n367231 );
buf ( n367233 , n367232 );
buf ( n367234 , n367233 );
nand ( n47047 , n367225 , n367234 );
buf ( n367236 , n47047 );
xor ( n47049 , n367220 , n367236 );
buf ( n367238 , n41835 );
not ( n367239 , n367238 );
buf ( n367240 , n366329 );
not ( n47053 , n367240 );
buf ( n367242 , n365760 );
not ( n47055 , n367242 );
or ( n367244 , n47053 , n47055 );
buf ( n367245 , n365757 );
buf ( n367246 , n364744 );
not ( n47059 , n367246 );
buf ( n367248 , n47059 );
buf ( n367249 , n367248 );
nand ( n47062 , n367245 , n367249 );
buf ( n47063 , n47062 );
buf ( n367252 , n47063 );
nand ( n47065 , n367244 , n367252 );
buf ( n367254 , n47065 );
buf ( n367255 , n367254 );
not ( n367256 , n367255 );
or ( n367257 , n367239 , n367256 );
buf ( n367258 , n46157 );
buf ( n367259 , n44591 );
nand ( n47072 , n367258 , n367259 );
buf ( n367261 , n47072 );
buf ( n367262 , n367261 );
nand ( n47075 , n367257 , n367262 );
buf ( n367264 , n47075 );
buf ( n367265 , n367264 );
not ( n47078 , n367265 );
buf ( n367267 , n47078 );
buf ( n367268 , n367267 );
buf ( n367269 , n366367 );
not ( n367270 , n367269 );
buf ( n367271 , n39207 );
not ( n367272 , n367271 );
buf ( n367273 , n367272 );
buf ( n367274 , n367273 );
not ( n367275 , n367274 );
or ( n367276 , n367270 , n367275 );
and ( n47089 , n35547 , n352212 );
nor ( n367278 , n352212 , n366356 );
nor ( n367279 , n47089 , n367278 );
buf ( n367280 , n367279 );
not ( n367281 , n367280 );
buf ( n367282 , n46582 );
nand ( n47095 , n367281 , n367282 );
buf ( n367284 , n47095 );
buf ( n367285 , n367284 );
nand ( n367286 , n367276 , n367285 );
buf ( n367287 , n367286 );
buf ( n367288 , n367287 );
not ( n367289 , n367288 );
buf ( n367290 , n367289 );
buf ( n367291 , n367290 );
xor ( n47104 , n367268 , n367291 );
buf ( n367293 , n47104 );
buf ( n47106 , n367293 );
buf ( n367295 , n45345 );
buf ( n367296 , n366474 );
and ( n367297 , n367295 , n367296 );
buf ( n367298 , n365440 );
not ( n367299 , n367298 );
buf ( n367300 , n360068 );
not ( n47113 , n367300 );
or ( n367302 , n367299 , n47113 );
buf ( n367303 , n363119 );
buf ( n367304 , n365452 );
nand ( n367305 , n367303 , n367304 );
buf ( n367306 , n367305 );
buf ( n367307 , n367306 );
nand ( n367308 , n367302 , n367307 );
buf ( n367309 , n367308 );
buf ( n367310 , n367309 );
not ( n367311 , n367310 );
buf ( n47124 , n360051 );
nor ( n47125 , n367311 , n47124 );
buf ( n47126 , n47125 );
buf ( n47127 , n47126 );
nor ( n47128 , n367297 , n47127 );
buf ( n47129 , n47128 );
buf ( n367318 , n47129 );
xor ( n47131 , n47106 , n367318 );
buf ( n367320 , n47131 );
xnor ( n47133 , n47049 , n367320 );
buf ( n367322 , n47133 );
buf ( n47135 , n367322 );
buf ( n367324 , n47135 );
buf ( n367325 , n367324 );
buf ( n367326 , n366654 );
not ( n367327 , n367326 );
buf ( n367328 , n367168 );
not ( n367329 , n367328 );
or ( n47142 , n367327 , n367329 );
buf ( n367331 , n367174 );
nand ( n367332 , n47142 , n367331 );
buf ( n367333 , n367332 );
buf ( n367334 , n367333 );
not ( n367335 , n367334 );
buf ( n367336 , n367184 );
not ( n47149 , n367336 );
or ( n367338 , n367335 , n47149 );
buf ( n367339 , n367184 );
buf ( n367340 , n367333 );
or ( n367341 , n367339 , n367340 );
buf ( n367342 , n367154 );
nand ( n47155 , n367341 , n367342 );
buf ( n367344 , n47155 );
buf ( n367345 , n367344 );
nand ( n47158 , n367338 , n367345 );
buf ( n367347 , n47158 );
buf ( n367348 , n43261 );
not ( n367349 , n367348 );
not ( n367350 , n22772 );
not ( n47163 , n366407 );
or ( n47164 , n367350 , n47163 );
not ( n47165 , n22772 );
nand ( n367354 , n47165 , n42149 );
nand ( n367355 , n47164 , n367354 );
buf ( n367356 , n367355 );
not ( n47169 , n367356 );
or ( n47170 , n367349 , n47169 );
buf ( n367359 , n365903 );
buf ( n367360 , n363429 );
nand ( n47173 , n367359 , n367360 );
buf ( n47174 , n47173 );
buf ( n367363 , n47174 );
nand ( n47176 , n47170 , n367363 );
buf ( n367365 , n47176 );
buf ( n47178 , n367365 );
xor ( n47179 , n46276 , n366481 );
and ( n367368 , n47179 , n366500 );
and ( n47181 , n46276 , n366481 );
or ( n47182 , n367368 , n47181 );
buf ( n367371 , n47182 );
xor ( n47184 , n47178 , n367371 );
buf ( n367373 , n46521 );
not ( n47186 , n367373 );
buf ( n367375 , n367168 );
not ( n47188 , n367375 );
or ( n47189 , n47186 , n47188 );
not ( n367378 , n360397 );
buf ( n47191 , n367378 );
not ( n47192 , n47191 );
buf ( n47193 , n47192 );
not ( n367382 , n47193 );
not ( n47195 , n46477 );
or ( n367384 , n367382 , n47195 );
buf ( n367385 , n366722 );
buf ( n367386 , n366683 );
nand ( n47199 , n367385 , n367386 );
buf ( n367388 , n47199 );
nand ( n47201 , n367384 , n367388 );
buf ( n367390 , n47201 );
buf ( n367391 , n366654 );
nand ( n47204 , n367390 , n367391 );
buf ( n47205 , n47204 );
buf ( n367394 , n47205 );
nand ( n47207 , n47189 , n367394 );
buf ( n367396 , n47207 );
buf ( n367397 , n367396 );
xor ( n47210 , n47184 , n367397 );
buf ( n367399 , n47210 );
buf ( n47212 , n367399 );
not ( n47213 , n47212 );
buf ( n367402 , n47213 );
and ( n367403 , n367347 , n367402 );
not ( n47216 , n367347 );
and ( n367405 , n47216 , n367399 );
or ( n47218 , n367403 , n367405 );
buf ( n367407 , n47218 );
xor ( n47220 , n367325 , n367407 );
buf ( n367409 , n47220 );
buf ( n47222 , n367409 );
nand ( n47223 , n367195 , n47222 );
buf ( n47224 , n47223 );
xor ( n367413 , n365089 , n44960 );
xor ( n47226 , n367413 , n44808 );
not ( n47227 , n47226 );
not ( n367416 , n47227 );
buf ( n367417 , n365980 );
not ( n367418 , n367417 );
buf ( n367419 , n364919 );
not ( n47232 , n367419 );
or ( n367421 , n367418 , n47232 );
buf ( n367422 , n44743 );
buf ( n367423 , n365989 );
nand ( n47236 , n367422 , n367423 );
buf ( n367425 , n47236 );
buf ( n367426 , n367425 );
nand ( n367427 , n367421 , n367426 );
buf ( n367428 , n367427 );
buf ( n367429 , n367428 );
not ( n47242 , n367429 );
buf ( n367431 , n47242 );
or ( n367432 , n364899 , n367431 );
and ( n47245 , n44737 , n364905 );
not ( n47246 , n44737 );
and ( n367435 , n47246 , n364909 );
nor ( n367436 , n47245 , n367435 );
not ( n47249 , n367436 );
buf ( n367438 , n359993 );
buf ( n47251 , n367438 );
buf ( n367440 , n47251 );
nand ( n47253 , n47249 , n367440 );
nand ( n47254 , n367432 , n47253 );
xor ( n47255 , n44629 , n44681 );
xor ( n367444 , n47255 , n44727 );
xor ( n47257 , n47254 , n367444 );
buf ( n367446 , n366434 );
not ( n47259 , n367446 );
buf ( n367448 , n367126 );
not ( n47261 , n367448 );
or ( n47262 , n47259 , n47261 );
buf ( n367451 , n22710 );
not ( n47264 , n367451 );
not ( n367453 , n361800 );
buf ( n367454 , n367453 );
not ( n367455 , n367454 );
or ( n47268 , n47264 , n367455 );
buf ( n367457 , n367453 );
not ( n367458 , n367457 );
buf ( n367459 , n367458 );
buf ( n367460 , n367459 );
buf ( n367461 , n342657 );
nand ( n367462 , n367460 , n367461 );
buf ( n367463 , n367462 );
buf ( n367464 , n367463 );
nand ( n367465 , n47268 , n367464 );
buf ( n367466 , n367465 );
buf ( n367467 , n367466 );
buf ( n367468 , n366402 );
nand ( n367469 , n367467 , n367468 );
buf ( n367470 , n367469 );
buf ( n367471 , n367470 );
nand ( n367472 , n47262 , n367471 );
buf ( n367473 , n367472 );
and ( n367474 , n47257 , n367473 );
and ( n47287 , n47254 , n367444 );
or ( n367476 , n367474 , n47287 );
not ( n47289 , n367476 );
not ( n47290 , n45021 );
not ( n367479 , n47290 );
buf ( n367480 , n22959 );
not ( n367481 , n367480 );
buf ( n367482 , n359976 );
not ( n47295 , n367482 );
or ( n367484 , n367481 , n47295 );
buf ( n367485 , n363171 );
buf ( n367486 , n342909 );
nand ( n367487 , n367485 , n367486 );
buf ( n367488 , n367487 );
buf ( n367489 , n367488 );
nand ( n367490 , n367484 , n367489 );
buf ( n367491 , n367490 );
not ( n367492 , n367491 );
or ( n47305 , n367479 , n367492 );
nand ( n367494 , n45005 , n365152 );
nand ( n367495 , n47305 , n367494 );
not ( n47308 , n367495 );
buf ( n367497 , n47308 );
buf ( n367498 , n42242 );
not ( n47311 , n367498 );
buf ( n367500 , n45747 );
not ( n47313 , n367500 );
or ( n367502 , n47311 , n47313 );
buf ( n367503 , n365915 );
not ( n47316 , n367503 );
buf ( n367505 , n362537 );
not ( n47318 , n367505 );
or ( n47319 , n47316 , n47318 );
buf ( n367508 , n46126 );
not ( n47321 , n367508 );
buf ( n367510 , n365918 );
nand ( n47323 , n47321 , n367510 );
buf ( n367512 , n47323 );
buf ( n367513 , n367512 );
nand ( n47326 , n47319 , n367513 );
buf ( n367515 , n47326 );
buf ( n367516 , n367515 );
buf ( n367517 , n42263 );
nand ( n47330 , n367516 , n367517 );
buf ( n47331 , n47330 );
buf ( n367520 , n47331 );
nand ( n47333 , n367502 , n367520 );
buf ( n367522 , n47333 );
buf ( n367523 , n367522 );
not ( n367524 , n367523 );
buf ( n367525 , n43261 );
not ( n47338 , n367525 );
buf ( n367527 , n364959 );
not ( n367528 , n367527 );
or ( n47341 , n47338 , n367528 );
buf ( n367530 , n44796 );
buf ( n367531 , n366903 );
nand ( n47344 , n367530 , n367531 );
buf ( n47345 , n47344 );
buf ( n367534 , n47345 );
nand ( n47347 , n47341 , n367534 );
buf ( n367536 , n47347 );
buf ( n47349 , n367536 );
not ( n367538 , n47349 );
buf ( n367539 , n367538 );
buf ( n367540 , n367539 );
nand ( n367541 , n367524 , n367540 );
buf ( n367542 , n367541 );
buf ( n367543 , n367542 );
not ( n47356 , n367543 );
buf ( n367545 , n42263 );
not ( n47358 , n367545 );
buf ( n367547 , n45595 );
not ( n47360 , n367547 );
buf ( n367549 , n32085 );
not ( n47362 , n367549 );
or ( n47363 , n47360 , n47362 );
buf ( n367552 , n364747 );
buf ( n367553 , n365773 );
nand ( n47366 , n367552 , n367553 );
buf ( n367555 , n47366 );
buf ( n47368 , n367555 );
nand ( n47369 , n47363 , n47368 );
buf ( n47370 , n47369 );
buf ( n367559 , n47370 );
not ( n47372 , n367559 );
or ( n367561 , n47358 , n47372 );
buf ( n367562 , n367515 );
buf ( n367563 , n42242 );
nand ( n367564 , n367562 , n367563 );
buf ( n367565 , n367564 );
buf ( n367566 , n367565 );
nand ( n47379 , n367561 , n367566 );
buf ( n367568 , n47379 );
buf ( n47381 , n367568 );
buf ( n367570 , n351107 );
not ( n367571 , n367570 );
buf ( n367572 , n366086 );
not ( n47385 , n367572 );
or ( n47386 , n367571 , n47385 );
not ( n367575 , n31072 );
not ( n367576 , n367575 );
buf ( n367577 , n367576 );
not ( n367578 , n367577 );
buf ( n367579 , n45908 );
nand ( n47392 , n367578 , n367579 );
buf ( n367581 , n47392 );
buf ( n367582 , n367581 );
nand ( n47395 , n47386 , n367582 );
buf ( n47396 , n47395 );
buf ( n367585 , n47396 );
not ( n47398 , n367585 );
buf ( n367587 , n361606 );
not ( n367588 , n367587 );
or ( n47401 , n47398 , n367588 );
not ( n367590 , n41481 );
nand ( n47403 , n367590 , n364876 );
buf ( n367592 , n47403 );
nand ( n367593 , n47401 , n367592 );
buf ( n367594 , n367593 );
buf ( n367595 , n367594 );
xor ( n47408 , n47381 , n367595 );
buf ( n367597 , n45376 );
buf ( n367598 , n351294 );
not ( n47411 , n367598 );
not ( n367600 , n365266 );
buf ( n367601 , n367600 );
not ( n47414 , n367601 );
or ( n367603 , n47411 , n47414 );
nand ( n367604 , n365474 , n45855 );
buf ( n367605 , n367604 );
nand ( n47418 , n367603 , n367605 );
buf ( n367607 , n47418 );
buf ( n367608 , n367607 );
not ( n47421 , n367608 );
buf ( n367610 , n47421 );
buf ( n367611 , n367610 );
or ( n47424 , n367597 , n367611 );
buf ( n367613 , n45384 );
buf ( n367614 , n365271 );
or ( n367615 , n367613 , n367614 );
nand ( n47428 , n47424 , n367615 );
buf ( n47429 , n47428 );
buf ( n367618 , n47429 );
and ( n47431 , n47408 , n367618 );
and ( n47432 , n47381 , n367595 );
or ( n47433 , n47431 , n47432 );
buf ( n367622 , n47433 );
buf ( n367623 , n367622 );
not ( n47436 , n367623 );
or ( n47437 , n47356 , n47436 );
buf ( n367626 , n367536 );
buf ( n367627 , n367522 );
nand ( n47440 , n367626 , n367627 );
buf ( n367629 , n47440 );
buf ( n367630 , n367629 );
nand ( n47443 , n47437 , n367630 );
buf ( n367632 , n47443 );
buf ( n367633 , n367632 );
not ( n47446 , n367633 );
buf ( n367635 , n47446 );
buf ( n47448 , n367635 );
nand ( n47449 , n367497 , n47448 );
buf ( n47450 , n47449 );
not ( n367639 , n47450 );
or ( n47452 , n47289 , n367639 );
not ( n367641 , n367635 );
nand ( n367642 , n367641 , n367495 );
nand ( n47455 , n47452 , n367642 );
not ( n367644 , n47455 );
or ( n47457 , n367416 , n367644 );
not ( n367646 , n47308 );
not ( n47459 , n367635 );
and ( n367648 , n367646 , n47459 );
and ( n47461 , n47450 , n367476 );
nor ( n47462 , n367648 , n47461 );
not ( n367651 , n47462 );
not ( n47464 , n47226 );
or ( n367653 , n367651 , n47464 );
not ( n47466 , n44913 );
not ( n47467 , n47466 );
buf ( n367656 , n365041 );
not ( n47469 , n367656 );
buf ( n367658 , n362179 );
not ( n47471 , n367658 );
or ( n47472 , n47469 , n47471 );
buf ( n367661 , n361617 );
buf ( n367662 , n365052 );
nand ( n47475 , n367661 , n367662 );
buf ( n367664 , n47475 );
buf ( n367665 , n367664 );
nand ( n367666 , n47472 , n367665 );
buf ( n367667 , n367666 );
not ( n47480 , n367667 );
or ( n367669 , n47467 , n47480 );
buf ( n47482 , n365058 );
buf ( n367671 , n44915 );
nand ( n367672 , n47482 , n367671 );
buf ( n367673 , n367672 );
nand ( n47486 , n367669 , n367673 );
not ( n47487 , n47486 );
not ( n47488 , n47487 );
not ( n47489 , n45075 );
not ( n47490 , n365208 );
or ( n367679 , n47489 , n47490 );
buf ( n367680 , n342881 );
not ( n367681 , n367680 );
buf ( n367682 , n362212 );
not ( n47495 , n367682 );
or ( n47496 , n367681 , n47495 );
buf ( n47497 , n359756 );
buf ( n367686 , n365202 );
nand ( n47499 , n47497 , n367686 );
buf ( n47500 , n47499 );
buf ( n367689 , n47500 );
nand ( n47502 , n47496 , n367689 );
buf ( n367691 , n47502 );
buf ( n47504 , n367691 );
buf ( n47505 , n45058 );
nand ( n47506 , n47504 , n47505 );
buf ( n47507 , n47506 );
nand ( n367696 , n367679 , n47507 );
not ( n47509 , n367696 );
not ( n367698 , n364968 );
not ( n47511 , n44766 );
and ( n367700 , n367698 , n47511 );
and ( n367701 , n44766 , n364968 );
nor ( n47514 , n367700 , n367701 );
not ( n367703 , n364895 );
xor ( n47516 , n47514 , n367703 );
not ( n367705 , n47516 );
nand ( n47518 , n47509 , n367705 );
nand ( n367707 , n47488 , n47518 );
nand ( n367708 , n367696 , n47516 );
nand ( n47521 , n367707 , n367708 );
nand ( n367710 , n367653 , n47521 );
nand ( n367711 , n47457 , n367710 );
and ( n47524 , n47224 , n367711 );
buf ( n367713 , n367191 );
not ( n367714 , n367713 );
buf ( n367715 , n367409 );
nor ( n367716 , n367714 , n367715 );
buf ( n367717 , n367716 );
nor ( n367718 , n47524 , n367717 );
not ( n47531 , n367718 );
not ( n47532 , n367236 );
buf ( n47533 , n366434 );
not ( n47534 , n47533 );
buf ( n47535 , n367209 );
not ( n47536 , n47535 );
or ( n47537 , n47534 , n47536 );
buf ( n367726 , n367216 );
nand ( n367727 , n47537 , n367726 );
buf ( n367728 , n367727 );
not ( n367729 , n367728 );
or ( n367730 , n47532 , n367729 );
buf ( n367731 , n367728 );
buf ( n367732 , n367236 );
nor ( n367733 , n367731 , n367732 );
buf ( n367734 , n367733 );
or ( n47547 , n367320 , n367734 );
nand ( n367736 , n367730 , n47547 );
buf ( n367737 , n367736 );
buf ( n367738 , n41835 );
not ( n367739 , n367738 );
buf ( n47552 , n41772 );
not ( n47553 , n47552 );
buf ( n47554 , n47553 );
buf ( n367743 , n47554 );
not ( n47556 , n367743 );
buf ( n367745 , n44783 );
not ( n47558 , n367745 );
or ( n47559 , n47556 , n47558 );
buf ( n367748 , n41607 );
buf ( n367749 , n41772 );
nand ( n47562 , n367748 , n367749 );
buf ( n367751 , n47562 );
buf ( n367752 , n367751 );
nand ( n47565 , n47559 , n367752 );
buf ( n367754 , n47565 );
buf ( n367755 , n367754 );
not ( n367756 , n367755 );
or ( n47569 , n367739 , n367756 );
buf ( n367758 , n367254 );
buf ( n367759 , n44591 );
buf ( n367760 , n367759 );
nand ( n47573 , n367758 , n367760 );
buf ( n367762 , n47573 );
buf ( n367763 , n367762 );
nand ( n367764 , n47569 , n367763 );
buf ( n367765 , n367764 );
buf ( n367766 , n367765 );
buf ( n367767 , n366145 );
not ( n367768 , n367767 );
buf ( n367769 , n367768 );
buf ( n367770 , n367769 );
not ( n47583 , n367770 );
buf ( n367772 , n45996 );
not ( n367773 , n367772 );
or ( n47586 , n47583 , n367773 );
buf ( n367775 , n366170 );
not ( n47588 , n367775 );
buf ( n367777 , n47588 );
buf ( n367778 , n367777 );
not ( n47591 , n367778 );
buf ( n367780 , n366145 );
not ( n367781 , n367780 );
or ( n47594 , n47591 , n367781 );
buf ( n367783 , n366199 );
nand ( n47596 , n47594 , n367783 );
buf ( n367785 , n47596 );
buf ( n367786 , n367785 );
nand ( n367787 , n47586 , n367786 );
buf ( n367788 , n367787 );
buf ( n367789 , n367788 );
xor ( n47602 , n367766 , n367789 );
buf ( n367791 , n366547 );
not ( n367792 , n367791 );
buf ( n367793 , n39701 );
not ( n367794 , n367793 );
or ( n47607 , n367792 , n367794 );
buf ( n367796 , n359685 );
buf ( n367797 , n367796 );
buf ( n367798 , n365490 );
not ( n367799 , n367798 );
buf ( n367800 , n366537 );
not ( n47613 , n367800 );
or ( n47614 , n367799 , n47613 );
buf ( n47615 , n39621 );
buf ( n47616 , n45336 );
nand ( n47617 , n47615 , n47616 );
buf ( n47618 , n47617 );
buf ( n367807 , n47618 );
nand ( n367808 , n47614 , n367807 );
buf ( n367809 , n367808 );
buf ( n367810 , n367809 );
nand ( n367811 , n367797 , n367810 );
buf ( n367812 , n367811 );
buf ( n367813 , n367812 );
nand ( n367814 , n47607 , n367813 );
buf ( n367815 , n367814 );
buf ( n367816 , n367815 );
not ( n47629 , n367816 );
buf ( n367818 , n47629 );
not ( n47631 , n367818 );
buf ( n367820 , n366193 );
not ( n367821 , n367820 );
buf ( n47634 , n45438 );
not ( n47635 , n47634 );
or ( n47636 , n367821 , n47635 );
buf ( n367825 , n45455 );
not ( n367826 , n367825 );
buf ( n367827 , n45915 );
not ( n367828 , n367827 );
or ( n367829 , n367826 , n367828 );
buf ( n367830 , n32084 );
buf ( n367831 , n44634 );
nand ( n367832 , n367830 , n367831 );
buf ( n367833 , n367832 );
buf ( n367834 , n367833 );
nand ( n367835 , n367829 , n367834 );
buf ( n367836 , n367835 );
buf ( n367837 , n367836 );
buf ( n367838 , n41915 );
nand ( n367839 , n367837 , n367838 );
buf ( n367840 , n367839 );
buf ( n367841 , n367840 );
nand ( n47654 , n47636 , n367841 );
buf ( n367843 , n47654 );
buf ( n367844 , n366137 );
not ( n47657 , n367844 );
buf ( n367846 , n366025 );
not ( n47659 , n367846 );
or ( n47660 , n47657 , n47659 );
buf ( n367849 , n40923 );
buf ( n367850 , n30912 );
not ( n47663 , n367850 );
buf ( n367852 , n367600 );
not ( n47665 , n367852 );
or ( n47666 , n47663 , n47665 );
buf ( n367855 , n45152 );
buf ( n367856 , n365569 );
nand ( n47669 , n367855 , n367856 );
buf ( n367858 , n47669 );
buf ( n367859 , n367858 );
nand ( n367860 , n47666 , n367859 );
buf ( n367861 , n367860 );
buf ( n367862 , n367861 );
nand ( n367863 , n367849 , n367862 );
buf ( n367864 , n367863 );
buf ( n367865 , n367864 );
nand ( n367866 , n47660 , n367865 );
buf ( n367867 , n367866 );
xor ( n367868 , n367843 , n367867 );
not ( n47681 , n367868 );
or ( n367870 , n47631 , n47681 );
or ( n47683 , n367818 , n367868 );
nand ( n47684 , n367870 , n47683 );
buf ( n367873 , n47684 );
xor ( n367874 , n47602 , n367873 );
buf ( n367875 , n367874 );
buf ( n367876 , n367875 );
xor ( n367877 , n367737 , n367876 );
not ( n47690 , n44796 );
not ( n367879 , n367355 );
or ( n367880 , n47690 , n367879 );
and ( n47693 , n360885 , n363444 );
not ( n367882 , n360885 );
and ( n47695 , n367882 , n22772 );
or ( n47696 , n47693 , n47695 );
buf ( n47697 , n47696 );
buf ( n47698 , n43261 );
nand ( n47699 , n47697 , n47698 );
buf ( n47700 , n47699 );
nand ( n367889 , n367880 , n47700 );
not ( n47702 , n366654 );
buf ( n367891 , n46477 );
not ( n367892 , n367891 );
buf ( n367893 , n45523 );
not ( n367894 , n367893 );
or ( n367895 , n367892 , n367894 );
buf ( n367896 , n40199 );
buf ( n367897 , n366683 );
nand ( n47710 , n367896 , n367897 );
buf ( n367899 , n47710 );
buf ( n367900 , n367899 );
nand ( n367901 , n367895 , n367900 );
buf ( n367902 , n367901 );
not ( n47715 , n367902 );
or ( n367904 , n47702 , n47715 );
nand ( n367905 , n47201 , n46521 );
nand ( n47718 , n367904 , n367905 );
xnor ( n367907 , n367889 , n47718 );
buf ( n367908 , n366434 );
not ( n47721 , n367908 );
buf ( n367910 , n22710 );
not ( n367911 , n367910 );
not ( n47724 , n40251 );
buf ( n367913 , n47724 );
not ( n367914 , n367913 );
or ( n47727 , n367911 , n367914 );
buf ( n367916 , n40251 );
buf ( n367917 , n342657 );
nand ( n47730 , n367916 , n367917 );
buf ( n47731 , n47730 );
buf ( n367920 , n47731 );
nand ( n367921 , n47727 , n367920 );
buf ( n367922 , n367921 );
buf ( n367923 , n367922 );
not ( n367924 , n367923 );
or ( n367925 , n47721 , n367924 );
buf ( n367926 , n366402 );
buf ( n367927 , n367209 );
nand ( n47733 , n367926 , n367927 );
buf ( n367929 , n47733 );
buf ( n367930 , n367929 );
nand ( n367931 , n367925 , n367930 );
buf ( n367932 , n367931 );
buf ( n367933 , n367932 );
not ( n367934 , n367933 );
buf ( n367935 , n367934 );
and ( n367936 , n367907 , n367935 );
not ( n47742 , n367907 );
and ( n47743 , n47742 , n367932 );
nor ( n47744 , n367936 , n47743 );
buf ( n367940 , n47744 );
xor ( n367941 , n367877 , n367940 );
buf ( n367942 , n367941 );
not ( n47748 , n367942 );
buf ( n367944 , n47133 );
not ( n47750 , n367944 );
buf ( n367946 , n47750 );
not ( n47752 , n367946 );
not ( n47753 , n367399 );
or ( n47754 , n47752 , n47753 );
not ( n47755 , n367402 );
not ( n47756 , n47133 );
or ( n367952 , n47755 , n47756 );
nand ( n47758 , n367952 , n367347 );
nand ( n47759 , n47754 , n47758 );
not ( n47760 , n47759 );
not ( n47761 , n47760 );
or ( n47762 , n47748 , n47761 );
not ( n47763 , n367942 );
not ( n47764 , n367946 );
not ( n47765 , n367399 );
or ( n47766 , n47764 , n47765 );
nand ( n47767 , n47766 , n47758 );
nand ( n47768 , n47763 , n47767 );
nand ( n367964 , n47762 , n47768 );
not ( n47770 , n365127 );
not ( n47771 , n365885 );
or ( n47772 , n47770 , n47771 );
buf ( n367968 , n365127 );
buf ( n47774 , n365885 );
nor ( n47775 , n367968 , n47774 );
buf ( n367971 , n47775 );
buf ( n367972 , n365656 );
not ( n367973 , n367972 );
buf ( n367974 , n367973 );
or ( n367975 , n367971 , n367974 );
nand ( n47781 , n47772 , n367975 );
and ( n47782 , n367964 , n47781 );
not ( n367978 , n367964 );
not ( n367979 , n47781 );
and ( n47785 , n367978 , n367979 );
nor ( n367981 , n47782 , n47785 );
and ( n367982 , n47531 , n367981 );
not ( n47788 , n47531 );
not ( n367984 , n367981 );
and ( n367985 , n47788 , n367984 );
nor ( n47791 , n367982 , n367985 );
not ( n47792 , n47791 );
not ( n367988 , n47792 );
buf ( n367989 , n366510 );
buf ( n367990 , n46432 );
nand ( n367991 , n367989 , n367990 );
buf ( n367992 , n367991 );
buf ( n367993 , n367992 );
buf ( n367994 , n366800 );
and ( n367995 , n367993 , n367994 );
buf ( n367996 , n46432 );
buf ( n367997 , n366510 );
nor ( n367998 , n367996 , n367997 );
buf ( n367999 , n367998 );
buf ( n368000 , n367999 );
nor ( n368001 , n367995 , n368000 );
buf ( n368002 , n368001 );
buf ( n368003 , n368002 );
not ( n47809 , n368003 );
not ( n47810 , n46393 );
nand ( n368006 , n366556 , n366522 );
not ( n47812 , n368006 );
or ( n368008 , n47810 , n47812 );
buf ( n368009 , n366553 );
buf ( n368010 , n46342 );
nand ( n368011 , n368009 , n368010 );
buf ( n368012 , n368011 );
nand ( n368013 , n368008 , n368012 );
buf ( n368014 , n365190 );
buf ( n368015 , n365155 );
nand ( n368016 , n368014 , n368015 );
buf ( n368017 , n368016 );
nand ( n368018 , n366586 , n368017 );
and ( n47824 , n368013 , n368018 );
not ( n368020 , n368013 );
not ( n368021 , n368018 );
and ( n47827 , n368020 , n368021 );
nor ( n368023 , n47824 , n47827 );
buf ( n368024 , n368023 );
not ( n47830 , n39217 );
and ( n47831 , n45113 , n35548 );
not ( n47832 , n45113 );
and ( n47833 , n47832 , n366356 );
nor ( n368029 , n47831 , n47833 );
not ( n47835 , n368029 );
or ( n368031 , n47830 , n47835 );
not ( n368032 , n367279 );
nand ( n368033 , n368032 , n45204 );
nand ( n47839 , n368031 , n368033 );
xor ( n47840 , n366522 , n47839 );
buf ( n47841 , n365801 );
not ( n47842 , n47841 );
buf ( n368038 , n47842 );
not ( n368039 , n368038 );
not ( n47845 , n44743 );
not ( n47846 , n365357 );
and ( n47847 , n47845 , n47846 );
and ( n47848 , n361762 , n365357 );
nor ( n47849 , n47847 , n47848 );
buf ( n368045 , n47849 );
not ( n368046 , n368045 );
buf ( n368047 , n368046 );
not ( n368048 , n368047 );
or ( n47854 , n368039 , n368048 );
not ( n47855 , n366245 );
not ( n368051 , n359913 );
nand ( n47857 , n47855 , n368051 );
nand ( n368053 , n47854 , n47857 );
xor ( n47859 , n47840 , n368053 );
buf ( n368055 , n47859 );
xnor ( n368056 , n368024 , n368055 );
buf ( n368057 , n368056 );
buf ( n368058 , n368057 );
not ( n47864 , n365876 );
not ( n47865 , n365734 );
and ( n47866 , n47864 , n47865 );
nor ( n47867 , n47866 , n365846 );
buf ( n368063 , n365876 );
buf ( n368064 , n365734 );
and ( n47870 , n368063 , n368064 );
buf ( n368066 , n47870 );
nor ( n47872 , n47867 , n368066 );
buf ( n368068 , n47872 );
xor ( n47874 , n368058 , n368068 );
xor ( n47875 , n366575 , n366589 );
and ( n47876 , n47875 , n366619 );
and ( n368072 , n366575 , n366589 );
or ( n47878 , n47876 , n368072 );
buf ( n368074 , n47878 );
xor ( n47880 , n47874 , n368074 );
buf ( n368076 , n47880 );
buf ( n47882 , n368076 );
not ( n368078 , n47882 );
buf ( n368079 , n368078 );
buf ( n368080 , n368079 );
not ( n368081 , n368080 );
or ( n47887 , n47809 , n368081 );
buf ( n368083 , n368002 );
not ( n47889 , n368083 );
buf ( n368085 , n47889 );
buf ( n368086 , n368085 );
buf ( n368087 , n368076 );
nand ( n368088 , n368086 , n368087 );
buf ( n368089 , n368088 );
buf ( n368090 , n368089 );
nand ( n368091 , n47887 , n368090 );
buf ( n368092 , n368091 );
buf ( n368093 , n368092 );
buf ( n368094 , n46089 );
not ( n47900 , n368094 );
buf ( n368096 , n47900 );
buf ( n368097 , n368096 );
not ( n368098 , n368097 );
buf ( n368099 , n366508 );
nand ( n368100 , n368098 , n368099 );
buf ( n368101 , n368100 );
buf ( n368102 , n368096 );
not ( n368103 , n368102 );
buf ( n368104 , n46322 );
not ( n47910 , n368104 );
or ( n368106 , n368103 , n47910 );
buf ( n47912 , n366113 );
buf ( n368108 , n47912 );
nand ( n368109 , n368106 , n368108 );
buf ( n368110 , n368109 );
nand ( n47916 , n368101 , n368110 );
not ( n368112 , n45075 );
not ( n368113 , n365202 );
not ( n47919 , n40899 );
or ( n368115 , n368113 , n47919 );
nand ( n368116 , n342881 , n40091 );
nand ( n47922 , n368115 , n368116 );
not ( n368118 , n47922 );
or ( n47924 , n368112 , n368118 );
buf ( n368120 , n45694 );
buf ( n368121 , n45058 );
nand ( n47927 , n368120 , n368121 );
buf ( n368123 , n47927 );
nand ( n47929 , n47924 , n368123 );
buf ( n368125 , n47929 );
not ( n47931 , n368125 );
buf ( n368127 , n365033 );
not ( n368128 , n368127 );
buf ( n368129 , n366610 );
not ( n47935 , n368129 );
or ( n368131 , n368128 , n47935 );
and ( n368132 , n44819 , n41907 );
not ( n47938 , n44819 );
and ( n368134 , n47938 , n39867 );
or ( n368135 , n368132 , n368134 );
buf ( n368136 , n368135 );
buf ( n368137 , n365118 );
nand ( n368138 , n368136 , n368137 );
buf ( n368139 , n368138 );
buf ( n368140 , n368139 );
nand ( n368141 , n368131 , n368140 );
buf ( n368142 , n368141 );
not ( n47948 , n368142 );
buf ( n368144 , n47948 );
not ( n368145 , n368144 );
or ( n47951 , n47931 , n368145 );
buf ( n368147 , n368142 );
not ( n47953 , n47929 );
buf ( n368149 , n47953 );
nand ( n368150 , n368147 , n368149 );
buf ( n368151 , n368150 );
buf ( n368152 , n368151 );
nand ( n368153 , n47951 , n368152 );
buf ( n368154 , n368153 );
buf ( n368155 , n366221 );
not ( n47961 , n368155 );
buf ( n368157 , n366251 );
nand ( n47963 , n47961 , n368157 );
buf ( n368159 , n47963 );
buf ( n368160 , n368159 );
not ( n47966 , n368160 );
not ( n368162 , n46025 );
buf ( n368163 , n368162 );
not ( n368164 , n368163 );
or ( n368165 , n47966 , n368164 );
buf ( n368166 , n366251 );
not ( n47972 , n368166 );
buf ( n368168 , n366221 );
nand ( n368169 , n47972 , n368168 );
buf ( n368170 , n368169 );
buf ( n368171 , n368170 );
nand ( n368172 , n368165 , n368171 );
buf ( n368173 , n368172 );
buf ( n368174 , n368173 );
not ( n368175 , n368174 );
buf ( n368176 , n368175 );
and ( n47982 , n368154 , n368176 );
not ( n368178 , n368154 );
and ( n368179 , n368178 , n368173 );
nor ( n47985 , n47982 , n368179 );
not ( n368181 , n47985 );
and ( n368182 , n47916 , n368181 );
not ( n47988 , n47916 );
and ( n47989 , n47988 , n47985 );
nor ( n368185 , n368182 , n47989 );
not ( n368186 , n45492 );
buf ( n368187 , n365676 );
not ( n368188 , n368187 );
buf ( n368189 , n362212 );
not ( n368190 , n368189 );
or ( n47996 , n368188 , n368190 );
buf ( n368192 , n359756 );
buf ( n368193 , n365673 );
nand ( n368194 , n368192 , n368193 );
buf ( n368195 , n368194 );
buf ( n368196 , n368195 );
nand ( n368197 , n47996 , n368196 );
buf ( n368198 , n368197 );
not ( n368199 , n368198 );
or ( n368200 , n368186 , n368199 );
buf ( n368201 , n365691 );
buf ( n368202 , n45553 );
nand ( n48008 , n368201 , n368202 );
buf ( n368204 , n48008 );
nand ( n368205 , n368200 , n368204 );
not ( n368206 , n368205 );
xor ( n48012 , n47178 , n367371 );
and ( n368208 , n48012 , n367397 );
and ( n368209 , n47178 , n367371 );
or ( n48015 , n368208 , n368209 );
buf ( n368211 , n48015 );
and ( n368212 , n368206 , n368211 );
not ( n48018 , n368206 );
not ( n48019 , n368211 );
and ( n368215 , n48018 , n48019 );
nor ( n368216 , n368212 , n368215 );
buf ( n368217 , n42242 );
not ( n368218 , n368217 );
buf ( n368219 , n366209 );
not ( n368220 , n368219 );
buf ( n368221 , n45718 );
not ( n48027 , n368221 );
or ( n368223 , n368220 , n48027 );
buf ( n368224 , n362133 );
buf ( n368225 , n366212 );
nand ( n368226 , n368224 , n368225 );
buf ( n368227 , n368226 );
buf ( n368228 , n368227 );
nand ( n368229 , n368223 , n368228 );
buf ( n368230 , n368229 );
buf ( n368231 , n368230 );
not ( n368232 , n368231 );
or ( n48038 , n368218 , n368232 );
buf ( n368234 , n46041 );
not ( n368235 , n368234 );
buf ( n48041 , n42263 );
buf ( n48042 , n48041 );
nand ( n48043 , n368235 , n48042 );
buf ( n48044 , n48043 );
buf ( n48045 , n48044 );
nand ( n48046 , n48038 , n48045 );
buf ( n48047 , n48046 );
and ( n368243 , n367268 , n367291 );
buf ( n368244 , n368243 );
or ( n48050 , n368244 , n47129 );
buf ( n368246 , n366367 );
not ( n368247 , n368246 );
buf ( n368248 , n45204 );
not ( n48054 , n368248 );
or ( n368250 , n368247 , n48054 );
buf ( n48056 , n367284 );
nand ( n48057 , n368250 , n48056 );
buf ( n48058 , n48057 );
buf ( n368254 , n48058 );
buf ( n368255 , n367264 );
nand ( n48061 , n368254 , n368255 );
buf ( n368257 , n48061 );
nand ( n368258 , n48050 , n368257 );
xor ( n368259 , n48047 , n368258 );
buf ( n368260 , n45993 );
not ( n48066 , n368260 );
buf ( n368262 , n366161 );
not ( n368263 , n368262 );
or ( n368264 , n48066 , n368263 );
buf ( n368265 , n364827 );
not ( n368266 , n368265 );
buf ( n368267 , n45270 );
not ( n48073 , n368267 );
or ( n48074 , n368266 , n48073 );
buf ( n48075 , n365471 );
buf ( n48076 , n44661 );
nand ( n48077 , n48075 , n48076 );
buf ( n48078 , n48077 );
buf ( n368274 , n48078 );
nand ( n368275 , n48074 , n368274 );
buf ( n368276 , n368275 );
buf ( n368277 , n368276 );
buf ( n48083 , n360574 );
nand ( n48084 , n368277 , n48083 );
buf ( n48085 , n48084 );
buf ( n368281 , n48085 );
nand ( n48087 , n368264 , n368281 );
buf ( n368283 , n48087 );
buf ( n368284 , n368283 );
buf ( n368285 , n367309 );
not ( n368286 , n368285 );
buf ( n368287 , n360164 );
buf ( n368288 , n360048 );
and ( n48094 , n368287 , n368288 );
buf ( n368290 , n48094 );
buf ( n368291 , n368290 );
not ( n48097 , n368291 );
or ( n48098 , n368286 , n48097 );
buf ( n368294 , n365486 );
buf ( n368295 , n45300 );
not ( n48101 , n368295 );
buf ( n368297 , n363116 );
not ( n368298 , n368297 );
or ( n48104 , n48101 , n368298 );
buf ( n368300 , n365495 );
buf ( n368301 , n365474 );
nand ( n368302 , n368300 , n368301 );
buf ( n368303 , n368302 );
buf ( n368304 , n368303 );
nand ( n368305 , n48104 , n368304 );
buf ( n368306 , n368305 );
buf ( n368307 , n368306 );
nand ( n368308 , n368294 , n368307 );
buf ( n368309 , n368308 );
buf ( n368310 , n368309 );
nand ( n48116 , n48098 , n368310 );
buf ( n48117 , n48116 );
buf ( n368313 , n48117 );
not ( n48119 , n368313 );
buf ( n368315 , n48119 );
buf ( n368316 , n368315 );
and ( n48122 , n368284 , n368316 );
not ( n48123 , n368284 );
buf ( n368319 , n48117 );
and ( n368320 , n48123 , n368319 );
nor ( n48126 , n48122 , n368320 );
buf ( n368322 , n48126 );
buf ( n368323 , n368322 );
buf ( n368324 , n366515 );
not ( n48130 , n368324 );
buf ( n368326 , n361606 );
not ( n48132 , n368326 );
or ( n48133 , n48130 , n48132 );
buf ( n368329 , n361531 );
not ( n368330 , n368329 );
buf ( n368331 , n363546 );
not ( n368332 , n368331 );
or ( n368333 , n368330 , n368332 );
buf ( n368334 , n361716 );
buf ( n368335 , n44717 );
nand ( n48141 , n368334 , n368335 );
buf ( n48142 , n48141 );
buf ( n368338 , n48142 );
nand ( n48144 , n368333 , n368338 );
buf ( n368340 , n48144 );
buf ( n368341 , n368340 );
buf ( n368342 , n361625 );
nand ( n48148 , n368341 , n368342 );
buf ( n48149 , n48148 );
buf ( n368345 , n48149 );
nand ( n48151 , n48133 , n368345 );
buf ( n48152 , n48151 );
buf ( n368348 , n48152 );
and ( n48154 , n368323 , n368348 );
not ( n48155 , n368323 );
buf ( n368351 , n48152 );
not ( n368352 , n368351 );
buf ( n368353 , n368352 );
buf ( n368354 , n368353 );
and ( n48160 , n48155 , n368354 );
nor ( n48161 , n48154 , n48160 );
buf ( n368357 , n48161 );
xnor ( n368358 , n368259 , n368357 );
and ( n48164 , n368216 , n368358 );
not ( n368360 , n368216 );
not ( n48166 , n368358 );
and ( n368362 , n368360 , n48166 );
nor ( n48168 , n48164 , n368362 );
and ( n368364 , n368185 , n48168 );
not ( n368365 , n368185 );
buf ( n368366 , n48168 );
not ( n368367 , n368366 );
buf ( n368368 , n368367 );
and ( n368369 , n368365 , n368368 );
nor ( n48175 , n368364 , n368369 );
buf ( n368371 , n48175 );
not ( n368372 , n368371 );
buf ( n368373 , n368372 );
buf ( n368374 , n368373 );
not ( n368375 , n368374 );
buf ( n368376 , n368375 );
buf ( n368377 , n368376 );
and ( n48183 , n368093 , n368377 );
not ( n368379 , n368093 );
buf ( n368380 , n368373 );
and ( n368381 , n368379 , n368380 );
nor ( n48187 , n48183 , n368381 );
buf ( n368383 , n48187 );
buf ( n368384 , n368383 );
not ( n368385 , n368384 );
buf ( n368386 , n368385 );
not ( n48192 , n368386 );
or ( n368388 , n367988 , n48192 );
buf ( n368389 , n368383 );
buf ( n368390 , n47791 );
nand ( n48196 , n368389 , n368390 );
buf ( n368392 , n48196 );
nand ( n48198 , n368388 , n368392 );
buf ( n368394 , n48198 );
xor ( n48200 , n367079 , n368394 );
and ( n48201 , n367409 , n367191 );
not ( n368397 , n367409 );
and ( n368398 , n368397 , n367194 );
or ( n368399 , n48201 , n368398 );
not ( n48205 , n367711 );
and ( n48206 , n368399 , n48205 );
not ( n48207 , n368399 );
not ( n368403 , n48205 );
and ( n48209 , n48207 , n368403 );
nor ( n48210 , n48206 , n48209 );
and ( n368406 , n47509 , n47487 );
not ( n368407 , n47509 );
and ( n48213 , n368407 , n47486 );
nor ( n368409 , n368406 , n48213 );
and ( n368410 , n368409 , n47516 );
not ( n48216 , n368409 );
and ( n48217 , n48216 , n367705 );
nor ( n368413 , n368410 , n48217 );
not ( n368414 , n368413 );
buf ( n368415 , n365428 );
not ( n368416 , n368415 );
buf ( n368417 , n359947 );
not ( n368418 , n368417 );
or ( n48224 , n368416 , n368418 );
buf ( n48225 , n361762 );
buf ( n368421 , n365422 );
nand ( n368422 , n48225 , n368421 );
buf ( n368423 , n368422 );
buf ( n368424 , n368423 );
nand ( n368425 , n48224 , n368424 );
buf ( n368426 , n368425 );
buf ( n368427 , n368426 );
not ( n368428 , n368427 );
buf ( n368429 , n366226 );
not ( n368430 , n368429 );
or ( n48236 , n368428 , n368430 );
buf ( n368432 , n359993 );
buf ( n368433 , n367428 );
nand ( n48239 , n368432 , n368433 );
buf ( n368435 , n48239 );
buf ( n368436 , n368435 );
nand ( n368437 , n48236 , n368436 );
buf ( n368438 , n368437 );
buf ( n368439 , n368438 );
not ( n368440 , n368439 );
buf ( n368441 , n366402 );
not ( n368442 , n368441 );
buf ( n48248 , n22710 );
not ( n48249 , n48248 );
buf ( n48250 , n44783 );
not ( n48251 , n48250 );
or ( n48252 , n48249 , n48251 );
buf ( n368448 , n41607 );
buf ( n368449 , n342657 );
nand ( n368450 , n368448 , n368449 );
buf ( n368451 , n368450 );
buf ( n368452 , n368451 );
nand ( n368453 , n48252 , n368452 );
buf ( n368454 , n368453 );
buf ( n368455 , n368454 );
not ( n368456 , n368455 );
or ( n48262 , n368442 , n368456 );
buf ( n368458 , n367466 );
buf ( n368459 , n366428 );
nand ( n368460 , n368458 , n368459 );
buf ( n368461 , n368460 );
buf ( n368462 , n368461 );
nand ( n48268 , n48262 , n368462 );
buf ( n368464 , n48268 );
buf ( n368465 , n368464 );
not ( n368466 , n368465 );
or ( n48272 , n368440 , n368466 );
or ( n48273 , n368464 , n368438 );
not ( n368469 , n45492 );
not ( n368470 , n366825 );
or ( n48276 , n368469 , n368470 );
buf ( n368472 , n360885 );
not ( n368473 , n368472 );
buf ( n368474 , n368473 );
and ( n48280 , n368474 , n365676 );
not ( n48281 , n368474 );
and ( n368477 , n48281 , n365673 );
or ( n368478 , n48280 , n368477 );
nand ( n48284 , n45553 , n368478 );
nand ( n48285 , n48276 , n48284 );
nand ( n48286 , n48273 , n48285 );
buf ( n368482 , n48286 );
nand ( n368483 , n48272 , n368482 );
buf ( n368484 , n368483 );
not ( n368485 , n368484 );
not ( n368486 , n368485 );
not ( n48292 , n368486 );
not ( n368488 , n367491 );
not ( n48294 , n365152 );
or ( n368490 , n368488 , n48294 );
buf ( n368491 , n342909 );
buf ( n368492 , n39830 );
and ( n48298 , n368491 , n368492 );
not ( n48299 , n368491 );
buf ( n48300 , n365206 );
and ( n368496 , n48299 , n48300 );
nor ( n48302 , n48298 , n368496 );
buf ( n48303 , n48302 );
not ( n368499 , n48303 );
nand ( n48305 , n368499 , n47290 );
nand ( n368501 , n368490 , n48305 );
not ( n368502 , n368501 );
or ( n48308 , n48292 , n368502 );
not ( n48309 , n368485 );
not ( n368505 , n368501 );
not ( n368506 , n368505 );
or ( n48312 , n48309 , n368506 );
buf ( n368508 , n44915 );
not ( n368509 , n368508 );
buf ( n368510 , n367667 );
not ( n368511 , n368510 );
or ( n48317 , n368509 , n368511 );
buf ( n368513 , n365041 );
not ( n48319 , n368513 );
buf ( n368515 , n363866 );
not ( n368516 , n368515 );
or ( n48322 , n48319 , n368516 );
buf ( n368518 , n365167 );
buf ( n368519 , n365052 );
nand ( n48325 , n368518 , n368519 );
buf ( n368521 , n48325 );
buf ( n368522 , n368521 );
nand ( n48328 , n48322 , n368522 );
buf ( n368524 , n48328 );
buf ( n368525 , n368524 );
buf ( n368526 , n47466 );
nand ( n368527 , n368525 , n368526 );
buf ( n368528 , n368527 );
buf ( n368529 , n368528 );
nand ( n368530 , n48317 , n368529 );
buf ( n368531 , n368530 );
buf ( n368532 , n368531 );
nand ( n368533 , n48312 , n368532 );
nand ( n368534 , n48308 , n368533 );
not ( n368535 , n368534 );
xor ( n368536 , n367632 , n47308 );
xor ( n368537 , n368536 , n367476 );
nand ( n368538 , n368535 , n368537 );
not ( n48338 , n368538 );
or ( n368540 , n368414 , n48338 );
not ( n368541 , n368537 );
nand ( n48341 , n368534 , n368541 );
nand ( n368543 , n368540 , n48341 );
not ( n48343 , n368543 );
not ( n48344 , n365047 );
buf ( n48345 , n48344 );
not ( n368547 , n48345 );
buf ( n368548 , n368547 );
buf ( n368549 , n23034 );
and ( n368550 , n368548 , n368549 );
not ( n48350 , n368548 );
buf ( n368552 , n368549 );
not ( n48352 , n368552 );
buf ( n368554 , n48352 );
and ( n48354 , n48350 , n368554 );
or ( n48355 , n368550 , n48354 );
xor ( n48356 , n22484 , n23034 );
buf ( n368558 , n48356 );
buf ( n368559 , n343193 );
not ( n48359 , n368559 );
buf ( n368561 , n48359 );
buf ( n368562 , n368561 );
not ( n368563 , n368562 );
buf ( n368564 , n368563 );
buf ( n368565 , n368564 );
not ( n368566 , n368565 );
buf ( n368567 , n22484 );
not ( n48367 , n368567 );
buf ( n368569 , n48367 );
buf ( n368570 , n368569 );
not ( n368571 , n368570 );
or ( n48371 , n368566 , n368571 );
buf ( n368573 , n22484 );
buf ( n368574 , n343179 );
buf ( n368575 , n343186 );
and ( n368576 , n368574 , n368575 );
not ( n368577 , n368574 );
buf ( n368578 , n343183 );
and ( n368579 , n368577 , n368578 );
nor ( n48379 , n368576 , n368579 );
buf ( n368581 , n48379 );
buf ( n368582 , n368581 );
not ( n48382 , n368582 );
buf ( n368584 , n48382 );
buf ( n368585 , n368584 );
nand ( n368586 , n368573 , n368585 );
buf ( n368587 , n368586 );
buf ( n368588 , n368587 );
nand ( n368589 , n48371 , n368588 );
buf ( n368590 , n368589 );
buf ( n368591 , n368590 );
not ( n368592 , n368591 );
buf ( n368593 , n368592 );
buf ( n368594 , n368593 );
nand ( n48394 , n368558 , n368594 );
buf ( n368596 , n48394 );
buf ( n48396 , n368596 );
not ( n368598 , n48396 );
buf ( n368599 , n368598 );
buf ( n368600 , n368599 );
buf ( n368601 , n368600 );
buf ( n368602 , n368601 );
buf ( n368603 , n368602 );
not ( n368604 , n368603 );
buf ( n368605 , n368604 );
buf ( n368606 , n368605 );
not ( n368607 , n368606 );
buf ( n368608 , n368607 );
buf ( n368609 , n368608 );
buf ( n368610 , n368609 );
buf ( n368611 , n368610 );
buf ( n368612 , n368611 );
not ( n368613 , n368612 );
buf ( n368614 , n368613 );
buf ( n368615 , n368614 );
not ( n48415 , n368564 );
not ( n368617 , n368569 );
or ( n48417 , n48415 , n368617 );
nand ( n48418 , n48417 , n368587 );
not ( n368620 , n48418 );
not ( n368621 , n368620 );
buf ( n368622 , n368621 );
not ( n368623 , n368622 );
buf ( n368624 , n368623 );
buf ( n368625 , n368624 );
nand ( n368626 , n368615 , n368625 );
buf ( n368627 , n368626 );
nand ( n48427 , n48355 , n368627 );
not ( n48428 , n48427 );
not ( n368630 , n365033 );
buf ( n368631 , n44819 );
not ( n48431 , n368631 );
buf ( n368633 , n366725 );
not ( n368634 , n368633 );
or ( n48434 , n48431 , n368634 );
buf ( n368636 , n364994 );
buf ( n368637 , n40275 );
nand ( n48437 , n368636 , n368637 );
buf ( n368639 , n48437 );
buf ( n368640 , n368639 );
nand ( n368641 , n48434 , n368640 );
buf ( n368642 , n368641 );
not ( n48442 , n368642 );
or ( n368644 , n368630 , n48442 );
nand ( n368645 , n46910 , n365118 );
nand ( n48445 , n368644 , n368645 );
not ( n368647 , n48445 );
or ( n368648 , n48428 , n368647 );
not ( n48448 , n48445 );
not ( n368650 , n48448 );
not ( n368651 , n48427 );
not ( n48451 , n368651 );
or ( n48452 , n368650 , n48451 );
buf ( n368654 , n352314 );
buf ( n368655 , n368654 );
buf ( n368656 , n368655 );
buf ( n368657 , n368656 );
not ( n48457 , n368657 );
buf ( n48458 , n48457 );
buf ( n48459 , n48458 );
buf ( n368661 , n48459 );
buf ( n368662 , n368661 );
buf ( n368663 , n368662 );
not ( n368664 , n368663 );
buf ( n368665 , n368664 );
buf ( n368666 , n368665 );
not ( n368667 , n368666 );
buf ( n368668 , n361631 );
not ( n48468 , n368668 );
or ( n368670 , n368667 , n48468 );
buf ( n368671 , n39621 );
buf ( n368672 , n368662 );
nand ( n368673 , n368671 , n368672 );
buf ( n368674 , n368673 );
buf ( n368675 , n368674 );
nand ( n48475 , n368670 , n368675 );
buf ( n368677 , n48475 );
buf ( n368678 , n368677 );
not ( n48478 , n368678 );
buf ( n368680 , n359809 );
not ( n368681 , n368680 );
or ( n368682 , n48478 , n368681 );
buf ( n368683 , n362521 );
buf ( n368684 , n45244 );
nand ( n368685 , n368683 , n368684 );
buf ( n368686 , n368685 );
buf ( n368687 , n368686 );
nand ( n368688 , n368682 , n368687 );
buf ( n368689 , n368688 );
not ( n368690 , n47370 );
not ( n48490 , n362385 );
not ( n368692 , n48490 );
or ( n48492 , n368690 , n368692 );
not ( n48493 , n365918 );
not ( n368695 , n364774 );
or ( n368696 , n48493 , n368695 );
not ( n48496 , n31728 );
buf ( n368698 , n48496 );
not ( n368699 , n368698 );
buf ( n368700 , n368699 );
or ( n368701 , n368700 , n362420 );
nand ( n368702 , n368696 , n368701 );
buf ( n48502 , n42259 );
buf ( n368704 , n48502 );
not ( n368705 , n368704 );
buf ( n368706 , n368705 );
nand ( n48506 , n368702 , n368706 );
nand ( n368708 , n48492 , n48506 );
not ( n368709 , n368708 );
buf ( n368710 , n364766 );
not ( n368711 , n368710 );
buf ( n368712 , n366131 );
not ( n48512 , n368712 );
and ( n368714 , n368711 , n48512 );
buf ( n368715 , n364744 );
buf ( n368716 , n364870 );
and ( n48516 , n368715 , n368716 );
nor ( n48517 , n368714 , n48516 );
buf ( n368719 , n48517 );
not ( n368720 , n368719 );
not ( n48520 , n361971 );
and ( n48521 , n368720 , n48520 );
buf ( n368723 , n365335 );
not ( n368724 , n366339 );
buf ( n368725 , n368724 );
and ( n368726 , n368723 , n368725 );
buf ( n368727 , n368726 );
nor ( n48527 , n48521 , n368727 );
not ( n368729 , n48527 );
not ( n368730 , n368729 );
or ( n48530 , n368709 , n368730 );
not ( n48531 , n368708 );
not ( n368733 , n48531 );
not ( n368734 , n48527 );
or ( n48534 , n368733 , n368734 );
buf ( n368736 , n365440 );
not ( n368737 , n368736 );
buf ( n368738 , n365290 );
not ( n48538 , n368738 );
or ( n368740 , n368737 , n48538 );
buf ( n368741 , n365569 );
buf ( n368742 , n365452 );
nand ( n48542 , n368741 , n368742 );
buf ( n368744 , n48542 );
buf ( n368745 , n368744 );
nand ( n368746 , n368740 , n368745 );
buf ( n368747 , n368746 );
not ( n368748 , n368747 );
not ( n368749 , n365279 );
or ( n48549 , n368748 , n368749 );
buf ( n368751 , n40923 );
buf ( n368752 , n367607 );
nand ( n48552 , n368751 , n368752 );
buf ( n48553 , n48552 );
nand ( n368755 , n48549 , n48553 );
nand ( n368756 , n48534 , n368755 );
nand ( n48556 , n48530 , n368756 );
xor ( n368758 , n368689 , n48556 );
not ( n48558 , n362385 );
not ( n368760 , n48558 );
not ( n368761 , n368702 );
or ( n48561 , n368760 , n368761 );
buf ( n368763 , n362417 );
not ( n48563 , n368763 );
buf ( n368765 , n48563 );
buf ( n368766 , n368765 );
buf ( n48566 , n365329 );
and ( n48567 , n368766 , n48566 );
not ( n48568 , n368766 );
buf ( n368770 , n45152 );
and ( n48570 , n48568 , n368770 );
nor ( n48571 , n48567 , n48570 );
buf ( n368773 , n48571 );
not ( n48573 , n368773 );
buf ( n368775 , n362405 );
not ( n368776 , n368775 );
buf ( n368777 , n368776 );
not ( n368778 , n368777 );
nand ( n368779 , n48573 , n368778 );
nand ( n48579 , n48561 , n368779 );
buf ( n368781 , n48579 );
buf ( n368782 , n352212 );
not ( n48582 , n368782 );
buf ( n368784 , n365626 );
not ( n368785 , n368784 );
or ( n48585 , n48582 , n368785 );
buf ( n368787 , n45455 );
buf ( n368788 , n365259 );
nand ( n368789 , n368787 , n368788 );
buf ( n368790 , n368789 );
buf ( n368791 , n368790 );
nand ( n368792 , n48585 , n368791 );
buf ( n368793 , n368792 );
buf ( n368794 , n368793 );
not ( n368795 , n368794 );
buf ( n368796 , n364797 );
not ( n368797 , n368796 );
or ( n48597 , n368795 , n368797 );
buf ( n368799 , n46678 );
buf ( n368800 , n41918 );
nand ( n48600 , n368799 , n368800 );
buf ( n368802 , n48600 );
buf ( n368803 , n368802 );
nand ( n48603 , n48597 , n368803 );
buf ( n48604 , n48603 );
buf ( n368806 , n48604 );
xor ( n48606 , n368781 , n368806 );
buf ( n368808 , n364852 );
buf ( n368809 , n365561 );
not ( n48609 , n368809 );
buf ( n368811 , n366086 );
not ( n368812 , n368811 );
or ( n368813 , n48609 , n368812 );
buf ( n368814 , n45414 );
buf ( n368815 , n351318 );
nand ( n368816 , n368814 , n368815 );
buf ( n368817 , n368816 );
buf ( n368818 , n368817 );
nand ( n368819 , n368813 , n368818 );
buf ( n368820 , n368819 );
buf ( n368821 , n368820 );
not ( n368822 , n368821 );
buf ( n368823 , n368822 );
buf ( n368824 , n368823 );
or ( n48624 , n368808 , n368824 );
buf ( n368826 , n47396 );
not ( n368827 , n368826 );
buf ( n368828 , n368827 );
buf ( n368829 , n368828 );
buf ( n368830 , n361626 );
or ( n48630 , n368829 , n368830 );
nand ( n48631 , n48624 , n48630 );
buf ( n368833 , n48631 );
buf ( n368834 , n368833 );
and ( n48634 , n48606 , n368834 );
and ( n368836 , n368781 , n368806 );
or ( n368837 , n48634 , n368836 );
buf ( n368838 , n368837 );
and ( n368839 , n368758 , n368838 );
and ( n368840 , n368689 , n48556 );
or ( n48640 , n368839 , n368840 );
nand ( n368842 , n48452 , n48640 );
nand ( n48642 , n368648 , n368842 );
buf ( n368844 , n46950 );
not ( n368845 , n368844 );
buf ( n368846 , n367133 );
not ( n48646 , n368846 );
and ( n368848 , n368845 , n48646 );
buf ( n48648 , n367133 );
buf ( n368850 , n46950 );
and ( n368851 , n48648 , n368850 );
nor ( n368852 , n368848 , n368851 );
buf ( n368853 , n368852 );
not ( n368854 , n367105 );
and ( n48654 , n368853 , n368854 );
not ( n368856 , n368853 );
and ( n48656 , n368856 , n367105 );
nor ( n368858 , n48654 , n48656 );
or ( n48658 , n48642 , n368858 );
buf ( n48659 , n366713 );
and ( n368861 , n48659 , n46548 );
not ( n368862 , n48659 );
and ( n48662 , n368862 , n46549 );
nor ( n368864 , n368861 , n48662 );
and ( n368865 , n368864 , n366779 );
not ( n48665 , n368864 );
not ( n368867 , n366779 );
and ( n368868 , n48665 , n368867 );
nor ( n48668 , n368865 , n368868 );
nand ( n48669 , n48658 , n48668 );
buf ( n48670 , n48669 );
nand ( n48671 , n48642 , n368858 );
buf ( n48672 , n48671 );
nand ( n48673 , n48670 , n48672 );
buf ( n48674 , n48673 );
not ( n368876 , n48674 );
xor ( n48676 , n367141 , n46960 );
xor ( n368878 , n48676 , n367187 );
buf ( n368879 , n368878 );
not ( n48679 , n368879 );
nand ( n48680 , n368876 , n48679 );
not ( n368882 , n48680 );
or ( n368883 , n48343 , n368882 );
nand ( n48683 , n48674 , n368879 );
nand ( n48684 , n368883 , n48683 );
not ( n368886 , n48684 );
nand ( n48686 , n48210 , n368886 );
buf ( n368888 , n48686 );
not ( n48688 , n368888 );
and ( n48689 , n46848 , n366846 );
not ( n368891 , n46848 );
and ( n368892 , n368891 , n366843 );
or ( n48692 , n48689 , n368892 );
and ( n368894 , n48692 , n366851 );
not ( n368895 , n48692 );
and ( n48695 , n368895 , n367044 );
nor ( n368897 , n368894 , n48695 );
not ( n48697 , n368897 );
xor ( n48698 , n367539 , n367522 );
not ( n48699 , n48698 );
not ( n48700 , n367622 );
not ( n48701 , n48700 );
and ( n48702 , n48699 , n48701 );
and ( n368904 , n48698 , n48700 );
nor ( n48704 , n48702 , n368904 );
not ( n368906 , n48704 );
buf ( n368907 , n45075 );
not ( n48707 , n368907 );
buf ( n368909 , n367691 );
not ( n368910 , n368909 );
or ( n48710 , n48707 , n368910 );
buf ( n368912 , n342881 );
not ( n48712 , n368912 );
buf ( n368914 , n365681 );
not ( n368915 , n368914 );
or ( n48715 , n48712 , n368915 );
buf ( n368917 , n359778 );
buf ( n368918 , n365202 );
nand ( n48718 , n368917 , n368918 );
buf ( n368920 , n48718 );
buf ( n368921 , n368920 );
nand ( n48721 , n48715 , n368921 );
buf ( n368923 , n48721 );
buf ( n368924 , n368923 );
buf ( n368925 , n45058 );
nand ( n48725 , n368924 , n368925 );
buf ( n368927 , n48725 );
buf ( n368928 , n368927 );
nand ( n368929 , n48710 , n368928 );
buf ( n368930 , n368929 );
not ( n48730 , n368930 );
or ( n368932 , n368906 , n48730 );
not ( n368933 , n48700 );
and ( n48733 , n48698 , n368933 );
not ( n48734 , n48698 );
and ( n48735 , n48734 , n48700 );
nor ( n48736 , n48733 , n48735 );
not ( n48737 , n48736 );
not ( n48738 , n368930 );
not ( n368940 , n48738 );
or ( n48740 , n48737 , n368940 );
buf ( n368942 , n365980 );
not ( n48742 , n368942 );
buf ( n368944 , n365945 );
not ( n368945 , n368944 );
or ( n48745 , n48742 , n368945 );
buf ( n368947 , n365507 );
buf ( n368948 , n365989 );
nand ( n368949 , n368947 , n368948 );
buf ( n368950 , n368949 );
buf ( n368951 , n368950 );
nand ( n368952 , n48745 , n368951 );
buf ( n368953 , n368952 );
buf ( n368954 , n368953 );
not ( n48754 , n368954 );
buf ( n368956 , n368290 );
not ( n368957 , n368956 );
or ( n368958 , n48754 , n368957 );
buf ( n368959 , n367013 );
buf ( n368960 , n365954 );
nand ( n368961 , n368959 , n368960 );
buf ( n368962 , n368961 );
buf ( n368963 , n368962 );
nand ( n368964 , n368958 , n368963 );
buf ( n368965 , n368964 );
buf ( n368966 , n368965 );
not ( n48766 , n368966 );
buf ( n368968 , n48766 );
not ( n48768 , n368968 );
not ( n48769 , n43261 );
not ( n368971 , n46701 );
or ( n48771 , n48769 , n368971 );
not ( n368973 , n342719 );
buf ( n368974 , n362534 );
not ( n48774 , n368974 );
buf ( n368976 , n48774 );
not ( n368977 , n368976 );
or ( n48777 , n368973 , n368977 );
buf ( n368979 , n362534 );
buf ( n368980 , n364953 );
nand ( n48780 , n368979 , n368980 );
buf ( n48781 , n48780 );
nand ( n368983 , n48777 , n48781 );
buf ( n368984 , n368983 );
buf ( n368985 , n44796 );
nand ( n368986 , n368984 , n368985 );
buf ( n368987 , n368986 );
nand ( n48787 , n48771 , n368987 );
not ( n368989 , n48787 );
not ( n368990 , n368989 );
or ( n48790 , n48768 , n368990 );
buf ( n48791 , n31009 );
not ( n48792 , n48791 );
buf ( n368994 , n48792 );
not ( n368995 , n368994 );
nand ( n48795 , n368995 , n366534 );
nand ( n368997 , n368994 , n361631 );
nand ( n368998 , n48795 , n368997 );
buf ( n368999 , n368998 );
not ( n369000 , n368999 );
buf ( n369001 , n359809 );
not ( n48801 , n369001 );
or ( n48802 , n369000 , n48801 );
buf ( n369004 , n362521 );
buf ( n369005 , n368677 );
nand ( n48805 , n369004 , n369005 );
buf ( n48806 , n48805 );
buf ( n369008 , n48806 );
nand ( n48808 , n48802 , n369008 );
buf ( n369010 , n48808 );
nand ( n48810 , n48790 , n369010 );
nand ( n369012 , n48787 , n368965 );
nand ( n48812 , n48810 , n369012 );
xor ( n48813 , n47381 , n367595 );
xor ( n369015 , n48813 , n367618 );
buf ( n369016 , n369015 );
xor ( n369017 , n48812 , n369016 );
buf ( n369018 , n365033 );
not ( n369019 , n369018 );
buf ( n369020 , n44819 );
not ( n48820 , n369020 );
not ( n369022 , n40251 );
buf ( n369023 , n369022 );
not ( n48823 , n369023 );
or ( n369025 , n48820 , n48823 );
buf ( n369026 , n364994 );
buf ( n369027 , n40251 );
nand ( n369028 , n369026 , n369027 );
buf ( n369029 , n369028 );
buf ( n369030 , n369029 );
nand ( n48830 , n369025 , n369030 );
buf ( n48831 , n48830 );
buf ( n369033 , n48831 );
not ( n48833 , n369033 );
or ( n369035 , n369019 , n48833 );
buf ( n369036 , n368642 );
buf ( n369037 , n365118 );
nand ( n369038 , n369036 , n369037 );
buf ( n369039 , n369038 );
buf ( n369040 , n369039 );
nand ( n369041 , n369035 , n369040 );
buf ( n369042 , n369041 );
and ( n48842 , n369017 , n369042 );
and ( n369044 , n48812 , n369016 );
or ( n369045 , n48842 , n369044 );
nand ( n369046 , n48740 , n369045 );
nand ( n48846 , n368932 , n369046 );
xor ( n369048 , n47254 , n367444 );
xor ( n48848 , n369048 , n367473 );
buf ( n369050 , n48848 );
not ( n369051 , n369050 );
buf ( n369052 , n369051 );
buf ( n369053 , n369052 );
not ( n369054 , n369053 );
buf ( n369055 , n46751 );
buf ( n369056 , n366964 );
xor ( n369057 , n369055 , n369056 );
buf ( n369058 , n367034 );
xor ( n369059 , n369057 , n369058 );
buf ( n369060 , n369059 );
buf ( n369061 , n369060 );
not ( n48861 , n369061 );
or ( n369063 , n369054 , n48861 );
buf ( n48863 , n365337 );
buf ( n369065 , n366994 );
xor ( n369066 , n48863 , n369065 );
buf ( n369067 , n367025 );
xnor ( n48867 , n369066 , n369067 );
buf ( n48868 , n48867 );
buf ( n48869 , n48868 );
xor ( n48870 , n366879 , n46721 );
xor ( n369072 , n48870 , n46747 );
buf ( n369073 , n369072 );
buf ( n369074 , n369073 );
xor ( n369075 , n48869 , n369074 );
buf ( n369076 , n366654 );
not ( n48876 , n369076 );
buf ( n369078 , n366954 );
not ( n369079 , n369078 );
or ( n369080 , n48876 , n369079 );
buf ( n369081 , n46477 );
not ( n369082 , n369081 );
buf ( n369083 , n362133 );
not ( n48883 , n369083 );
buf ( n369085 , n48883 );
buf ( n369086 , n369085 );
not ( n369087 , n369086 );
or ( n48887 , n369082 , n369087 );
buf ( n369089 , n362136 );
buf ( n369090 , n366683 );
nand ( n369091 , n369089 , n369090 );
buf ( n369092 , n369091 );
buf ( n369093 , n369092 );
nand ( n369094 , n48887 , n369093 );
buf ( n369095 , n369094 );
buf ( n369096 , n369095 );
buf ( n369097 , n46521 );
nand ( n369098 , n369096 , n369097 );
buf ( n369099 , n369098 );
buf ( n369100 , n369099 );
nand ( n369101 , n369080 , n369100 );
buf ( n369102 , n369101 );
buf ( n369103 , n369102 );
and ( n369104 , n369075 , n369103 );
and ( n48904 , n48869 , n369074 );
or ( n48905 , n369104 , n48904 );
buf ( n369107 , n48905 );
buf ( n369108 , n369107 );
nand ( n369109 , n369063 , n369108 );
buf ( n369110 , n369109 );
buf ( n369111 , n369060 );
not ( n48911 , n369111 );
buf ( n369113 , n48911 );
buf ( n48913 , n369113 );
buf ( n48914 , n48848 );
nand ( n48915 , n48913 , n48914 );
buf ( n48916 , n48915 );
nand ( n369118 , n369110 , n48916 );
nand ( n48918 , n48846 , n369118 );
not ( n369120 , n48918 );
or ( n369121 , n48697 , n369120 );
not ( n369122 , n369118 );
not ( n48922 , n48846 );
nand ( n369124 , n369122 , n48922 );
nand ( n48924 , n369121 , n369124 );
buf ( n369126 , n48924 );
not ( n48926 , n369126 );
buf ( n369128 , n48926 );
not ( n48928 , n369128 );
not ( n369130 , n47462 );
not ( n48930 , n47227 );
or ( n48931 , n369130 , n48930 );
nand ( n369133 , n47226 , n47455 );
nand ( n48933 , n48931 , n369133 );
not ( n369135 , n47521 );
and ( n48935 , n48933 , n369135 );
not ( n48936 , n48933 );
and ( n48937 , n48936 , n47521 );
nor ( n369139 , n48935 , n48937 );
not ( n48939 , n369139 );
not ( n369141 , n48939 );
or ( n48941 , n48928 , n369141 );
not ( n48942 , n369139 );
not ( n369144 , n48924 );
or ( n369145 , n48942 , n369144 );
xor ( n48945 , n366810 , n367051 );
xor ( n369147 , n48945 , n367069 );
buf ( n369148 , n369147 );
nand ( n48948 , n369145 , n369148 );
nand ( n369150 , n48941 , n48948 );
buf ( n369151 , n369150 );
not ( n48951 , n369151 );
or ( n369153 , n48688 , n48951 );
not ( n369154 , n48210 );
nand ( n48954 , n369154 , n48684 );
buf ( n369156 , n48954 );
nand ( n369157 , n369153 , n369156 );
buf ( n369158 , n369157 );
buf ( n369159 , n369158 );
not ( n369160 , n369159 );
buf ( n369161 , n369160 );
buf ( n369162 , n369161 );
xnor ( n369163 , n48200 , n369162 );
buf ( n369164 , n369163 );
xor ( n369165 , n365887 , n366805 );
xor ( n369166 , n369165 , n367074 );
buf ( n369167 , n369166 );
buf ( n369168 , n369167 );
not ( n48968 , n368879 );
not ( n48969 , n368876 );
or ( n48970 , n48968 , n48969 );
nand ( n48971 , n48679 , n48674 );
nand ( n48972 , n48970 , n48971 );
not ( n369174 , n368543 );
and ( n48974 , n48972 , n369174 );
not ( n369176 , n48972 );
and ( n48976 , n369176 , n368543 );
nor ( n48977 , n48974 , n48976 );
not ( n369179 , n44915 );
not ( n48979 , n368524 );
or ( n48980 , n369179 , n48979 );
not ( n369182 , n44913 );
not ( n369183 , n342965 );
not ( n48983 , n369183 );
and ( n369185 , n39860 , n48983 );
not ( n369186 , n39860 );
not ( n48986 , n365041 );
and ( n369188 , n369186 , n48986 );
or ( n48988 , n369185 , n369188 );
and ( n48989 , n359966 , n48988 );
not ( n369191 , n359966 );
not ( n369192 , n369183 );
and ( n48992 , n39863 , n369192 );
not ( n48993 , n39863 );
not ( n369195 , n365041 );
and ( n369196 , n48993 , n369195 );
or ( n48996 , n48992 , n369196 );
and ( n369198 , n369191 , n48996 );
or ( n369199 , n48989 , n369198 );
nand ( n48999 , n369182 , n369199 );
nand ( n49000 , n48980 , n48999 );
not ( n369202 , n49000 );
not ( n369203 , n45075 );
not ( n49003 , n368923 );
or ( n369205 , n369203 , n49003 );
buf ( n369206 , n342881 );
not ( n369207 , n369206 );
buf ( n369208 , n46902 );
not ( n369209 , n369208 );
or ( n49009 , n369207 , n369209 );
buf ( n369211 , n40199 );
buf ( n49011 , n365202 );
nand ( n49012 , n369211 , n49011 );
buf ( n49013 , n49012 );
buf ( n369215 , n49013 );
nand ( n49015 , n49009 , n369215 );
buf ( n369217 , n49015 );
buf ( n369218 , n369217 );
buf ( n369219 , n45058 );
nand ( n369220 , n369218 , n369219 );
buf ( n369221 , n369220 );
nand ( n49021 , n369205 , n369221 );
not ( n369223 , n49021 );
or ( n369224 , n369202 , n369223 );
nor ( n49024 , n49000 , n49021 );
not ( n369226 , n351229 );
not ( n49026 , n365471 );
or ( n49027 , n369226 , n49026 );
nand ( n49028 , n360613 , n31197 );
nand ( n369230 , n49027 , n49028 );
buf ( n369231 , n369230 );
not ( n49031 , n369231 );
buf ( n369233 , n40475 );
not ( n49033 , n369233 );
or ( n49034 , n49031 , n49033 );
buf ( n369236 , n366922 );
buf ( n369237 , n360574 );
nand ( n49037 , n369236 , n369237 );
buf ( n369239 , n49037 );
buf ( n369240 , n369239 );
nand ( n49040 , n49034 , n369240 );
buf ( n369242 , n49040 );
buf ( n369243 , n369242 );
buf ( n369244 , n351160 );
not ( n49044 , n369244 );
buf ( n369246 , n365368 );
not ( n49046 , n369246 );
or ( n49047 , n49044 , n49046 );
buf ( n369249 , n35548 );
buf ( n369250 , n364915 );
nand ( n49050 , n369249 , n369250 );
buf ( n369252 , n49050 );
buf ( n369253 , n369252 );
nand ( n369254 , n49047 , n369253 );
buf ( n369255 , n369254 );
buf ( n369256 , n369255 );
not ( n49056 , n369256 );
buf ( n369258 , n39207 );
not ( n49058 , n369258 );
buf ( n369260 , n49058 );
buf ( n369261 , n369260 );
not ( n49061 , n369261 );
or ( n49062 , n49056 , n49061 );
buf ( n369264 , n46582 );
buf ( n369265 , n366981 );
nand ( n49065 , n369264 , n369265 );
buf ( n369267 , n49065 );
buf ( n369268 , n369267 );
nand ( n49068 , n49062 , n369268 );
buf ( n369270 , n49068 );
buf ( n369271 , n369270 );
xor ( n49071 , n369243 , n369271 );
buf ( n369273 , n366434 );
not ( n369274 , n369273 );
buf ( n369275 , n368454 );
not ( n49075 , n369275 );
or ( n369277 , n369274 , n49075 );
buf ( n369278 , n22710 );
not ( n49078 , n369278 );
buf ( n369280 , n41528 );
not ( n49080 , n369280 );
buf ( n369282 , n49080 );
buf ( n369283 , n369282 );
not ( n49083 , n369283 );
or ( n49084 , n49078 , n49083 );
buf ( n369286 , n41528 );
buf ( n369287 , n342657 );
nand ( n49087 , n369286 , n369287 );
buf ( n369289 , n49087 );
buf ( n369290 , n369289 );
nand ( n49090 , n49084 , n369290 );
buf ( n369292 , n49090 );
buf ( n369293 , n369292 );
buf ( n369294 , n366402 );
nand ( n369295 , n369293 , n369294 );
buf ( n369296 , n369295 );
buf ( n369297 , n369296 );
nand ( n49097 , n369277 , n369297 );
buf ( n369299 , n49097 );
buf ( n369300 , n369299 );
and ( n49100 , n49071 , n369300 );
and ( n49101 , n369243 , n369271 );
or ( n49102 , n49100 , n49101 );
buf ( n369304 , n49102 );
buf ( n369305 , n369304 );
not ( n49105 , n369305 );
buf ( n369307 , n49105 );
or ( n49107 , n49024 , n369307 );
nand ( n49108 , n369224 , n49107 );
xor ( n369310 , n366831 , n366835 );
xor ( n49110 , n369310 , n366839 );
buf ( n369312 , n49110 );
xor ( n49112 , n49108 , n369312 );
xor ( n369314 , n368689 , n48556 );
xor ( n49114 , n369314 , n368838 );
not ( n369316 , n49114 );
buf ( n369317 , n368438 );
buf ( n369318 , n368464 );
xor ( n369319 , n369317 , n369318 );
buf ( n369320 , n48285 );
xnor ( n49120 , n369319 , n369320 );
buf ( n369322 , n49120 );
nand ( n49122 , n369316 , n369322 );
not ( n369324 , n49122 );
and ( n369325 , n48531 , n368729 );
not ( n49125 , n48531 );
and ( n49126 , n49125 , n48527 );
nor ( n49127 , n369325 , n49126 );
not ( n369329 , n368755 );
and ( n49129 , n49127 , n369329 );
not ( n369331 , n49127 );
and ( n49131 , n369331 , n368755 );
nor ( n49132 , n49129 , n49131 );
buf ( n369334 , n366654 );
not ( n49134 , n369334 );
buf ( n369336 , n369095 );
not ( n49136 , n369336 );
or ( n369338 , n49134 , n49136 );
buf ( n369339 , n46477 );
not ( n49139 , n369339 );
buf ( n369341 , n46031 );
not ( n49141 , n369341 );
buf ( n369343 , n49141 );
buf ( n369344 , n369343 );
not ( n49144 , n369344 );
or ( n49145 , n49139 , n49144 );
buf ( n369347 , n367453 );
buf ( n49147 , n369347 );
buf ( n369349 , n49147 );
buf ( n369350 , n369349 );
not ( n49150 , n369350 );
buf ( n369352 , n49150 );
buf ( n369353 , n369352 );
buf ( n49153 , n366683 );
nand ( n49154 , n369353 , n49153 );
buf ( n369356 , n49154 );
buf ( n369357 , n369356 );
nand ( n49157 , n49145 , n369357 );
buf ( n369359 , n49157 );
buf ( n369360 , n369359 );
buf ( n369361 , n46521 );
nand ( n49161 , n369360 , n369361 );
buf ( n369363 , n49161 );
buf ( n369364 , n369363 );
nand ( n369365 , n369338 , n369364 );
buf ( n369366 , n369365 );
xor ( n49166 , n49132 , n369366 );
not ( n49167 , n39592 );
not ( n49168 , n368998 );
or ( n369370 , n49167 , n49168 );
not ( n369371 , n42886 );
not ( n369372 , n352353 );
not ( n49172 , n369372 );
buf ( n369374 , n49172 );
not ( n49174 , n369374 );
not ( n369376 , n45231 );
or ( n49176 , n49174 , n369376 );
buf ( n369378 , n39621 );
not ( n49178 , n369374 );
buf ( n369380 , n49178 );
nand ( n369381 , n369378 , n369380 );
buf ( n369382 , n369381 );
nand ( n49182 , n49176 , n369382 );
nand ( n369384 , n369371 , n49182 );
nand ( n369385 , n369370 , n369384 );
buf ( n369386 , n45345 );
not ( n369387 , n369386 );
buf ( n369388 , n365428 );
not ( n49188 , n369388 );
buf ( n369390 , n363116 );
not ( n369391 , n369390 );
or ( n369392 , n49188 , n369391 );
buf ( n369393 , n363119 );
buf ( n369394 , n365422 );
nand ( n369395 , n369393 , n369394 );
buf ( n369396 , n369395 );
buf ( n369397 , n369396 );
nand ( n369398 , n369392 , n369397 );
buf ( n369399 , n369398 );
buf ( n369400 , n369399 );
not ( n49200 , n369400 );
or ( n49201 , n369387 , n49200 );
buf ( n369403 , n39949 );
buf ( n49203 , n368953 );
nand ( n49204 , n369403 , n49203 );
buf ( n369406 , n49204 );
buf ( n369407 , n369406 );
nand ( n49207 , n49201 , n369407 );
buf ( n369409 , n49207 );
xor ( n49209 , n369385 , n369409 );
not ( n49210 , n366356 );
not ( n369412 , n46303 );
or ( n369413 , n49210 , n369412 );
buf ( n369414 , n365353 );
buf ( n369415 , n44737 );
nand ( n369416 , n369414 , n369415 );
buf ( n369417 , n369416 );
nand ( n49217 , n369413 , n369417 );
not ( n369419 , n49217 );
not ( n369420 , n45204 );
or ( n49218 , n369419 , n369420 );
buf ( n369422 , n39217 );
buf ( n369423 , n369255 );
nand ( n369424 , n369422 , n369423 );
buf ( n369425 , n369424 );
nand ( n49223 , n49218 , n369425 );
and ( n369427 , n49209 , n49223 );
and ( n369428 , n369385 , n369409 );
or ( n369429 , n369427 , n369428 );
and ( n49227 , n49166 , n369429 );
and ( n369431 , n49132 , n369366 );
or ( n369432 , n49227 , n369431 );
not ( n49230 , n369432 );
or ( n49231 , n369324 , n49230 );
buf ( n49232 , n369322 );
not ( n49233 , n49232 );
buf ( n369437 , n49233 );
nand ( n369438 , n369437 , n49114 );
nand ( n369439 , n49231 , n369438 );
and ( n49237 , n49112 , n369439 );
and ( n369441 , n49108 , n369312 );
or ( n369442 , n49237 , n369441 );
buf ( n369443 , n369442 );
not ( n369444 , n368620 );
not ( n369445 , n369444 );
not ( n49243 , n48355 );
or ( n369447 , n369445 , n49243 );
and ( n369448 , n40090 , n368554 );
not ( n369449 , n40090 );
and ( n49247 , n369449 , n368549 );
or ( n369451 , n369448 , n49247 );
nand ( n49249 , n368611 , n369451 );
nand ( n49250 , n369447 , n49249 );
buf ( n369454 , n49250 );
not ( n369455 , n369454 );
buf ( n369456 , n365155 );
not ( n369457 , n369456 );
buf ( n369458 , n48303 );
not ( n49256 , n369458 );
and ( n369460 , n369457 , n49256 );
buf ( n369461 , n22959 );
not ( n49259 , n369461 );
buf ( n369463 , n362208 );
not ( n369464 , n369463 );
or ( n49262 , n49259 , n369464 );
buf ( n369466 , n342909 );
buf ( n49264 , n359756 );
nand ( n49265 , n369466 , n49264 );
buf ( n49266 , n49265 );
buf ( n49267 , n49266 );
nand ( n49268 , n49262 , n49267 );
buf ( n49269 , n49268 );
buf ( n369473 , n49269 );
buf ( n369474 , n47290 );
and ( n369475 , n369473 , n369474 );
nor ( n49273 , n369460 , n369475 );
buf ( n369477 , n49273 );
buf ( n369478 , n369477 );
not ( n49276 , n369478 );
buf ( n369480 , n49276 );
buf ( n369481 , n369480 );
not ( n49279 , n369481 );
or ( n369483 , n369455 , n49279 );
buf ( n369484 , n49250 );
not ( n369485 , n369484 );
buf ( n369486 , n369485 );
buf ( n369487 , n369486 );
not ( n49285 , n369487 );
buf ( n369489 , n369477 );
not ( n369490 , n369489 );
or ( n369491 , n49285 , n369490 );
buf ( n369492 , n368983 );
buf ( n369493 , n43261 );
nand ( n369494 , n369492 , n369493 );
buf ( n369495 , n369494 );
buf ( n369496 , n369495 );
buf ( n369497 , n46693 );
buf ( n369498 , n369497 );
not ( n49296 , n369498 );
buf ( n369500 , n32085 );
not ( n369501 , n369500 );
or ( n49299 , n49296 , n369501 );
not ( n369503 , n369497 );
nand ( n369504 , n369503 , n32084 );
buf ( n369505 , n369504 );
nand ( n369506 , n49299 , n369505 );
buf ( n369507 , n369506 );
nand ( n369508 , n363429 , n369507 );
buf ( n49306 , n369508 );
nand ( n369510 , n369496 , n49306 , n48579 );
not ( n49308 , n369510 );
buf ( n369512 , n45177 );
not ( n49310 , n369512 );
buf ( n369514 , n40891 );
not ( n49312 , n369514 );
or ( n49313 , n49310 , n49312 );
buf ( n369517 , n365293 );
buf ( n49315 , n365344 );
buf ( n49316 , n49315 );
nand ( n49317 , n369517 , n49316 );
buf ( n49318 , n49317 );
buf ( n49319 , n49318 );
nand ( n49320 , n49313 , n49319 );
buf ( n49321 , n49320 );
not ( n369525 , n49321 );
not ( n49323 , n361013 );
or ( n369527 , n369525 , n49323 );
buf ( n369528 , n40923 );
buf ( n369529 , n368747 );
nand ( n369530 , n369528 , n369529 );
buf ( n369531 , n369530 );
nand ( n369532 , n369527 , n369531 );
not ( n49330 , n369532 );
or ( n49331 , n49308 , n49330 );
not ( n369535 , n369508 );
not ( n49333 , n369495 );
or ( n369537 , n369535 , n49333 );
not ( n49335 , n48579 );
nand ( n369539 , n369537 , n49335 );
nand ( n369540 , n49331 , n369539 );
not ( n49338 , n369540 );
not ( n49339 , n366229 );
not ( n369543 , n49339 );
buf ( n369544 , n365408 );
buf ( n369545 , n366243 );
and ( n369546 , n369544 , n369545 );
not ( n369547 , n369544 );
buf ( n369548 , n41623 );
and ( n369549 , n369547 , n369548 );
nor ( n369550 , n369546 , n369549 );
buf ( n369551 , n369550 );
not ( n49349 , n369551 );
not ( n369553 , n49349 );
or ( n369554 , n369543 , n369553 );
buf ( n369555 , n368426 );
not ( n369556 , n369555 );
buf ( n369557 , n359996 );
nor ( n49355 , n369556 , n369557 );
buf ( n369559 , n49355 );
not ( n369560 , n369559 );
nand ( n369561 , n369554 , n369560 );
not ( n49359 , n369561 );
or ( n369563 , n49338 , n49359 );
and ( n49361 , n49339 , n49349 );
nor ( n49362 , n49361 , n369559 );
not ( n49363 , n49362 );
not ( n49364 , n369540 );
not ( n49365 , n49364 );
or ( n49366 , n49363 , n49365 );
buf ( n369570 , n45113 );
not ( n369571 , n369570 );
buf ( n369572 , n44717 );
not ( n369573 , n369572 );
or ( n369574 , n369571 , n369573 );
buf ( n369575 , n41386 );
not ( n369576 , n369575 );
buf ( n369577 , n369576 );
buf ( n369578 , n369577 );
buf ( n369579 , n45125 );
nand ( n369580 , n369578 , n369579 );
buf ( n369581 , n369580 );
buf ( n369582 , n369581 );
nand ( n369583 , n369574 , n369582 );
buf ( n369584 , n369583 );
buf ( n369585 , n369584 );
not ( n369586 , n369585 );
buf ( n369587 , n361603 );
not ( n369588 , n369587 );
buf ( n369589 , n369588 );
buf ( n369590 , n369589 );
not ( n49388 , n369590 );
or ( n369592 , n369586 , n49388 );
buf ( n369593 , n368820 );
buf ( n369594 , n366518 );
nand ( n369595 , n369593 , n369594 );
buf ( n369596 , n369595 );
buf ( n369597 , n369596 );
nand ( n369598 , n369592 , n369597 );
buf ( n369599 , n369598 );
not ( n369600 , n369599 );
and ( n49398 , n364827 , n41772 );
not ( n49399 , n364827 );
and ( n369603 , n49399 , n44570 );
nor ( n369604 , n49398 , n369603 );
or ( n369605 , n366317 , n369604 );
or ( n49403 , n365312 , n368719 );
nand ( n369607 , n369605 , n49403 );
not ( n49405 , n369607 );
or ( n49406 , n369600 , n49405 );
buf ( n369610 , n369599 );
buf ( n369611 , n369607 );
or ( n49409 , n369610 , n369611 );
buf ( n369613 , n45300 );
not ( n49411 , n369613 );
buf ( n369615 , n364832 );
not ( n49413 , n369615 );
or ( n49414 , n49411 , n49413 );
buf ( n369618 , n45455 );
buf ( n369619 , n365464 );
nand ( n369620 , n369618 , n369619 );
buf ( n369621 , n369620 );
buf ( n369622 , n369621 );
nand ( n369623 , n49414 , n369622 );
buf ( n369624 , n369623 );
buf ( n369625 , n369624 );
not ( n369626 , n369625 );
buf ( n369627 , n362027 );
not ( n369628 , n369627 );
or ( n369629 , n369626 , n369628 );
buf ( n369630 , n364824 );
buf ( n369631 , n368793 );
nand ( n369632 , n369630 , n369631 );
buf ( n369633 , n369632 );
buf ( n369634 , n369633 );
nand ( n369635 , n369629 , n369634 );
buf ( n369636 , n369635 );
buf ( n369637 , n369636 );
nand ( n369638 , n49409 , n369637 );
buf ( n369639 , n369638 );
nand ( n49437 , n49406 , n369639 );
nand ( n369641 , n49366 , n49437 );
nand ( n369642 , n369563 , n369641 );
buf ( n369643 , n369642 );
nand ( n49441 , n369491 , n369643 );
buf ( n49442 , n49441 );
buf ( n369646 , n49442 );
nand ( n49444 , n369483 , n369646 );
buf ( n369648 , n49444 );
not ( n369649 , n369648 );
xor ( n49447 , n48427 , n48448 );
xor ( n369651 , n49447 , n48640 );
nand ( n369652 , n369649 , n369651 );
not ( n49450 , n369652 );
not ( n369654 , n48738 );
not ( n369655 , n48704 );
or ( n49453 , n369654 , n369655 );
nand ( n49454 , n48736 , n368930 );
nand ( n49455 , n49453 , n49454 );
and ( n49456 , n49455 , n369045 );
not ( n49457 , n49455 );
not ( n369661 , n369045 );
and ( n369662 , n49457 , n369661 );
nor ( n49460 , n49456 , n369662 );
not ( n369664 , n49460 );
or ( n49462 , n49450 , n369664 );
not ( n369666 , n369651 );
nand ( n49464 , n369666 , n369648 );
nand ( n369668 , n49462 , n49464 );
buf ( n369669 , n369668 );
xor ( n49467 , n369443 , n369669 );
xor ( n49468 , n48642 , n48668 );
xor ( n49469 , n49468 , n368858 );
buf ( n369673 , n49469 );
and ( n369674 , n49467 , n369673 );
and ( n49472 , n369443 , n369669 );
or ( n369676 , n369674 , n49472 );
buf ( n369677 , n369676 );
buf ( n369678 , n369677 );
not ( n49476 , n369678 );
buf ( n369680 , n49476 );
nand ( n369681 , n48977 , n369680 );
not ( n49479 , n369681 );
not ( n369683 , n368413 );
and ( n49481 , n368537 , n368534 );
not ( n49482 , n368537 );
not ( n369686 , n368534 );
and ( n369687 , n49482 , n369686 );
nor ( n49485 , n49481 , n369687 );
xor ( n369689 , n369683 , n49485 );
buf ( n369690 , n369689 );
not ( n49488 , n369690 );
buf ( n49489 , n49488 );
not ( n369693 , n49489 );
not ( n369694 , n368897 );
not ( n49492 , n369694 );
not ( n369696 , n48922 );
not ( n49494 , n369118 );
or ( n49495 , n369696 , n49494 );
or ( n49496 , n48922 , n369118 );
nand ( n49497 , n49495 , n49496 );
not ( n49498 , n49497 );
or ( n49499 , n49492 , n49498 );
or ( n369703 , n369694 , n49497 );
nand ( n49501 , n49499 , n369703 );
not ( n369705 , n49501 );
or ( n49503 , n369693 , n369705 );
xor ( n49504 , n368484 , n368501 );
xor ( n369708 , n49504 , n368532 );
not ( n369709 , n368989 );
not ( n49507 , n368968 );
or ( n369711 , n369709 , n49507 );
nand ( n369712 , n369711 , n369012 );
xor ( n49510 , n369712 , n369010 );
buf ( n369714 , n49510 );
not ( n49512 , n369714 );
buf ( n369716 , n49512 );
not ( n49514 , n369716 );
buf ( n369718 , n44819 );
not ( n49516 , n369718 );
buf ( n369720 , n360845 );
not ( n49518 , n369720 );
buf ( n369722 , n49518 );
buf ( n369723 , n369722 );
not ( n369724 , n369723 );
or ( n369725 , n49516 , n369724 );
buf ( n369726 , n362458 );
buf ( n369727 , n364994 );
nand ( n369728 , n369726 , n369727 );
buf ( n369729 , n369728 );
buf ( n369730 , n369729 );
nand ( n49528 , n369725 , n369730 );
buf ( n369732 , n49528 );
buf ( n369733 , n369732 );
buf ( n369734 , n365033 );
nand ( n49532 , n369733 , n369734 );
buf ( n369736 , n49532 );
buf ( n369737 , n369736 );
buf ( n49535 , n48831 );
buf ( n369739 , n365118 );
nand ( n49537 , n49535 , n369739 );
buf ( n369741 , n49537 );
buf ( n369742 , n369741 );
and ( n369743 , n369737 , n369742 );
buf ( n369744 , n369743 );
not ( n49542 , n369744 );
not ( n369746 , n49542 );
or ( n49544 , n49514 , n369746 );
not ( n369748 , n49510 );
not ( n49546 , n369744 );
or ( n49547 , n369748 , n49546 );
xor ( n369751 , n368781 , n368806 );
xor ( n49549 , n369751 , n368834 );
buf ( n369753 , n49549 );
nand ( n49551 , n49547 , n369753 );
nand ( n49552 , n49544 , n49551 );
buf ( n369756 , n49552 );
xor ( n49554 , n48812 , n369016 );
xor ( n369758 , n49554 , n369042 );
buf ( n369759 , n369758 );
xor ( n49557 , n369756 , n369759 );
buf ( n369761 , n368584 );
buf ( n369762 , n369761 );
buf ( n369763 , n369762 );
buf ( n369764 , n369763 );
buf ( n49562 , n369764 );
buf ( n369766 , n49562 );
buf ( n369767 , n369766 );
not ( n49565 , n369767 );
buf ( n369769 , n49565 );
not ( n49567 , n369769 );
not ( n49568 , n363439 );
or ( n49569 , n49567 , n49568 );
buf ( n369773 , n359144 );
buf ( n369774 , n369766 );
nand ( n369775 , n369773 , n369774 );
buf ( n369776 , n369775 );
nand ( n369777 , n49569 , n369776 );
buf ( n369778 , n369777 );
and ( n369779 , n343031 , n343034 );
not ( n49577 , n343031 );
and ( n49578 , n49577 , n23069 );
nor ( n49579 , n369779 , n49578 );
buf ( n369783 , n49579 );
buf ( n49581 , n369783 );
buf ( n49582 , n49581 );
not ( n369786 , n49582 );
and ( n49584 , n369786 , n343053 );
not ( n49585 , n369786 );
not ( n369789 , n343053 );
and ( n369790 , n49585 , n369789 );
nor ( n49588 , n49584 , n369790 );
buf ( n369792 , n49588 );
nand ( n369793 , n368581 , n343053 );
buf ( n369794 , n369793 );
nand ( n369795 , n369789 , n368584 );
buf ( n369796 , n369795 );
nand ( n49594 , n369792 , n369794 , n369796 );
buf ( n369798 , n49594 );
buf ( n49596 , n369798 );
not ( n369800 , n49596 );
buf ( n369801 , n369800 );
buf ( n369802 , n369801 );
buf ( n49600 , n369802 );
buf ( n369804 , n49600 );
buf ( n369805 , n369804 );
not ( n49603 , n369805 );
buf ( n49604 , n49603 );
buf ( n49605 , n49604 );
not ( n369809 , n49588 );
buf ( n369810 , n369809 );
buf ( n49608 , n369810 );
buf ( n49609 , n49608 );
not ( n369813 , n49609 );
buf ( n369814 , n369813 );
nand ( n369815 , n49605 , n369814 );
buf ( n369816 , n369815 );
buf ( n369817 , n369816 );
nand ( n49615 , n369778 , n369817 );
buf ( n369819 , n49615 );
buf ( n369820 , n369819 );
buf ( n369821 , n366428 );
not ( n369822 , n369821 );
buf ( n369823 , n369292 );
not ( n369824 , n369823 );
or ( n49622 , n369822 , n369824 );
buf ( n369826 , n342656 );
not ( n49624 , n369826 );
buf ( n369828 , n43377 );
not ( n369829 , n369828 );
or ( n49627 , n49624 , n369829 );
buf ( n369831 , n361716 );
buf ( n369832 , n342657 );
nand ( n49630 , n369831 , n369832 );
buf ( n369834 , n49630 );
buf ( n369835 , n369834 );
nand ( n49633 , n49627 , n369835 );
buf ( n49634 , n49633 );
buf ( n369838 , n49634 );
buf ( n369839 , n366402 );
nand ( n369840 , n369838 , n369839 );
buf ( n369841 , n369840 );
buf ( n369842 , n369841 );
nand ( n49640 , n49622 , n369842 );
buf ( n49641 , n49640 );
buf ( n369845 , n49641 );
buf ( n369846 , n365490 );
not ( n369847 , n369846 );
buf ( n369848 , n360613 );
not ( n49646 , n369848 );
or ( n49647 , n369847 , n49646 );
buf ( n369851 , n362452 );
buf ( n369852 , n45336 );
nand ( n49650 , n369851 , n369852 );
buf ( n369854 , n49650 );
buf ( n369855 , n369854 );
nand ( n49653 , n49647 , n369855 );
buf ( n369857 , n49653 );
buf ( n49655 , n369857 );
not ( n49656 , n49655 );
buf ( n369860 , n46557 );
not ( n49658 , n369860 );
or ( n49659 , n49656 , n49658 );
buf ( n369863 , n369230 );
buf ( n369864 , n366757 );
nand ( n49662 , n369863 , n369864 );
buf ( n369866 , n49662 );
buf ( n369867 , n369866 );
nand ( n369868 , n49659 , n369867 );
buf ( n369869 , n369868 );
buf ( n369870 , n369869 );
xor ( n369871 , n369845 , n369870 );
not ( n49669 , n48502 );
not ( n369873 , n49669 );
not ( n49671 , n364855 );
not ( n49672 , n45595 );
or ( n49673 , n49671 , n49672 );
buf ( n369877 , n365773 );
buf ( n369878 , n364858 );
nand ( n369879 , n369877 , n369878 );
buf ( n369880 , n369879 );
nand ( n369881 , n49673 , n369880 );
not ( n49679 , n369881 );
or ( n369883 , n369873 , n49679 );
buf ( n369884 , n368773 );
not ( n49682 , n369884 );
buf ( n369886 , n48490 );
nand ( n49684 , n49682 , n369886 );
buf ( n369888 , n49684 );
nand ( n49686 , n369883 , n369888 );
buf ( n369890 , n49686 );
buf ( n369891 , n366317 );
xor ( n49689 , n364744 , n31286 );
buf ( n369893 , n49689 );
or ( n369894 , n369891 , n369893 );
not ( n49692 , n41834 );
buf ( n369896 , n49692 );
buf ( n369897 , n369896 );
buf ( n369898 , n369604 );
or ( n49696 , n369897 , n369898 );
nand ( n369900 , n369894 , n49696 );
buf ( n369901 , n369900 );
buf ( n369902 , n369901 );
xor ( n49700 , n369890 , n369902 );
buf ( n369904 , n364852 );
buf ( n369905 , n352212 );
not ( n369906 , n369905 );
buf ( n369907 , n44717 );
not ( n369908 , n369907 );
or ( n369909 , n369906 , n369908 );
buf ( n369910 , n366096 );
buf ( n369911 , n365259 );
nand ( n369912 , n369910 , n369911 );
buf ( n369913 , n369912 );
buf ( n369914 , n369913 );
nand ( n49712 , n369909 , n369914 );
buf ( n369916 , n49712 );
buf ( n369917 , n369916 );
not ( n49715 , n369917 );
buf ( n369919 , n49715 );
buf ( n369920 , n369919 );
or ( n49718 , n369904 , n369920 );
buf ( n369922 , n369584 );
not ( n49720 , n369922 );
buf ( n369924 , n49720 );
buf ( n369925 , n369924 );
not ( n49723 , n366518 );
buf ( n369927 , n49723 );
or ( n49725 , n369925 , n369927 );
nand ( n369929 , n49718 , n49725 );
buf ( n369930 , n369929 );
buf ( n369931 , n369930 );
and ( n49729 , n49700 , n369931 );
and ( n369933 , n369890 , n369902 );
or ( n49731 , n49729 , n369933 );
buf ( n369935 , n49731 );
buf ( n369936 , n369935 );
and ( n369937 , n369871 , n369936 );
and ( n49735 , n369845 , n369870 );
or ( n369939 , n369937 , n49735 );
buf ( n369940 , n369939 );
buf ( n369941 , n369940 );
xor ( n369942 , n369820 , n369941 );
buf ( n369943 , n368051 );
not ( n49741 , n369943 );
buf ( n369945 , n49741 );
not ( n49743 , n369945 );
buf ( n369947 , n368662 );
buf ( n369948 , n359950 );
and ( n49746 , n369947 , n369948 );
not ( n369950 , n369947 );
buf ( n369951 , n364919 );
and ( n369952 , n369950 , n369951 );
nor ( n369953 , n49746 , n369952 );
buf ( n369954 , n369953 );
not ( n369955 , n369954 );
and ( n369956 , n49743 , n369955 );
buf ( n369957 , n367440 );
not ( n369958 , n369957 );
buf ( n369959 , n369958 );
buf ( n369960 , n369959 );
buf ( n369961 , n369551 );
nor ( n49759 , n369960 , n369961 );
buf ( n369963 , n49759 );
nor ( n369964 , n369956 , n369963 );
not ( n49762 , n369964 );
buf ( n369966 , n46521 );
not ( n369967 , n369966 );
buf ( n369968 , n46477 );
not ( n369969 , n369968 );
buf ( n369970 , n44783 );
not ( n49768 , n369970 );
or ( n369972 , n369969 , n49768 );
buf ( n369973 , n41607 );
buf ( n369974 , n366683 );
nand ( n49772 , n369973 , n369974 );
buf ( n369976 , n49772 );
buf ( n49774 , n369976 );
nand ( n49775 , n369972 , n49774 );
buf ( n49776 , n49775 );
buf ( n49777 , n49776 );
not ( n49778 , n49777 );
or ( n49779 , n369967 , n49778 );
buf ( n369983 , n369359 );
buf ( n369984 , n366654 );
nand ( n49782 , n369983 , n369984 );
buf ( n369986 , n49782 );
buf ( n369987 , n369986 );
nand ( n369988 , n49779 , n369987 );
buf ( n369989 , n369988 );
not ( n369990 , n369989 );
not ( n369991 , n369990 );
or ( n49789 , n49762 , n369991 );
buf ( n369993 , n43261 );
not ( n369994 , n369993 );
buf ( n369995 , n369497 );
not ( n49793 , n369995 );
buf ( n369997 , n364777 );
not ( n369998 , n369997 );
or ( n49796 , n49793 , n369998 );
buf ( n370000 , n364774 );
buf ( n370001 , n342718 );
nand ( n370002 , n370000 , n370001 );
buf ( n370003 , n370002 );
buf ( n370004 , n370003 );
nand ( n370005 , n49796 , n370004 );
buf ( n370006 , n370005 );
buf ( n370007 , n370006 );
not ( n370008 , n370007 );
or ( n370009 , n369994 , n370008 );
buf ( n370010 , n46693 );
not ( n370011 , n370010 );
buf ( n370012 , n45152 );
not ( n49810 , n370012 );
or ( n370014 , n370011 , n49810 );
buf ( n370015 , n30912 );
buf ( n370016 , n342718 );
nand ( n49814 , n370015 , n370016 );
buf ( n370018 , n49814 );
buf ( n370019 , n370018 );
nand ( n370020 , n370014 , n370019 );
buf ( n370021 , n370020 );
buf ( n370022 , n370021 );
buf ( n370023 , n363429 );
nand ( n370024 , n370022 , n370023 );
buf ( n370025 , n370024 );
buf ( n370026 , n370025 );
nand ( n370027 , n370009 , n370026 );
buf ( n370028 , n370027 );
buf ( n49826 , n370028 );
not ( n49827 , n49826 );
buf ( n49828 , n49827 );
buf ( n370032 , n49828 );
not ( n49830 , n370032 );
buf ( n370034 , n49830 );
buf ( n370035 , n370034 );
not ( n370036 , n370035 );
and ( n49834 , n369507 , n43261 );
not ( n370038 , n370006 );
nor ( n49836 , n370038 , n43274 );
nor ( n370040 , n49834 , n49836 );
not ( n370041 , n370040 );
buf ( n370042 , n370041 );
not ( n370043 , n370042 );
or ( n370044 , n370036 , n370043 );
not ( n49842 , n370040 );
not ( n370046 , n49828 );
or ( n49844 , n49842 , n370046 );
buf ( n370048 , n365303 );
not ( n49846 , n370048 );
buf ( n370050 , n49846 );
buf ( n370051 , n49321 );
not ( n49849 , n370051 );
buf ( n370053 , n49849 );
or ( n370054 , n370050 , n370053 );
not ( n49852 , n31197 );
not ( n370056 , n45855 );
or ( n370057 , n49852 , n370056 );
or ( n49855 , n365293 , n31197 );
nand ( n370059 , n370057 , n49855 );
buf ( n370060 , n40878 );
or ( n49858 , n370059 , n370060 );
nand ( n49859 , n370054 , n49858 );
nand ( n370063 , n49844 , n49859 );
buf ( n370064 , n370063 );
nand ( n370065 , n370044 , n370064 );
buf ( n370066 , n370065 );
nand ( n370067 , n49789 , n370066 );
buf ( n370068 , n370067 );
not ( n49866 , n369964 );
nand ( n370070 , n49866 , n369989 );
buf ( n370071 , n370070 );
nand ( n370072 , n370068 , n370071 );
buf ( n370073 , n370072 );
buf ( n370074 , n370073 );
and ( n370075 , n369942 , n370074 );
and ( n370076 , n369820 , n369941 );
or ( n370077 , n370075 , n370076 );
buf ( n370078 , n370077 );
buf ( n370079 , n370078 );
and ( n370080 , n49557 , n370079 );
and ( n49878 , n369756 , n369759 );
or ( n370082 , n370080 , n49878 );
buf ( n370083 , n370082 );
xor ( n49881 , n369708 , n370083 );
buf ( n370085 , n369107 );
buf ( n370086 , n48848 );
and ( n49884 , n370085 , n370086 );
not ( n49885 , n370085 );
buf ( n370089 , n369052 );
and ( n370090 , n49885 , n370089 );
nor ( n370091 , n49884 , n370090 );
buf ( n370092 , n370091 );
buf ( n370093 , n370092 );
buf ( n370094 , n369113 );
and ( n49892 , n370093 , n370094 );
not ( n370096 , n370093 );
buf ( n370097 , n369060 );
and ( n49895 , n370096 , n370097 );
nor ( n370099 , n49892 , n49895 );
buf ( n370100 , n370099 );
and ( n49898 , n49881 , n370100 );
and ( n370102 , n369708 , n370083 );
or ( n49900 , n49898 , n370102 );
nand ( n49901 , n49503 , n49900 );
buf ( n370105 , n49501 );
not ( n370106 , n370105 );
buf ( n370107 , n370106 );
buf ( n370108 , n369689 );
nand ( n49906 , n370107 , n370108 );
nand ( n370110 , n49901 , n49906 );
not ( n49908 , n370110 );
or ( n370112 , n49479 , n49908 );
not ( n49910 , n48977 );
buf ( n370114 , n369677 );
nand ( n49912 , n49910 , n370114 );
nand ( n370116 , n370112 , n49912 );
buf ( n370117 , n370116 );
xor ( n370118 , n369168 , n370117 );
and ( n49916 , n369154 , n368886 );
not ( n49917 , n369154 );
and ( n370121 , n49917 , n48684 );
nor ( n370122 , n49916 , n370121 );
not ( n49920 , n369150 );
and ( n370124 , n370122 , n49920 );
not ( n370125 , n370122 );
and ( n49923 , n370125 , n369150 );
nor ( n370127 , n370124 , n49923 );
buf ( n370128 , n370127 );
and ( n49926 , n370118 , n370128 );
and ( n49927 , n369168 , n370117 );
or ( n370131 , n49926 , n49927 );
buf ( n370132 , n370131 );
or ( n49930 , n369164 , n370132 );
buf ( n370134 , n368021 );
not ( n370135 , n370134 );
buf ( n370136 , n47859 );
not ( n370137 , n370136 );
buf ( n370138 , n370137 );
buf ( n370139 , n370138 );
not ( n370140 , n370139 );
or ( n370141 , n370135 , n370140 );
not ( n49939 , n46393 );
not ( n49940 , n368006 );
or ( n49941 , n49939 , n49940 );
nand ( n49942 , n49941 , n368012 );
buf ( n370146 , n49942 );
nand ( n49944 , n370141 , n370146 );
buf ( n370148 , n49944 );
buf ( n370149 , n370148 );
buf ( n370150 , n47859 );
buf ( n370151 , n368018 );
nand ( n370152 , n370150 , n370151 );
buf ( n370153 , n370152 );
buf ( n370154 , n370153 );
nand ( n370155 , n370149 , n370154 );
buf ( n370156 , n370155 );
buf ( n370157 , n370156 );
buf ( n370158 , n368340 );
not ( n49956 , n370158 );
buf ( n370160 , n361606 );
not ( n49958 , n370160 );
or ( n370162 , n49956 , n49958 );
buf ( n370163 , n361531 );
not ( n49961 , n370163 );
buf ( n370165 , n365760 );
not ( n370166 , n370165 );
or ( n49964 , n49961 , n370166 );
buf ( n370168 , n365757 );
buf ( n370169 , n44717 );
nand ( n49967 , n370168 , n370169 );
buf ( n49968 , n49967 );
buf ( n370172 , n49968 );
nand ( n370173 , n49964 , n370172 );
buf ( n370174 , n370173 );
buf ( n370175 , n370174 );
buf ( n370176 , n366518 );
nand ( n49974 , n370175 , n370176 );
buf ( n49975 , n49974 );
buf ( n370179 , n49975 );
nand ( n49977 , n370162 , n370179 );
buf ( n370181 , n49977 );
buf ( n370182 , n370181 );
buf ( n370183 , n367861 );
not ( n370184 , n370183 );
buf ( n370185 , n361013 );
not ( n49983 , n370185 );
or ( n370187 , n370184 , n49983 );
buf ( n370188 , n40923 );
buf ( n49986 , n364777 );
buf ( n49987 , n49986 );
buf ( n49988 , n49987 );
not ( n370192 , n49988 );
not ( n49990 , n365293 );
or ( n49991 , n370192 , n49990 );
nand ( n49992 , n45116 , n42911 );
nand ( n49993 , n49991 , n49992 );
buf ( n370197 , n49993 );
nand ( n49995 , n370188 , n370197 );
buf ( n370199 , n49995 );
buf ( n370200 , n370199 );
nand ( n370201 , n370187 , n370200 );
buf ( n370202 , n370201 );
buf ( n370203 , n370202 );
and ( n50001 , n370182 , n370203 );
not ( n50002 , n370182 );
buf ( n370206 , n370202 );
not ( n50004 , n370206 );
buf ( n370208 , n50004 );
buf ( n370209 , n370208 );
and ( n370210 , n50002 , n370209 );
nor ( n370211 , n50001 , n370210 );
buf ( n370212 , n370211 );
buf ( n370213 , n370212 );
buf ( n370214 , n368306 );
not ( n50012 , n370214 );
buf ( n370216 , n45345 );
not ( n370217 , n370216 );
or ( n370218 , n50012 , n370217 );
buf ( n370219 , n352212 );
not ( n370220 , n370219 );
buf ( n370221 , n365945 );
not ( n50019 , n370221 );
or ( n370223 , n370220 , n50019 );
buf ( n370224 , n363119 );
buf ( n370225 , n365259 );
nand ( n50023 , n370224 , n370225 );
buf ( n370227 , n50023 );
buf ( n370228 , n370227 );
nand ( n50026 , n370223 , n370228 );
buf ( n370230 , n50026 );
buf ( n370231 , n370230 );
buf ( n370232 , n365486 );
nand ( n50030 , n370231 , n370232 );
buf ( n370234 , n50030 );
buf ( n370235 , n370234 );
nand ( n370236 , n370218 , n370235 );
buf ( n370237 , n370236 );
buf ( n370238 , n370237 );
and ( n50036 , n370213 , n370238 );
not ( n50037 , n370213 );
buf ( n50038 , n370237 );
not ( n50039 , n50038 );
buf ( n50040 , n50039 );
buf ( n50041 , n50040 );
and ( n50042 , n50037 , n50041 );
nor ( n370246 , n50036 , n50042 );
buf ( n370247 , n370246 );
buf ( n370248 , n370247 );
xor ( n370249 , n366522 , n47839 );
and ( n50047 , n370249 , n368053 );
and ( n370251 , n366522 , n47839 );
or ( n370252 , n50047 , n370251 );
buf ( n370253 , n370252 );
xor ( n370254 , n370248 , n370253 );
buf ( n370255 , n366654 );
not ( n50053 , n370255 );
not ( n370257 , n359778 );
not ( n370258 , n370257 );
xor ( n50056 , n46477 , n370258 );
buf ( n370260 , n50056 );
not ( n370261 , n370260 );
or ( n50059 , n50053 , n370261 );
buf ( n370263 , n367902 );
buf ( n370264 , n46521 );
nand ( n50062 , n370263 , n370264 );
buf ( n370266 , n50062 );
buf ( n370267 , n370266 );
nand ( n50065 , n50059 , n370267 );
buf ( n370269 , n50065 );
buf ( n370270 , n370269 );
xor ( n370271 , n370254 , n370270 );
buf ( n370272 , n370271 );
buf ( n370273 , n370272 );
xor ( n370274 , n370157 , n370273 );
buf ( n370275 , n47929 );
not ( n370276 , n370275 );
buf ( n370277 , n368142 );
not ( n370278 , n370277 );
or ( n370279 , n370276 , n370278 );
buf ( n370280 , n47953 );
not ( n370281 , n370280 );
buf ( n370282 , n47948 );
not ( n370283 , n370282 );
or ( n50076 , n370281 , n370283 );
buf ( n370285 , n368173 );
nand ( n370286 , n50076 , n370285 );
buf ( n370287 , n370286 );
buf ( n370288 , n370287 );
nand ( n370289 , n370279 , n370288 );
buf ( n370290 , n370289 );
buf ( n370291 , n370290 );
xor ( n50084 , n370274 , n370291 );
buf ( n370293 , n50084 );
buf ( n370294 , n370293 );
nand ( n50087 , n48019 , n368206 );
nand ( n370296 , n368358 , n50087 );
nand ( n370297 , n368205 , n368211 );
nand ( n50090 , n370296 , n370297 );
xor ( n370299 , n367766 , n367789 );
and ( n370300 , n370299 , n367873 );
and ( n50093 , n367766 , n367789 );
or ( n370302 , n370300 , n50093 );
buf ( n370303 , n370302 );
buf ( n370304 , n370303 );
not ( n370305 , n366046 );
not ( n370306 , n367836 );
or ( n50099 , n370305 , n370306 );
buf ( n370308 , n368976 );
not ( n50101 , n370308 );
buf ( n370310 , n50101 );
not ( n370311 , n365626 );
or ( n50104 , n370310 , n370311 );
nand ( n370313 , n370311 , n362534 );
nand ( n50106 , n50104 , n370313 );
not ( n370315 , n50106 );
nand ( n370316 , n370315 , n364824 );
nand ( n50109 , n50099 , n370316 );
not ( n370318 , n50109 );
buf ( n370319 , n370318 );
buf ( n370320 , n367759 );
not ( n370321 , n370320 );
buf ( n370322 , n367754 );
not ( n370323 , n370322 );
or ( n50116 , n370321 , n370323 );
buf ( n370325 , n47554 );
not ( n370326 , n370325 );
buf ( n370327 , n369349 );
not ( n50120 , n370327 );
or ( n370329 , n370326 , n50120 );
buf ( n370330 , n46031 );
buf ( n370331 , n41772 );
nand ( n370332 , n370330 , n370331 );
buf ( n370333 , n370332 );
buf ( n370334 , n370333 );
nand ( n50127 , n370329 , n370334 );
buf ( n50128 , n50127 );
buf ( n370337 , n50128 );
buf ( n370338 , n41835 );
nand ( n370339 , n370337 , n370338 );
buf ( n370340 , n370339 );
buf ( n370341 , n370340 );
nand ( n370342 , n50116 , n370341 );
buf ( n370343 , n370342 );
buf ( n370344 , n370343 );
xor ( n370345 , n370319 , n370344 );
buf ( n370346 , n368047 );
not ( n50139 , n370346 );
buf ( n370348 , n363291 );
not ( n370349 , n370348 );
buf ( n370350 , n370349 );
buf ( n370351 , n370350 );
not ( n370352 , n370351 );
or ( n50145 , n50139 , n370352 );
buf ( n370354 , n367440 );
buf ( n50147 , n365440 );
not ( n50148 , n50147 );
buf ( n50149 , n42455 );
not ( n50150 , n50149 );
or ( n50151 , n50148 , n50150 );
buf ( n370360 , n364905 );
buf ( n370361 , n365452 );
nand ( n50154 , n370360 , n370361 );
buf ( n370363 , n50154 );
buf ( n370364 , n370363 );
nand ( n50157 , n50151 , n370364 );
buf ( n370366 , n50157 );
buf ( n370367 , n370366 );
nand ( n50160 , n370354 , n370367 );
buf ( n370369 , n50160 );
buf ( n370370 , n370369 );
nand ( n50163 , n50145 , n370370 );
buf ( n370372 , n50163 );
buf ( n370373 , n370372 );
xnor ( n370374 , n370345 , n370373 );
buf ( n370375 , n370374 );
buf ( n50168 , n370375 );
xor ( n50169 , n370304 , n50168 );
not ( n370378 , n367889 );
nand ( n50171 , n370378 , n367935 );
buf ( n370380 , n50171 );
buf ( n370381 , n47718 );
and ( n370382 , n370380 , n370381 );
not ( n370383 , n367889 );
nor ( n50176 , n370383 , n367935 );
buf ( n370385 , n50176 );
nor ( n370386 , n370382 , n370385 );
buf ( n370387 , n370386 );
buf ( n370388 , n370387 );
xnor ( n50181 , n50169 , n370388 );
buf ( n370390 , n50181 );
buf ( n370391 , n365118 );
not ( n50184 , n370391 );
buf ( n370393 , n44819 );
not ( n370394 , n370393 );
buf ( n370395 , n363866 );
not ( n370396 , n370395 );
or ( n370397 , n370394 , n370396 );
buf ( n370398 , n41406 );
buf ( n370399 , n364997 );
nand ( n370400 , n370398 , n370399 );
buf ( n370401 , n370400 );
buf ( n370402 , n370401 );
nand ( n370403 , n370397 , n370402 );
buf ( n370404 , n370403 );
buf ( n370405 , n370404 );
not ( n50198 , n370405 );
or ( n50199 , n50184 , n50198 );
buf ( n370408 , n368135 );
buf ( n370409 , n365033 );
nand ( n50202 , n370408 , n370409 );
buf ( n370411 , n50202 );
buf ( n370412 , n370411 );
nand ( n50205 , n50199 , n370412 );
buf ( n370414 , n50205 );
buf ( n370415 , n370414 );
buf ( n370416 , n45058 );
not ( n50209 , n370416 );
buf ( n370418 , n47922 );
not ( n50211 , n370418 );
or ( n50212 , n50209 , n50211 );
buf ( n370421 , n342881 );
not ( n370422 , n370421 );
buf ( n370423 , n368548 );
not ( n50216 , n370423 );
or ( n50217 , n370422 , n50216 );
buf ( n370426 , n48344 );
buf ( n370427 , n365202 );
nand ( n50220 , n370426 , n370427 );
buf ( n370429 , n50220 );
buf ( n370430 , n370429 );
nand ( n50223 , n50217 , n370430 );
buf ( n50224 , n50223 );
buf ( n370433 , n50224 );
buf ( n370434 , n45075 );
nand ( n50227 , n370433 , n370434 );
buf ( n370436 , n50227 );
buf ( n370437 , n370436 );
nand ( n50230 , n50212 , n370437 );
buf ( n370439 , n50230 );
buf ( n370440 , n370439 );
xor ( n50233 , n370415 , n370440 );
buf ( n370442 , n45553 );
not ( n50235 , n370442 );
buf ( n370444 , n368198 );
not ( n370445 , n370444 );
or ( n370446 , n50235 , n370445 );
and ( n50239 , n39830 , n365673 );
not ( n50240 , n39830 );
and ( n50241 , n50240 , n365676 );
or ( n370450 , n50239 , n50241 );
buf ( n370451 , n370450 );
buf ( n370452 , n45492 );
nand ( n50245 , n370451 , n370452 );
buf ( n370454 , n50245 );
buf ( n370455 , n370454 );
nand ( n370456 , n370446 , n370455 );
buf ( n370457 , n370456 );
buf ( n370458 , n370457 );
xor ( n370459 , n50233 , n370458 );
buf ( n370460 , n370459 );
xnor ( n50253 , n370390 , n370460 );
xor ( n370462 , n50090 , n50253 );
buf ( n370463 , n370462 );
xor ( n50256 , n370294 , n370463 );
buf ( n370465 , n47985 );
not ( n370466 , n370465 );
buf ( n370467 , n48168 );
not ( n50260 , n370467 );
or ( n370469 , n370466 , n50260 );
buf ( n370470 , n47916 );
nand ( n370471 , n370469 , n370470 );
buf ( n370472 , n370471 );
buf ( n370473 , n370472 );
buf ( n370474 , n47985 );
not ( n50267 , n370474 );
buf ( n370476 , n368368 );
nand ( n370477 , n50267 , n370476 );
buf ( n370478 , n370477 );
buf ( n370479 , n370478 );
nand ( n50272 , n370473 , n370479 );
buf ( n370481 , n50272 );
buf ( n370482 , n370481 );
and ( n50275 , n50256 , n370482 );
and ( n370484 , n370294 , n370463 );
or ( n50277 , n50275 , n370484 );
buf ( n370486 , n50277 );
buf ( n370487 , n370486 );
not ( n50280 , n367867 );
not ( n370489 , n367843 );
or ( n50282 , n50280 , n370489 );
buf ( n370491 , n367867 );
buf ( n370492 , n367843 );
nor ( n50285 , n370491 , n370492 );
buf ( n50286 , n50285 );
or ( n370495 , n367818 , n50286 );
nand ( n370496 , n50282 , n370495 );
buf ( n370497 , n43261 );
not ( n370498 , n370497 );
buf ( n370499 , n22772 );
not ( n50292 , n370499 );
buf ( n370501 , n366673 );
not ( n50294 , n370501 );
or ( n50295 , n50292 , n50294 );
buf ( n370504 , n360845 );
buf ( n370505 , n363444 );
nand ( n370506 , n370504 , n370505 );
buf ( n370507 , n370506 );
buf ( n370508 , n370507 );
nand ( n50301 , n50295 , n370508 );
buf ( n370510 , n50301 );
buf ( n370511 , n370510 );
not ( n370512 , n370511 );
or ( n50305 , n370498 , n370512 );
buf ( n370514 , n47696 );
buf ( n370515 , n363429 );
nand ( n50308 , n370514 , n370515 );
buf ( n370517 , n50308 );
buf ( n370518 , n370517 );
nand ( n50311 , n50305 , n370518 );
buf ( n370520 , n50311 );
not ( n50313 , n370520 );
xor ( n50314 , n370496 , n50313 );
buf ( n370523 , n368315 );
not ( n50316 , n370523 );
buf ( n370525 , n50316 );
buf ( n370526 , n370525 );
not ( n50319 , n370526 );
buf ( n370528 , n48152 );
not ( n50321 , n370528 );
or ( n50322 , n50319 , n50321 );
buf ( n370531 , n370525 );
buf ( n370532 , n48152 );
or ( n370533 , n370531 , n370532 );
buf ( n370534 , n368283 );
nand ( n50327 , n370533 , n370534 );
buf ( n370536 , n50327 );
buf ( n370537 , n370536 );
nand ( n370538 , n50322 , n370537 );
buf ( n370539 , n370538 );
xor ( n370540 , n50314 , n370539 );
buf ( n370541 , n370540 );
buf ( n370542 , n48047 );
not ( n50335 , n370542 );
buf ( n370544 , n368357 );
nand ( n50337 , n50335 , n370544 );
buf ( n370546 , n50337 );
buf ( n370547 , n370546 );
buf ( n370548 , n368258 );
and ( n50341 , n370547 , n370548 );
buf ( n370550 , n48047 );
not ( n370551 , n370550 );
buf ( n370552 , n368357 );
nor ( n370553 , n370551 , n370552 );
buf ( n370554 , n370553 );
buf ( n370555 , n370554 );
nor ( n50348 , n50341 , n370555 );
buf ( n370557 , n50348 );
buf ( n50350 , n370557 );
xor ( n50351 , n370541 , n50350 );
not ( n370560 , n42242 );
not ( n370561 , n42149 );
not ( n50354 , n362435 );
or ( n370563 , n370561 , n50354 );
buf ( n370564 , n362285 );
not ( n50357 , n370564 );
buf ( n370566 , n50357 );
nand ( n50359 , n370566 , n362426 );
nand ( n370568 , n370563 , n50359 );
not ( n370569 , n370568 );
or ( n50362 , n370560 , n370569 );
buf ( n370571 , n368230 );
buf ( n370572 , n363210 );
nand ( n370573 , n370571 , n370572 );
buf ( n370574 , n370573 );
nand ( n50367 , n50362 , n370574 );
buf ( n370576 , n366402 );
not ( n50369 , n370576 );
buf ( n370578 , n367922 );
not ( n50371 , n370578 );
or ( n370580 , n50369 , n50371 );
buf ( n370581 , n342657 );
buf ( n370582 , n366722 );
xor ( n370583 , n370581 , n370582 );
buf ( n370584 , n370583 );
buf ( n370585 , n370584 );
not ( n370586 , n370585 );
buf ( n50379 , n366434 );
nand ( n50380 , n370586 , n50379 );
buf ( n50381 , n50380 );
buf ( n50382 , n50381 );
nand ( n50383 , n370580 , n50382 );
buf ( n50384 , n50383 );
xor ( n370593 , n50367 , n50384 );
buf ( n370594 , n367809 );
not ( n370595 , n370594 );
buf ( n370596 , n45795 );
not ( n370597 , n370596 );
or ( n50390 , n370595 , n370597 );
buf ( n370599 , n362521 );
buf ( n50392 , n31197 );
not ( n50393 , n50392 );
buf ( n50394 , n45231 );
not ( n50395 , n50394 );
or ( n50396 , n50393 , n50395 );
buf ( n50397 , n366534 );
buf ( n50398 , n351229 );
nand ( n50399 , n50397 , n50398 );
buf ( n50400 , n50399 );
buf ( n50401 , n50400 );
nand ( n50402 , n50396 , n50401 );
buf ( n50403 , n50402 );
buf ( n370612 , n50403 );
nand ( n370613 , n370599 , n370612 );
buf ( n370614 , n370613 );
buf ( n370615 , n370614 );
nand ( n370616 , n50390 , n370615 );
buf ( n370617 , n370616 );
buf ( n370618 , n370617 );
buf ( n370619 , n368276 );
not ( n50412 , n370619 );
buf ( n370621 , n46113 );
not ( n50414 , n370621 );
or ( n370623 , n50412 , n50414 );
buf ( n370624 , n364858 );
not ( n50417 , n370624 );
buf ( n370626 , n365468 );
not ( n370627 , n370626 );
or ( n370628 , n50417 , n370627 );
buf ( n370629 , n362452 );
buf ( n370630 , n364870 );
nand ( n50423 , n370629 , n370630 );
buf ( n370632 , n50423 );
buf ( n370633 , n370632 );
nand ( n370634 , n370628 , n370633 );
buf ( n370635 , n370634 );
buf ( n370636 , n370635 );
buf ( n370637 , n366757 );
nand ( n50430 , n370636 , n370637 );
buf ( n370639 , n50430 );
buf ( n370640 , n370639 );
nand ( n370641 , n370623 , n370640 );
buf ( n370642 , n370641 );
buf ( n370643 , n370642 );
xor ( n370644 , n370618 , n370643 );
buf ( n370645 , n368029 );
not ( n370646 , n370645 );
buf ( n370647 , n45204 );
not ( n50440 , n370647 );
or ( n370649 , n370646 , n50440 );
buf ( n370650 , n365353 );
not ( n50443 , n370650 );
not ( n370652 , n364808 );
buf ( n370653 , n370652 );
not ( n50446 , n370653 );
and ( n370655 , n50443 , n50446 );
buf ( n370656 , n35548 );
buf ( n370657 , n31286 );
and ( n50450 , n370656 , n370657 );
nor ( n370659 , n370655 , n50450 );
buf ( n370660 , n370659 );
buf ( n370661 , n370660 );
not ( n370662 , n370661 );
buf ( n370663 , n39217 );
nand ( n370664 , n370662 , n370663 );
buf ( n370665 , n370664 );
buf ( n370666 , n370665 );
nand ( n50459 , n370649 , n370666 );
buf ( n370668 , n50459 );
buf ( n370669 , n370668 );
xor ( n50462 , n370644 , n370669 );
buf ( n370671 , n50462 );
xor ( n370672 , n370593 , n370671 );
buf ( n370673 , n370672 );
xnor ( n50466 , n50351 , n370673 );
buf ( n50467 , n50466 );
xor ( n370676 , n367737 , n367876 );
and ( n50469 , n370676 , n367940 );
and ( n370678 , n367737 , n367876 );
or ( n370679 , n50469 , n370678 );
buf ( n370680 , n370679 );
and ( n50473 , n50467 , n370680 );
not ( n370682 , n50467 );
not ( n370683 , n370680 );
and ( n50476 , n370682 , n370683 );
nor ( n370685 , n50473 , n50476 );
xor ( n370686 , n368058 , n368068 );
and ( n50479 , n370686 , n368074 );
and ( n370688 , n368058 , n368068 );
or ( n370689 , n50479 , n370688 );
buf ( n370690 , n370689 );
and ( n370691 , n370685 , n370690 );
not ( n50484 , n370685 );
not ( n50485 , n370690 );
and ( n370694 , n50484 , n50485 );
nor ( n370695 , n370691 , n370694 );
not ( n50488 , n370695 );
buf ( n370697 , n50488 );
not ( n370698 , n47781 );
not ( n50491 , n47767 );
nand ( n50492 , n50491 , n47763 );
not ( n370701 , n50492 );
or ( n370702 , n370698 , n370701 );
not ( n50495 , n47763 );
nand ( n370704 , n50495 , n47767 );
nand ( n50497 , n370702 , n370704 );
not ( n50498 , n50497 );
buf ( n370707 , n50498 );
nand ( n370708 , n370697 , n370707 );
buf ( n370709 , n370708 );
buf ( n370710 , n370709 );
not ( n370711 , n370710 );
not ( n50504 , n368373 );
not ( n370713 , n368079 );
or ( n50506 , n50504 , n370713 );
not ( n50507 , n368076 );
not ( n370716 , n48175 );
or ( n50509 , n50507 , n370716 );
nand ( n370718 , n50509 , n368085 );
nand ( n50511 , n50506 , n370718 );
buf ( n50512 , n50511 );
not ( n50513 , n50512 );
or ( n50514 , n370711 , n50513 );
not ( n370723 , n50498 );
nand ( n370724 , n370723 , n370695 );
buf ( n370725 , n370724 );
nand ( n370726 , n50514 , n370725 );
buf ( n370727 , n370726 );
buf ( n370728 , n370727 );
xor ( n370729 , n370487 , n370728 );
not ( n370730 , n50485 );
buf ( n370731 , n50467 );
buf ( n370732 , n370731 );
buf ( n370733 , n370732 );
nand ( n50526 , n370733 , n370683 );
not ( n370735 , n50526 );
or ( n370736 , n370730 , n370735 );
buf ( n370737 , n370733 );
not ( n370738 , n370737 );
buf ( n370739 , n370680 );
nand ( n50532 , n370738 , n370739 );
buf ( n50533 , n50532 );
nand ( n370742 , n370736 , n50533 );
not ( n50535 , n370557 );
not ( n50536 , n370672 );
buf ( n370745 , n370540 );
nand ( n50538 , n50536 , n370745 );
nand ( n370747 , n50535 , n50538 );
buf ( n370748 , n370747 );
buf ( n370749 , n370745 );
not ( n370750 , n370749 );
buf ( n370751 , n370672 );
nand ( n50544 , n370750 , n370751 );
buf ( n370753 , n50544 );
buf ( n370754 , n370753 );
nand ( n370755 , n370748 , n370754 );
buf ( n370756 , n370755 );
buf ( n370757 , n370756 );
xor ( n370758 , n50367 , n50384 );
and ( n370759 , n370758 , n370671 );
and ( n50552 , n50367 , n50384 );
or ( n370761 , n370759 , n50552 );
not ( n370762 , n370237 );
not ( n50555 , n370181 );
nand ( n370764 , n50555 , n370208 );
not ( n370765 , n370764 );
or ( n50558 , n370762 , n370765 );
buf ( n370767 , n370181 );
buf ( n370768 , n370202 );
nand ( n50561 , n370767 , n370768 );
buf ( n370770 , n50561 );
nand ( n50563 , n50558 , n370770 );
buf ( n370772 , n50563 );
buf ( n370773 , n41835 );
not ( n370774 , n370773 );
buf ( n370775 , n47554 );
not ( n50568 , n370775 );
buf ( n370777 , n362145 );
not ( n50570 , n370777 );
or ( n50571 , n50568 , n50570 );
buf ( n370780 , n45718 );
not ( n370781 , n370780 );
buf ( n370782 , n370781 );
buf ( n370783 , n370782 );
buf ( n370784 , n41772 );
nand ( n50577 , n370783 , n370784 );
buf ( n50578 , n50577 );
buf ( n370787 , n50578 );
nand ( n50580 , n50571 , n370787 );
buf ( n370789 , n50580 );
buf ( n370790 , n370789 );
not ( n370791 , n370790 );
or ( n370792 , n370774 , n370791 );
buf ( n370793 , n50128 );
buf ( n370794 , n41830 );
nand ( n370795 , n370793 , n370794 );
buf ( n370796 , n370795 );
buf ( n370797 , n370796 );
nand ( n50590 , n370792 , n370797 );
buf ( n370799 , n50590 );
buf ( n370800 , n370799 );
xor ( n50593 , n370772 , n370800 );
xor ( n370802 , n370618 , n370643 );
and ( n50595 , n370802 , n370669 );
and ( n50596 , n370618 , n370643 );
or ( n370805 , n50595 , n50596 );
buf ( n370806 , n370805 );
buf ( n370807 , n370806 );
xnor ( n370808 , n50593 , n370807 );
buf ( n370809 , n370808 );
xor ( n370810 , n370761 , n370809 );
buf ( n370811 , n363210 );
not ( n50604 , n370811 );
buf ( n370813 , n370568 );
not ( n370814 , n370813 );
or ( n50607 , n50604 , n370814 );
buf ( n370816 , n362426 );
not ( n50609 , n370816 );
buf ( n370818 , n368474 );
not ( n370819 , n370818 );
or ( n370820 , n50609 , n370819 );
buf ( n370821 , n360885 );
buf ( n370822 , n366212 );
nand ( n50615 , n370821 , n370822 );
buf ( n370824 , n50615 );
buf ( n370825 , n370824 );
nand ( n370826 , n370820 , n370825 );
buf ( n370827 , n370826 );
buf ( n370828 , n370827 );
buf ( n50621 , n42242 );
nand ( n50622 , n370828 , n50621 );
buf ( n370831 , n50622 );
buf ( n370832 , n370831 );
nand ( n370833 , n50607 , n370832 );
buf ( n370834 , n370833 );
buf ( n370835 , n370834 );
buf ( n370836 , n370230 );
not ( n50629 , n370836 );
buf ( n370838 , n45345 );
not ( n370839 , n370838 );
or ( n50632 , n50629 , n370839 );
buf ( n370841 , n45113 );
not ( n370842 , n370841 );
buf ( n370843 , n365495 );
not ( n370844 , n370843 );
buf ( n370845 , n370844 );
buf ( n370846 , n370845 );
not ( n370847 , n370846 );
or ( n370848 , n370842 , n370847 );
buf ( n370849 , n363119 );
buf ( n370850 , n352194 );
nand ( n50643 , n370849 , n370850 );
buf ( n50644 , n50643 );
buf ( n50645 , n50644 );
nand ( n370854 , n370848 , n50645 );
buf ( n370855 , n370854 );
buf ( n370856 , n370855 );
buf ( n370857 , n365954 );
nand ( n370858 , n370856 , n370857 );
buf ( n370859 , n370858 );
buf ( n370860 , n370859 );
nand ( n50653 , n50632 , n370860 );
buf ( n370862 , n50653 );
buf ( n370863 , n370862 );
not ( n50656 , n370863 );
buf ( n370865 , n50656 );
buf ( n370866 , n370865 );
not ( n50659 , n370866 );
buf ( n370868 , n50403 );
not ( n370869 , n370868 );
buf ( n370870 , n39701 );
not ( n370871 , n370870 );
or ( n370872 , n370869 , n370871 );
buf ( n370873 , n39592 );
buf ( n370874 , n45177 );
not ( n370875 , n370874 );
buf ( n370876 , n45231 );
not ( n370877 , n370876 );
or ( n50670 , n370875 , n370877 );
buf ( n370879 , n39621 );
buf ( n370880 , n365357 );
nand ( n50673 , n370879 , n370880 );
buf ( n370882 , n50673 );
buf ( n370883 , n370882 );
nand ( n370884 , n50670 , n370883 );
buf ( n370885 , n370884 );
buf ( n370886 , n370885 );
nand ( n370887 , n370873 , n370886 );
buf ( n370888 , n370887 );
buf ( n370889 , n370888 );
nand ( n50682 , n370872 , n370889 );
buf ( n370891 , n50682 );
buf ( n370892 , n370635 );
not ( n50685 , n370892 );
buf ( n370894 , n46113 );
not ( n370895 , n370894 );
or ( n50688 , n50685 , n370895 );
buf ( n370897 , n30912 );
not ( n370898 , n370897 );
buf ( n370899 , n45270 );
not ( n370900 , n370899 );
or ( n50693 , n370898 , n370900 );
buf ( n370902 , n366151 );
buf ( n370903 , n45152 );
nand ( n370904 , n370902 , n370903 );
buf ( n370905 , n370904 );
buf ( n370906 , n370905 );
nand ( n50699 , n50693 , n370906 );
buf ( n370908 , n50699 );
buf ( n370909 , n370908 );
buf ( n370910 , n360574 );
nand ( n50703 , n370909 , n370910 );
buf ( n370912 , n50703 );
buf ( n370913 , n370912 );
nand ( n50706 , n50688 , n370913 );
buf ( n370915 , n50706 );
xor ( n370916 , n370891 , n370915 );
buf ( n370917 , n370916 );
not ( n370918 , n370917 );
or ( n50711 , n50659 , n370918 );
buf ( n370920 , n370916 );
buf ( n370921 , n370865 );
or ( n50714 , n370920 , n370921 );
nand ( n370923 , n50711 , n50714 );
buf ( n370924 , n370923 );
buf ( n370925 , n370924 );
xor ( n370926 , n370835 , n370925 );
buf ( n370927 , n370318 );
not ( n370928 , n370927 );
buf ( n370929 , n370343 );
not ( n50722 , n370929 );
or ( n50723 , n370928 , n50722 );
buf ( n370932 , n50109 );
not ( n50725 , n370932 );
buf ( n370934 , n370343 );
not ( n370935 , n370934 );
buf ( n370936 , n370935 );
buf ( n370937 , n370936 );
not ( n50730 , n370937 );
or ( n370939 , n50725 , n50730 );
buf ( n370940 , n370372 );
nand ( n50733 , n370939 , n370940 );
buf ( n370942 , n50733 );
buf ( n370943 , n370942 );
nand ( n50736 , n50723 , n370943 );
buf ( n370945 , n50736 );
buf ( n370946 , n370945 );
xor ( n370947 , n370926 , n370946 );
buf ( n370948 , n370947 );
xnor ( n370949 , n370810 , n370948 );
buf ( n370950 , n370949 );
xor ( n50743 , n370757 , n370950 );
xor ( n50744 , n370248 , n370253 );
and ( n50745 , n50744 , n370270 );
and ( n50746 , n370248 , n370253 );
or ( n370955 , n50745 , n50746 );
buf ( n370956 , n370955 );
buf ( n370957 , n370956 );
not ( n370958 , n370510 );
not ( n370959 , n370958 );
not ( n50752 , n43274 );
and ( n370961 , n370959 , n50752 );
buf ( n370962 , n22772 );
not ( n50755 , n370962 );
buf ( n370964 , n362803 );
not ( n370965 , n370964 );
or ( n50758 , n50755 , n370965 );
buf ( n370967 , n40251 );
buf ( n370968 , n363444 );
nand ( n50761 , n370967 , n370968 );
buf ( n50762 , n50761 );
buf ( n370971 , n50762 );
nand ( n50764 , n50758 , n370971 );
buf ( n370973 , n50764 );
and ( n50766 , n370973 , n43261 );
nor ( n50767 , n370961 , n50766 );
buf ( n370976 , n50767 );
not ( n370977 , n370976 );
buf ( n370978 , n370977 );
buf ( n370979 , n370584 );
not ( n370980 , n370979 );
buf ( n370981 , n342654 );
buf ( n370982 , n342759 );
nor ( n50775 , n370981 , n370982 );
buf ( n370984 , n50775 );
not ( n50777 , n370984 );
not ( n370986 , n366393 );
not ( n50779 , n46204 );
nor ( n50780 , n370986 , n50779 );
nand ( n370989 , n50777 , n50780 );
buf ( n50782 , n370989 );
buf ( n370991 , n50782 );
not ( n370992 , n370991 );
and ( n370993 , n370980 , n370992 );
buf ( n370994 , n22710 );
not ( n370995 , n370994 );
buf ( n370996 , n46902 );
not ( n50789 , n370996 );
or ( n370998 , n370995 , n50789 );
buf ( n370999 , n45523 );
not ( n50792 , n370999 );
buf ( n371001 , n342657 );
nand ( n371002 , n50792 , n371001 );
buf ( n371003 , n371002 );
buf ( n371004 , n371003 );
nand ( n371005 , n370998 , n371004 );
buf ( n371006 , n371005 );
buf ( n371007 , n371006 );
buf ( n371008 , n366434 );
and ( n371009 , n371007 , n371008 );
nor ( n50802 , n370993 , n371009 );
buf ( n371011 , n50802 );
xor ( n50804 , n370978 , n371011 );
buf ( n371013 , n39207 );
buf ( n371014 , n370660 );
or ( n50807 , n371013 , n371014 );
buf ( n371016 , n39218 );
buf ( n371017 , n367576 );
not ( n50810 , n371017 );
buf ( n371019 , n35547 );
not ( n50812 , n371019 );
or ( n50813 , n50810 , n50812 );
buf ( n371022 , n366360 );
buf ( n371023 , n367575 );
buf ( n371024 , n371023 );
nand ( n50817 , n371022 , n371024 );
buf ( n371026 , n50817 );
buf ( n371027 , n371026 );
nand ( n371028 , n50813 , n371027 );
buf ( n371029 , n371028 );
buf ( n371030 , n371029 );
not ( n50823 , n371030 );
buf ( n371032 , n50823 );
buf ( n371033 , n371032 );
or ( n50826 , n371016 , n371033 );
nand ( n50827 , n50807 , n50826 );
buf ( n371036 , n50827 );
buf ( n371037 , n371036 );
not ( n50830 , n371037 );
buf ( n371039 , n50830 );
buf ( n371040 , n371039 );
not ( n50833 , n371040 );
buf ( n371042 , n50106 );
not ( n50835 , n371042 );
buf ( n371044 , n41882 );
not ( n50837 , n371044 );
and ( n50838 , n50835 , n50837 );
buf ( n371047 , n41892 );
not ( n50840 , n371047 );
buf ( n371049 , n43377 );
not ( n50842 , n371049 );
or ( n371051 , n50840 , n50842 );
buf ( n371052 , n45455 );
not ( n50845 , n371052 );
buf ( n371054 , n361716 );
nand ( n50847 , n50845 , n371054 );
buf ( n371056 , n50847 );
buf ( n371057 , n371056 );
nand ( n50850 , n371051 , n371057 );
buf ( n371059 , n50850 );
buf ( n371060 , n371059 );
buf ( n371061 , n365619 );
not ( n50854 , n371061 );
buf ( n371063 , n50854 );
buf ( n371064 , n371063 );
and ( n371065 , n371060 , n371064 );
nor ( n371066 , n50838 , n371065 );
buf ( n371067 , n371066 );
buf ( n371068 , n371067 );
not ( n50861 , n371068 );
buf ( n371070 , n365279 );
not ( n371071 , n371070 );
buf ( n371072 , n49993 );
not ( n50865 , n371072 );
or ( n371074 , n371071 , n50865 );
not ( n50867 , n40891 );
not ( n371076 , n50867 );
not ( n50869 , n44573 );
or ( n50870 , n371076 , n50869 );
not ( n50871 , n32085 );
buf ( n371080 , n50871 );
buf ( n371081 , n365267 );
nand ( n371082 , n371080 , n371081 );
buf ( n371083 , n371082 );
nand ( n50876 , n50870 , n371083 );
buf ( n371085 , n50876 );
buf ( n371086 , n40923 );
nand ( n371087 , n371085 , n371086 );
buf ( n371088 , n371087 );
buf ( n371089 , n371088 );
nand ( n50882 , n371074 , n371089 );
buf ( n371091 , n50882 );
buf ( n371092 , n371091 );
not ( n371093 , n371092 );
or ( n50886 , n50861 , n371093 );
buf ( n371095 , n371067 );
buf ( n371096 , n371091 );
or ( n50889 , n371095 , n371096 );
nand ( n371098 , n50886 , n50889 );
buf ( n371099 , n371098 );
buf ( n371100 , n371099 );
not ( n371101 , n371100 );
or ( n371102 , n50833 , n371101 );
buf ( n371103 , n371099 );
buf ( n371104 , n371039 );
or ( n50897 , n371103 , n371104 );
nand ( n50898 , n371102 , n50897 );
buf ( n371107 , n50898 );
xnor ( n50900 , n50804 , n371107 );
buf ( n371109 , n50900 );
xor ( n371110 , n370957 , n371109 );
xor ( n50903 , n370415 , n370440 );
and ( n50904 , n50903 , n370458 );
and ( n371113 , n370415 , n370440 );
or ( n371114 , n50904 , n371113 );
buf ( n371115 , n371114 );
buf ( n371116 , n371115 );
xor ( n371117 , n371110 , n371116 );
buf ( n371118 , n371117 );
buf ( n371119 , n371118 );
xor ( n50912 , n50743 , n371119 );
buf ( n371121 , n50912 );
xor ( n50914 , n370742 , n371121 );
xor ( n50915 , n370157 , n370273 );
and ( n371124 , n50915 , n370291 );
and ( n50917 , n370157 , n370273 );
or ( n371126 , n371124 , n50917 );
buf ( n371127 , n371126 );
buf ( n371128 , n371127 );
buf ( n50921 , n50090 );
not ( n50922 , n50921 );
buf ( n371131 , n370460 );
not ( n50924 , n371131 );
or ( n371133 , n50922 , n50924 );
not ( n371134 , n370296 );
not ( n50927 , n370297 );
nor ( n50928 , n50927 , n370460 );
not ( n371137 , n50928 );
or ( n371138 , n371134 , n371137 );
buf ( n371139 , n370390 );
not ( n371140 , n371139 );
buf ( n371141 , n371140 );
nand ( n50934 , n371138 , n371141 );
buf ( n371143 , n50934 );
nand ( n371144 , n371133 , n371143 );
buf ( n371145 , n371144 );
buf ( n371146 , n371145 );
xor ( n371147 , n371128 , n371146 );
buf ( n371148 , n50224 );
not ( n50941 , n45075 );
nand ( n371150 , n50941 , n365227 );
buf ( n371151 , n371150 );
nand ( n371152 , n371148 , n371151 );
buf ( n371153 , n371152 );
buf ( n371154 , n371153 );
buf ( n371155 , n365118 );
not ( n50948 , n371155 );
buf ( n371157 , n44819 );
not ( n371158 , n371157 );
buf ( n371159 , n40091 );
not ( n371160 , n371159 );
or ( n50953 , n371158 , n371160 );
buf ( n371162 , n40899 );
buf ( n371163 , n364997 );
nand ( n50956 , n371162 , n371163 );
buf ( n50957 , n50956 );
buf ( n371166 , n50957 );
nand ( n50959 , n50953 , n371166 );
buf ( n371168 , n50959 );
buf ( n371169 , n371168 );
not ( n50962 , n371169 );
or ( n371171 , n50948 , n50962 );
buf ( n371172 , n370404 );
buf ( n371173 , n365033 );
nand ( n371174 , n371172 , n371173 );
buf ( n371175 , n371174 );
buf ( n371176 , n371175 );
nand ( n50969 , n371171 , n371176 );
buf ( n371178 , n50969 );
buf ( n371179 , n371178 );
xor ( n371180 , n371154 , n371179 );
buf ( n371181 , n370318 );
buf ( n371182 , n361531 );
not ( n371183 , n371182 );
buf ( n371184 , n41615 );
not ( n371185 , n371184 );
or ( n371186 , n371183 , n371185 );
buf ( n371187 , n41607 );
buf ( n371188 , n361534 );
nand ( n50981 , n371187 , n371188 );
buf ( n50982 , n50981 );
buf ( n371191 , n50982 );
nand ( n50984 , n371186 , n371191 );
buf ( n50985 , n50984 );
not ( n371194 , n50985 );
not ( n50987 , n41482 );
not ( n371196 , n50987 );
or ( n371197 , n371194 , n371196 );
not ( n371198 , n364852 );
nand ( n50991 , n371198 , n370174 );
nand ( n371200 , n371197 , n50991 );
buf ( n371201 , n371200 );
xor ( n50994 , n371181 , n371201 );
buf ( n371203 , n370366 );
not ( n371204 , n371203 );
buf ( n371205 , n359916 );
not ( n371206 , n371205 );
or ( n371207 , n371204 , n371206 );
buf ( n371208 , n368038 );
buf ( n371209 , n351294 );
not ( n371210 , n371209 );
buf ( n371211 , n42455 );
not ( n371212 , n371211 );
or ( n371213 , n371210 , n371212 );
buf ( n371214 , n366243 );
buf ( n371215 , n365464 );
nand ( n51008 , n371214 , n371215 );
buf ( n371217 , n51008 );
buf ( n371218 , n371217 );
nand ( n371219 , n371213 , n371218 );
buf ( n371220 , n371219 );
buf ( n371221 , n371220 );
nand ( n371222 , n371208 , n371221 );
buf ( n371223 , n371222 );
buf ( n371224 , n371223 );
nand ( n371225 , n371207 , n371224 );
buf ( n371226 , n371225 );
buf ( n371227 , n371226 );
xnor ( n371228 , n50994 , n371227 );
buf ( n371229 , n371228 );
buf ( n371230 , n371229 );
xor ( n371231 , n371180 , n371230 );
buf ( n371232 , n371231 );
buf ( n371233 , n371232 );
buf ( n371234 , n370375 );
not ( n51022 , n371234 );
buf ( n371236 , n370387 );
not ( n371237 , n371236 );
or ( n51025 , n51022 , n371237 );
buf ( n371239 , n370303 );
nand ( n51027 , n51025 , n371239 );
buf ( n371241 , n51027 );
buf ( n371242 , n371241 );
buf ( n371243 , n370387 );
buf ( n371244 , n370375 );
or ( n51032 , n371243 , n371244 );
buf ( n371246 , n51032 );
buf ( n371247 , n371246 );
nand ( n371248 , n371242 , n371247 );
buf ( n371249 , n371248 );
buf ( n371250 , n371249 );
xor ( n371251 , n371233 , n371250 );
buf ( n371252 , n365676 );
not ( n51040 , n371252 );
not ( n371254 , n359974 );
buf ( n371255 , n371254 );
not ( n51043 , n371255 );
or ( n371257 , n51040 , n51043 );
buf ( n371258 , n359974 );
buf ( n371259 , n365673 );
nand ( n51047 , n371258 , n371259 );
buf ( n371261 , n51047 );
buf ( n371262 , n371261 );
nand ( n51050 , n371257 , n371262 );
buf ( n371264 , n51050 );
buf ( n51052 , n371264 );
not ( n51053 , n51052 );
buf ( n51054 , n51053 );
buf ( n371268 , n51054 );
not ( n51056 , n371268 );
buf ( n371270 , n45492 );
not ( n371271 , n371270 );
buf ( n371272 , n371271 );
buf ( n371273 , n371272 );
not ( n51061 , n371273 );
and ( n371275 , n51056 , n51061 );
buf ( n371276 , n370450 );
buf ( n371277 , n45553 );
and ( n371278 , n371276 , n371277 );
nor ( n371279 , n371275 , n371278 );
buf ( n371280 , n371279 );
buf ( n371281 , n366654 );
not ( n51069 , n371281 );
buf ( n371283 , n46477 );
not ( n371284 , n371283 );
buf ( n371285 , n44925 );
not ( n371286 , n371285 );
or ( n51074 , n371284 , n371286 );
buf ( n51075 , n44926 );
buf ( n51076 , n366683 );
nand ( n51077 , n51075 , n51076 );
buf ( n371291 , n51077 );
buf ( n371292 , n371291 );
nand ( n371293 , n51074 , n371292 );
buf ( n371294 , n371293 );
buf ( n371295 , n371294 );
not ( n51083 , n371295 );
or ( n371297 , n51069 , n51083 );
buf ( n371298 , n46521 );
not ( n371299 , n371298 );
buf ( n371300 , n371299 );
buf ( n371301 , n371300 );
not ( n371302 , n371301 );
buf ( n371303 , n50056 );
nand ( n51091 , n371302 , n371303 );
buf ( n371305 , n51091 );
buf ( n371306 , n371305 );
nand ( n371307 , n371297 , n371306 );
buf ( n371308 , n371307 );
xor ( n371309 , n371280 , n371308 );
buf ( n371310 , n370539 );
not ( n51098 , n371310 );
buf ( n371312 , n370520 );
not ( n51100 , n371312 );
or ( n51101 , n51098 , n51100 );
or ( n371315 , n370539 , n370520 );
nand ( n51103 , n371315 , n370496 );
buf ( n371317 , n51103 );
nand ( n51105 , n51101 , n371317 );
buf ( n371319 , n51105 );
xor ( n51107 , n371309 , n371319 );
buf ( n371321 , n51107 );
xnor ( n371322 , n371251 , n371321 );
buf ( n371323 , n371322 );
buf ( n371324 , n371323 );
xor ( n51112 , n371147 , n371324 );
buf ( n371326 , n51112 );
xor ( n51114 , n50914 , n371326 );
buf ( n371328 , n51114 );
xor ( n51116 , n370729 , n371328 );
buf ( n371330 , n51116 );
buf ( n371331 , n371330 );
xor ( n371332 , n370294 , n370463 );
xor ( n51120 , n371332 , n370482 );
buf ( n371334 , n51120 );
buf ( n371335 , n371334 );
and ( n371336 , n50497 , n370695 );
not ( n371337 , n50497 );
and ( n51125 , n371337 , n50488 );
nor ( n371339 , n371336 , n51125 );
and ( n371340 , n371339 , n50511 );
not ( n51128 , n371339 );
not ( n371342 , n50511 );
and ( n371343 , n51128 , n371342 );
nor ( n51131 , n371340 , n371343 );
buf ( n371345 , n51131 );
xor ( n51133 , n371335 , n371345 );
buf ( n371347 , n367981 );
not ( n51135 , n371347 );
buf ( n51136 , n367718 );
buf ( n371350 , n51136 );
buf ( n371351 , n371350 );
buf ( n371352 , n371351 );
nand ( n371353 , n51135 , n371352 );
buf ( n371354 , n371353 );
buf ( n371355 , n371354 );
not ( n371356 , n371355 );
buf ( n371357 , n368386 );
not ( n51145 , n371357 );
or ( n371359 , n371356 , n51145 );
buf ( n371360 , n371351 );
not ( n371361 , n371360 );
buf ( n371362 , n367981 );
nand ( n51150 , n371361 , n371362 );
buf ( n371364 , n51150 );
buf ( n371365 , n371364 );
nand ( n51153 , n371359 , n371365 );
buf ( n51154 , n51153 );
buf ( n371368 , n51154 );
and ( n51156 , n51133 , n371368 );
and ( n371370 , n371335 , n371345 );
or ( n51158 , n51156 , n371370 );
buf ( n371372 , n51158 );
buf ( n371373 , n371372 );
nor ( n371374 , n371331 , n371373 );
buf ( n371375 , n371374 );
buf ( n371376 , n371375 );
not ( n371377 , n371376 );
buf ( n371378 , n371377 );
xor ( n51166 , n371128 , n371146 );
and ( n371380 , n51166 , n371324 );
and ( n371381 , n371128 , n371146 );
or ( n371382 , n371380 , n371381 );
buf ( n371383 , n371382 );
buf ( n371384 , n371383 );
xor ( n371385 , n370742 , n371121 );
and ( n51173 , n371385 , n371326 );
and ( n371387 , n370742 , n371121 );
or ( n371388 , n51173 , n371387 );
buf ( n371389 , n371388 );
xor ( n371390 , n371384 , n371389 );
not ( n51178 , n370948 );
not ( n51179 , n370761 );
nand ( n51180 , n51179 , n370809 );
not ( n51181 , n51180 );
or ( n371395 , n51178 , n51181 );
buf ( n371396 , n50563 );
buf ( n371397 , n370799 );
xor ( n371398 , n371396 , n371397 );
buf ( n371399 , n370806 );
xnor ( n371400 , n371398 , n371399 );
buf ( n371401 , n371400 );
buf ( n371402 , n371401 );
not ( n51190 , n371402 );
buf ( n371404 , n370761 );
nand ( n371405 , n51190 , n371404 );
buf ( n371406 , n371405 );
nand ( n51194 , n371395 , n371406 );
not ( n51195 , n51194 );
buf ( n371409 , n366654 );
not ( n371410 , n371409 );
buf ( n371411 , n46477 );
not ( n371412 , n371411 );
buf ( n371413 , n366600 );
not ( n371414 , n371413 );
or ( n51202 , n371412 , n371414 );
not ( n371416 , n366600 );
buf ( n51204 , n371416 );
buf ( n51205 , n366683 );
nand ( n51206 , n51204 , n51205 );
buf ( n51207 , n51206 );
buf ( n371421 , n51207 );
nand ( n51209 , n51202 , n371421 );
buf ( n51210 , n51209 );
buf ( n51211 , n51210 );
not ( n51212 , n51211 );
or ( n51213 , n371410 , n51212 );
buf ( n51214 , n371294 );
buf ( n371428 , n46521 );
nand ( n371429 , n51214 , n371428 );
buf ( n371430 , n371429 );
buf ( n371431 , n371430 );
nand ( n51219 , n51213 , n371431 );
buf ( n371433 , n51219 );
buf ( n371434 , n371433 );
buf ( n371435 , n371011 );
not ( n371436 , n371435 );
buf ( n371437 , n371436 );
not ( n371438 , n371437 );
not ( n51226 , n370978 );
or ( n51227 , n371438 , n51226 );
not ( n371441 , n371011 );
not ( n371442 , n50767 );
or ( n51230 , n371441 , n371442 );
nand ( n51231 , n51230 , n371107 );
nand ( n371445 , n51227 , n51231 );
buf ( n371446 , n371445 );
xor ( n371447 , n371434 , n371446 );
buf ( n371448 , n42242 );
not ( n371449 , n371448 );
buf ( n371450 , n366209 );
not ( n51238 , n371450 );
buf ( n371452 , n366673 );
not ( n371453 , n371452 );
or ( n51241 , n51238 , n371453 );
buf ( n371455 , n362458 );
buf ( n371456 , n366212 );
nand ( n51244 , n371455 , n371456 );
buf ( n371458 , n51244 );
buf ( n371459 , n371458 );
nand ( n51247 , n51241 , n371459 );
buf ( n371461 , n51247 );
buf ( n371462 , n371461 );
not ( n51250 , n371462 );
or ( n371464 , n371449 , n51250 );
buf ( n371465 , n370827 );
buf ( n371466 , n42263 );
nand ( n371467 , n371465 , n371466 );
buf ( n371468 , n371467 );
buf ( n371469 , n371468 );
nand ( n371470 , n371464 , n371469 );
buf ( n371471 , n371470 );
buf ( n371472 , n371471 );
not ( n371473 , n370891 );
buf ( n371474 , n370915 );
not ( n371475 , n371474 );
buf ( n371476 , n370865 );
nand ( n371477 , n371475 , n371476 );
buf ( n371478 , n371477 );
not ( n51266 , n371478 );
or ( n51267 , n371473 , n51266 );
buf ( n371481 , n370862 );
buf ( n371482 , n370915 );
nand ( n51270 , n371481 , n371482 );
buf ( n371484 , n51270 );
nand ( n51272 , n51267 , n371484 );
buf ( n371486 , n51272 );
xor ( n371487 , n371472 , n371486 );
buf ( n371488 , n41835 );
not ( n51276 , n371488 );
buf ( n371490 , n47554 );
not ( n371491 , n371490 );
buf ( n371492 , n366407 );
not ( n371493 , n371492 );
or ( n51281 , n371491 , n371493 );
buf ( n371495 , n362285 );
buf ( n371496 , n41772 );
nand ( n51284 , n371495 , n371496 );
buf ( n371498 , n51284 );
buf ( n371499 , n371498 );
nand ( n371500 , n51281 , n371499 );
buf ( n371501 , n371500 );
buf ( n371502 , n371501 );
not ( n51290 , n371502 );
or ( n371504 , n51276 , n51290 );
buf ( n371505 , n370789 );
buf ( n371506 , n41830 );
nand ( n51294 , n371505 , n371506 );
buf ( n371508 , n51294 );
buf ( n371509 , n371508 );
nand ( n51297 , n371504 , n371509 );
buf ( n371511 , n51297 );
buf ( n371512 , n371511 );
not ( n371513 , n371512 );
buf ( n371514 , n371513 );
buf ( n371515 , n371514 );
xnor ( n371516 , n371487 , n371515 );
buf ( n371517 , n371516 );
buf ( n371518 , n371517 );
xor ( n371519 , n371447 , n371518 );
buf ( n371520 , n371519 );
not ( n51308 , n371520 );
not ( n371522 , n51308 );
and ( n51310 , n51195 , n371522 );
and ( n51311 , n51194 , n51308 );
nor ( n371525 , n51310 , n51311 );
xor ( n371526 , n370835 , n370925 );
and ( n51314 , n371526 , n370946 );
and ( n371528 , n370835 , n370925 );
or ( n51316 , n51314 , n371528 );
buf ( n371530 , n51316 );
buf ( n371531 , n371530 );
buf ( n371532 , n45492 );
not ( n51320 , n371532 );
and ( n51321 , n40005 , n365673 );
not ( n51322 , n40005 );
and ( n371536 , n51322 , n365676 );
or ( n371537 , n51321 , n371536 );
buf ( n371538 , n371537 );
not ( n371539 , n371538 );
or ( n51327 , n51320 , n371539 );
buf ( n371541 , n371264 );
buf ( n371542 , n45553 );
nand ( n371543 , n371541 , n371542 );
buf ( n371544 , n371543 );
buf ( n371545 , n371544 );
nand ( n51333 , n51327 , n371545 );
buf ( n371547 , n51333 );
buf ( n371548 , n371547 );
not ( n371549 , n371200 );
not ( n51337 , n50109 );
or ( n51338 , n371549 , n51337 );
not ( n371552 , n370318 );
buf ( n371553 , n50985 );
buf ( n371554 , n50987 );
and ( n371555 , n371553 , n371554 );
buf ( n371556 , n370174 );
not ( n51344 , n371556 );
buf ( n371558 , n364852 );
nor ( n371559 , n51344 , n371558 );
buf ( n371560 , n371559 );
buf ( n371561 , n371560 );
nor ( n371562 , n371555 , n371561 );
buf ( n371563 , n371562 );
not ( n371564 , n371563 );
or ( n51352 , n371552 , n371564 );
nand ( n51353 , n51352 , n371226 );
nand ( n51354 , n51338 , n51353 );
buf ( n371568 , n51354 );
xor ( n371569 , n371548 , n371568 );
buf ( n371570 , n366402 );
not ( n371571 , n371570 );
buf ( n371572 , n371006 );
not ( n51360 , n371572 );
or ( n51361 , n371571 , n51360 );
buf ( n371575 , n22710 );
not ( n51363 , n371575 );
buf ( n371577 , n370257 );
not ( n371578 , n371577 );
or ( n51366 , n51363 , n371578 );
buf ( n371580 , n359778 );
buf ( n371581 , n342657 );
nand ( n51369 , n371580 , n371581 );
buf ( n371583 , n51369 );
buf ( n371584 , n371583 );
nand ( n371585 , n51366 , n371584 );
buf ( n371586 , n371585 );
buf ( n371587 , n371586 );
buf ( n371588 , n366434 );
nand ( n51376 , n371587 , n371588 );
buf ( n371590 , n51376 );
buf ( n371591 , n371590 );
nand ( n371592 , n51361 , n371591 );
buf ( n371593 , n371592 );
buf ( n371594 , n371593 );
xor ( n371595 , n371569 , n371594 );
buf ( n371596 , n371595 );
buf ( n371597 , n371596 );
xor ( n371598 , n371531 , n371597 );
not ( n51386 , n363429 );
not ( n371600 , n370973 );
or ( n51388 , n51386 , n371600 );
and ( n51389 , n367378 , n363444 );
not ( n371603 , n367378 );
and ( n51391 , n371603 , n22772 );
or ( n371605 , n51389 , n51391 );
nand ( n51393 , n371605 , n43261 );
nand ( n371607 , n51388 , n51393 );
buf ( n371608 , n50876 );
not ( n371609 , n371608 );
buf ( n371610 , n361013 );
not ( n371611 , n371610 );
or ( n371612 , n371609 , n371611 );
buf ( n371613 , n365293 );
not ( n371614 , n371613 );
buf ( n371615 , n46126 );
not ( n371616 , n371615 );
or ( n371617 , n371614 , n371616 );
buf ( n371618 , n40891 );
buf ( n371619 , n362534 );
nand ( n51407 , n371618 , n371619 );
buf ( n371621 , n51407 );
buf ( n371622 , n371621 );
nand ( n51410 , n371617 , n371622 );
buf ( n371624 , n51410 );
buf ( n371625 , n371624 );
buf ( n371626 , n40923 );
nand ( n371627 , n371625 , n371626 );
buf ( n371628 , n371627 );
buf ( n371629 , n371628 );
nand ( n51417 , n371612 , n371629 );
buf ( n371631 , n51417 );
buf ( n371632 , n371631 );
not ( n371633 , n371632 );
buf ( n371634 , n371633 );
buf ( n371635 , n371634 );
buf ( n371636 , n370885 );
not ( n51424 , n371636 );
buf ( n371638 , n45795 );
not ( n371639 , n371638 );
or ( n371640 , n51424 , n371639 );
buf ( n371641 , n367796 );
buf ( n371642 , n365440 );
not ( n371643 , n371642 );
buf ( n371644 , n45231 );
not ( n51432 , n371644 );
or ( n371646 , n371643 , n51432 );
buf ( n371647 , n45234 );
buf ( n371648 , n365452 );
nand ( n371649 , n371647 , n371648 );
buf ( n371650 , n371649 );
buf ( n371651 , n371650 );
nand ( n51439 , n371646 , n371651 );
buf ( n371653 , n51439 );
buf ( n371654 , n371653 );
nand ( n51442 , n371641 , n371654 );
buf ( n371656 , n51442 );
buf ( n371657 , n371656 );
nand ( n51445 , n371640 , n371657 );
buf ( n51446 , n51445 );
buf ( n371660 , n51446 );
xor ( n51448 , n371635 , n371660 );
buf ( n371662 , n371029 );
not ( n371663 , n371662 );
buf ( n371664 , n45204 );
not ( n371665 , n371664 );
or ( n51453 , n371663 , n371665 );
buf ( n371667 , n364870 );
not ( n371668 , n371667 );
buf ( n371669 , n371668 );
and ( n371670 , n371669 , n366356 );
not ( n51458 , n371669 );
and ( n51459 , n51458 , n366360 );
nor ( n371673 , n371670 , n51459 );
buf ( n371674 , n371673 );
not ( n371675 , n371674 );
buf ( n371676 , n359312 );
nand ( n371677 , n371675 , n371676 );
buf ( n371678 , n371677 );
buf ( n371679 , n371678 );
nand ( n371680 , n51453 , n371679 );
buf ( n371681 , n371680 );
buf ( n371682 , n371681 );
xor ( n371683 , n51448 , n371682 );
buf ( n371684 , n371683 );
xor ( n371685 , n371607 , n371684 );
buf ( n371686 , n362027 );
not ( n371687 , n371686 );
buf ( n371688 , n371059 );
not ( n371689 , n371688 );
or ( n371690 , n371687 , n371689 );
buf ( n371691 , n45455 );
not ( n371692 , n371691 );
buf ( n371693 , n365760 );
not ( n371694 , n371693 );
or ( n371695 , n371692 , n371694 );
buf ( n371696 , n41528 );
buf ( n371697 , n364832 );
nand ( n371698 , n371696 , n371697 );
buf ( n371699 , n371698 );
buf ( n371700 , n371699 );
nand ( n51468 , n371695 , n371700 );
buf ( n371702 , n51468 );
buf ( n371703 , n371702 );
buf ( n371704 , n365622 );
nand ( n371705 , n371703 , n371704 );
buf ( n371706 , n371705 );
buf ( n371707 , n371706 );
nand ( n51471 , n371690 , n371707 );
buf ( n371709 , n51471 );
buf ( n371710 , n371709 );
buf ( n51474 , n370908 );
not ( n51475 , n51474 );
buf ( n371713 , n40475 );
not ( n51477 , n371713 );
or ( n51478 , n51475 , n51477 );
buf ( n371716 , n351762 );
not ( n51480 , n371716 );
buf ( n371718 , n45270 );
not ( n51482 , n371718 );
or ( n51483 , n51480 , n51482 );
buf ( n371721 , n42911 );
not ( n51485 , n371721 );
buf ( n371723 , n365471 );
nand ( n51487 , n51485 , n371723 );
buf ( n371725 , n51487 );
buf ( n371726 , n371725 );
nand ( n371727 , n51483 , n371726 );
buf ( n371728 , n371727 );
buf ( n371729 , n371728 );
buf ( n371730 , n360583 );
not ( n371731 , n371730 );
buf ( n371732 , n371731 );
buf ( n371733 , n371732 );
nand ( n371734 , n371729 , n371733 );
buf ( n371735 , n371734 );
buf ( n371736 , n371735 );
nand ( n51500 , n51478 , n371736 );
buf ( n371738 , n51500 );
buf ( n371739 , n371738 );
xor ( n371740 , n371710 , n371739 );
buf ( n371741 , n370855 );
not ( n371742 , n371741 );
buf ( n371743 , n40058 );
not ( n51507 , n371743 );
or ( n371745 , n371742 , n51507 );
and ( n371746 , n351320 , n363122 );
not ( n51510 , n351320 );
and ( n371748 , n51510 , n363119 );
or ( n51512 , n371746 , n371748 );
nand ( n51513 , n39946 , n51512 );
buf ( n371751 , n51513 );
nand ( n51515 , n371745 , n371751 );
buf ( n371753 , n51515 );
buf ( n371754 , n371753 );
xor ( n371755 , n371740 , n371754 );
buf ( n371756 , n371755 );
xor ( n371757 , n371685 , n371756 );
buf ( n371758 , n371757 );
xor ( n371759 , n371598 , n371758 );
buf ( n371760 , n371759 );
and ( n51524 , n371525 , n371760 );
not ( n371762 , n371525 );
buf ( n371763 , n371760 );
not ( n371764 , n371763 );
buf ( n371765 , n371764 );
and ( n51529 , n371762 , n371765 );
nor ( n371767 , n51524 , n51529 );
not ( n371768 , n371767 );
xor ( n51532 , n370757 , n370950 );
and ( n51533 , n51532 , n371119 );
and ( n371771 , n370757 , n370950 );
or ( n51535 , n51533 , n371771 );
buf ( n371773 , n51535 );
not ( n371774 , n371773 );
and ( n51538 , n371768 , n371774 );
not ( n371776 , n371768 );
and ( n51540 , n371776 , n371773 );
nor ( n51541 , n51538 , n51540 );
xor ( n51542 , n371154 , n371179 );
and ( n51543 , n51542 , n371230 );
and ( n371781 , n371154 , n371179 );
or ( n371782 , n51543 , n371781 );
buf ( n371783 , n371782 );
buf ( n371784 , n371783 );
buf ( n371785 , n371280 );
not ( n51549 , n371785 );
buf ( n51550 , n51549 );
buf ( n371788 , n51550 );
not ( n51552 , n371788 );
buf ( n371790 , n371308 );
not ( n51554 , n371790 );
or ( n371792 , n51552 , n51554 );
buf ( n371793 , n371308 );
buf ( n371794 , n51550 );
or ( n51558 , n371793 , n371794 );
buf ( n371796 , n371319 );
nand ( n371797 , n51558 , n371796 );
buf ( n371798 , n371797 );
buf ( n371799 , n371798 );
nand ( n371800 , n371792 , n371799 );
buf ( n371801 , n371800 );
buf ( n371802 , n371801 );
xor ( n371803 , n371784 , n371802 );
buf ( n371804 , n365033 );
not ( n51568 , n371804 );
buf ( n371806 , n371168 );
not ( n371807 , n371806 );
or ( n51571 , n51568 , n371807 );
buf ( n371809 , n44819 );
not ( n371810 , n371809 );
buf ( n371811 , n363439 );
not ( n371812 , n371811 );
or ( n371813 , n371810 , n371812 );
buf ( n371814 , n363442 );
buf ( n371815 , n364997 );
nand ( n371816 , n371814 , n371815 );
buf ( n371817 , n371816 );
buf ( n371818 , n371817 );
nand ( n51582 , n371813 , n371818 );
buf ( n371820 , n51582 );
buf ( n371821 , n371820 );
buf ( n371822 , n365118 );
nand ( n371823 , n371821 , n371822 );
buf ( n371824 , n371823 );
buf ( n371825 , n371824 );
nand ( n51589 , n51571 , n371825 );
buf ( n371827 , n51589 );
buf ( n371828 , n371827 );
buf ( n371829 , n371220 );
not ( n51593 , n371829 );
buf ( n371831 , n368051 );
not ( n51595 , n371831 );
or ( n51596 , n51593 , n51595 );
buf ( n371834 , n352212 );
buf ( n371835 , n364909 );
and ( n51599 , n371834 , n371835 );
not ( n51600 , n371834 );
buf ( n371838 , n366243 );
and ( n371839 , n51600 , n371838 );
nor ( n371840 , n51599 , n371839 );
buf ( n371841 , n371840 );
buf ( n371842 , n371841 );
not ( n51606 , n371842 );
buf ( n371844 , n366237 );
not ( n51608 , n371844 );
buf ( n371846 , n51608 );
buf ( n371847 , n371846 );
nand ( n371848 , n51606 , n371847 );
buf ( n371849 , n371848 );
buf ( n371850 , n371849 );
nand ( n371851 , n51596 , n371850 );
buf ( n371852 , n371851 );
buf ( n371853 , n371852 );
buf ( n371854 , n363603 );
not ( n51618 , n371854 );
buf ( n371856 , n363317 );
not ( n371857 , n371856 );
or ( n51621 , n51618 , n371857 );
buf ( n371859 , n41663 );
buf ( n371860 , n361534 );
nand ( n51624 , n371859 , n371860 );
buf ( n371862 , n51624 );
buf ( n371863 , n371862 );
nand ( n51627 , n51621 , n371863 );
buf ( n371865 , n51627 );
not ( n371866 , n371865 );
not ( n51630 , n41485 );
or ( n371868 , n371866 , n51630 );
nand ( n371869 , n50985 , n361606 );
nand ( n51633 , n371868 , n371869 );
buf ( n371871 , n51633 );
xor ( n371872 , n371853 , n371871 );
buf ( n371873 , n371091 );
not ( n51637 , n371873 );
buf ( n371875 , n51637 );
buf ( n371876 , n371875 );
not ( n371877 , n371876 );
buf ( n371878 , n371067 );
not ( n371879 , n371878 );
or ( n51643 , n371877 , n371879 );
buf ( n371881 , n371036 );
nand ( n51645 , n51643 , n371881 );
buf ( n371883 , n51645 );
buf ( n51647 , n371883 );
buf ( n371885 , n371067 );
buf ( n371886 , n371875 );
or ( n371887 , n371885 , n371886 );
buf ( n371888 , n371887 );
buf ( n371889 , n371888 );
nand ( n371890 , n51647 , n371889 );
buf ( n371891 , n371890 );
buf ( n371892 , n371891 );
xor ( n371893 , n371872 , n371892 );
buf ( n371894 , n371893 );
buf ( n371895 , n371894 );
xor ( n51659 , n371828 , n371895 );
buf ( n371897 , n50563 );
not ( n51661 , n371897 );
buf ( n51662 , n370799 );
not ( n51663 , n51662 );
or ( n51664 , n51661 , n51663 );
or ( n371902 , n50563 , n370799 );
nand ( n51666 , n371902 , n370806 );
buf ( n371904 , n51666 );
nand ( n51668 , n51664 , n371904 );
buf ( n371906 , n51668 );
buf ( n371907 , n371906 );
xor ( n51671 , n51659 , n371907 );
buf ( n371909 , n51671 );
buf ( n371910 , n371909 );
xnor ( n51674 , n371803 , n371910 );
buf ( n371912 , n51674 );
not ( n371913 , n371912 );
not ( n51677 , n371913 );
xor ( n371915 , n370957 , n371109 );
and ( n371916 , n371915 , n371116 );
and ( n51680 , n370957 , n371109 );
or ( n371918 , n371916 , n51680 );
buf ( n371919 , n371918 );
buf ( n371920 , n371919 );
not ( n51684 , n371920 );
buf ( n51685 , n51684 );
buf ( n371923 , n51685 );
not ( n51687 , n371923 );
buf ( n371925 , n371232 );
not ( n371926 , n371925 );
buf ( n371927 , n51107 );
nand ( n371928 , n371926 , n371927 );
buf ( n371929 , n371928 );
buf ( n371930 , n371929 );
buf ( n371931 , n371249 );
and ( n51695 , n371930 , n371931 );
buf ( n371933 , n371232 );
not ( n51697 , n371933 );
buf ( n51698 , n51107 );
nor ( n51699 , n51697 , n51698 );
buf ( n51700 , n51699 );
buf ( n371938 , n51700 );
nor ( n51702 , n51695 , n371938 );
buf ( n51703 , n51702 );
buf ( n371941 , n51703 );
not ( n51705 , n371941 );
buf ( n371943 , n51705 );
buf ( n371944 , n371943 );
not ( n371945 , n371944 );
or ( n51709 , n51687 , n371945 );
buf ( n371947 , n51703 );
buf ( n371948 , n371919 );
nand ( n371949 , n371947 , n371948 );
buf ( n371950 , n371949 );
buf ( n371951 , n371950 );
nand ( n371952 , n51709 , n371951 );
buf ( n371953 , n371952 );
not ( n51717 , n371953 );
or ( n371955 , n51677 , n51717 );
or ( n51719 , n371953 , n371913 );
nand ( n371957 , n371955 , n51719 );
buf ( n371958 , n371957 );
not ( n51722 , n371958 );
buf ( n371960 , n51722 );
and ( n371961 , n51541 , n371960 );
not ( n51725 , n51541 );
buf ( n371963 , n371957 );
and ( n371964 , n51725 , n371963 );
nor ( n51728 , n371961 , n371964 );
buf ( n371966 , n51728 );
xnor ( n371967 , n371390 , n371966 );
buf ( n371968 , n371967 );
xor ( n51732 , n370487 , n370728 );
and ( n371970 , n51732 , n371328 );
and ( n371971 , n370487 , n370728 );
or ( n51735 , n371970 , n371971 );
buf ( n371973 , n51735 );
nor ( n371974 , n371968 , n371973 );
not ( n51738 , n371974 );
xor ( n371976 , n371335 , n371345 );
xor ( n371977 , n371976 , n371368 );
buf ( n371978 , n371977 );
buf ( n371979 , n371978 );
not ( n51743 , n371979 );
buf ( n371981 , n51743 );
buf ( n51745 , n371981 );
buf ( n371983 , n367078 );
not ( n51747 , n371983 );
buf ( n51748 , n51747 );
not ( n371986 , n51748 );
buf ( n371987 , n48198 );
not ( n371988 , n371987 );
buf ( n371989 , n371988 );
not ( n51753 , n371989 );
and ( n371991 , n371986 , n51753 );
buf ( n371992 , n371989 );
buf ( n371993 , n51748 );
nand ( n51757 , n371992 , n371993 );
buf ( n371995 , n51757 );
and ( n51759 , n371995 , n369158 );
nor ( n371997 , n371991 , n51759 );
buf ( n371998 , n371997 );
nand ( n371999 , n51745 , n371998 );
buf ( n372000 , n371999 );
and ( n372001 , n49930 , n371378 , n51738 , n372000 );
buf ( n372002 , n371757 );
not ( n372003 , n372002 );
buf ( n372004 , n371596 );
not ( n51768 , n372004 );
or ( n372006 , n372003 , n51768 );
buf ( n372007 , n371596 );
buf ( n372008 , n371757 );
or ( n372009 , n372007 , n372008 );
buf ( n51773 , n371530 );
nand ( n51774 , n372009 , n51773 );
buf ( n51775 , n51774 );
buf ( n372013 , n51775 );
nand ( n51777 , n372006 , n372013 );
buf ( n372015 , n51777 );
buf ( n372016 , n372015 );
not ( n51780 , n372016 );
buf ( n372018 , n51780 );
not ( n372019 , n372018 );
buf ( n372020 , n366434 );
not ( n372021 , n372020 );
buf ( n372022 , n22710 );
not ( n51786 , n372022 );
buf ( n372024 , n362212 );
not ( n372025 , n372024 );
or ( n51789 , n51786 , n372025 );
buf ( n372027 , n359756 );
buf ( n372028 , n342657 );
nand ( n372029 , n372027 , n372028 );
buf ( n372030 , n372029 );
buf ( n372031 , n372030 );
nand ( n51795 , n51789 , n372031 );
buf ( n372033 , n51795 );
buf ( n372034 , n372033 );
not ( n372035 , n372034 );
or ( n51799 , n372021 , n372035 );
buf ( n372037 , n371586 );
buf ( n372038 , n366402 );
nand ( n372039 , n372037 , n372038 );
buf ( n372040 , n372039 );
buf ( n372041 , n372040 );
nand ( n372042 , n51799 , n372041 );
buf ( n372043 , n372042 );
buf ( n372044 , n372043 );
not ( n51808 , n371471 );
nand ( n372046 , n51808 , n371514 );
and ( n372047 , n372046 , n51272 );
and ( n51811 , n371511 , n371471 );
nor ( n372049 , n372047 , n51811 );
buf ( n372050 , n372049 );
not ( n51814 , n372050 );
buf ( n51815 , n51814 );
buf ( n372053 , n51815 );
xor ( n51817 , n372044 , n372053 );
buf ( n372055 , n371607 );
buf ( n372056 , n371684 );
or ( n372057 , n372055 , n372056 );
buf ( n372058 , n371756 );
nand ( n51822 , n372057 , n372058 );
buf ( n372060 , n51822 );
buf ( n372061 , n372060 );
buf ( n372062 , n371607 );
buf ( n51826 , n371684 );
nand ( n51827 , n372062 , n51826 );
buf ( n372065 , n51827 );
buf ( n372066 , n372065 );
nand ( n372067 , n372061 , n372066 );
buf ( n372068 , n372067 );
buf ( n372069 , n372068 );
xnor ( n372070 , n51817 , n372069 );
buf ( n372071 , n372070 );
buf ( n372072 , n372071 );
not ( n51836 , n372072 );
buf ( n372074 , n51836 );
not ( n51838 , n372074 );
xor ( n51839 , n371434 , n371446 );
and ( n372077 , n51839 , n371518 );
and ( n372078 , n371434 , n371446 );
or ( n51842 , n372077 , n372078 );
buf ( n372080 , n51842 );
buf ( n51844 , n372080 );
not ( n372082 , n51844 );
buf ( n372083 , n372082 );
not ( n372084 , n372083 );
or ( n372085 , n51838 , n372084 );
buf ( n372086 , n372071 );
buf ( n372087 , n372080 );
nand ( n372088 , n372086 , n372087 );
buf ( n372089 , n372088 );
nand ( n51853 , n372085 , n372089 );
not ( n51854 , n51853 );
or ( n372092 , n372019 , n51854 );
or ( n372093 , n372018 , n51853 );
nand ( n51857 , n372092 , n372093 );
buf ( n372095 , n371520 );
not ( n51859 , n372095 );
buf ( n372097 , n371760 );
not ( n51861 , n372097 );
or ( n372099 , n51859 , n51861 );
buf ( n372100 , n371760 );
buf ( n372101 , n371520 );
or ( n372102 , n372100 , n372101 );
buf ( n372103 , n51194 );
nand ( n372104 , n372102 , n372103 );
buf ( n372105 , n372104 );
buf ( n372106 , n372105 );
nand ( n372107 , n372099 , n372106 );
buf ( n372108 , n372107 );
xor ( n372109 , n51857 , n372108 );
not ( n372110 , n371913 );
not ( n372111 , n371919 );
or ( n51875 , n372110 , n372111 );
not ( n372113 , n51685 );
not ( n372114 , n371912 );
or ( n51878 , n372113 , n372114 );
nand ( n372116 , n51878 , n371943 );
nand ( n51880 , n51875 , n372116 );
and ( n51881 , n372109 , n51880 );
and ( n372119 , n51857 , n372108 );
or ( n372120 , n51881 , n372119 );
buf ( n372121 , n372120 );
not ( n372122 , n372121 );
buf ( n372123 , n372071 );
not ( n372124 , n372123 );
buf ( n372125 , n372083 );
not ( n51889 , n372125 );
or ( n372127 , n372124 , n51889 );
buf ( n372128 , n372015 );
nand ( n51892 , n372127 , n372128 );
buf ( n372130 , n51892 );
buf ( n372131 , n372074 );
buf ( n372132 , n372080 );
nand ( n372133 , n372131 , n372132 );
buf ( n372134 , n372133 );
nand ( n372135 , n372130 , n372134 );
not ( n51899 , n372135 );
not ( n51900 , n51899 );
not ( n51901 , n372043 );
nand ( n372139 , n51901 , n372049 );
not ( n372140 , n372139 );
not ( n51904 , n372068 );
or ( n372142 , n372140 , n51904 );
buf ( n372143 , n51815 );
buf ( n372144 , n372043 );
nand ( n372145 , n372143 , n372144 );
buf ( n372146 , n372145 );
nand ( n372147 , n372142 , n372146 );
xor ( n51911 , n371548 , n371568 );
and ( n372149 , n51911 , n371594 );
and ( n51913 , n371548 , n371568 );
or ( n51914 , n372149 , n51913 );
buf ( n372152 , n51914 );
buf ( n372153 , n372152 );
not ( n51917 , n372153 );
buf ( n372155 , n44796 );
not ( n51919 , n372155 );
buf ( n372157 , n371605 );
not ( n372158 , n372157 );
or ( n51922 , n51919 , n372158 );
and ( n372160 , n40199 , n363444 );
not ( n51924 , n40199 );
and ( n51925 , n51924 , n22772 );
or ( n372163 , n372160 , n51925 );
buf ( n372164 , n372163 );
buf ( n372165 , n43261 );
nand ( n372166 , n372164 , n372165 );
buf ( n372167 , n372166 );
buf ( n372168 , n372167 );
nand ( n372169 , n51922 , n372168 );
buf ( n372170 , n372169 );
buf ( n372171 , n372170 );
xor ( n372172 , n371710 , n371739 );
and ( n51936 , n372172 , n371754 );
and ( n372174 , n371710 , n371739 );
or ( n372175 , n51936 , n372174 );
buf ( n372176 , n372175 );
buf ( n372177 , n372176 );
xor ( n372178 , n372171 , n372177 );
not ( n372179 , n45345 );
not ( n51943 , n51512 );
or ( n372181 , n372179 , n51943 );
buf ( n372182 , n367576 );
not ( n51946 , n372182 );
buf ( n372184 , n365945 );
not ( n51948 , n372184 );
or ( n51949 , n51946 , n51948 );
buf ( n372187 , n365507 );
buf ( n372188 , n44661 );
nand ( n51952 , n372187 , n372188 );
buf ( n51953 , n51952 );
buf ( n51954 , n51953 );
nand ( n51955 , n51949 , n51954 );
buf ( n51956 , n51955 );
buf ( n372194 , n51956 );
buf ( n372195 , n365954 );
nand ( n372196 , n372194 , n372195 );
buf ( n372197 , n372196 );
nand ( n372198 , n372181 , n372197 );
xor ( n372199 , n371631 , n372198 );
not ( n51963 , n46582 );
not ( n372201 , n30912 );
not ( n372202 , n372201 );
not ( n51966 , n366356 );
not ( n372204 , n51966 );
or ( n372205 , n372202 , n372204 );
or ( n51969 , n45152 , n365367 );
nand ( n372207 , n372205 , n51969 );
not ( n372208 , n372207 );
or ( n51972 , n51963 , n372208 );
or ( n372210 , n371673 , n39207 );
nand ( n372211 , n51972 , n372210 );
xor ( n51975 , n372199 , n372211 );
buf ( n372213 , n51975 );
xor ( n372214 , n372178 , n372213 );
buf ( n372215 , n372214 );
buf ( n372216 , n372215 );
not ( n51980 , n372216 );
or ( n372218 , n51917 , n51980 );
buf ( n372219 , n372215 );
buf ( n372220 , n372152 );
or ( n51984 , n372219 , n372220 );
xor ( n51985 , n371635 , n371660 );
and ( n51986 , n51985 , n371682 );
and ( n372224 , n371635 , n371660 );
or ( n51988 , n51986 , n372224 );
buf ( n372226 , n51988 );
buf ( n372227 , n372226 );
buf ( n372228 , n40923 );
not ( n51992 , n372228 );
not ( n372230 , n45116 );
buf ( n372231 , n372230 );
not ( n51995 , n372231 );
not ( n51996 , n361716 );
buf ( n372234 , n51996 );
not ( n51998 , n372234 );
or ( n51999 , n51995 , n51998 );
buf ( n372237 , n361716 );
buf ( n372238 , n367600 );
nand ( n52002 , n372237 , n372238 );
buf ( n372240 , n52002 );
buf ( n372241 , n372240 );
nand ( n372242 , n51999 , n372241 );
buf ( n372243 , n372242 );
buf ( n372244 , n372243 );
not ( n52008 , n372244 );
or ( n372246 , n51992 , n52008 );
not ( n372247 , n40878 );
buf ( n372248 , n372247 );
buf ( n372249 , n371624 );
nand ( n372250 , n372248 , n372249 );
buf ( n372251 , n372250 );
buf ( n372252 , n372251 );
nand ( n372253 , n372246 , n372252 );
buf ( n372254 , n372253 );
buf ( n372255 , n372254 );
buf ( n372256 , n371728 );
not ( n372257 , n372256 );
buf ( n372258 , n40475 );
not ( n52022 , n372258 );
or ( n372260 , n372257 , n52022 );
buf ( n372261 , n42355 );
not ( n52025 , n372261 );
buf ( n372263 , n45270 );
not ( n52027 , n372263 );
or ( n52028 , n52025 , n52027 );
not ( n52029 , n366078 );
buf ( n372267 , n52029 );
buf ( n372268 , n365471 );
nand ( n52032 , n372267 , n372268 );
buf ( n372270 , n52032 );
buf ( n372271 , n372270 );
nand ( n52035 , n52028 , n372271 );
buf ( n372273 , n52035 );
buf ( n52037 , n372273 );
buf ( n372275 , n360574 );
nand ( n372276 , n52037 , n372275 );
buf ( n372277 , n372276 );
buf ( n372278 , n372277 );
nand ( n52042 , n372260 , n372278 );
buf ( n372280 , n52042 );
buf ( n372281 , n372280 );
xor ( n52045 , n372255 , n372281 );
buf ( n372283 , n371653 );
not ( n52047 , n372283 );
buf ( n372285 , n359809 );
not ( n372286 , n372285 );
or ( n372287 , n52047 , n372286 );
buf ( n372288 , n362521 );
buf ( n372289 , n45300 );
not ( n372290 , n372289 );
buf ( n372291 , n361631 );
not ( n372292 , n372291 );
or ( n372293 , n372290 , n372292 );
buf ( n372294 , n366534 );
buf ( n372295 , n365464 );
nand ( n372296 , n372294 , n372295 );
buf ( n372297 , n372296 );
buf ( n372298 , n372297 );
nand ( n372299 , n372293 , n372298 );
buf ( n372300 , n372299 );
buf ( n372301 , n372300 );
nand ( n52065 , n372288 , n372301 );
buf ( n372303 , n52065 );
buf ( n372304 , n372303 );
nand ( n52068 , n372287 , n372304 );
buf ( n372306 , n52068 );
buf ( n372307 , n372306 );
xor ( n52071 , n52045 , n372307 );
buf ( n372309 , n52071 );
buf ( n372310 , n372309 );
xor ( n52074 , n372227 , n372310 );
buf ( n372312 , n42242 );
not ( n52076 , n372312 );
buf ( n372314 , n362426 );
not ( n372315 , n372314 );
buf ( n372316 , n47724 );
not ( n372317 , n372316 );
or ( n52081 , n372315 , n372317 );
buf ( n372319 , n40251 );
buf ( n372320 , n362435 );
nand ( n52084 , n372319 , n372320 );
buf ( n372322 , n52084 );
buf ( n372323 , n372322 );
nand ( n52087 , n52081 , n372323 );
buf ( n372325 , n52087 );
buf ( n372326 , n372325 );
not ( n52090 , n372326 );
or ( n52091 , n52076 , n52090 );
buf ( n372329 , n371461 );
buf ( n372330 , n363210 );
nand ( n52094 , n372329 , n372330 );
buf ( n372332 , n52094 );
buf ( n372333 , n372332 );
nand ( n52097 , n52091 , n372333 );
buf ( n372335 , n52097 );
buf ( n372336 , n372335 );
xor ( n52100 , n52074 , n372336 );
buf ( n372338 , n52100 );
buf ( n372339 , n372338 );
nand ( n372340 , n51984 , n372339 );
buf ( n372341 , n372340 );
buf ( n372342 , n372341 );
nand ( n372343 , n372218 , n372342 );
buf ( n372344 , n372343 );
xor ( n372345 , n372147 , n372344 );
buf ( n372346 , n362066 );
not ( n372347 , n372346 );
buf ( n372348 , n41892 );
not ( n372349 , n372348 );
buf ( n372350 , n41615 );
not ( n52108 , n372350 );
or ( n372352 , n372349 , n52108 );
buf ( n52110 , n41607 );
buf ( n372354 , n44634 );
nand ( n52112 , n52110 , n372354 );
buf ( n372356 , n52112 );
buf ( n372357 , n372356 );
nand ( n52115 , n372352 , n372357 );
buf ( n372359 , n52115 );
buf ( n372360 , n372359 );
not ( n52118 , n372360 );
or ( n52119 , n372347 , n52118 );
buf ( n372363 , n362030 );
buf ( n372364 , n371702 );
buf ( n52122 , n372364 );
nand ( n52123 , n372363 , n52122 );
buf ( n52124 , n52123 );
buf ( n52125 , n52124 );
nand ( n52126 , n52119 , n52125 );
buf ( n52127 , n52126 );
buf ( n372371 , n52127 );
buf ( n372372 , n371841 );
not ( n372373 , n372372 );
buf ( n372374 , n372373 );
buf ( n372375 , n372374 );
not ( n372376 , n372375 );
buf ( n372377 , n359916 );
not ( n52135 , n372377 );
or ( n372379 , n372376 , n52135 );
buf ( n372380 , n44743 );
not ( n52138 , n372380 );
not ( n372382 , n45113 );
buf ( n52140 , n372382 );
not ( n52141 , n52140 );
and ( n52142 , n52138 , n52141 );
buf ( n372386 , n44743 );
buf ( n372387 , n372382 );
and ( n52145 , n372386 , n372387 );
nor ( n372389 , n52142 , n52145 );
buf ( n372390 , n372389 );
buf ( n372391 , n372390 );
not ( n372392 , n372391 );
buf ( n372393 , n367440 );
nand ( n372394 , n372392 , n372393 );
buf ( n372395 , n372394 );
buf ( n372396 , n372395 );
nand ( n52154 , n372379 , n372396 );
buf ( n372398 , n52154 );
buf ( n372399 , n372398 );
xor ( n52157 , n372371 , n372399 );
buf ( n372401 , n41485 );
not ( n372402 , n372401 );
buf ( n372403 , n361531 );
not ( n372404 , n372403 );
buf ( n372405 , n362145 );
not ( n52163 , n372405 );
or ( n372407 , n372404 , n52163 );
buf ( n372408 , n45718 );
not ( n52166 , n372408 );
buf ( n372410 , n361534 );
nand ( n372411 , n52166 , n372410 );
buf ( n372412 , n372411 );
buf ( n372413 , n372412 );
nand ( n372414 , n372407 , n372413 );
buf ( n372415 , n372414 );
buf ( n372416 , n372415 );
not ( n372417 , n372416 );
or ( n372418 , n372402 , n372417 );
buf ( n372419 , n371865 );
buf ( n372420 , n361606 );
nand ( n372421 , n372419 , n372420 );
buf ( n372422 , n372421 );
buf ( n372423 , n372422 );
nand ( n372424 , n372418 , n372423 );
buf ( n372425 , n372424 );
buf ( n372426 , n372425 );
and ( n52184 , n52157 , n372426 );
and ( n372428 , n372371 , n372399 );
or ( n52186 , n52184 , n372428 );
buf ( n372430 , n52186 );
buf ( n372431 , n372430 );
xor ( n52189 , n372171 , n372177 );
and ( n372433 , n52189 , n372213 );
and ( n372434 , n372171 , n372177 );
or ( n52192 , n372433 , n372434 );
buf ( n372436 , n52192 );
buf ( n372437 , n372436 );
xor ( n52195 , n372431 , n372437 );
xor ( n372439 , n372227 , n372310 );
and ( n372440 , n372439 , n372336 );
and ( n52198 , n372227 , n372310 );
or ( n52199 , n372440 , n52198 );
buf ( n372443 , n52199 );
buf ( n372444 , n372443 );
xor ( n52202 , n52195 , n372444 );
buf ( n372446 , n52202 );
xor ( n372447 , n372345 , n372446 );
not ( n52205 , n372447 );
or ( n52206 , n51900 , n52205 );
not ( n52207 , n372447 );
nand ( n372451 , n52207 , n372135 );
nand ( n372452 , n52206 , n372451 );
buf ( n372453 , n51210 );
buf ( n372454 , n46521 );
and ( n52212 , n372453 , n372454 );
buf ( n372456 , n46477 );
not ( n52214 , n372456 );
not ( n372458 , n359974 );
buf ( n372459 , n372458 );
not ( n372460 , n372459 );
or ( n52218 , n52214 , n372460 );
buf ( n372462 , n363171 );
buf ( n372463 , n366683 );
nand ( n52221 , n372462 , n372463 );
buf ( n372465 , n52221 );
buf ( n372466 , n372465 );
nand ( n372467 , n52218 , n372466 );
buf ( n372468 , n372467 );
buf ( n372469 , n372468 );
not ( n372470 , n372469 );
buf ( n372471 , n366654 );
not ( n372472 , n372471 );
buf ( n372473 , n372472 );
buf ( n372474 , n372473 );
nor ( n372475 , n372470 , n372474 );
buf ( n372476 , n372475 );
buf ( n372477 , n372476 );
nor ( n372478 , n52212 , n372477 );
buf ( n372479 , n372478 );
buf ( n372480 , n372479 );
not ( n52238 , n372480 );
and ( n52239 , n47554 , n360886 );
not ( n52240 , n47554 );
and ( n52241 , n52240 , n360893 );
or ( n372485 , n52239 , n52241 );
and ( n52243 , n372485 , n41835 );
and ( n372487 , n371501 , n367759 );
nor ( n52245 , n52243 , n372487 );
buf ( n372489 , n52245 );
not ( n372490 , n372489 );
buf ( n372491 , n366615 );
not ( n52249 , n372491 );
buf ( n372493 , n365036 );
not ( n372494 , n372493 );
or ( n52252 , n52249 , n372494 );
buf ( n372496 , n371820 );
nand ( n372497 , n52252 , n372496 );
buf ( n372498 , n372497 );
buf ( n52256 , n372498 );
not ( n52257 , n52256 );
or ( n52258 , n372490 , n52257 );
buf ( n372502 , n366615 );
not ( n372503 , n372502 );
buf ( n372504 , n365036 );
not ( n372505 , n372504 );
or ( n372506 , n372503 , n372505 );
buf ( n372507 , n371820 );
nand ( n372508 , n372506 , n372507 );
buf ( n372509 , n372508 );
buf ( n372510 , n372509 );
buf ( n372511 , n52245 );
or ( n372512 , n372510 , n372511 );
nand ( n52270 , n52258 , n372512 );
buf ( n372514 , n52270 );
buf ( n372515 , n372514 );
not ( n52273 , n372515 );
or ( n52274 , n52238 , n52273 );
buf ( n372518 , n372479 );
buf ( n372519 , n372514 );
or ( n52277 , n372518 , n372519 );
nand ( n372521 , n52274 , n52277 );
buf ( n372522 , n372521 );
buf ( n372523 , n372522 );
xor ( n372524 , n371828 , n371895 );
and ( n52282 , n372524 , n371907 );
and ( n52283 , n371828 , n371895 );
or ( n52284 , n52282 , n52283 );
buf ( n372528 , n52284 );
buf ( n372529 , n372528 );
xor ( n52287 , n372523 , n372529 );
xor ( n52288 , n371853 , n371871 );
and ( n372532 , n52288 , n371892 );
and ( n52290 , n371853 , n371871 );
or ( n372534 , n372532 , n52290 );
buf ( n372535 , n372534 );
buf ( n372536 , n372535 );
buf ( n372537 , n45492 );
not ( n372538 , n372537 );
buf ( n372539 , n365676 );
not ( n372540 , n372539 );
buf ( n372541 , n362179 );
not ( n52299 , n372541 );
or ( n372543 , n372540 , n52299 );
buf ( n372544 , n40899 );
buf ( n372545 , n365673 );
nand ( n52303 , n372544 , n372545 );
buf ( n372547 , n52303 );
buf ( n372548 , n372547 );
nand ( n52306 , n372543 , n372548 );
buf ( n372550 , n52306 );
buf ( n52308 , n372550 );
not ( n52309 , n52308 );
or ( n52310 , n372538 , n52309 );
buf ( n52311 , n371537 );
buf ( n372555 , n45553 );
nand ( n372556 , n52311 , n372555 );
buf ( n372557 , n372556 );
buf ( n372558 , n372557 );
nand ( n372559 , n52310 , n372558 );
buf ( n372560 , n372559 );
buf ( n372561 , n372560 );
xor ( n372562 , n372536 , n372561 );
xor ( n52320 , n372371 , n372399 );
xor ( n52321 , n52320 , n372426 );
buf ( n372565 , n52321 );
buf ( n372566 , n372565 );
xor ( n52324 , n372562 , n372566 );
buf ( n372568 , n52324 );
buf ( n372569 , n372568 );
xor ( n52327 , n52287 , n372569 );
buf ( n372571 , n52327 );
buf ( n372572 , n371801 );
buf ( n372573 , n371783 );
or ( n52331 , n372572 , n372573 );
buf ( n372575 , n371909 );
nand ( n372576 , n52331 , n372575 );
buf ( n372577 , n372576 );
buf ( n372578 , n372577 );
buf ( n372579 , n371801 );
buf ( n372580 , n371783 );
nand ( n372581 , n372579 , n372580 );
buf ( n372582 , n372581 );
buf ( n372583 , n372582 );
nand ( n372584 , n372578 , n372583 );
buf ( n372585 , n372584 );
or ( n372586 , n372571 , n372585 );
buf ( n52344 , n372152 );
xor ( n372588 , n372338 , n52344 );
buf ( n372589 , n372215 );
buf ( n372590 , n372589 );
buf ( n372591 , n372590 );
xor ( n52349 , n372588 , n372591 );
nand ( n372593 , n372586 , n52349 );
nand ( n372594 , n372571 , n372585 );
nand ( n52352 , n372593 , n372594 );
buf ( n52353 , n52352 );
not ( n372597 , n52353 );
buf ( n372598 , n372597 );
and ( n372599 , n372452 , n372598 );
not ( n372600 , n372452 );
and ( n52358 , n372600 , n52352 );
nor ( n372602 , n372599 , n52358 );
buf ( n372603 , n362030 );
not ( n52361 , n372603 );
buf ( n372605 , n372359 );
not ( n52363 , n372605 );
or ( n52364 , n52361 , n52363 );
buf ( n52365 , n41892 );
not ( n52366 , n52365 );
buf ( n52367 , n363317 );
not ( n52368 , n52367 );
or ( n52369 , n52366 , n52368 );
buf ( n372613 , n41663 );
buf ( n372614 , n365626 );
nand ( n372615 , n372613 , n372614 );
buf ( n372616 , n372615 );
buf ( n372617 , n372616 );
nand ( n372618 , n52369 , n372617 );
buf ( n372619 , n372618 );
buf ( n372620 , n372619 );
buf ( n372621 , n362066 );
nand ( n372622 , n372620 , n372621 );
buf ( n372623 , n372622 );
buf ( n372624 , n372623 );
nand ( n372625 , n52364 , n372624 );
buf ( n372626 , n372625 );
buf ( n372627 , n372626 );
buf ( n372628 , n41835 );
not ( n52386 , n372628 );
buf ( n372630 , n44570 );
not ( n372631 , n372630 );
buf ( n372632 , n362461 );
not ( n52390 , n372632 );
or ( n372634 , n372631 , n52390 );
buf ( n372635 , n46491 );
buf ( n372636 , n41772 );
nand ( n372637 , n372635 , n372636 );
buf ( n372638 , n372637 );
buf ( n372639 , n372638 );
nand ( n372640 , n372634 , n372639 );
buf ( n372641 , n372640 );
buf ( n372642 , n372641 );
not ( n52400 , n372642 );
or ( n52401 , n52386 , n52400 );
buf ( n372645 , n47554 );
not ( n52403 , n372645 );
buf ( n372647 , n360886 );
not ( n52405 , n372647 );
or ( n52406 , n52403 , n52405 );
buf ( n372650 , n360893 );
buf ( n372651 , n41772 );
nand ( n52409 , n372650 , n372651 );
buf ( n372653 , n52409 );
buf ( n372654 , n372653 );
nand ( n52412 , n52406 , n372654 );
buf ( n372656 , n52412 );
buf ( n372657 , n372656 );
buf ( n372658 , n367759 );
nand ( n372659 , n372657 , n372658 );
buf ( n372660 , n372659 );
buf ( n372661 , n372660 );
nand ( n52419 , n52401 , n372661 );
buf ( n372663 , n52419 );
buf ( n372664 , n372663 );
xor ( n52422 , n372627 , n372664 );
xor ( n52423 , n372255 , n372281 );
and ( n52424 , n52423 , n372307 );
and ( n52425 , n372255 , n372281 );
or ( n52426 , n52424 , n52425 );
buf ( n372670 , n52426 );
buf ( n372671 , n372670 );
xor ( n372672 , n52422 , n372671 );
buf ( n372673 , n372672 );
buf ( n372674 , n372673 );
xor ( n372675 , n371631 , n372198 );
and ( n52433 , n372675 , n372211 );
and ( n372677 , n371631 , n372198 );
or ( n372678 , n52433 , n372677 );
buf ( n372679 , n372678 );
buf ( n52437 , n41485 );
not ( n52438 , n52437 );
and ( n372682 , n363603 , n366407 );
not ( n52440 , n363603 );
and ( n52441 , n52440 , n42149 );
or ( n372685 , n372682 , n52441 );
buf ( n372686 , n372685 );
not ( n372687 , n372686 );
or ( n372688 , n52438 , n372687 );
buf ( n372689 , n372415 );
buf ( n372690 , n361606 );
nand ( n372691 , n372689 , n372690 );
buf ( n372692 , n372691 );
buf ( n372693 , n372692 );
nand ( n372694 , n372688 , n372693 );
buf ( n372695 , n372694 );
buf ( n372696 , n372695 );
xor ( n52454 , n372679 , n372696 );
buf ( n372698 , n363210 );
not ( n52456 , n372698 );
buf ( n372700 , n372325 );
not ( n52458 , n372700 );
or ( n372702 , n52456 , n52458 );
not ( n372703 , n362426 );
not ( n52461 , n363391 );
or ( n372705 , n372703 , n52461 );
nand ( n372706 , n40275 , n362435 );
nand ( n52464 , n372705 , n372706 );
buf ( n372708 , n52464 );
buf ( n52466 , n42242 );
nand ( n52467 , n372708 , n52466 );
buf ( n372711 , n52467 );
buf ( n372712 , n372711 );
nand ( n372713 , n372702 , n372712 );
buf ( n372714 , n372713 );
buf ( n372715 , n372714 );
xor ( n52473 , n52454 , n372715 );
buf ( n372717 , n52473 );
buf ( n372718 , n372717 );
xor ( n52476 , n372674 , n372718 );
buf ( n372720 , n372509 );
not ( n372721 , n372720 );
buf ( n372722 , n52245 );
nand ( n372723 , n372721 , n372722 );
buf ( n372724 , n372723 );
buf ( n372725 , n372724 );
not ( n372726 , n372725 );
buf ( n372727 , n372479 );
not ( n372728 , n372727 );
buf ( n372729 , n372728 );
buf ( n372730 , n372729 );
not ( n52488 , n372730 );
or ( n372732 , n372726 , n52488 );
buf ( n372733 , n52245 );
not ( n372734 , n372733 );
buf ( n372735 , n372509 );
nand ( n372736 , n372734 , n372735 );
buf ( n372737 , n372736 );
buf ( n372738 , n372737 );
nand ( n52496 , n372732 , n372738 );
buf ( n372740 , n52496 );
buf ( n372741 , n372740 );
xnor ( n372742 , n52476 , n372741 );
buf ( n372743 , n372742 );
buf ( n372744 , n372743 );
xor ( n52502 , n372523 , n372529 );
and ( n372746 , n52502 , n372569 );
and ( n52504 , n372523 , n372529 );
or ( n372748 , n372746 , n52504 );
buf ( n372749 , n372748 );
buf ( n372750 , n372749 );
xor ( n372751 , n372744 , n372750 );
buf ( n372752 , n43261 );
not ( n52510 , n372752 );
buf ( n372754 , n22772 );
not ( n372755 , n372754 );
buf ( n372756 , n364987 );
not ( n372757 , n372756 );
or ( n372758 , n372755 , n372757 );
buf ( n372759 , n359778 );
buf ( n372760 , n363444 );
nand ( n372761 , n372759 , n372760 );
buf ( n372762 , n372761 );
buf ( n372763 , n372762 );
nand ( n372764 , n372758 , n372763 );
buf ( n372765 , n372764 );
buf ( n52523 , n372765 );
not ( n52524 , n52523 );
or ( n52525 , n52510 , n52524 );
buf ( n52526 , n363429 );
buf ( n52527 , n372163 );
nand ( n52528 , n52526 , n52527 );
buf ( n52529 , n52528 );
buf ( n52530 , n52529 );
nand ( n52531 , n52525 , n52530 );
buf ( n52532 , n52531 );
buf ( n52533 , n366654 );
not ( n52534 , n52533 );
buf ( n372778 , n46477 );
not ( n52536 , n372778 );
buf ( n372780 , n363866 );
not ( n372781 , n372780 );
or ( n52539 , n52536 , n372781 );
buf ( n372783 , n365170 );
buf ( n372784 , n366683 );
nand ( n372785 , n372783 , n372784 );
buf ( n372786 , n372785 );
buf ( n372787 , n372786 );
nand ( n372788 , n52539 , n372787 );
buf ( n372789 , n372788 );
buf ( n372790 , n372789 );
not ( n52548 , n372790 );
or ( n372792 , n52534 , n52548 );
buf ( n372793 , n372468 );
buf ( n372794 , n46521 );
nand ( n372795 , n372793 , n372794 );
buf ( n372796 , n372795 );
buf ( n372797 , n372796 );
nand ( n52555 , n372792 , n372797 );
buf ( n372799 , n52555 );
xor ( n52557 , n52532 , n372799 );
buf ( n372801 , n51956 );
not ( n372802 , n372801 );
buf ( n372803 , n40059 );
not ( n372804 , n372803 );
or ( n52562 , n372802 , n372804 );
buf ( n372806 , n371669 );
not ( n372807 , n372806 );
buf ( n372808 , n363122 );
not ( n52566 , n372808 );
or ( n372810 , n372807 , n52566 );
buf ( n372811 , n363119 );
buf ( n372812 , n364870 );
nand ( n372813 , n372811 , n372812 );
buf ( n372814 , n372813 );
buf ( n372815 , n372814 );
nand ( n372816 , n372810 , n372815 );
buf ( n372817 , n372816 );
buf ( n372818 , n372817 );
buf ( n372819 , n39949 );
nand ( n52577 , n372818 , n372819 );
buf ( n372821 , n52577 );
buf ( n372822 , n372821 );
nand ( n52580 , n52562 , n372822 );
buf ( n372824 , n52580 );
buf ( n372825 , n372273 );
not ( n52583 , n372825 );
buf ( n372827 , n40475 );
not ( n372828 , n372827 );
or ( n52586 , n52583 , n372828 );
buf ( n372830 , n362540 );
not ( n372831 , n372830 );
buf ( n372832 , n366277 );
not ( n372833 , n372832 );
or ( n52591 , n372831 , n372833 );
buf ( n372835 , n362452 );
buf ( n372836 , n362552 );
nand ( n52594 , n372835 , n372836 );
buf ( n372838 , n52594 );
buf ( n372839 , n372838 );
nand ( n52597 , n52591 , n372839 );
buf ( n52598 , n52597 );
buf ( n372842 , n52598 );
buf ( n372843 , n360577 );
nand ( n372844 , n372842 , n372843 );
buf ( n372845 , n372844 );
buf ( n372846 , n372845 );
nand ( n372847 , n52586 , n372846 );
buf ( n372848 , n372847 );
xor ( n52606 , n372824 , n372848 );
buf ( n372850 , n52606 );
buf ( n372851 , n372300 );
not ( n372852 , n372851 );
buf ( n372853 , n359809 );
not ( n372854 , n372853 );
or ( n372855 , n372852 , n372854 );
buf ( n372856 , n39592 );
and ( n52614 , n352212 , n361631 );
not ( n372858 , n352212 );
and ( n52616 , n372858 , n39621 );
or ( n52617 , n52614 , n52616 );
buf ( n372861 , n52617 );
nand ( n372862 , n372856 , n372861 );
buf ( n372863 , n372862 );
buf ( n372864 , n372863 );
nand ( n372865 , n372855 , n372864 );
buf ( n372866 , n372865 );
buf ( n372867 , n372866 );
xor ( n372868 , n372850 , n372867 );
buf ( n372869 , n372868 );
xnor ( n52627 , n52557 , n372869 );
buf ( n372871 , n52627 );
not ( n52629 , n372871 );
buf ( n372873 , n52629 );
not ( n52631 , n372873 );
buf ( n372875 , n365279 );
not ( n52633 , n372875 );
buf ( n372877 , n372243 );
not ( n52635 , n372877 );
or ( n372879 , n52633 , n52635 );
buf ( n372880 , n365293 );
not ( n52638 , n372880 );
buf ( n372882 , n52638 );
buf ( n372883 , n372882 );
buf ( n372884 , n365760 );
and ( n372885 , n372883 , n372884 );
not ( n52643 , n372883 );
buf ( n372887 , n361664 );
not ( n52645 , n372887 );
buf ( n372889 , n52645 );
buf ( n52647 , n372889 );
and ( n372891 , n52643 , n52647 );
nor ( n52649 , n372885 , n372891 );
buf ( n52650 , n52649 );
buf ( n372894 , n52650 );
buf ( n372895 , n365303 );
nand ( n372896 , n372894 , n372895 );
buf ( n372897 , n372896 );
buf ( n372898 , n372897 );
nand ( n52656 , n372879 , n372898 );
buf ( n52657 , n52656 );
not ( n372901 , n366989 );
not ( n52659 , n372207 );
or ( n372903 , n372901 , n52659 );
buf ( n372904 , n42911 );
not ( n52662 , n372904 );
buf ( n372906 , n365368 );
not ( n52664 , n372906 );
or ( n372908 , n52662 , n52664 );
buf ( n372909 , n51966 );
buf ( n372910 , n49988 );
nand ( n372911 , n372909 , n372910 );
buf ( n372912 , n372911 );
buf ( n372913 , n372912 );
nand ( n372914 , n372908 , n372913 );
buf ( n372915 , n372914 );
nand ( n372916 , n372915 , n46582 );
nand ( n52674 , n372903 , n372916 );
not ( n52675 , n52674 );
xor ( n52676 , n52657 , n52675 );
buf ( n372920 , n369945 );
buf ( n372921 , n372390 );
or ( n372922 , n372920 , n372921 );
buf ( n372923 , n359996 );
buf ( n372924 , n31286 );
buf ( n372925 , n361762 );
and ( n372926 , n372924 , n372925 );
not ( n52684 , n372924 );
buf ( n372928 , n359947 );
and ( n372929 , n52684 , n372928 );
nor ( n372930 , n372926 , n372929 );
buf ( n372931 , n372930 );
buf ( n372932 , n372931 );
or ( n52690 , n372923 , n372932 );
nand ( n52691 , n372922 , n52690 );
buf ( n372935 , n52691 );
xor ( n372936 , n52676 , n372935 );
buf ( n372937 , n372936 );
buf ( n372938 , n45553 );
not ( n372939 , n372938 );
buf ( n372940 , n372550 );
not ( n372941 , n372940 );
or ( n372942 , n372939 , n372941 );
nand ( n52700 , n365676 , n359147 );
not ( n372944 , n52700 );
buf ( n372945 , n363442 );
buf ( n372946 , n365673 );
nand ( n372947 , n372945 , n372946 );
buf ( n372948 , n372947 );
not ( n52706 , n372948 );
or ( n372950 , n372944 , n52706 );
nand ( n372951 , n372950 , n45492 );
buf ( n372952 , n372951 );
nand ( n372953 , n372942 , n372952 );
buf ( n372954 , n372953 );
buf ( n372955 , n372954 );
xor ( n372956 , n372937 , n372955 );
buf ( n372957 , n366402 );
not ( n372958 , n372957 );
buf ( n372959 , n372033 );
not ( n52717 , n372959 );
or ( n372961 , n372958 , n52717 );
and ( n52719 , n22710 , n359939 );
not ( n372963 , n22710 );
and ( n52721 , n372963 , n40943 );
or ( n52722 , n52719 , n52721 );
buf ( n52723 , n52722 );
buf ( n372967 , n366434 );
nand ( n52725 , n52723 , n372967 );
buf ( n372969 , n52725 );
buf ( n372970 , n372969 );
nand ( n372971 , n372961 , n372970 );
buf ( n372972 , n372971 );
buf ( n372973 , n372972 );
xor ( n372974 , n372956 , n372973 );
buf ( n372975 , n372974 );
buf ( n372976 , n372975 );
not ( n52734 , n372976 );
buf ( n52735 , n52734 );
not ( n372979 , n52735 );
or ( n52737 , n52631 , n372979 );
buf ( n372981 , n372975 );
buf ( n372982 , n52627 );
nand ( n52740 , n372981 , n372982 );
buf ( n52741 , n52740 );
nand ( n372985 , n52737 , n52741 );
xor ( n372986 , n372536 , n372561 );
and ( n372987 , n372986 , n372566 );
and ( n52745 , n372536 , n372561 );
or ( n372989 , n372987 , n52745 );
buf ( n372990 , n372989 );
xnor ( n52748 , n372985 , n372990 );
buf ( n372992 , n52748 );
xor ( n372993 , n372751 , n372992 );
buf ( n372994 , n372993 );
and ( n372995 , n372602 , n372994 );
not ( n52753 , n372602 );
not ( n52754 , n372994 );
and ( n372998 , n52753 , n52754 );
nor ( n372999 , n372995 , n372998 );
buf ( n373000 , n372999 );
not ( n373001 , n373000 );
or ( n373002 , n372122 , n373001 );
buf ( n373003 , n372999 );
buf ( n373004 , n372120 );
or ( n373005 , n373003 , n373004 );
nand ( n52763 , n373002 , n373005 );
buf ( n373007 , n52763 );
buf ( n373008 , n373007 );
not ( n52766 , n373008 );
xor ( n373010 , n52349 , n372585 );
buf ( n373011 , n373010 );
buf ( n373012 , n372571 );
buf ( n373013 , n373012 );
buf ( n373014 , n373013 );
buf ( n373015 , n373014 );
and ( n373016 , n373011 , n373015 );
not ( n52774 , n373011 );
buf ( n373018 , n373014 );
not ( n52776 , n373018 );
buf ( n373020 , n52776 );
buf ( n52778 , n373020 );
and ( n52779 , n52774 , n52778 );
nor ( n373023 , n373016 , n52779 );
buf ( n373024 , n373023 );
buf ( n373025 , n373024 );
not ( n373026 , n373025 );
not ( n52784 , n371960 );
not ( n52785 , n371768 );
or ( n373029 , n52784 , n52785 );
not ( n373030 , n371767 );
not ( n52788 , n371957 );
or ( n373032 , n373030 , n52788 );
nand ( n373033 , n373032 , n371773 );
nand ( n52791 , n373029 , n373033 );
not ( n373035 , n52791 );
buf ( n373036 , n373035 );
nand ( n52794 , n373026 , n373036 );
buf ( n52795 , n52794 );
buf ( n373039 , n52795 );
xor ( n373040 , n51857 , n372108 );
xor ( n373041 , n373040 , n51880 );
buf ( n373042 , n373041 );
buf ( n373043 , n373042 );
buf ( n373044 , n373043 );
buf ( n373045 , n373044 );
and ( n52798 , n373039 , n373045 );
buf ( n373047 , n52791 );
buf ( n373048 , n373024 );
and ( n52801 , n373047 , n373048 );
buf ( n373050 , n52801 );
buf ( n373051 , n373050 );
nor ( n373052 , n52798 , n373051 );
buf ( n373053 , n373052 );
buf ( n373054 , n373053 );
nand ( n52807 , n52766 , n373054 );
buf ( n373056 , n52807 );
buf ( n373057 , n373056 );
not ( n52810 , n373024 );
and ( n52811 , n373041 , n52810 );
not ( n373060 , n373041 );
and ( n52813 , n373060 , n373024 );
nor ( n373062 , n52811 , n52813 );
and ( n373063 , n373062 , n52791 );
not ( n52816 , n373062 );
and ( n373065 , n52816 , n373035 );
nor ( n52818 , n373063 , n373065 );
buf ( n52819 , n52818 );
not ( n373068 , n51728 );
buf ( n373069 , n371383 );
not ( n373070 , n373069 );
buf ( n373071 , n373070 );
not ( n373072 , n373071 );
and ( n52825 , n373068 , n373072 );
buf ( n373074 , n51728 );
buf ( n373075 , n373071 );
nand ( n52828 , n373074 , n373075 );
buf ( n373077 , n52828 );
buf ( n52830 , n371388 );
and ( n373079 , n373077 , n52830 );
nor ( n373080 , n52825 , n373079 );
buf ( n373081 , n373080 );
nand ( n373082 , n52819 , n373081 );
buf ( n373083 , n373082 );
buf ( n373084 , n373083 );
buf ( n373085 , n372673 );
not ( n52838 , n373085 );
buf ( n373087 , n372717 );
not ( n373088 , n373087 );
or ( n52841 , n52838 , n373088 );
or ( n52842 , n372717 , n372673 );
nand ( n373091 , n52842 , n372740 );
buf ( n373092 , n373091 );
nand ( n373093 , n52841 , n373092 );
buf ( n373094 , n373093 );
not ( n373095 , n372873 );
not ( n373096 , n372975 );
or ( n52849 , n373095 , n373096 );
buf ( n373098 , n52735 );
not ( n52851 , n373098 );
buf ( n373100 , n52627 );
not ( n373101 , n373100 );
or ( n52854 , n52851 , n373101 );
buf ( n373103 , n372990 );
nand ( n52856 , n52854 , n373103 );
buf ( n373105 , n52856 );
nand ( n52858 , n52849 , n373105 );
not ( n52859 , n52858 );
xor ( n52860 , n373094 , n52859 );
xor ( n373109 , n52657 , n52675 );
and ( n373110 , n373109 , n372935 );
and ( n373111 , n52657 , n52675 );
or ( n52864 , n373110 , n373111 );
buf ( n373113 , n52864 );
not ( n373114 , n372948 );
not ( n52867 , n52700 );
or ( n52868 , n373114 , n52867 );
buf ( n373117 , n45553 );
not ( n52870 , n373117 );
buf ( n373119 , n371272 );
nand ( n373120 , n52870 , n373119 );
buf ( n373121 , n373120 );
nand ( n373122 , n52868 , n373121 );
buf ( n373123 , n373122 );
xor ( n373124 , n373113 , n373123 );
buf ( n52877 , n52598 );
not ( n52878 , n52877 );
buf ( n373127 , n46557 );
not ( n52880 , n373127 );
or ( n52881 , n52878 , n52880 );
not ( n373130 , n51996 );
nand ( n52883 , n373130 , n365468 );
nand ( n52884 , n361712 , n360610 );
nand ( n373133 , n52883 , n52884 );
nand ( n52886 , n360577 , n373133 );
buf ( n373135 , n52886 );
nand ( n52888 , n52881 , n373135 );
buf ( n373137 , n52888 );
buf ( n373138 , n372915 );
not ( n52891 , n373138 );
buf ( n373140 , n39208 );
not ( n373141 , n373140 );
or ( n52894 , n52891 , n373141 );
buf ( n373143 , n39217 );
buf ( n373144 , n51966 );
not ( n52897 , n373144 );
buf ( n373146 , n366077 );
not ( n52899 , n373146 );
or ( n373148 , n52897 , n52899 );
buf ( n52901 , n366078 );
buf ( n373150 , n359297 );
buf ( n373151 , n373150 );
nand ( n373152 , n52901 , n373151 );
buf ( n373153 , n373152 );
buf ( n373154 , n373153 );
nand ( n373155 , n373148 , n373154 );
buf ( n373156 , n373155 );
buf ( n373157 , n373156 );
nand ( n52910 , n373143 , n373157 );
buf ( n373159 , n52910 );
buf ( n373160 , n373159 );
nand ( n373161 , n52894 , n373160 );
buf ( n373162 , n373161 );
xor ( n373163 , n373137 , n373162 );
buf ( n373164 , n372817 );
not ( n52917 , n373164 );
buf ( n373166 , n40059 );
not ( n373167 , n373166 );
or ( n373168 , n52917 , n373167 );
buf ( n373169 , n30912 );
not ( n373170 , n373169 );
buf ( n373171 , n365945 );
not ( n52924 , n373171 );
or ( n373173 , n373170 , n52924 );
buf ( n373174 , n363107 );
buf ( n373175 , n42898 );
nand ( n52928 , n373174 , n373175 );
buf ( n373177 , n52928 );
buf ( n373178 , n373177 );
nand ( n373179 , n373173 , n373178 );
buf ( n373180 , n373179 );
buf ( n373181 , n373180 );
buf ( n373182 , n39949 );
nand ( n373183 , n373181 , n373182 );
buf ( n373184 , n373183 );
buf ( n373185 , n373184 );
nand ( n52938 , n373168 , n373185 );
buf ( n373187 , n52938 );
xor ( n52940 , n373163 , n373187 );
buf ( n373189 , n52940 );
xor ( n52942 , n373124 , n373189 );
buf ( n373191 , n52942 );
buf ( n52944 , n373191 );
xor ( n373193 , n372937 , n372955 );
and ( n52946 , n373193 , n372973 );
and ( n373195 , n372937 , n372955 );
or ( n373196 , n52946 , n373195 );
buf ( n373197 , n373196 );
buf ( n373198 , n373197 );
xor ( n373199 , n52944 , n373198 );
xor ( n52952 , n372431 , n372437 );
and ( n52953 , n52952 , n372444 );
and ( n373202 , n372431 , n372437 );
or ( n373203 , n52953 , n373202 );
buf ( n373204 , n373203 );
buf ( n373205 , n373204 );
xor ( n373206 , n373199 , n373205 );
buf ( n373207 , n373206 );
xor ( n373208 , n52860 , n373207 );
buf ( n373209 , n372135 );
not ( n52962 , n373209 );
not ( n373211 , n52207 );
buf ( n373212 , n373211 );
not ( n52965 , n373212 );
or ( n52966 , n52962 , n52965 );
not ( n373215 , n372594 );
not ( n52968 , n372593 );
or ( n52969 , n373215 , n52968 );
or ( n373218 , n372135 , n372447 );
nand ( n373219 , n52969 , n373218 );
buf ( n373220 , n373219 );
nand ( n373221 , n52966 , n373220 );
buf ( n373222 , n373221 );
xor ( n52975 , n373208 , n373222 );
buf ( n373224 , n372344 );
buf ( n52977 , n373224 );
buf ( n373226 , n52977 );
buf ( n373227 , n373226 );
buf ( n373228 , n372446 );
or ( n52981 , n373227 , n373228 );
buf ( n373230 , n372147 );
nand ( n373231 , n52981 , n373230 );
buf ( n373232 , n373231 );
buf ( n373233 , n373232 );
buf ( n52986 , n372446 );
buf ( n373235 , n373226 );
nand ( n373236 , n52986 , n373235 );
buf ( n373237 , n373236 );
buf ( n373238 , n373237 );
nand ( n52991 , n373233 , n373238 );
buf ( n373240 , n52991 );
buf ( n373241 , n366402 );
not ( n373242 , n373241 );
buf ( n373243 , n52722 );
not ( n52996 , n373243 );
or ( n373245 , n373242 , n52996 );
buf ( n373246 , n22710 );
not ( n52999 , n373246 );
buf ( n373248 , n363172 );
not ( n373249 , n373248 );
or ( n53002 , n52999 , n373249 );
buf ( n373251 , n42606 );
buf ( n373252 , n342657 );
nand ( n53005 , n373251 , n373252 );
buf ( n373254 , n53005 );
buf ( n373255 , n373254 );
nand ( n53008 , n53002 , n373255 );
buf ( n53009 , n53008 );
buf ( n373258 , n53009 );
buf ( n373259 , n366434 );
nand ( n373260 , n373258 , n373259 );
buf ( n373261 , n373260 );
buf ( n373262 , n373261 );
nand ( n53015 , n373245 , n373262 );
buf ( n373264 , n53015 );
buf ( n373265 , n43261 );
not ( n373266 , n373265 );
and ( n53019 , n44925 , n22772 );
not ( n373268 , n44925 );
and ( n373269 , n373268 , n363444 );
or ( n373270 , n53019 , n373269 );
buf ( n373271 , n373270 );
not ( n53024 , n373271 );
or ( n373273 , n373266 , n53024 );
buf ( n373274 , n372765 );
buf ( n373275 , n44796 );
nand ( n373276 , n373274 , n373275 );
buf ( n373277 , n373276 );
buf ( n373278 , n373277 );
nand ( n53031 , n373273 , n373278 );
buf ( n373280 , n53031 );
or ( n53033 , n373264 , n373280 );
buf ( n373282 , n373264 );
not ( n53035 , n373282 );
buf ( n373284 , n53035 );
not ( n53037 , n373280 );
or ( n373286 , n373284 , n53037 );
not ( n373287 , n366654 );
not ( n53040 , n46477 );
not ( n53041 , n41472 );
or ( n373290 , n53040 , n53041 );
nand ( n53043 , n40899 , n46474 );
nand ( n373292 , n373290 , n53043 );
not ( n373293 , n373292 );
or ( n53046 , n373287 , n373293 );
buf ( n373295 , n372789 );
buf ( n373296 , n46521 );
nand ( n53049 , n373295 , n373296 );
buf ( n373298 , n53049 );
nand ( n373299 , n53046 , n373298 );
nand ( n53052 , n53033 , n373286 , n373299 );
not ( n53053 , n373299 );
not ( n53054 , n373284 );
not ( n373303 , n53037 );
or ( n373304 , n53054 , n373303 );
nand ( n53057 , n373280 , n373264 );
nand ( n53058 , n373304 , n53057 );
nand ( n53059 , n53053 , n53058 );
nand ( n373308 , n53052 , n53059 );
buf ( n373309 , n52617 );
not ( n53062 , n373309 );
buf ( n373311 , n363038 );
not ( n53064 , n373311 );
or ( n373313 , n53062 , n53064 );
buf ( n373314 , n362521 );
buf ( n373315 , n352195 );
not ( n373316 , n373315 );
buf ( n373317 , n361631 );
not ( n53070 , n373317 );
or ( n373319 , n373316 , n53070 );
buf ( n53072 , n39621 );
buf ( n373321 , n352194 );
nand ( n373322 , n53072 , n373321 );
buf ( n373323 , n373322 );
buf ( n373324 , n373323 );
nand ( n373325 , n373319 , n373324 );
buf ( n373326 , n373325 );
buf ( n373327 , n373326 );
nand ( n373328 , n373314 , n373327 );
buf ( n373329 , n373328 );
buf ( n373330 , n373329 );
nand ( n373331 , n373313 , n373330 );
buf ( n373332 , n373331 );
buf ( n373333 , n373332 );
buf ( n373334 , n42171 );
not ( n53087 , n373334 );
buf ( n373336 , n41615 );
not ( n373337 , n373336 );
or ( n53090 , n53087 , n373337 );
buf ( n373339 , n41607 );
buf ( n373340 , n361026 );
nand ( n53093 , n373339 , n373340 );
buf ( n373342 , n53093 );
buf ( n373343 , n373342 );
nand ( n373344 , n53090 , n373343 );
buf ( n373345 , n373344 );
and ( n53098 , n373345 , n361060 );
and ( n373347 , n52650 , n361019 );
nor ( n53100 , n53098 , n373347 );
buf ( n373349 , n53100 );
not ( n53102 , n373349 );
buf ( n373351 , n53102 );
buf ( n373352 , n373351 );
xor ( n373353 , n373333 , n373352 );
buf ( n373354 , n369945 );
not ( n373355 , n373354 );
buf ( n373356 , n372931 );
not ( n53109 , n373356 );
and ( n53110 , n373355 , n53109 );
buf ( n373359 , n365801 );
xor ( n53112 , n44743 , n31073 );
buf ( n373361 , n53112 );
nor ( n53114 , n373359 , n373361 );
buf ( n373363 , n53114 );
buf ( n373364 , n373363 );
nor ( n53117 , n53110 , n373364 );
buf ( n373366 , n53117 );
buf ( n373367 , n373366 );
not ( n53120 , n373367 );
buf ( n373369 , n53120 );
buf ( n373370 , n373369 );
xor ( n53123 , n373353 , n373370 );
buf ( n373372 , n53123 );
buf ( n373373 , n373372 );
xor ( n373374 , n372627 , n372664 );
and ( n53127 , n373374 , n372671 );
and ( n53128 , n372627 , n372664 );
or ( n53129 , n53127 , n53128 );
buf ( n53130 , n53129 );
buf ( n373379 , n53130 );
xor ( n53132 , n373373 , n373379 );
buf ( n373381 , n41892 );
not ( n373382 , n373381 );
buf ( n373383 , n367116 );
not ( n53136 , n373383 );
or ( n373385 , n373382 , n53136 );
buf ( n373386 , n362136 );
buf ( n373387 , n362037 );
nand ( n53140 , n373386 , n373387 );
buf ( n373389 , n53140 );
buf ( n373390 , n373389 );
nand ( n53143 , n373385 , n373390 );
buf ( n373392 , n53143 );
buf ( n373393 , n373392 );
buf ( n373394 , n362066 );
and ( n373395 , n373393 , n373394 );
buf ( n373396 , n372619 );
buf ( n373397 , n362030 );
and ( n373398 , n373396 , n373397 );
buf ( n373399 , n373398 );
buf ( n373400 , n373399 );
nor ( n373401 , n373395 , n373400 );
buf ( n373402 , n373401 );
buf ( n373403 , n373402 );
not ( n53156 , n373403 );
buf ( n373405 , n53156 );
xor ( n373406 , n52674 , n373405 );
buf ( n373407 , n372848 );
buf ( n373408 , n372824 );
or ( n373409 , n373407 , n373408 );
buf ( n373410 , n372866 );
nand ( n373411 , n373409 , n373410 );
buf ( n373412 , n373411 );
buf ( n373413 , n373412 );
buf ( n373414 , n372824 );
buf ( n373415 , n372848 );
nand ( n373416 , n373414 , n373415 );
buf ( n373417 , n373416 );
buf ( n373418 , n373417 );
nand ( n373419 , n373413 , n373418 );
buf ( n373420 , n373419 );
xnor ( n373421 , n373406 , n373420 );
buf ( n373422 , n373421 );
not ( n373423 , n373422 );
buf ( n373424 , n373423 );
buf ( n373425 , n373424 );
xnor ( n373426 , n53132 , n373425 );
buf ( n373427 , n373426 );
xor ( n373428 , n373308 , n373427 );
xor ( n373429 , n372679 , n372696 );
and ( n373430 , n373429 , n372715 );
and ( n373431 , n372679 , n372696 );
or ( n373432 , n373430 , n373431 );
buf ( n373433 , n373432 );
buf ( n373434 , n373433 );
buf ( n373435 , n363210 );
not ( n373436 , n373435 );
buf ( n373437 , n52464 );
not ( n373438 , n373437 );
or ( n373439 , n373436 , n373438 );
and ( n373440 , n360308 , n362426 );
not ( n373441 , n360308 );
and ( n373442 , n373441 , n362435 );
or ( n373443 , n373440 , n373442 );
buf ( n373444 , n373443 );
buf ( n373445 , n42242 );
nand ( n373446 , n373444 , n373445 );
buf ( n373447 , n373446 );
buf ( n373448 , n373447 );
nand ( n373449 , n373439 , n373448 );
buf ( n373450 , n373449 );
buf ( n373451 , n361606 );
not ( n373452 , n373451 );
buf ( n373453 , n372685 );
not ( n373454 , n373453 );
or ( n373455 , n373452 , n373454 );
buf ( n373456 , n363603 );
not ( n373457 , n373456 );
buf ( n373458 , n46236 );
not ( n373459 , n373458 );
or ( n373460 , n373457 , n373459 );
buf ( n373461 , n360885 );
not ( n373462 , n373461 );
buf ( n373463 , n373462 );
buf ( n373464 , n373463 );
not ( n373465 , n373464 );
buf ( n373466 , n361534 );
nand ( n373467 , n373465 , n373466 );
buf ( n373468 , n373467 );
buf ( n373469 , n373468 );
nand ( n373470 , n373460 , n373469 );
buf ( n373471 , n373470 );
buf ( n373472 , n373471 );
buf ( n373473 , n41485 );
nand ( n373474 , n373472 , n373473 );
buf ( n373475 , n373474 );
buf ( n373476 , n373475 );
nand ( n373477 , n373455 , n373476 );
buf ( n373478 , n373477 );
xor ( n373479 , n373450 , n373478 );
not ( n373480 , n372641 );
nor ( n373481 , n373480 , n41831 );
buf ( n373482 , n47554 );
not ( n373483 , n373482 );
buf ( n373484 , n362803 );
not ( n53161 , n373484 );
or ( n373486 , n373483 , n53161 );
buf ( n373487 , n40251 );
buf ( n373488 , n41772 );
nand ( n53162 , n373487 , n373488 );
buf ( n373490 , n53162 );
buf ( n373491 , n373490 );
nand ( n53165 , n373486 , n373491 );
buf ( n373493 , n53165 );
not ( n53167 , n373493 );
nor ( n53168 , n53167 , n41836 );
nor ( n53169 , n373481 , n53168 );
and ( n53170 , n373479 , n53169 );
not ( n53171 , n373479 );
not ( n53172 , n53169 );
and ( n53173 , n53171 , n53172 );
or ( n373501 , n53170 , n53173 );
buf ( n373502 , n373501 );
xor ( n373503 , n373434 , n373502 );
buf ( n373504 , n52532 );
not ( n53178 , n373504 );
buf ( n373506 , n372799 );
buf ( n373507 , n373506 );
not ( n53181 , n373507 );
or ( n373509 , n53178 , n53181 );
buf ( n373510 , n372799 );
buf ( n373511 , n52532 );
or ( n373512 , n373510 , n373511 );
buf ( n373513 , n372869 );
nand ( n373514 , n373512 , n373513 );
buf ( n373515 , n373514 );
buf ( n373516 , n373515 );
nand ( n53190 , n373509 , n373516 );
buf ( n373518 , n53190 );
buf ( n373519 , n373518 );
xnor ( n373520 , n373503 , n373519 );
buf ( n373521 , n373520 );
xor ( n53195 , n373428 , n373521 );
not ( n53196 , n53195 );
xor ( n53197 , n373240 , n53196 );
not ( n53198 , n372743 );
nand ( n373526 , n53198 , n372749 );
not ( n53200 , n373526 );
not ( n53201 , n52748 );
or ( n53202 , n53200 , n53201 );
not ( n53203 , n372749 );
nand ( n53204 , n53203 , n372743 );
nand ( n53205 , n53202 , n53204 );
buf ( n373533 , n53205 );
not ( n53207 , n373533 );
buf ( n373535 , n53207 );
xnor ( n53209 , n53197 , n373535 );
xnor ( n373537 , n52975 , n53209 );
buf ( n53211 , n373537 );
buf ( n373539 , n372994 );
not ( n53213 , n373539 );
buf ( n373541 , n372602 );
buf ( n373542 , n373541 );
buf ( n373543 , n373542 );
buf ( n373544 , n373543 );
nand ( n373545 , n53213 , n373544 );
buf ( n373546 , n373545 );
buf ( n373547 , n373546 );
buf ( n373548 , n372120 );
and ( n53222 , n373547 , n373548 );
buf ( n373550 , n372994 );
not ( n373551 , n373550 );
buf ( n373552 , n373543 );
nor ( n373553 , n373551 , n373552 );
buf ( n373554 , n373553 );
buf ( n373555 , n373554 );
nor ( n373556 , n53222 , n373555 );
buf ( n373557 , n373556 );
buf ( n373558 , n373557 );
nand ( n373559 , n53211 , n373558 );
buf ( n373560 , n373559 );
buf ( n373561 , n373560 );
nand ( n53235 , n373057 , n373084 , n373561 );
buf ( n373563 , n53235 );
buf ( n373564 , n373563 );
not ( n53238 , n373564 );
nand ( n373566 , n53209 , n373208 );
not ( n373567 , n373566 );
not ( n53241 , n373222 );
or ( n373569 , n373567 , n53241 );
or ( n373570 , n53209 , n373208 );
nand ( n53244 , n373569 , n373570 );
not ( n373572 , n53244 );
buf ( n373573 , n373572 );
xor ( n53247 , n373113 , n373123 );
and ( n373575 , n53247 , n373189 );
and ( n53249 , n373113 , n373123 );
or ( n53250 , n373575 , n53249 );
buf ( n373578 , n53250 );
buf ( n373579 , n373450 );
not ( n53253 , n373579 );
buf ( n373581 , n53172 );
not ( n373582 , n373581 );
or ( n373583 , n53253 , n373582 );
buf ( n373584 , n53169 );
not ( n373585 , n373584 );
buf ( n373586 , n373450 );
not ( n53260 , n373586 );
buf ( n373588 , n53260 );
buf ( n373589 , n373588 );
not ( n373590 , n373589 );
or ( n53264 , n373585 , n373590 );
buf ( n373592 , n373478 );
nand ( n373593 , n53264 , n373592 );
buf ( n373594 , n373593 );
buf ( n373595 , n373594 );
nand ( n53269 , n373583 , n373595 );
buf ( n53270 , n53269 );
buf ( n373598 , n53270 );
not ( n53272 , n373598 );
buf ( n373600 , n41485 );
not ( n53274 , n373600 );
buf ( n373602 , n363603 );
not ( n373603 , n373602 );
buf ( n373604 , n366673 );
not ( n373605 , n373604 );
or ( n373606 , n373603 , n373605 );
buf ( n373607 , n362458 );
buf ( n373608 , n361534 );
nand ( n53282 , n373607 , n373608 );
buf ( n373610 , n53282 );
buf ( n373611 , n373610 );
nand ( n53285 , n373606 , n373611 );
buf ( n373613 , n53285 );
buf ( n373614 , n373613 );
not ( n53288 , n373614 );
or ( n373616 , n53274 , n53288 );
buf ( n373617 , n373471 );
buf ( n373618 , n361606 );
nand ( n373619 , n373617 , n373618 );
buf ( n373620 , n373619 );
buf ( n373621 , n373620 );
nand ( n373622 , n373616 , n373621 );
buf ( n373623 , n373622 );
buf ( n373624 , n373623 );
buf ( n373625 , n41835 );
not ( n373626 , n373625 );
buf ( n373627 , n44570 );
not ( n373628 , n373627 );
buf ( n373629 , n47193 );
not ( n53303 , n373629 );
or ( n53304 , n373628 , n53303 );
buf ( n373632 , n363388 );
buf ( n373633 , n361917 );
nand ( n373634 , n373632 , n373633 );
buf ( n373635 , n373634 );
buf ( n373636 , n373635 );
nand ( n53310 , n53304 , n373636 );
buf ( n373638 , n53310 );
buf ( n373639 , n373638 );
not ( n53313 , n373639 );
or ( n53314 , n373626 , n53313 );
buf ( n373642 , n373493 );
buf ( n373643 , n41830 );
nand ( n53317 , n373642 , n373643 );
buf ( n373645 , n53317 );
buf ( n373646 , n373645 );
nand ( n53320 , n53314 , n373646 );
buf ( n373648 , n53320 );
buf ( n53322 , n373648 );
xor ( n53323 , n373624 , n53322 );
buf ( n373651 , n373137 );
not ( n373652 , n373651 );
buf ( n373653 , n373162 );
not ( n53327 , n373653 );
or ( n373655 , n373652 , n53327 );
buf ( n373656 , n373162 );
buf ( n373657 , n373137 );
or ( n53331 , n373656 , n373657 );
buf ( n373659 , n373187 );
nand ( n53333 , n53331 , n373659 );
buf ( n373661 , n53333 );
buf ( n373662 , n373661 );
nand ( n53336 , n373655 , n373662 );
buf ( n373664 , n53336 );
buf ( n373665 , n373664 );
xnor ( n53339 , n53323 , n373665 );
buf ( n373667 , n53339 );
buf ( n373668 , n373667 );
not ( n53342 , n373668 );
or ( n373670 , n53272 , n53342 );
buf ( n373671 , n53270 );
buf ( n373672 , n373667 );
or ( n53346 , n373671 , n373672 );
nand ( n373674 , n373670 , n53346 );
buf ( n373675 , n373674 );
xor ( n53349 , n373578 , n373675 );
buf ( n373677 , n53349 );
xor ( n53351 , n52944 , n373198 );
and ( n373679 , n53351 , n373205 );
and ( n373680 , n52944 , n373198 );
or ( n53354 , n373679 , n373680 );
buf ( n373682 , n53354 );
buf ( n53356 , n373682 );
xor ( n53357 , n373677 , n53356 );
not ( n373685 , n362066 );
buf ( n373686 , n41892 );
not ( n53360 , n373686 );
buf ( n53361 , n363362 );
not ( n53362 , n53361 );
or ( n53363 , n53360 , n53362 );
buf ( n373691 , n362285 );
buf ( n373692 , n362037 );
nand ( n53366 , n373691 , n373692 );
buf ( n373694 , n53366 );
buf ( n373695 , n373694 );
nand ( n373696 , n53363 , n373695 );
buf ( n373697 , n373696 );
not ( n53371 , n373697 );
or ( n53372 , n373685 , n53371 );
buf ( n373700 , n373392 );
buf ( n373701 , n362030 );
nand ( n53375 , n373700 , n373701 );
buf ( n53376 , n53375 );
nand ( n53377 , n53372 , n53376 );
buf ( n373705 , n373180 );
not ( n53379 , n373705 );
buf ( n373707 , n40059 );
not ( n53381 , n373707 );
or ( n53382 , n53379 , n53381 );
buf ( n373710 , n39946 );
buf ( n373711 , n42911 );
not ( n53385 , n373711 );
buf ( n373713 , n365504 );
not ( n53387 , n373713 );
or ( n53388 , n53385 , n53387 );
buf ( n373716 , n363119 );
buf ( n373717 , n364771 );
nand ( n53391 , n373716 , n373717 );
buf ( n373719 , n53391 );
buf ( n373720 , n373719 );
nand ( n373721 , n53388 , n373720 );
buf ( n373722 , n373721 );
buf ( n373723 , n373722 );
nand ( n53397 , n373710 , n373723 );
buf ( n53398 , n53397 );
buf ( n373726 , n53398 );
nand ( n373727 , n53382 , n373726 );
buf ( n373728 , n373727 );
buf ( n373729 , n373728 );
buf ( n373730 , n373326 );
not ( n53404 , n373730 );
buf ( n373732 , n359809 );
not ( n373733 , n373732 );
or ( n53407 , n53404 , n373733 );
buf ( n373735 , n39592 );
buf ( n373736 , n351320 );
not ( n373737 , n373736 );
buf ( n373738 , n361631 );
not ( n53412 , n373738 );
or ( n373740 , n373737 , n53412 );
buf ( n373741 , n45234 );
buf ( n373742 , n31286 );
nand ( n373743 , n373741 , n373742 );
buf ( n373744 , n373743 );
buf ( n373745 , n373744 );
nand ( n373746 , n373740 , n373745 );
buf ( n373747 , n373746 );
buf ( n373748 , n373747 );
nand ( n53422 , n373735 , n373748 );
buf ( n373750 , n53422 );
buf ( n373751 , n373750 );
nand ( n373752 , n53407 , n373751 );
buf ( n373753 , n373752 );
buf ( n373754 , n373753 );
xor ( n53428 , n373729 , n373754 );
buf ( n373756 , n373156 );
not ( n53430 , n373756 );
buf ( n373758 , n359307 );
not ( n53432 , n373758 );
or ( n53433 , n53430 , n53432 );
buf ( n373761 , n39217 );
buf ( n373762 , n368976 );
buf ( n53436 , n373762 );
buf ( n373764 , n53436 );
and ( n53438 , n373764 , n35548 );
not ( n53439 , n373764 );
and ( n373767 , n53439 , n361851 );
or ( n53441 , n53438 , n373767 );
buf ( n373769 , n53441 );
nand ( n373770 , n373761 , n373769 );
buf ( n373771 , n373770 );
buf ( n373772 , n373771 );
nand ( n53446 , n53433 , n373772 );
buf ( n373774 , n53446 );
buf ( n373775 , n373774 );
xor ( n53449 , n53428 , n373775 );
buf ( n373777 , n53449 );
xor ( n53451 , n53377 , n373777 );
buf ( n373779 , n366434 );
not ( n373780 , n373779 );
buf ( n373781 , n342657 );
buf ( n53455 , n363866 );
and ( n53456 , n373781 , n53455 );
not ( n53457 , n373781 );
buf ( n53458 , n41406 );
and ( n53459 , n53457 , n53458 );
nor ( n53460 , n53456 , n53459 );
buf ( n53461 , n53460 );
buf ( n373789 , n53461 );
not ( n53463 , n373789 );
or ( n53464 , n373780 , n53463 );
buf ( n373792 , n53009 );
buf ( n373793 , n366402 );
nand ( n53467 , n373792 , n373793 );
buf ( n373795 , n53467 );
buf ( n373796 , n373795 );
nand ( n53470 , n53464 , n373796 );
buf ( n373798 , n53470 );
xor ( n53472 , n53451 , n373798 );
buf ( n373800 , n53472 );
not ( n53474 , n373264 );
not ( n53475 , n373280 );
or ( n373803 , n53474 , n53475 );
not ( n373804 , n53037 );
not ( n53478 , n373284 );
or ( n53479 , n373804 , n53478 );
nand ( n373807 , n53479 , n373299 );
nand ( n53481 , n373803 , n373807 );
buf ( n373809 , n53481 );
xor ( n373810 , n373800 , n373809 );
not ( n53484 , n373369 );
not ( n373812 , n373351 );
or ( n53486 , n53484 , n373812 );
not ( n373814 , n373366 );
not ( n53488 , n53100 );
or ( n53489 , n373814 , n53488 );
nand ( n373817 , n53489 , n373332 );
nand ( n53491 , n53486 , n373817 );
buf ( n373819 , n53491 );
not ( n373820 , n42242 );
not ( n53494 , n359781 );
not ( n373822 , n363218 );
and ( n53496 , n53494 , n373822 );
nor ( n53497 , n370257 , n362438 );
nor ( n373825 , n53496 , n53497 );
not ( n373826 , n373825 );
or ( n53500 , n373820 , n373826 );
buf ( n373828 , n373443 );
buf ( n373829 , n363210 );
nand ( n53503 , n373828 , n373829 );
buf ( n53504 , n53503 );
nand ( n373832 , n53500 , n53504 );
buf ( n53506 , n373832 );
xor ( n53507 , n373819 , n53506 );
buf ( n373835 , n46521 );
not ( n373836 , n373835 );
buf ( n373837 , n373292 );
not ( n373838 , n373837 );
or ( n373839 , n373836 , n373838 );
or ( n53513 , n46477 , n363442 );
not ( n53514 , n40083 );
not ( n53515 , n39039 );
or ( n373843 , n53514 , n53515 );
not ( n53517 , n359141 );
nand ( n373845 , n373843 , n53517 );
not ( n53519 , n373845 );
nand ( n53520 , n53519 , n46477 );
nand ( n373848 , n53513 , n53520 );
buf ( n373849 , n373848 );
not ( n53523 , n373849 );
buf ( n373851 , n366654 );
nand ( n373852 , n53523 , n373851 );
buf ( n373853 , n373852 );
buf ( n373854 , n373853 );
nand ( n373855 , n373839 , n373854 );
buf ( n373856 , n373855 );
buf ( n373857 , n373856 );
xor ( n373858 , n53507 , n373857 );
buf ( n373859 , n373858 );
buf ( n373860 , n373859 );
xor ( n53534 , n373810 , n373860 );
buf ( n373862 , n53534 );
buf ( n373863 , n373862 );
xor ( n373864 , n53357 , n373863 );
buf ( n373865 , n373864 );
buf ( n373866 , n373865 );
buf ( n53540 , n53196 );
not ( n53541 , n53540 );
buf ( n53542 , n373535 );
not ( n53543 , n53542 );
or ( n53544 , n53541 , n53543 );
buf ( n373872 , n53195 );
not ( n373873 , n373872 );
buf ( n373874 , n53205 );
not ( n373875 , n373874 );
or ( n373876 , n373873 , n373875 );
buf ( n373877 , n373240 );
nand ( n373878 , n373876 , n373877 );
buf ( n373879 , n373878 );
buf ( n373880 , n373879 );
nand ( n373881 , n53544 , n373880 );
buf ( n373882 , n373881 );
buf ( n373883 , n373882 );
xor ( n373884 , n373866 , n373883 );
xor ( n373885 , n373308 , n373427 );
and ( n373886 , n373885 , n373521 );
and ( n53557 , n373308 , n373427 );
or ( n373888 , n373886 , n53557 );
not ( n53559 , n373501 );
buf ( n373890 , n373433 );
not ( n53561 , n373890 );
buf ( n373892 , n53561 );
nand ( n53563 , n53559 , n373892 );
not ( n53564 , n53563 );
not ( n53565 , n373518 );
or ( n53566 , n53564 , n53565 );
buf ( n373897 , n373892 );
not ( n53568 , n373897 );
buf ( n373899 , n373501 );
nand ( n53570 , n53568 , n373899 );
buf ( n373901 , n53570 );
nand ( n53572 , n53566 , n373901 );
buf ( n373903 , n373372 );
not ( n373904 , n373903 );
buf ( n373905 , n373904 );
buf ( n373906 , n373905 );
not ( n373907 , n373906 );
buf ( n373908 , n373421 );
not ( n53579 , n373908 );
or ( n373910 , n373907 , n53579 );
buf ( n373911 , n53130 );
nand ( n53582 , n373910 , n373911 );
buf ( n373913 , n53582 );
buf ( n373914 , n373913 );
buf ( n373915 , n373424 );
buf ( n373916 , n373372 );
nand ( n373917 , n373915 , n373916 );
buf ( n373918 , n373917 );
buf ( n373919 , n373918 );
nand ( n373920 , n373914 , n373919 );
buf ( n373921 , n373920 );
buf ( n373922 , n373921 );
not ( n373923 , n373922 );
not ( n373924 , n50867 );
buf ( n373925 , n373924 );
buf ( n373926 , n361802 );
and ( n373927 , n373925 , n373926 );
not ( n53598 , n373925 );
buf ( n373929 , n369349 );
and ( n373930 , n53598 , n373929 );
nor ( n373931 , n373927 , n373930 );
buf ( n373932 , n373931 );
buf ( n373933 , n373932 );
not ( n53604 , n373933 );
buf ( n373935 , n45384 );
not ( n373936 , n373935 );
and ( n373937 , n53604 , n373936 );
buf ( n373938 , n373345 );
buf ( n373939 , n372247 );
and ( n373940 , n373938 , n373939 );
nor ( n53611 , n373937 , n373940 );
buf ( n53612 , n53611 );
not ( n373943 , n360574 );
buf ( n373944 , n362452 );
not ( n373945 , n373944 );
buf ( n373946 , n369282 );
not ( n53617 , n373946 );
or ( n373948 , n373945 , n53617 );
buf ( n373949 , n41528 );
buf ( n53620 , n365468 );
nand ( n53621 , n373949 , n53620 );
buf ( n53622 , n53621 );
buf ( n53623 , n53622 );
nand ( n53624 , n373948 , n53623 );
buf ( n53625 , n53624 );
not ( n373956 , n53625 );
or ( n53627 , n373943 , n373956 );
not ( n53628 , n52884 );
not ( n373959 , n52883 );
or ( n53630 , n53628 , n373959 );
nand ( n373961 , n53630 , n40475 );
nand ( n53632 , n53627 , n373961 );
buf ( n373963 , n53632 );
not ( n53634 , n373963 );
buf ( n373965 , n53634 );
and ( n373966 , n53612 , n373965 );
not ( n373967 , n53612 );
and ( n53638 , n373967 , n53632 );
or ( n373969 , n373966 , n53638 );
or ( n373970 , n364899 , n53112 );
buf ( n373971 , n371669 );
buf ( n373972 , n364909 );
and ( n373973 , n373971 , n373972 );
not ( n53644 , n373971 );
buf ( n373975 , n364922 );
and ( n373976 , n53644 , n373975 );
nor ( n373977 , n373973 , n373976 );
buf ( n373978 , n373977 );
not ( n373979 , n373978 );
nand ( n373980 , n373979 , n368038 );
nand ( n53651 , n373970 , n373980 );
and ( n373982 , n373969 , n53651 );
not ( n373983 , n373969 );
not ( n53654 , n53651 );
and ( n373985 , n373983 , n53654 );
nor ( n373986 , n373982 , n373985 );
buf ( n373987 , n43261 );
not ( n373988 , n373987 );
buf ( n373989 , n22772 );
not ( n373990 , n373989 );
buf ( n373991 , n361073 );
not ( n53662 , n373991 );
or ( n373993 , n373990 , n53662 );
buf ( n373994 , n39832 );
buf ( n373995 , n363444 );
nand ( n373996 , n373994 , n373995 );
buf ( n373997 , n373996 );
buf ( n373998 , n373997 );
nand ( n53669 , n373993 , n373998 );
buf ( n374000 , n53669 );
buf ( n374001 , n374000 );
not ( n53672 , n374001 );
or ( n53673 , n373988 , n53672 );
buf ( n374004 , n373270 );
buf ( n374005 , n44796 );
nand ( n374006 , n374004 , n374005 );
buf ( n374007 , n374006 );
buf ( n374008 , n374007 );
nand ( n374009 , n53673 , n374008 );
buf ( n374010 , n374009 );
xor ( n53681 , n373986 , n374010 );
not ( n374012 , n373420 );
not ( n53683 , n52674 );
nand ( n374014 , n53683 , n373402 );
not ( n53685 , n374014 );
or ( n374016 , n374012 , n53685 );
nand ( n374017 , n373405 , n52674 );
nand ( n53688 , n374016 , n374017 );
xor ( n374019 , n53681 , n53688 );
buf ( n374020 , n374019 );
not ( n53691 , n374020 );
buf ( n374022 , n53691 );
buf ( n374023 , n374022 );
not ( n374024 , n374023 );
or ( n53695 , n373923 , n374024 );
buf ( n374026 , n374019 );
buf ( n53697 , n373921 );
not ( n374028 , n53697 );
buf ( n374029 , n374028 );
buf ( n374030 , n374029 );
nand ( n374031 , n374026 , n374030 );
buf ( n374032 , n374031 );
buf ( n374033 , n374032 );
nand ( n374034 , n53695 , n374033 );
buf ( n374035 , n374034 );
xor ( n374036 , n53572 , n374035 );
xor ( n53707 , n373888 , n374036 );
not ( n53708 , n373094 );
nand ( n374039 , n53708 , n52859 );
and ( n374040 , n374039 , n373207 );
and ( n53711 , n52858 , n373094 );
nor ( n374042 , n374040 , n53711 );
xnor ( n374043 , n53707 , n374042 );
buf ( n374044 , n374043 );
xnor ( n374045 , n373884 , n374044 );
buf ( n374046 , n374045 );
buf ( n374047 , n374046 );
not ( n53718 , n374047 );
buf ( n374049 , n53718 );
buf ( n374050 , n374049 );
nand ( n374051 , n373573 , n374050 );
buf ( n374052 , n374051 );
buf ( n374053 , n374052 );
nand ( n53724 , n53238 , n374053 );
buf ( n374055 , n53724 );
buf ( n374056 , n374055 );
not ( n374057 , n374056 );
buf ( n374058 , n374057 );
nand ( n53729 , n372001 , n374058 );
not ( n374060 , n53729 );
buf ( n374061 , n359307 );
not ( n53732 , n374061 );
buf ( n374063 , n355582 );
not ( n374064 , n374063 );
buf ( n374065 , n361751 );
not ( n374066 , n374065 );
or ( n374067 , n374064 , n374066 );
buf ( n374068 , n41946 );
buf ( n374069 , n361851 );
nand ( n374070 , n374068 , n374069 );
buf ( n374071 , n374070 );
buf ( n374072 , n374071 );
nand ( n374073 , n374067 , n374072 );
buf ( n374074 , n374073 );
buf ( n374075 , n374074 );
not ( n374076 , n374075 );
or ( n374077 , n53732 , n374076 );
buf ( n374078 , n363327 );
buf ( n374079 , n39217 );
nand ( n53750 , n374078 , n374079 );
buf ( n374081 , n53750 );
buf ( n374082 , n374081 );
nand ( n53753 , n374077 , n374082 );
buf ( n374084 , n53753 );
buf ( n374085 , n374084 );
buf ( n374086 , n361060 );
not ( n53757 , n374086 );
buf ( n374088 , n363344 );
not ( n374089 , n374088 );
or ( n53760 , n53757 , n374089 );
buf ( n374091 , n42171 );
not ( n53762 , n374091 );
buf ( n374093 , n360893 );
not ( n374094 , n374093 );
buf ( n374095 , n374094 );
buf ( n374096 , n374095 );
not ( n53767 , n374096 );
or ( n374098 , n53762 , n53767 );
buf ( n374099 , n360893 );
buf ( n374100 , n361026 );
nand ( n374101 , n374099 , n374100 );
buf ( n374102 , n374101 );
buf ( n374103 , n374102 );
nand ( n53774 , n374098 , n374103 );
buf ( n53775 , n53774 );
buf ( n374106 , n53775 );
buf ( n374107 , n361022 );
nand ( n374108 , n374106 , n374107 );
buf ( n374109 , n374108 );
buf ( n374110 , n374109 );
nand ( n53781 , n53760 , n374110 );
buf ( n374112 , n53781 );
buf ( n374113 , n374112 );
xor ( n374114 , n374085 , n374113 );
buf ( n374115 , n362066 );
not ( n53786 , n374115 );
buf ( n374117 , n363395 );
not ( n374118 , n374117 );
or ( n374119 , n53786 , n374118 );
buf ( n374120 , n41892 );
not ( n53791 , n374120 );
buf ( n374122 , n40252 );
not ( n374123 , n374122 );
or ( n374124 , n53791 , n374123 );
buf ( n374125 , n42659 );
buf ( n374126 , n362037 );
nand ( n53797 , n374125 , n374126 );
buf ( n374128 , n53797 );
buf ( n374129 , n374128 );
nand ( n374130 , n374124 , n374129 );
buf ( n374131 , n374130 );
buf ( n374132 , n374131 );
buf ( n374133 , n362030 );
nand ( n53804 , n374132 , n374133 );
buf ( n374135 , n53804 );
buf ( n374136 , n374135 );
nand ( n53807 , n374119 , n374136 );
buf ( n53808 , n53807 );
buf ( n374139 , n53808 );
xor ( n53810 , n374114 , n374139 );
buf ( n374141 , n53810 );
buf ( n374142 , n374141 );
not ( n374143 , n374142 );
buf ( n374144 , n42911 );
not ( n374145 , n374144 );
buf ( n374146 , n41623 );
not ( n374147 , n374146 );
or ( n53818 , n374145 , n374147 );
buf ( n374149 , n359950 );
buf ( n374150 , n363071 );
nand ( n53821 , n374149 , n374150 );
buf ( n53822 , n53821 );
buf ( n374153 , n53822 );
nand ( n374154 , n53818 , n374153 );
buf ( n374155 , n374154 );
buf ( n374156 , n374155 );
not ( n374157 , n374156 );
buf ( n374158 , n370350 );
not ( n374159 , n374158 );
or ( n374160 , n374157 , n374159 );
buf ( n374161 , n39891 );
buf ( n374162 , n363581 );
nand ( n53833 , n374161 , n374162 );
buf ( n374164 , n53833 );
buf ( n374165 , n374164 );
nand ( n53836 , n374160 , n374165 );
buf ( n374167 , n53836 );
buf ( n374168 , n374167 );
not ( n53839 , n374168 );
buf ( n374170 , n53839 );
buf ( n374171 , n374170 );
not ( n53842 , n374171 );
not ( n374173 , n360616 );
not ( n53844 , n369349 );
or ( n374175 , n374173 , n53844 );
buf ( n374176 , n363317 );
not ( n53847 , n374176 );
buf ( n374178 , n53847 );
nand ( n374179 , n374178 , n362489 );
nand ( n53850 , n374175 , n374179 );
not ( n374181 , n53850 );
not ( n374182 , n374181 );
buf ( n53853 , n40474 );
buf ( n374184 , n53853 );
not ( n53855 , n374184 );
and ( n53856 , n374182 , n53855 );
buf ( n374187 , n360616 );
not ( n53858 , n374187 );
buf ( n374189 , n362139 );
not ( n53860 , n374189 );
or ( n374191 , n53858 , n53860 );
buf ( n374192 , n362133 );
buf ( n374193 , n362471 );
nand ( n53864 , n374192 , n374193 );
buf ( n374195 , n53864 );
buf ( n374196 , n374195 );
nand ( n53867 , n374191 , n374196 );
buf ( n374198 , n53867 );
and ( n374199 , n374198 , n360577 );
nor ( n53870 , n53856 , n374199 );
buf ( n374201 , n53870 );
not ( n53872 , n374201 );
or ( n374203 , n53842 , n53872 );
buf ( n374204 , n359809 );
buf ( n374205 , n367576 );
not ( n53876 , n374205 );
buf ( n374207 , n45231 );
not ( n53878 , n374207 );
or ( n374209 , n53876 , n53878 );
buf ( n374210 , n39621 );
buf ( n374211 , n44661 );
nand ( n374212 , n374210 , n374211 );
buf ( n374213 , n374212 );
buf ( n374214 , n374213 );
nand ( n53885 , n374209 , n374214 );
buf ( n374216 , n53885 );
buf ( n374217 , n374216 );
and ( n374218 , n374204 , n374217 );
buf ( n374219 , n39592 );
buf ( n374220 , n45459 );
not ( n374221 , n374220 );
buf ( n374222 , n45234 );
not ( n53893 , n374222 );
or ( n374224 , n374221 , n53893 );
buf ( n53895 , n39621 );
buf ( n374226 , n364870 );
or ( n374227 , n53895 , n374226 );
nand ( n53898 , n374224 , n374227 );
buf ( n374229 , n53898 );
buf ( n374230 , n374229 );
and ( n374231 , n374219 , n374230 );
buf ( n374232 , n374231 );
buf ( n374233 , n374232 );
nor ( n53904 , n374218 , n374233 );
buf ( n374235 , n53904 );
buf ( n374236 , n374235 );
not ( n374237 , n374236 );
buf ( n374238 , n374237 );
buf ( n53909 , n374238 );
nand ( n53910 , n374203 , n53909 );
buf ( n53911 , n53910 );
buf ( n374242 , n53911 );
buf ( n374243 , n53870 );
not ( n53914 , n374243 );
buf ( n374245 , n53914 );
buf ( n374246 , n374245 );
buf ( n374247 , n374167 );
nand ( n53918 , n374246 , n374247 );
buf ( n374249 , n53918 );
buf ( n374250 , n374249 );
and ( n53921 , n374242 , n374250 );
buf ( n374252 , n53921 );
buf ( n374253 , n374252 );
not ( n53924 , n374253 );
buf ( n53925 , n53924 );
buf ( n374256 , n53925 );
not ( n53927 , n374256 );
buf ( n374258 , n43283 );
not ( n374259 , n374258 );
buf ( n374260 , n363420 );
not ( n374261 , n374260 );
and ( n53932 , n374259 , n374261 );
and ( n53933 , n41472 , n22772 );
not ( n53934 , n41472 );
and ( n53935 , n53934 , n363444 );
or ( n374266 , n53933 , n53935 );
buf ( n374267 , n374266 );
buf ( n374268 , n44796 );
and ( n53939 , n374267 , n374268 );
nor ( n374270 , n53932 , n53939 );
buf ( n374271 , n374270 );
buf ( n374272 , n374271 );
not ( n53943 , n374272 );
and ( n374274 , n53927 , n53943 );
buf ( n374275 , n374271 );
buf ( n374276 , n53925 );
and ( n53947 , n374275 , n374276 );
nor ( n53948 , n374274 , n53947 );
buf ( n374279 , n53948 );
buf ( n374280 , n374279 );
not ( n53951 , n374280 );
or ( n53952 , n374143 , n53951 );
buf ( n53953 , n374279 );
buf ( n374284 , n374141 );
or ( n374285 , n53953 , n374284 );
nand ( n374286 , n53952 , n374285 );
buf ( n374287 , n374286 );
buf ( n374288 , n374287 );
buf ( n53959 , n361022 );
not ( n53960 , n53959 );
buf ( n374291 , n40893 );
not ( n53962 , n374291 );
buf ( n374293 , n363362 );
not ( n374294 , n374293 );
or ( n374295 , n53962 , n374294 );
buf ( n374296 , n362285 );
buf ( n374297 , n361026 );
nand ( n374298 , n374296 , n374297 );
buf ( n374299 , n374298 );
buf ( n374300 , n374299 );
nand ( n374301 , n374295 , n374300 );
buf ( n374302 , n374301 );
buf ( n53973 , n374302 );
not ( n53974 , n53973 );
or ( n53975 , n53960 , n53974 );
buf ( n53976 , n53775 );
buf ( n53977 , n361060 );
nand ( n53978 , n53976 , n53977 );
buf ( n53979 , n53978 );
buf ( n53980 , n53979 );
nand ( n53981 , n53975 , n53980 );
buf ( n53982 , n53981 );
not ( n374313 , n361609 );
buf ( n374314 , n366725 );
not ( n53985 , n374314 );
buf ( n374316 , n361537 );
nand ( n53987 , n53985 , n374316 );
buf ( n374318 , n53987 );
nand ( n53989 , n363391 , n363603 );
nand ( n53990 , n374318 , n53989 );
not ( n53991 , n53990 );
or ( n374322 , n374313 , n53991 );
buf ( n374323 , n361540 );
not ( n53994 , n374323 );
buf ( n374325 , n46902 );
not ( n53996 , n374325 );
or ( n374327 , n53994 , n53996 );
buf ( n374328 , n40201 );
buf ( n374329 , n361537 );
nand ( n374330 , n374328 , n374329 );
buf ( n374331 , n374330 );
buf ( n374332 , n374331 );
nand ( n374333 , n374327 , n374332 );
buf ( n374334 , n374333 );
nand ( n374335 , n41485 , n374334 );
nand ( n54006 , n374322 , n374335 );
xor ( n54007 , n53982 , n54006 );
buf ( n374338 , n362066 );
not ( n374339 , n374338 );
buf ( n374340 , n374131 );
not ( n374341 , n374340 );
or ( n374342 , n374339 , n374341 );
buf ( n374343 , n41892 );
not ( n374344 , n374343 );
buf ( n374345 , n362461 );
not ( n54016 , n374345 );
or ( n374347 , n374344 , n54016 );
buf ( n374348 , n362467 );
buf ( n374349 , n362037 );
nand ( n374350 , n374348 , n374349 );
buf ( n374351 , n374350 );
buf ( n374352 , n374351 );
nand ( n374353 , n374347 , n374352 );
buf ( n374354 , n374353 );
buf ( n374355 , n374354 );
buf ( n374356 , n362030 );
nand ( n374357 , n374355 , n374356 );
buf ( n374358 , n374357 );
buf ( n374359 , n374358 );
nand ( n54030 , n374342 , n374359 );
buf ( n374361 , n54030 );
xor ( n54032 , n54007 , n374361 );
buf ( n374363 , n54032 );
buf ( n54034 , n53632 );
buf ( n374365 , n360577 );
not ( n54036 , n374365 );
buf ( n374367 , n362452 );
not ( n374368 , n374367 );
buf ( n374369 , n41615 );
not ( n374370 , n374369 );
or ( n374371 , n374368 , n374370 );
buf ( n374372 , n361750 );
buf ( n374373 , n360613 );
nand ( n54044 , n374372 , n374373 );
buf ( n374375 , n54044 );
buf ( n374376 , n374375 );
nand ( n374377 , n374371 , n374376 );
buf ( n374378 , n374377 );
buf ( n374379 , n374378 );
not ( n374380 , n374379 );
or ( n54051 , n54036 , n374380 );
buf ( n374382 , n46557 );
buf ( n374383 , n53625 );
nand ( n54054 , n374382 , n374383 );
buf ( n374385 , n54054 );
buf ( n374386 , n374385 );
nand ( n374387 , n54051 , n374386 );
buf ( n374388 , n374387 );
buf ( n374389 , n374388 );
xor ( n54060 , n54034 , n374389 );
buf ( n374391 , n363291 );
buf ( n374392 , n373978 );
or ( n54063 , n374391 , n374392 );
buf ( n374394 , n369959 );
buf ( n374395 , n42898 );
buf ( n374396 , n359950 );
and ( n54067 , n374395 , n374396 );
not ( n54068 , n374395 );
buf ( n374399 , n42455 );
and ( n54070 , n54068 , n374399 );
nor ( n54071 , n54067 , n54070 );
buf ( n374402 , n54071 );
buf ( n374403 , n374402 );
or ( n374404 , n374394 , n374403 );
nand ( n374405 , n54063 , n374404 );
buf ( n374406 , n374405 );
buf ( n374407 , n374406 );
and ( n374408 , n54060 , n374407 );
and ( n54079 , n54034 , n374389 );
or ( n374410 , n374408 , n54079 );
buf ( n374411 , n374410 );
buf ( n374412 , n374411 );
buf ( n374413 , n41835 );
not ( n374414 , n374413 );
buf ( n374415 , n41778 );
not ( n374416 , n374415 );
buf ( n374417 , n359784 );
not ( n374418 , n374417 );
or ( n374419 , n374416 , n374418 );
buf ( n374420 , n365681 );
not ( n374421 , n374420 );
buf ( n374422 , n374421 );
buf ( n374423 , n374422 );
buf ( n374424 , n361917 );
nand ( n54095 , n374423 , n374424 );
buf ( n374426 , n54095 );
buf ( n374427 , n374426 );
nand ( n374428 , n374419 , n374427 );
buf ( n374429 , n374428 );
buf ( n374430 , n374429 );
not ( n374431 , n374430 );
or ( n54102 , n374414 , n374431 );
buf ( n374433 , n41778 );
not ( n54104 , n374433 );
buf ( n374435 , n360308 );
not ( n54106 , n374435 );
or ( n54107 , n54104 , n54106 );
buf ( n374438 , n40199 );
buf ( n374439 , n361917 );
nand ( n374440 , n374438 , n374439 );
buf ( n374441 , n374440 );
buf ( n374442 , n374441 );
nand ( n374443 , n54107 , n374442 );
buf ( n374444 , n374443 );
buf ( n374445 , n374444 );
buf ( n374446 , n41830 );
nand ( n54117 , n374445 , n374446 );
buf ( n374448 , n54117 );
buf ( n374449 , n374448 );
nand ( n374450 , n54102 , n374449 );
buf ( n374451 , n374450 );
buf ( n54122 , n374451 );
xor ( n54123 , n374412 , n54122 );
buf ( n374454 , n44796 );
not ( n54125 , n374454 );
buf ( n374456 , n22772 );
not ( n374457 , n374456 );
buf ( n374458 , n362752 );
not ( n54129 , n374458 );
or ( n374460 , n374457 , n54129 );
buf ( n374461 , n42606 );
buf ( n374462 , n363444 );
nand ( n374463 , n374461 , n374462 );
buf ( n374464 , n374463 );
buf ( n374465 , n374464 );
nand ( n54136 , n374460 , n374465 );
buf ( n374467 , n54136 );
buf ( n374468 , n374467 );
not ( n54139 , n374468 );
or ( n54140 , n54125 , n54139 );
buf ( n374471 , n22772 );
buf ( n374472 , n363869 );
and ( n54143 , n374471 , n374472 );
not ( n54144 , n374471 );
buf ( n374475 , n360116 );
and ( n54146 , n54144 , n374475 );
nor ( n54147 , n54143 , n54146 );
buf ( n374478 , n54147 );
buf ( n374479 , n374478 );
buf ( n374480 , n43261 );
nand ( n54151 , n374479 , n374480 );
buf ( n374482 , n54151 );
buf ( n374483 , n374482 );
nand ( n54154 , n54140 , n374483 );
buf ( n374485 , n54154 );
buf ( n374486 , n374485 );
and ( n54157 , n54123 , n374486 );
and ( n54158 , n374412 , n54122 );
or ( n54159 , n54157 , n54158 );
buf ( n374490 , n54159 );
buf ( n374491 , n374490 );
xor ( n54162 , n374363 , n374491 );
buf ( n374493 , n366431 );
not ( n54164 , n374493 );
buf ( n374495 , n50782 );
not ( n54166 , n374495 );
or ( n54167 , n54164 , n54166 );
buf ( n374498 , n22710 );
not ( n54169 , n374498 );
buf ( n374500 , n363439 );
not ( n54171 , n374500 );
or ( n54172 , n54169 , n54171 );
buf ( n374503 , n363442 );
buf ( n374504 , n342657 );
nand ( n54175 , n374503 , n374504 );
buf ( n374506 , n54175 );
buf ( n374507 , n374506 );
nand ( n54178 , n54172 , n374507 );
buf ( n374509 , n54178 );
buf ( n374510 , n374509 );
nand ( n54181 , n54167 , n374510 );
buf ( n374512 , n54181 );
buf ( n374513 , n374512 );
not ( n54184 , n39949 );
xor ( n54185 , n362552 , n365945 );
not ( n54186 , n54185 );
or ( n54187 , n54184 , n54186 );
not ( n54188 , n42355 );
not ( n54189 , n363122 );
or ( n54190 , n54188 , n54189 );
buf ( n374521 , n352119 );
buf ( n374522 , n365507 );
nand ( n54193 , n374521 , n374522 );
buf ( n374524 , n54193 );
nand ( n54195 , n54190 , n374524 );
nand ( n54196 , n54195 , n40059 );
nand ( n54197 , n54187 , n54196 );
buf ( n374528 , n355582 );
not ( n54199 , n374528 );
buf ( n374530 , n361712 );
not ( n54201 , n374530 );
or ( n54202 , n54199 , n54201 );
buf ( n374533 , n361717 );
buf ( n374534 , n361851 );
nand ( n54205 , n374533 , n374534 );
buf ( n374536 , n54205 );
buf ( n374537 , n374536 );
nand ( n54208 , n54202 , n374537 );
buf ( n374539 , n54208 );
buf ( n374540 , n374539 );
not ( n54211 , n374540 );
buf ( n374542 , n359307 );
not ( n54213 , n374542 );
or ( n54214 , n54211 , n54213 );
buf ( n374545 , n41528 );
not ( n54216 , n374545 );
buf ( n374547 , n54216 );
and ( n54218 , n355582 , n374547 );
not ( n54219 , n355582 );
and ( n54220 , n54219 , n361673 );
or ( n54221 , n54218 , n54220 );
buf ( n374552 , n54221 );
buf ( n374553 , n39217 );
nand ( n54224 , n374552 , n374553 );
buf ( n374555 , n54224 );
buf ( n374556 , n374555 );
nand ( n54227 , n54214 , n374556 );
buf ( n374558 , n54227 );
xor ( n54229 , n54197 , n374558 );
buf ( n374560 , n360601 );
not ( n54231 , n374560 );
buf ( n374562 , n374378 );
not ( n54233 , n374562 );
or ( n54234 , n54231 , n54233 );
nand ( n54235 , n53850 , n360577 );
buf ( n374566 , n54235 );
nand ( n54237 , n54234 , n374566 );
buf ( n374568 , n54237 );
and ( n54239 , n54229 , n374568 );
and ( n54240 , n54197 , n374558 );
or ( n54241 , n54239 , n54240 );
buf ( n374572 , n54241 );
xor ( n54243 , n374513 , n374572 );
buf ( n374574 , n54185 );
not ( n54245 , n374574 );
buf ( n374576 , n40059 );
not ( n54247 , n374576 );
or ( n54248 , n54245 , n54247 );
buf ( n374579 , n43389 );
buf ( n374580 , n39949 );
nand ( n54251 , n374579 , n374580 );
buf ( n374582 , n54251 );
buf ( n374583 , n374582 );
nand ( n54254 , n54248 , n374583 );
buf ( n374585 , n54254 );
buf ( n374586 , n374585 );
buf ( n374587 , n374229 );
not ( n54258 , n374587 );
buf ( n374589 , n359809 );
not ( n54260 , n374589 );
or ( n54261 , n54258 , n54260 );
buf ( n374592 , n362521 );
buf ( n374593 , n363055 );
nand ( n54264 , n374592 , n374593 );
buf ( n374595 , n54264 );
buf ( n374596 , n374595 );
nand ( n54267 , n54261 , n374596 );
buf ( n374598 , n54267 );
buf ( n374599 , n374598 );
xor ( n54270 , n374586 , n374599 );
buf ( n374601 , n39217 );
not ( n54272 , n374601 );
buf ( n374603 , n374074 );
not ( n54274 , n374603 );
or ( n54275 , n54272 , n54274 );
buf ( n374606 , n359307 );
buf ( n374607 , n54221 );
nand ( n54278 , n374606 , n374607 );
buf ( n374609 , n54278 );
buf ( n374610 , n374609 );
nand ( n54281 , n54275 , n374610 );
buf ( n374612 , n54281 );
buf ( n374613 , n374612 );
xor ( n54284 , n54270 , n374613 );
buf ( n374615 , n54284 );
buf ( n374616 , n374615 );
xor ( n54287 , n54243 , n374616 );
buf ( n374618 , n54287 );
buf ( n374619 , n374618 );
and ( n54290 , n54162 , n374619 );
and ( n54291 , n374363 , n374491 );
or ( n54292 , n54290 , n54291 );
buf ( n374623 , n54292 );
buf ( n374624 , n374623 );
xor ( n54295 , n374288 , n374624 );
xor ( n54296 , n53982 , n54006 );
and ( n54297 , n54296 , n374361 );
and ( n54298 , n53982 , n54006 );
or ( n54299 , n54297 , n54298 );
buf ( n374630 , n54299 );
xor ( n54301 , n374513 , n374572 );
and ( n54302 , n54301 , n374616 );
and ( n54303 , n374513 , n374572 );
or ( n54304 , n54302 , n54303 );
buf ( n374635 , n54304 );
buf ( n374636 , n374635 );
xor ( n54307 , n374630 , n374636 );
buf ( n374638 , n374235 );
buf ( n374639 , n374167 );
xor ( n54310 , n374638 , n374639 );
buf ( n374641 , n374245 );
xnor ( n54312 , n54310 , n374641 );
buf ( n374643 , n54312 );
buf ( n374644 , n374643 );
buf ( n374645 , n41835 );
not ( n54316 , n374645 );
buf ( n374647 , n41778 );
not ( n54318 , n374647 );
buf ( n374649 , n40999 );
not ( n54320 , n374649 );
or ( n54321 , n54318 , n54320 );
buf ( n374652 , n359756 );
buf ( n374653 , n361917 );
nand ( n54324 , n374652 , n374653 );
buf ( n374655 , n54324 );
buf ( n374656 , n374655 );
nand ( n54327 , n54321 , n374656 );
buf ( n374658 , n54327 );
buf ( n374659 , n374658 );
not ( n54330 , n374659 );
or ( n54331 , n54316 , n54330 );
buf ( n374662 , n374429 );
buf ( n374663 , n41830 );
nand ( n54334 , n374662 , n374663 );
buf ( n374665 , n54334 );
buf ( n374666 , n374665 );
nand ( n54337 , n54331 , n374666 );
buf ( n374668 , n54337 );
buf ( n374669 , n374668 );
xor ( n54340 , n374644 , n374669 );
buf ( n374671 , n374402 );
not ( n54342 , n374671 );
buf ( n374673 , n54342 );
buf ( n374674 , n374673 );
not ( n54345 , n374674 );
buf ( n374676 , n359919 );
not ( n54347 , n374676 );
or ( n54348 , n54345 , n54347 );
buf ( n374679 , n39891 );
buf ( n374680 , n374155 );
nand ( n54351 , n374679 , n374680 );
buf ( n374682 , n54351 );
buf ( n374683 , n374682 );
nand ( n54354 , n54348 , n374683 );
buf ( n374685 , n54354 );
xor ( n54356 , n374235 , n374685 );
not ( n54357 , n362066 );
not ( n54358 , n374354 );
or ( n54359 , n54357 , n54358 );
buf ( n374690 , n41892 );
not ( n54361 , n374690 );
buf ( n374692 , n374095 );
not ( n54363 , n374692 );
or ( n54364 , n54361 , n54363 );
buf ( n374695 , n360893 );
buf ( n374696 , n362037 );
nand ( n54367 , n374695 , n374696 );
buf ( n374698 , n54367 );
buf ( n374699 , n374698 );
nand ( n54370 , n54364 , n374699 );
buf ( n374701 , n54370 );
buf ( n374702 , n374701 );
buf ( n374703 , n362030 );
nand ( n54374 , n374702 , n374703 );
buf ( n374705 , n54374 );
nand ( n54376 , n54359 , n374705 );
and ( n54377 , n54356 , n54376 );
and ( n54378 , n374235 , n374685 );
or ( n54379 , n54377 , n54378 );
buf ( n374710 , n54379 );
and ( n54381 , n54340 , n374710 );
and ( n54382 , n374644 , n374669 );
or ( n54383 , n54381 , n54382 );
buf ( n374714 , n54383 );
buf ( n374715 , n374714 );
xor ( n54386 , n54307 , n374715 );
buf ( n374717 , n54386 );
buf ( n374718 , n374717 );
xor ( n54389 , n54295 , n374718 );
buf ( n374720 , n54389 );
buf ( n374721 , n374720 );
xor ( n54392 , n54197 , n374558 );
xor ( n54393 , n54392 , n374568 );
buf ( n374724 , n54393 );
buf ( n374725 , n42242 );
not ( n54396 , n374725 );
buf ( n374727 , n363218 );
not ( n54398 , n374727 );
buf ( n374729 , n366600 );
not ( n54400 , n374729 );
or ( n54401 , n54398 , n54400 );
buf ( n374732 , n40943 );
buf ( n374733 , n362438 );
nand ( n54404 , n374732 , n374733 );
buf ( n374735 , n54404 );
buf ( n374736 , n374735 );
nand ( n54407 , n54401 , n374736 );
buf ( n374738 , n54407 );
buf ( n374739 , n374738 );
not ( n54410 , n374739 );
or ( n54411 , n54396 , n54410 );
and ( n54412 , n44925 , n362426 );
not ( n54413 , n44925 );
and ( n54414 , n54413 , n362435 );
or ( n54415 , n54412 , n54414 );
buf ( n374746 , n54415 );
buf ( n374747 , n363210 );
nand ( n54418 , n374746 , n374747 );
buf ( n374749 , n54418 );
buf ( n374750 , n374749 );
nand ( n54421 , n54411 , n374750 );
buf ( n374752 , n54421 );
buf ( n374753 , n374752 );
xor ( n54424 , n374724 , n374753 );
xor ( n54425 , n374235 , n374685 );
xor ( n54426 , n54425 , n54376 );
buf ( n374757 , n54426 );
and ( n54428 , n54424 , n374757 );
and ( n54429 , n374724 , n374753 );
or ( n54430 , n54428 , n54429 );
buf ( n374761 , n54430 );
buf ( n374762 , n374761 );
buf ( n374763 , n366402 );
not ( n54434 , n374763 );
buf ( n374765 , n22710 );
not ( n54436 , n374765 );
buf ( n374767 , n40091 );
not ( n54438 , n374767 );
or ( n54439 , n54436 , n54438 );
buf ( n374770 , n40899 );
buf ( n374771 , n342657 );
nand ( n54442 , n374770 , n374771 );
buf ( n374773 , n54442 );
buf ( n374774 , n374773 );
nand ( n54445 , n54439 , n374774 );
buf ( n374776 , n54445 );
buf ( n374777 , n374776 );
not ( n54448 , n374777 );
or ( n54449 , n54434 , n54448 );
buf ( n374780 , n366434 );
buf ( n374781 , n374509 );
nand ( n54452 , n374780 , n374781 );
buf ( n374783 , n54452 );
buf ( n374784 , n374783 );
nand ( n54455 , n54449 , n374784 );
buf ( n374786 , n54455 );
buf ( n54457 , n374786 );
buf ( n374788 , n54457 );
not ( n54459 , n374788 );
buf ( n374790 , n361060 );
not ( n54461 , n374790 );
buf ( n374792 , n42171 );
not ( n54463 , n374792 );
buf ( n374794 , n45718 );
not ( n54465 , n374794 );
or ( n54466 , n54463 , n54465 );
buf ( n374797 , n362133 );
buf ( n374798 , n361026 );
nand ( n54469 , n374797 , n374798 );
buf ( n374800 , n54469 );
buf ( n374801 , n374800 );
nand ( n54472 , n54466 , n374801 );
buf ( n374803 , n54472 );
buf ( n374804 , n374803 );
not ( n54475 , n374804 );
or ( n54476 , n54461 , n54475 );
buf ( n374807 , n373932 );
not ( n54478 , n374807 );
buf ( n374809 , n361022 );
nand ( n54480 , n54478 , n374809 );
buf ( n374811 , n54480 );
buf ( n374812 , n374811 );
nand ( n54483 , n54476 , n374812 );
buf ( n374814 , n54483 );
not ( n54485 , n374814 );
buf ( n374816 , n363603 );
not ( n54487 , n374816 );
buf ( n374818 , n54487 );
buf ( n374819 , n374818 );
not ( n54490 , n374819 );
not ( n54491 , n367158 );
buf ( n374822 , n54491 );
not ( n54493 , n374822 );
or ( n54494 , n54490 , n54493 );
buf ( n374825 , n40251 );
not ( n54496 , n374825 );
buf ( n374827 , n363603 );
nand ( n54498 , n54496 , n374827 );
buf ( n374829 , n54498 );
buf ( n374830 , n374829 );
nand ( n54501 , n54494 , n374830 );
buf ( n374832 , n54501 );
buf ( n374833 , n374832 );
buf ( n374834 , n41485 );
and ( n54505 , n374833 , n374834 );
buf ( n374836 , n373613 );
not ( n54507 , n374836 );
buf ( n374838 , n361603 );
nor ( n54509 , n54507 , n374838 );
buf ( n374840 , n54509 );
buf ( n374841 , n374840 );
nor ( n54512 , n54505 , n374841 );
buf ( n374843 , n54512 );
nand ( n54514 , n54485 , n374843 );
not ( n54515 , n54514 );
xor ( n54516 , n373729 , n373754 );
and ( n54517 , n54516 , n373775 );
and ( n54518 , n373729 , n373754 );
or ( n54519 , n54517 , n54518 );
buf ( n374850 , n54519 );
not ( n54521 , n374850 );
or ( n54522 , n54515 , n54521 );
buf ( n374853 , n374843 );
not ( n54524 , n374853 );
buf ( n374855 , n54524 );
buf ( n374856 , n374855 );
buf ( n374857 , n374814 );
nand ( n54528 , n374856 , n374857 );
buf ( n374859 , n54528 );
nand ( n54530 , n54522 , n374859 );
buf ( n374861 , n54530 );
not ( n54532 , n374861 );
or ( n54533 , n54459 , n54532 );
buf ( n374864 , n374786 );
buf ( n374865 , n54530 );
or ( n54536 , n374864 , n374865 );
buf ( n374867 , n362030 );
not ( n54538 , n374867 );
buf ( n374869 , n373697 );
not ( n54540 , n374869 );
or ( n54541 , n54538 , n54540 );
buf ( n374872 , n374701 );
buf ( n374873 , n362066 );
nand ( n54544 , n374872 , n374873 );
buf ( n374875 , n54544 );
buf ( n374876 , n374875 );
nand ( n54547 , n54541 , n374876 );
buf ( n374878 , n54547 );
buf ( n374879 , n374878 );
not ( n54550 , n374879 );
buf ( n374881 , n367759 );
not ( n54552 , n374881 );
buf ( n374883 , n373638 );
not ( n54554 , n374883 );
or ( n54555 , n54552 , n54554 );
buf ( n374886 , n374444 );
buf ( n374887 , n41835 );
nand ( n54558 , n374886 , n374887 );
buf ( n374889 , n54558 );
buf ( n374890 , n374889 );
nand ( n54561 , n54555 , n374890 );
buf ( n374892 , n54561 );
buf ( n374893 , n374892 );
not ( n54564 , n374893 );
or ( n54565 , n54550 , n54564 );
buf ( n374896 , n374892 );
buf ( n374897 , n374878 );
or ( n54568 , n374896 , n374897 );
buf ( n374899 , n373747 );
not ( n54570 , n374899 );
buf ( n374901 , n45795 );
not ( n54572 , n374901 );
or ( n54573 , n54570 , n54572 );
buf ( n374904 , n362521 );
buf ( n374905 , n374216 );
nand ( n54576 , n374904 , n374905 );
buf ( n374907 , n54576 );
buf ( n374908 , n374907 );
nand ( n54579 , n54573 , n374908 );
buf ( n374910 , n54579 );
buf ( n374911 , n373722 );
not ( n54582 , n374911 );
buf ( n374913 , n40058 );
not ( n54584 , n374913 );
or ( n54585 , n54582 , n54584 );
nand ( n54586 , n54195 , n39949 );
buf ( n374917 , n54586 );
nand ( n54588 , n54585 , n374917 );
buf ( n374919 , n54588 );
xor ( n54590 , n374910 , n374919 );
buf ( n374921 , n53441 );
not ( n54592 , n374921 );
buf ( n374923 , n45204 );
not ( n54594 , n374923 );
or ( n54595 , n54592 , n54594 );
buf ( n374926 , n374539 );
buf ( n374927 , n39217 );
nand ( n54598 , n374926 , n374927 );
buf ( n374929 , n54598 );
buf ( n374930 , n374929 );
nand ( n54601 , n54595 , n374930 );
buf ( n374932 , n54601 );
xor ( n54603 , n54590 , n374932 );
buf ( n374934 , n54603 );
nand ( n54605 , n54568 , n374934 );
buf ( n374936 , n54605 );
buf ( n374937 , n374936 );
nand ( n54608 , n54565 , n374937 );
buf ( n374939 , n54608 );
buf ( n374940 , n374939 );
nand ( n54611 , n54536 , n374940 );
buf ( n374942 , n54611 );
buf ( n374943 , n374942 );
nand ( n54614 , n54533 , n374943 );
buf ( n374945 , n54614 );
buf ( n374946 , n374945 );
xor ( n54617 , n374762 , n374946 );
buf ( n374948 , n43261 );
not ( n54619 , n374948 );
buf ( n374950 , n374266 );
not ( n54621 , n374950 );
or ( n54622 , n54619 , n54621 );
buf ( n374953 , n374478 );
buf ( n374954 , n44796 );
nand ( n54625 , n374953 , n374954 );
buf ( n374956 , n54625 );
buf ( n374957 , n374956 );
nand ( n54628 , n54622 , n374957 );
buf ( n374959 , n54628 );
buf ( n374960 , n374959 );
buf ( n374961 , n363218 );
not ( n54632 , n374961 );
buf ( n374963 , n363172 );
not ( n54634 , n374963 );
or ( n54635 , n54632 , n54634 );
buf ( n374966 , n42606 );
buf ( n374967 , n362438 );
nand ( n54638 , n374966 , n374967 );
buf ( n374969 , n54638 );
buf ( n374970 , n374969 );
nand ( n54641 , n54635 , n374970 );
buf ( n374972 , n54641 );
not ( n54643 , n374972 );
not ( n54644 , n42242 );
or ( n54645 , n54643 , n54644 );
buf ( n374976 , n374738 );
not ( n54647 , n374976 );
buf ( n374978 , n54647 );
or ( n54649 , n374978 , n42266 );
nand ( n54650 , n54645 , n54649 );
buf ( n374981 , n54650 );
xor ( n54652 , n374960 , n374981 );
buf ( n374983 , n361060 );
not ( n54654 , n374983 );
buf ( n374985 , n374302 );
not ( n54656 , n374985 );
or ( n54657 , n54654 , n54656 );
buf ( n374988 , n374803 );
buf ( n374989 , n361022 );
nand ( n54660 , n374988 , n374989 );
buf ( n374991 , n54660 );
buf ( n374992 , n374991 );
nand ( n54663 , n54657 , n374992 );
buf ( n374994 , n54663 );
buf ( n374995 , n374994 );
xor ( n54666 , n374910 , n374919 );
and ( n54667 , n54666 , n374932 );
and ( n54668 , n374910 , n374919 );
or ( n54669 , n54667 , n54668 );
buf ( n375000 , n54669 );
xor ( n54671 , n374995 , n375000 );
buf ( n375002 , n41485 );
not ( n54673 , n375002 );
buf ( n375004 , n53990 );
not ( n54675 , n375004 );
or ( n54676 , n54673 , n54675 );
buf ( n375007 , n374832 );
buf ( n375008 , n361609 );
nand ( n54679 , n375007 , n375008 );
buf ( n375010 , n54679 );
buf ( n375011 , n375010 );
nand ( n54682 , n54676 , n375011 );
buf ( n375013 , n54682 );
buf ( n375014 , n375013 );
and ( n54685 , n54671 , n375014 );
and ( n54686 , n374995 , n375000 );
or ( n54687 , n54685 , n54686 );
buf ( n375018 , n54687 );
buf ( n375019 , n375018 );
xor ( n54690 , n54652 , n375019 );
buf ( n375021 , n54690 );
buf ( n375022 , n375021 );
and ( n54693 , n54617 , n375022 );
and ( n54694 , n374762 , n374946 );
or ( n54695 , n54693 , n54694 );
buf ( n375026 , n54695 );
buf ( n375027 , n375026 );
buf ( n375028 , n360577 );
not ( n54699 , n375028 );
buf ( n375030 , n363372 );
not ( n54701 , n375030 );
or ( n54702 , n54699 , n54701 );
buf ( n375033 , n374198 );
buf ( n375034 , n360601 );
nand ( n54705 , n375033 , n375034 );
buf ( n375036 , n54705 );
buf ( n375037 , n375036 );
nand ( n54708 , n54702 , n375037 );
buf ( n375039 , n54708 );
buf ( n375040 , n375039 );
buf ( n375041 , n41485 );
not ( n54712 , n375041 );
buf ( n375043 , n363607 );
not ( n54714 , n375043 );
or ( n54715 , n54712 , n54714 );
buf ( n375046 , n374334 );
buf ( n375047 , n361609 );
nand ( n54718 , n375046 , n375047 );
buf ( n375049 , n54718 );
buf ( n375050 , n375049 );
nand ( n54721 , n54715 , n375050 );
buf ( n375052 , n54721 );
buf ( n375053 , n375052 );
xor ( n54724 , n375040 , n375053 );
buf ( n375055 , n42242 );
not ( n54726 , n375055 );
buf ( n375057 , n363505 );
not ( n54728 , n375057 );
or ( n54729 , n54726 , n54728 );
buf ( n375060 , n374972 );
buf ( n375061 , n363210 );
nand ( n54732 , n375060 , n375061 );
buf ( n375063 , n54732 );
buf ( n375064 , n375063 );
nand ( n54735 , n54729 , n375064 );
buf ( n375066 , n54735 );
buf ( n375067 , n375066 );
xor ( n54738 , n54724 , n375067 );
buf ( n375069 , n54738 );
buf ( n375070 , n375069 );
xor ( n54741 , n374960 , n374981 );
and ( n54742 , n54741 , n375019 );
and ( n54743 , n374960 , n374981 );
or ( n54744 , n54742 , n54743 );
buf ( n375075 , n54744 );
buf ( n375076 , n375075 );
xor ( n54747 , n375070 , n375076 );
xor ( n54748 , n374586 , n374599 );
and ( n54749 , n54748 , n374613 );
and ( n54750 , n374586 , n374599 );
or ( n54751 , n54749 , n54750 );
buf ( n375082 , n54751 );
buf ( n375083 , n375082 );
xor ( n54754 , n363539 , n363567 );
xor ( n54755 , n54754 , n363592 );
buf ( n375086 , n54755 );
buf ( n375087 , n375086 );
xor ( n54758 , n375083 , n375087 );
not ( n54759 , n41835 );
not ( n54760 , n363517 );
or ( n54761 , n54759 , n54760 );
buf ( n375092 , n374658 );
not ( n54763 , n375092 );
buf ( n375094 , n54763 );
or ( n54765 , n375094 , n41831 );
nand ( n54766 , n54761 , n54765 );
buf ( n375097 , n54766 );
xor ( n54768 , n54758 , n375097 );
buf ( n375099 , n54768 );
buf ( n375100 , n375099 );
xor ( n54771 , n54747 , n375100 );
buf ( n375102 , n54771 );
buf ( n375103 , n375102 );
xor ( n54774 , n375027 , n375103 );
xor ( n54775 , n374644 , n374669 );
xor ( n54776 , n54775 , n374710 );
buf ( n375107 , n54776 );
buf ( n375108 , n375107 );
xor ( n54779 , n374995 , n375000 );
xor ( n54780 , n54779 , n375014 );
buf ( n375111 , n54780 );
buf ( n375112 , n375111 );
and ( n54783 , n371300 , n372473 );
nor ( n54784 , n54783 , n373848 );
not ( n54785 , n54784 );
not ( n54786 , n54785 );
not ( n54787 , n42242 );
not ( n54788 , n54415 );
or ( n54789 , n54787 , n54788 );
not ( n54790 , n42266 );
nand ( n54791 , n54790 , n373825 );
nand ( n54792 , n54789 , n54791 );
not ( n54793 , n54792 );
or ( n54794 , n54786 , n54793 );
or ( n54795 , n54792 , n54785 );
not ( n54796 , n53632 );
not ( n54797 , n53612 );
or ( n54798 , n54796 , n54797 );
nand ( n54799 , n54798 , n53651 );
buf ( n375130 , n54799 );
buf ( n375131 , n53612 );
not ( n54802 , n375131 );
buf ( n375133 , n373965 );
nand ( n54804 , n54802 , n375133 );
buf ( n375135 , n54804 );
buf ( n375136 , n375135 );
nand ( n54807 , n375130 , n375136 );
buf ( n375138 , n54807 );
nand ( n54809 , n54795 , n375138 );
nand ( n54810 , n54794 , n54809 );
buf ( n375141 , n54810 );
xor ( n54812 , n375112 , n375141 );
xor ( n54813 , n374412 , n54122 );
xor ( n54814 , n54813 , n374486 );
buf ( n375145 , n54814 );
buf ( n375146 , n375145 );
and ( n54817 , n54812 , n375146 );
and ( n54818 , n375112 , n375141 );
or ( n54819 , n54817 , n54818 );
buf ( n375150 , n54819 );
buf ( n375151 , n375150 );
xor ( n54822 , n375108 , n375151 );
xor ( n54823 , n374363 , n374491 );
xor ( n54824 , n54823 , n374619 );
buf ( n375155 , n54824 );
buf ( n375156 , n375155 );
and ( n54827 , n54822 , n375156 );
and ( n54828 , n375108 , n375151 );
or ( n54829 , n54827 , n54828 );
buf ( n375160 , n54829 );
buf ( n375161 , n375160 );
xor ( n54832 , n54774 , n375161 );
buf ( n375163 , n54832 );
buf ( n375164 , n375163 );
xor ( n54835 , n374721 , n375164 );
buf ( n375166 , n366434 );
not ( n54837 , n375166 );
buf ( n375168 , n374776 );
not ( n54839 , n375168 );
or ( n54840 , n54837 , n54839 );
buf ( n375171 , n53461 );
buf ( n375172 , n366402 );
nand ( n54843 , n375171 , n375172 );
buf ( n375174 , n54843 );
buf ( n375175 , n375174 );
nand ( n54846 , n54840 , n375175 );
buf ( n375177 , n54846 );
buf ( n375178 , n375177 );
xor ( n54849 , n54034 , n374389 );
xor ( n54850 , n54849 , n374407 );
buf ( n375181 , n54850 );
buf ( n375182 , n375181 );
xor ( n54853 , n375178 , n375182 );
buf ( n375184 , n44796 );
not ( n54855 , n375184 );
buf ( n375186 , n374000 );
not ( n54857 , n375186 );
or ( n54858 , n54855 , n54857 );
buf ( n375189 , n374467 );
buf ( n375190 , n43261 );
nand ( n54861 , n375189 , n375190 );
buf ( n375192 , n54861 );
buf ( n375193 , n375192 );
nand ( n54864 , n54858 , n375193 );
buf ( n375195 , n54864 );
buf ( n375196 , n375195 );
and ( n54867 , n54853 , n375196 );
and ( n54868 , n375178 , n375182 );
or ( n54869 , n54867 , n54868 );
buf ( n375200 , n54869 );
buf ( n375201 , n375200 );
xor ( n54872 , n374724 , n374753 );
xor ( n54873 , n54872 , n374757 );
buf ( n375204 , n54873 );
buf ( n375205 , n375204 );
xor ( n54876 , n375201 , n375205 );
buf ( n375207 , n373623 );
not ( n54878 , n375207 );
buf ( n375209 , n373648 );
not ( n54880 , n375209 );
or ( n54881 , n54878 , n54880 );
buf ( n375212 , n373648 );
buf ( n375213 , n373623 );
or ( n54884 , n375212 , n375213 );
buf ( n375215 , n373664 );
nand ( n54886 , n54884 , n375215 );
buf ( n375217 , n54886 );
buf ( n375218 , n375217 );
nand ( n54889 , n54881 , n375218 );
buf ( n375220 , n54889 );
buf ( n375221 , n375220 );
not ( n54892 , n375221 );
buf ( n375223 , n54892 );
buf ( n375224 , n375223 );
not ( n54895 , n375224 );
buf ( n375226 , n374814 );
buf ( n375227 , n374855 );
xor ( n54898 , n375226 , n375227 );
buf ( n375229 , n374850 );
xnor ( n54900 , n54898 , n375229 );
buf ( n375231 , n54900 );
buf ( n375232 , n375231 );
not ( n54903 , n375232 );
or ( n54904 , n54895 , n54903 );
xor ( n54905 , n53377 , n373777 );
and ( n54906 , n54905 , n373798 );
and ( n54907 , n53377 , n373777 );
or ( n54908 , n54906 , n54907 );
buf ( n375239 , n54908 );
nand ( n54910 , n54904 , n375239 );
buf ( n375241 , n54910 );
buf ( n375242 , n375241 );
buf ( n375243 , n375231 );
not ( n54914 , n375243 );
buf ( n375245 , n54914 );
buf ( n375246 , n375245 );
buf ( n375247 , n375220 );
nand ( n54918 , n375246 , n375247 );
buf ( n375249 , n54918 );
buf ( n375250 , n375249 );
nand ( n54921 , n375242 , n375250 );
buf ( n375252 , n54921 );
buf ( n375253 , n375252 );
and ( n54924 , n54876 , n375253 );
and ( n54925 , n375201 , n375205 );
or ( n54926 , n54924 , n54925 );
buf ( n375257 , n54926 );
buf ( n375258 , n375257 );
xor ( n54929 , n374762 , n374946 );
xor ( n54930 , n54929 , n375022 );
buf ( n375261 , n54930 );
buf ( n375262 , n375261 );
xor ( n54933 , n375258 , n375262 );
xor ( n54934 , n375108 , n375151 );
xor ( n54935 , n54934 , n375156 );
buf ( n375266 , n54935 );
buf ( n375267 , n375266 );
and ( n54938 , n54933 , n375267 );
and ( n54939 , n375258 , n375262 );
or ( n54940 , n54938 , n54939 );
buf ( n375271 , n54940 );
buf ( n375272 , n375271 );
xnor ( n54943 , n54835 , n375272 );
buf ( n375274 , n54943 );
buf ( n375275 , n375274 );
xor ( n54946 , n375258 , n375262 );
xor ( n54947 , n54946 , n375267 );
buf ( n375278 , n54947 );
not ( n54949 , n375278 );
xor ( n54950 , n375112 , n375141 );
xor ( n54951 , n54950 , n375146 );
buf ( n375282 , n54951 );
buf ( n375283 , n375282 );
not ( n54954 , n375283 );
buf ( n375285 , n54954 );
not ( n54956 , n375285 );
buf ( n375287 , n374786 );
buf ( n375288 , n374939 );
xor ( n54959 , n375287 , n375288 );
buf ( n375290 , n54530 );
xnor ( n54961 , n54959 , n375290 );
buf ( n375292 , n54961 );
not ( n54963 , n375292 );
and ( n54964 , n54956 , n54963 );
buf ( n375295 , n375285 );
buf ( n375296 , n375292 );
nand ( n54967 , n375295 , n375296 );
buf ( n375298 , n54967 );
xor ( n54969 , n374892 , n374878 );
buf ( n54970 , n54603 );
and ( n54971 , n54969 , n54970 );
not ( n54972 , n54969 );
not ( n54973 , n54970 );
and ( n54974 , n54972 , n54973 );
nor ( n54975 , n54971 , n54974 );
not ( n54976 , n54975 );
buf ( n375307 , n375138 );
not ( n54978 , n375307 );
buf ( n375309 , n54784 );
not ( n54980 , n375309 );
and ( n54981 , n54978 , n54980 );
buf ( n375312 , n54784 );
buf ( n375313 , n375138 );
and ( n54984 , n375312 , n375313 );
nor ( n54985 , n54981 , n54984 );
buf ( n375316 , n54985 );
not ( n54987 , n54792 );
and ( n54988 , n375316 , n54987 );
not ( n54989 , n375316 );
and ( n54990 , n54989 , n54792 );
nor ( n54991 , n54988 , n54990 );
not ( n54992 , n54991 );
nand ( n54993 , n54976 , n54992 );
not ( n54994 , n54993 );
xor ( n54995 , n373986 , n374010 );
and ( n54996 , n54995 , n53688 );
and ( n54997 , n373986 , n374010 );
or ( n54998 , n54996 , n54997 );
not ( n54999 , n54998 );
or ( n55000 , n54994 , n54999 );
buf ( n375331 , n54991 );
buf ( n375332 , n54975 );
nand ( n55003 , n375331 , n375332 );
buf ( n375334 , n55003 );
nand ( n55005 , n55000 , n375334 );
and ( n55006 , n375298 , n55005 );
nor ( n55007 , n54964 , n55006 );
nand ( n55008 , n54949 , n55007 );
xor ( n55009 , n373819 , n53506 );
and ( n55010 , n55009 , n373857 );
and ( n55011 , n373819 , n53506 );
or ( n55012 , n55010 , n55011 );
buf ( n375343 , n55012 );
buf ( n375344 , n375343 );
xor ( n55015 , n375178 , n375182 );
xor ( n55016 , n55015 , n375196 );
buf ( n375347 , n55016 );
buf ( n375348 , n375347 );
xor ( n55019 , n375344 , n375348 );
buf ( n375350 , n53270 );
not ( n55021 , n375350 );
buf ( n375352 , n55021 );
buf ( n375353 , n375352 );
not ( n55024 , n375353 );
buf ( n375355 , n373667 );
not ( n55026 , n375355 );
or ( n55027 , n55024 , n55026 );
buf ( n375358 , n373578 );
nand ( n55029 , n55027 , n375358 );
buf ( n375360 , n55029 );
buf ( n375361 , n375360 );
buf ( n375362 , n373667 );
not ( n55033 , n375362 );
buf ( n375364 , n53270 );
nand ( n55035 , n55033 , n375364 );
buf ( n375366 , n55035 );
buf ( n375367 , n375366 );
nand ( n55038 , n375361 , n375367 );
buf ( n375369 , n55038 );
buf ( n375370 , n375369 );
and ( n55041 , n55019 , n375370 );
and ( n55042 , n375344 , n375348 );
or ( n55043 , n55041 , n55042 );
buf ( n375374 , n55043 );
buf ( n375375 , n375374 );
xor ( n55046 , n375201 , n375205 );
xor ( n55047 , n55046 , n375253 );
buf ( n375378 , n55047 );
buf ( n375379 , n375378 );
xor ( n55050 , n375375 , n375379 );
buf ( n375381 , n375292 );
buf ( n375382 , n55005 );
xor ( n55053 , n375381 , n375382 );
buf ( n375384 , n375282 );
xnor ( n55055 , n55053 , n375384 );
buf ( n375386 , n55055 );
buf ( n375387 , n375386 );
and ( n55058 , n55050 , n375387 );
and ( n55059 , n375375 , n375379 );
or ( n55060 , n55058 , n55059 );
buf ( n375391 , n55060 );
and ( n55062 , n55008 , n375391 );
not ( n55063 , n375278 );
nor ( n55064 , n55063 , n55007 );
nor ( n55065 , n55062 , n55064 );
buf ( n375396 , n55065 );
nand ( n55067 , n375275 , n375396 );
buf ( n375398 , n55067 );
xor ( n55069 , n375391 , n375278 );
xnor ( n55070 , n55069 , n55007 );
buf ( n375401 , n55070 );
buf ( n375402 , n375223 );
not ( n55073 , n375402 );
buf ( n375404 , n375245 );
not ( n55075 , n375404 );
or ( n55076 , n55073 , n55075 );
buf ( n375407 , n375231 );
buf ( n375408 , n375220 );
nand ( n55079 , n375407 , n375408 );
buf ( n375410 , n55079 );
buf ( n375411 , n375410 );
nand ( n55082 , n55076 , n375411 );
buf ( n375413 , n55082 );
buf ( n375414 , n375413 );
buf ( n375415 , n54908 );
not ( n55086 , n375415 );
buf ( n375417 , n55086 );
buf ( n375418 , n375417 );
and ( n55089 , n375414 , n375418 );
not ( n55090 , n375414 );
buf ( n375421 , n54908 );
and ( n55092 , n55090 , n375421 );
nor ( n55093 , n55089 , n55092 );
buf ( n375424 , n55093 );
buf ( n375425 , n375424 );
not ( n55096 , n375425 );
buf ( n375427 , n55096 );
buf ( n375428 , n375427 );
not ( n55099 , n375428 );
buf ( n55100 , n54975 );
xor ( n55101 , n54998 , n55100 );
xnor ( n55102 , n55101 , n54992 );
buf ( n375433 , n55102 );
not ( n55104 , n375433 );
or ( n55105 , n55099 , n55104 );
buf ( n375436 , n55102 );
buf ( n375437 , n375427 );
or ( n55108 , n375436 , n375437 );
xor ( n55109 , n373800 , n373809 );
and ( n55110 , n55109 , n373860 );
and ( n55111 , n373800 , n373809 );
or ( n55112 , n55110 , n55111 );
buf ( n375443 , n55112 );
buf ( n375444 , n375443 );
nand ( n375445 , n55108 , n375444 );
buf ( n375446 , n375445 );
buf ( n375447 , n375446 );
nand ( n375448 , n55105 , n375447 );
buf ( n375449 , n375448 );
buf ( n375450 , n375449 );
xor ( n55121 , n375375 , n375379 );
xor ( n375452 , n55121 , n375387 );
buf ( n375453 , n375452 );
buf ( n375454 , n375453 );
or ( n375455 , n375450 , n375454 );
xor ( n375456 , n375344 , n375348 );
xor ( n375457 , n375456 , n375370 );
buf ( n375458 , n375457 );
buf ( n375459 , n375458 );
not ( n375460 , n375459 );
not ( n55131 , n374022 );
not ( n375462 , n374029 );
and ( n375463 , n55131 , n375462 );
buf ( n375464 , n374022 );
buf ( n375465 , n374029 );
nand ( n55136 , n375464 , n375465 );
buf ( n375467 , n55136 );
and ( n55138 , n375467 , n53572 );
nor ( n55139 , n375463 , n55138 );
buf ( n375470 , n55139 );
nand ( n55141 , n375460 , n375470 );
buf ( n375472 , n55141 );
buf ( n375473 , n375472 );
not ( n55144 , n375473 );
xor ( n55145 , n373677 , n53356 );
and ( n55146 , n55145 , n373863 );
and ( n55147 , n373677 , n53356 );
or ( n55148 , n55146 , n55147 );
buf ( n375479 , n55148 );
buf ( n375480 , n375479 );
not ( n55151 , n375480 );
or ( n55152 , n55144 , n55151 );
buf ( n375483 , n55139 );
not ( n375484 , n375483 );
buf ( n375485 , n375458 );
nand ( n375486 , n375484 , n375485 );
buf ( n375487 , n375486 );
buf ( n375488 , n375487 );
nand ( n55159 , n55152 , n375488 );
buf ( n55160 , n55159 );
buf ( n375491 , n55160 );
nand ( n55162 , n375455 , n375491 );
buf ( n375493 , n55162 );
buf ( n375494 , n375493 );
buf ( n375495 , n375453 );
buf ( n375496 , n375449 );
nand ( n375497 , n375495 , n375496 );
buf ( n375498 , n375497 );
buf ( n375499 , n375498 );
nand ( n375500 , n375494 , n375499 );
buf ( n375501 , n375500 );
buf ( n375502 , n375501 );
nor ( n375503 , n375401 , n375502 );
buf ( n375504 , n375503 );
buf ( n375505 , n375504 );
not ( n55176 , n375505 );
buf ( n55177 , n55176 );
nand ( n375508 , n375398 , n55177 );
not ( n55179 , n374043 );
buf ( n375510 , n373865 );
not ( n375511 , n375510 );
buf ( n375512 , n375511 );
not ( n55183 , n375512 );
and ( n375514 , n55179 , n55183 );
buf ( n375515 , n374043 );
buf ( n375516 , n375512 );
nand ( n375517 , n375515 , n375516 );
buf ( n375518 , n375517 );
and ( n55189 , n375518 , n373882 );
nor ( n375520 , n375514 , n55189 );
xor ( n375521 , n375424 , n375443 );
xor ( n55192 , n375521 , n55102 );
not ( n375523 , n374042 );
not ( n55194 , n373888 );
nand ( n375525 , n374036 , n55194 );
not ( n375526 , n375525 );
or ( n55197 , n375523 , n375526 );
not ( n375528 , n374036 );
not ( n375529 , n55194 );
nand ( n55200 , n375528 , n375529 );
nand ( n375531 , n55197 , n55200 );
xor ( n375532 , n55192 , n375531 );
xor ( n375533 , n375458 , n55139 );
xor ( n55204 , n375533 , n375479 );
xor ( n375535 , n375532 , n55204 );
nand ( n375536 , n375520 , n375535 );
buf ( n375537 , n375449 );
buf ( n375538 , n375453 );
xor ( n375539 , n375537 , n375538 );
buf ( n375540 , n55160 );
xnor ( n55211 , n375539 , n375540 );
buf ( n55212 , n55211 );
xor ( n375543 , n55192 , n375531 );
and ( n55214 , n375543 , n55204 );
and ( n375545 , n55192 , n375531 );
or ( n375546 , n55214 , n375545 );
nand ( n375547 , n55212 , n375546 );
nand ( n55218 , n375536 , n375547 );
nor ( n375549 , n375508 , n55218 );
buf ( n375550 , n375549 );
xor ( n375551 , n363511 , n363520 );
xor ( n375552 , n375551 , n363525 );
buf ( n375553 , n375552 );
buf ( n375554 , n375553 );
xor ( n55225 , n374630 , n374636 );
and ( n55226 , n55225 , n374715 );
and ( n55227 , n374630 , n374636 );
or ( n55228 , n55226 , n55227 );
buf ( n375559 , n55228 );
buf ( n375560 , n375559 );
xor ( n55231 , n375554 , n375560 );
xor ( n55232 , n374085 , n374113 );
and ( n55233 , n55232 , n374139 );
and ( n55234 , n374085 , n374113 );
or ( n55235 , n55233 , n55234 );
buf ( n375566 , n55235 );
buf ( n375567 , n375566 );
buf ( n375568 , n363380 );
not ( n55239 , n375568 );
buf ( n375570 , n363402 );
not ( n55241 , n375570 );
or ( n55242 , n55239 , n55241 );
buf ( n375573 , n363402 );
buf ( n375574 , n363380 );
or ( n55245 , n375573 , n375574 );
nand ( n55246 , n55242 , n55245 );
buf ( n375577 , n55246 );
xor ( n55248 , n363454 , n375577 );
buf ( n375579 , n55248 );
xor ( n375580 , n375567 , n375579 );
xor ( n375581 , n375040 , n375053 );
and ( n55252 , n375581 , n375067 );
and ( n375583 , n375040 , n375053 );
or ( n375584 , n55252 , n375583 );
buf ( n375585 , n375584 );
buf ( n375586 , n375585 );
xor ( n375587 , n375580 , n375586 );
buf ( n375588 , n375587 );
buf ( n375589 , n375588 );
xor ( n375590 , n55231 , n375589 );
buf ( n375591 , n375590 );
xor ( n55262 , n375070 , n375076 );
and ( n375593 , n55262 , n375100 );
and ( n375594 , n375070 , n375076 );
or ( n55265 , n375593 , n375594 );
buf ( n375596 , n55265 );
buf ( n375597 , n375596 );
not ( n375598 , n374141 );
buf ( n55269 , n374271 );
buf ( n375600 , n374252 );
nand ( n375601 , n55269 , n375600 );
buf ( n375602 , n375601 );
not ( n375603 , n375602 );
or ( n375604 , n375598 , n375603 );
buf ( n375605 , n374271 );
not ( n375606 , n375605 );
buf ( n375607 , n53925 );
nand ( n55278 , n375606 , n375607 );
buf ( n375609 , n55278 );
nand ( n55280 , n375604 , n375609 );
buf ( n375611 , n55280 );
xor ( n375612 , n375083 , n375087 );
and ( n375613 , n375612 , n375097 );
and ( n55284 , n375083 , n375087 );
or ( n55285 , n375613 , n55284 );
buf ( n375616 , n55285 );
buf ( n375617 , n375616 );
xor ( n55288 , n375611 , n375617 );
xor ( n375619 , n363535 , n363597 );
xor ( n375620 , n375619 , n363618 );
buf ( n375621 , n375620 );
buf ( n375622 , n375621 );
xor ( n55293 , n55288 , n375622 );
buf ( n375624 , n55293 );
buf ( n375625 , n375624 );
xor ( n375626 , n375597 , n375625 );
xor ( n55297 , n374288 , n374624 );
and ( n55298 , n55297 , n374718 );
and ( n375629 , n374288 , n374624 );
or ( n375630 , n55298 , n375629 );
buf ( n375631 , n375630 );
buf ( n375632 , n375631 );
xor ( n55303 , n375626 , n375632 );
buf ( n375634 , n55303 );
xor ( n375635 , n375591 , n375634 );
xor ( n375636 , n375027 , n375103 );
and ( n55307 , n375636 , n375161 );
and ( n375638 , n375027 , n375103 );
or ( n55309 , n55307 , n375638 );
buf ( n375640 , n55309 );
not ( n375641 , n375640 );
and ( n55312 , n375635 , n375641 );
not ( n375643 , n375635 );
and ( n55314 , n375643 , n375640 );
nor ( n55315 , n55312 , n55314 );
buf ( n375646 , n375163 );
buf ( n375647 , n374720 );
or ( n55318 , n375646 , n375647 );
buf ( n375649 , n375271 );
nand ( n375650 , n55318 , n375649 );
buf ( n375651 , n375650 );
buf ( n375652 , n375651 );
buf ( n55323 , n375163 );
buf ( n55324 , n374720 );
nand ( n55325 , n55323 , n55324 );
buf ( n55326 , n55325 );
buf ( n375657 , n55326 );
nand ( n55328 , n375652 , n375657 );
buf ( n55329 , n55328 );
not ( n375660 , n55329 );
nand ( n55331 , n55315 , n375660 );
buf ( n375662 , n55331 );
xor ( n375663 , n43051 , n363231 );
xor ( n55334 , n375663 , n363257 );
buf ( n375665 , n55334 );
buf ( n375666 , n375665 );
not ( n55337 , n375666 );
xor ( n55338 , n363357 , n363467 );
xor ( n375669 , n55338 , n363471 );
buf ( n375670 , n375669 );
buf ( n375671 , n375670 );
not ( n375672 , n375671 );
or ( n55343 , n55337 , n375672 );
buf ( n375674 , n375665 );
buf ( n375675 , n375670 );
or ( n55346 , n375674 , n375675 );
xor ( n375677 , n375567 , n375579 );
and ( n55348 , n375677 , n375586 );
and ( n375679 , n375567 , n375579 );
or ( n375680 , n55348 , n375679 );
buf ( n375681 , n375680 );
buf ( n375682 , n375681 );
nand ( n375683 , n55346 , n375682 );
buf ( n375684 , n375683 );
buf ( n375685 , n375684 );
nand ( n55356 , n55343 , n375685 );
buf ( n375687 , n55356 );
buf ( n375688 , n375687 );
not ( n55359 , n375688 );
buf ( n375690 , n55359 );
buf ( n375691 , n375690 );
not ( n55362 , n375691 );
xor ( n55363 , n43463 , n363632 );
xor ( n375694 , n55363 , n363637 );
buf ( n375695 , n375694 );
buf ( n375696 , n375695 );
not ( n55367 , n375696 );
or ( n375698 , n55362 , n55367 );
buf ( n375699 , n375695 );
not ( n375700 , n375699 );
buf ( n375701 , n375700 );
buf ( n375702 , n375701 );
buf ( n375703 , n375687 );
nand ( n55374 , n375702 , n375703 );
buf ( n375705 , n55374 );
buf ( n375706 , n375705 );
nand ( n375707 , n375698 , n375706 );
buf ( n375708 , n375707 );
buf ( n375709 , n375708 );
buf ( n375710 , n375616 );
buf ( n375711 , n375621 );
or ( n55382 , n375710 , n375711 );
buf ( n375713 , n55280 );
nand ( n375714 , n55382 , n375713 );
buf ( n375715 , n375714 );
buf ( n375716 , n375715 );
buf ( n375717 , n375616 );
buf ( n375718 , n375621 );
nand ( n55389 , n375717 , n375718 );
buf ( n55390 , n55389 );
buf ( n375721 , n55390 );
and ( n55392 , n375716 , n375721 );
buf ( n375723 , n55392 );
buf ( n375724 , n375723 );
not ( n375725 , n375724 );
buf ( n375726 , n375725 );
buf ( n375727 , n375726 );
not ( n375728 , n375727 );
xor ( n375729 , n363490 , n363530 );
xor ( n55400 , n375729 , n363623 );
buf ( n375731 , n55400 );
buf ( n375732 , n375731 );
not ( n55403 , n375732 );
or ( n55404 , n375728 , n55403 );
xor ( n375735 , n375554 , n375560 );
and ( n55406 , n375735 , n375589 );
and ( n55407 , n375554 , n375560 );
or ( n55408 , n55406 , n55407 );
buf ( n375739 , n55408 );
buf ( n375740 , n375739 );
buf ( n375741 , n375731 );
not ( n55412 , n375741 );
buf ( n375743 , n375723 );
nand ( n375744 , n55412 , n375743 );
buf ( n375745 , n375744 );
buf ( n375746 , n375745 );
nand ( n55417 , n375740 , n375746 );
buf ( n375748 , n55417 );
buf ( n375749 , n375748 );
nand ( n55420 , n55404 , n375749 );
buf ( n375751 , n55420 );
buf ( n375752 , n375751 );
xnor ( n55423 , n375709 , n375752 );
buf ( n375754 , n55423 );
buf ( n375755 , n375754 );
buf ( n375756 , n375665 );
buf ( n375757 , n375681 );
xor ( n55428 , n375756 , n375757 );
buf ( n375759 , n375670 );
xnor ( n55430 , n55428 , n375759 );
buf ( n375761 , n55430 );
buf ( n375762 , n375761 );
xor ( n55433 , n375597 , n375625 );
and ( n375764 , n55433 , n375632 );
and ( n375765 , n375597 , n375625 );
or ( n55436 , n375764 , n375765 );
buf ( n375767 , n55436 );
buf ( n375768 , n375767 );
not ( n375769 , n375768 );
buf ( n375770 , n375769 );
buf ( n375771 , n375770 );
xor ( n375772 , n375762 , n375771 );
buf ( n375773 , n375723 );
not ( n55444 , n375773 );
buf ( n375775 , n375731 );
not ( n375776 , n375775 );
or ( n55447 , n55444 , n375776 );
buf ( n375778 , n375723 );
buf ( n375779 , n375731 );
or ( n375780 , n375778 , n375779 );
nand ( n375781 , n55447 , n375780 );
buf ( n375782 , n375781 );
buf ( n375783 , n375782 );
buf ( n375784 , n375739 );
not ( n55455 , n375784 );
buf ( n375786 , n55455 );
buf ( n375787 , n375786 );
and ( n55458 , n375783 , n375787 );
not ( n55459 , n375783 );
buf ( n375790 , n375739 );
and ( n55461 , n55459 , n375790 );
nor ( n55462 , n55458 , n55461 );
buf ( n375793 , n55462 );
buf ( n375794 , n375793 );
and ( n55465 , n375772 , n375794 );
and ( n55466 , n375762 , n375771 );
or ( n375797 , n55465 , n55466 );
buf ( n375798 , n375797 );
buf ( n375799 , n375798 );
nand ( n55470 , n375755 , n375799 );
buf ( n375801 , n55470 );
buf ( n375802 , n375801 );
xor ( n375803 , n375762 , n375771 );
xor ( n55474 , n375803 , n375794 );
buf ( n375805 , n55474 );
buf ( n55476 , n375805 );
buf ( n375807 , n375634 );
buf ( n55478 , n375591 );
or ( n55479 , n375807 , n55478 );
buf ( n375810 , n55479 );
and ( n375811 , n375810 , n375640 );
and ( n55482 , n375591 , n375634 );
nor ( n55483 , n375811 , n55482 );
buf ( n375814 , n55483 );
nand ( n55485 , n55476 , n375814 );
buf ( n375816 , n55485 );
buf ( n375817 , n375816 );
nand ( n55488 , n375662 , n375802 , n375817 );
buf ( n375819 , n55488 );
buf ( n375820 , n375819 );
buf ( n375821 , n375690 );
not ( n55492 , n375821 );
buf ( n375823 , n375701 );
not ( n55494 , n375823 );
or ( n375825 , n55492 , n55494 );
buf ( n375826 , n375751 );
nand ( n55497 , n375825 , n375826 );
buf ( n375828 , n55497 );
buf ( n375829 , n375828 );
buf ( n375830 , n375695 );
buf ( n375831 , n375687 );
nand ( n55502 , n375830 , n375831 );
buf ( n375833 , n55502 );
buf ( n375834 , n375833 );
nand ( n55505 , n375829 , n375834 );
buf ( n375836 , n55505 );
buf ( n375837 , n375836 );
xor ( n375838 , n363486 , n363642 );
xor ( n55509 , n375838 , n363647 );
buf ( n375840 , n55509 );
buf ( n55511 , n375840 );
nor ( n55512 , n375837 , n55511 );
buf ( n375843 , n55512 );
buf ( n375844 , n375843 );
nor ( n375845 , n375820 , n375844 );
buf ( n375846 , n375845 );
buf ( n375847 , n375846 );
and ( n375848 , n375550 , n375847 );
buf ( n375849 , n375848 );
nand ( n55520 , n374060 , n375849 );
not ( n55521 , n55520 );
not ( n375852 , n55521 );
xnor ( n375853 , n360885 , n369769 );
not ( n375854 , n375853 );
not ( n55525 , n49604 );
and ( n375856 , n375854 , n55525 );
not ( n55527 , n369769 );
not ( n375858 , n360848 );
or ( n55529 , n55527 , n375858 );
buf ( n375860 , n362458 );
buf ( n375861 , n369766 );
nand ( n375862 , n375860 , n375861 );
buf ( n375863 , n375862 );
nand ( n375864 , n55529 , n375863 );
and ( n375865 , n375864 , n49609 );
nor ( n55536 , n375856 , n375865 );
buf ( n375867 , n55536 );
not ( n375868 , n375867 );
not ( n55539 , n362376 );
buf ( n375870 , n55539 );
buf ( n55541 , n31231 );
not ( n375872 , n55541 );
buf ( n375873 , n375872 );
buf ( n375874 , n375873 );
nand ( n375875 , n375870 , n375874 );
buf ( n375876 , n375875 );
nand ( n375877 , n31231 , n362376 );
nand ( n375878 , n375876 , n375877 );
not ( n375879 , n375878 );
not ( n375880 , n363428 );
or ( n375881 , n375879 , n375880 );
not ( n375882 , n363416 );
not ( n375883 , n55539 );
buf ( n375884 , n32202 );
not ( n375885 , n375884 );
buf ( n375886 , n375885 );
not ( n375887 , n375886 );
or ( n375888 , n375883 , n375887 );
nand ( n375889 , n32202 , n362376 );
nand ( n375890 , n375888 , n375889 );
nand ( n375891 , n375882 , n375890 );
nand ( n375892 , n375881 , n375891 );
buf ( n375893 , n375892 );
buf ( n375894 , n366708 );
not ( n375895 , n375894 );
buf ( n375896 , n375895 );
buf ( n375897 , n375896 );
not ( n375898 , n375897 );
buf ( n375899 , n342617 );
buf ( n375900 , n375899 );
buf ( n375901 , n375900 );
or ( n375902 , n32160 , n375901 );
not ( n375903 , n352192 );
nand ( n375904 , n375903 , n375901 );
nand ( n375905 , n375902 , n375904 );
buf ( n375906 , n375905 );
not ( n375907 , n375906 );
or ( n375908 , n375898 , n375907 );
not ( n375909 , n375901 );
not ( n55551 , n31283 );
or ( n375911 , n375909 , n55551 );
buf ( n375912 , n366659 );
not ( n375913 , n375912 );
buf ( n375914 , n375913 );
not ( n55556 , n375914 );
nand ( n375916 , n55556 , n351310 , n351315 );
nand ( n55558 , n375911 , n375916 );
buf ( n375918 , n366649 );
not ( n55560 , n375918 );
buf ( n375920 , n55560 );
nand ( n375921 , n55558 , n375920 );
buf ( n375922 , n375921 );
nand ( n55564 , n375908 , n375922 );
buf ( n55565 , n55564 );
buf ( n375925 , n55565 );
xor ( n55567 , n375893 , n375925 );
not ( n375927 , n342635 );
not ( n375928 , n22698 );
or ( n375929 , n375927 , n375928 );
nand ( n55571 , n375929 , n22704 );
not ( n375931 , n55571 );
not ( n375932 , n375931 );
not ( n55574 , n375932 );
not ( n375934 , n32202 );
or ( n375935 , n55574 , n375934 );
or ( n55577 , n32202 , n375932 );
nand ( n375937 , n375935 , n55577 );
not ( n55578 , n375937 );
nand ( n375939 , n366399 , n55578 );
buf ( n375940 , n375939 );
not ( n55581 , n351291 );
not ( n55582 , n55581 );
not ( n55583 , n342654 );
buf ( n375944 , n55583 );
not ( n55585 , n375944 );
or ( n55586 , n55582 , n55585 );
or ( n55587 , n55581 , n375944 );
nand ( n375948 , n55586 , n55587 );
buf ( n375949 , n375948 );
not ( n375950 , n375949 );
buf ( n375951 , n375950 );
buf ( n375952 , n375951 );
buf ( n375953 , n366428 );
nand ( n55594 , n375952 , n375953 );
buf ( n375955 , n55594 );
buf ( n375956 , n375955 );
and ( n55597 , n608 , n618 );
and ( n55598 , n610 , n616 );
xor ( n375959 , n55597 , n55598 );
and ( n375960 , n610 , n617 );
and ( n55601 , n612 , n615 );
xor ( n55602 , n375960 , n55601 );
and ( n375963 , n609 , n618 );
and ( n375964 , n55602 , n375963 );
and ( n55605 , n375960 , n55601 );
or ( n55606 , n375964 , n55605 );
and ( n55607 , n375959 , n55606 );
and ( n375968 , n55597 , n55598 );
or ( n375969 , n55607 , n375968 );
and ( n55610 , n612 , n614 );
and ( n55611 , n611 , n615 );
xor ( n55612 , n55610 , n55611 );
and ( n55613 , n609 , n617 );
and ( n55614 , n55612 , n55613 );
and ( n55615 , n55610 , n55611 );
or ( n55616 , n55614 , n55615 );
and ( n55617 , n612 , n613 );
xor ( n55618 , n612 , n55617 );
and ( n55619 , n610 , n615 );
xor ( n55620 , n55618 , n55619 );
xor ( n55621 , n55616 , n55620 );
and ( n55622 , n609 , n616 );
and ( n55623 , n611 , n614 );
xor ( n375984 , n55622 , n55623 );
and ( n55625 , n608 , n617 );
xor ( n55626 , n375984 , n55625 );
xor ( n55627 , n55621 , n55626 );
xor ( n375988 , n375969 , n55627 );
and ( n55629 , n613 , n614 );
xor ( n375990 , n613 , n55629 );
and ( n55631 , n611 , n616 );
and ( n55632 , n375990 , n55631 );
and ( n55633 , n613 , n55629 );
or ( n55634 , n55632 , n55633 );
xor ( n55635 , n55610 , n55611 );
xor ( n375996 , n55635 , n55613 );
xor ( n55637 , n55634 , n375996 );
and ( n375998 , n608 , n619 );
and ( n55639 , n613 , n615 );
and ( n55640 , n612 , n616 );
xor ( n376001 , n55639 , n55640 );
and ( n376002 , n610 , n618 );
and ( n55643 , n376001 , n376002 );
and ( n376004 , n55639 , n55640 );
or ( n376005 , n55643 , n376004 );
xor ( n55646 , n375998 , n376005 );
and ( n376007 , n609 , n619 );
and ( n376008 , n611 , n617 );
xor ( n376009 , n376007 , n376008 );
and ( n55650 , n608 , n620 );
and ( n376011 , n376009 , n55650 );
and ( n55652 , n376007 , n376008 );
or ( n376013 , n376011 , n55652 );
and ( n376014 , n55646 , n376013 );
and ( n55655 , n375998 , n376005 );
or ( n376016 , n376014 , n55655 );
and ( n55657 , n55637 , n376016 );
and ( n55658 , n55634 , n375996 );
or ( n55659 , n55657 , n55658 );
and ( n376020 , n375988 , n55659 );
and ( n55661 , n375969 , n55627 );
or ( n376022 , n376020 , n55661 );
and ( n55663 , n611 , n613 );
and ( n376024 , n610 , n614 );
xor ( n376025 , n55663 , n376024 );
and ( n55666 , n608 , n616 );
xor ( n376027 , n376025 , n55666 );
and ( n376028 , n609 , n615 );
xor ( n55669 , n612 , n55617 );
and ( n376030 , n55669 , n55619 );
and ( n376031 , n612 , n55617 );
or ( n55672 , n376030 , n376031 );
xor ( n376033 , n376028 , n55672 );
xor ( n55674 , n55622 , n55623 );
and ( n376035 , n55674 , n55625 );
and ( n55676 , n55622 , n55623 );
or ( n55677 , n376035 , n55676 );
xor ( n55678 , n376033 , n55677 );
xor ( n55679 , n376027 , n55678 );
xor ( n55680 , n55616 , n55620 );
and ( n376041 , n55680 , n55626 );
and ( n55682 , n55616 , n55620 );
or ( n376043 , n376041 , n55682 );
xor ( n55684 , n55679 , n376043 );
or ( n55685 , n376022 , n55684 );
xor ( n376046 , n376027 , n55678 );
and ( n376047 , n376046 , n376043 );
and ( n55688 , n376027 , n55678 );
or ( n376049 , n376047 , n55688 );
and ( n376050 , n611 , n612 );
xor ( n55691 , n611 , n376050 );
and ( n376052 , n609 , n614 );
xor ( n376053 , n55691 , n376052 );
and ( n376054 , n608 , n615 );
and ( n55695 , n610 , n613 );
xor ( n376056 , n376054 , n55695 );
xor ( n55697 , n55663 , n376024 );
and ( n55698 , n55697 , n55666 );
and ( n55699 , n55663 , n376024 );
or ( n55700 , n55698 , n55699 );
xor ( n55701 , n376056 , n55700 );
xor ( n55702 , n376053 , n55701 );
xor ( n55703 , n376028 , n55672 );
and ( n55704 , n55703 , n55677 );
and ( n55705 , n376028 , n55672 );
or ( n55706 , n55704 , n55705 );
xor ( n376067 , n55702 , n55706 );
nor ( n55708 , n376049 , n376067 );
xor ( n55709 , n376053 , n55701 );
and ( n55710 , n55709 , n55706 );
and ( n55711 , n376053 , n55701 );
or ( n55712 , n55710 , n55711 );
xor ( n55713 , n611 , n376050 );
and ( n55714 , n55713 , n376052 );
and ( n55715 , n611 , n376050 );
or ( n55716 , n55714 , n55715 );
and ( n55717 , n610 , n612 );
and ( n55718 , n609 , n613 );
xor ( n376079 , n55717 , n55718 );
and ( n55720 , n608 , n614 );
xor ( n376081 , n376079 , n55720 );
xor ( n376082 , n55716 , n376081 );
xor ( n55723 , n376054 , n55695 );
and ( n376084 , n55723 , n55700 );
and ( n55725 , n376054 , n55695 );
or ( n376086 , n376084 , n55725 );
xor ( n55727 , n376082 , n376086 );
nor ( n55728 , n55712 , n55727 );
nor ( n55729 , n55708 , n55728 );
xor ( n55730 , n55716 , n376081 );
and ( n55731 , n55730 , n376086 );
and ( n55732 , n55716 , n376081 );
or ( n376093 , n55731 , n55732 );
not ( n376094 , n376093 );
and ( n55735 , n609 , n612 );
xor ( n376096 , n55717 , n55718 );
and ( n55737 , n376096 , n55720 );
and ( n55738 , n55717 , n55718 );
or ( n55739 , n55737 , n55738 );
xor ( n55740 , n55735 , n55739 );
and ( n376101 , n610 , n611 );
xor ( n55742 , n610 , n376101 );
and ( n55743 , n608 , n613 );
xor ( n376104 , n55742 , n55743 );
xor ( n55745 , n55740 , n376104 );
not ( n55746 , n55745 );
nand ( n376107 , n376094 , n55746 );
xor ( n376108 , n55735 , n55739 );
and ( n55749 , n376108 , n376104 );
and ( n376110 , n55735 , n55739 );
or ( n376111 , n55749 , n376110 );
and ( n55752 , n609 , n611 );
and ( n376113 , n608 , n612 );
xor ( n376114 , n55752 , n376113 );
xor ( n55755 , n610 , n376101 );
and ( n376116 , n55755 , n55743 );
and ( n55757 , n610 , n376101 );
or ( n55758 , n376116 , n55757 );
xor ( n376119 , n376114 , n55758 );
or ( n376120 , n376111 , n376119 );
nand ( n55761 , n376107 , n376120 );
xor ( n376122 , n55752 , n376113 );
and ( n376123 , n376122 , n55758 );
and ( n55764 , n55752 , n376113 );
or ( n376125 , n376123 , n55764 );
not ( n55766 , n376125 );
and ( n55767 , n609 , n610 );
xor ( n55768 , n609 , n55767 );
and ( n376129 , n608 , n611 );
xor ( n55770 , n55768 , n376129 );
not ( n55771 , n55770 );
nand ( n55772 , n55766 , n55771 );
xor ( n376133 , n609 , n55767 );
and ( n55774 , n376133 , n376129 );
and ( n55775 , n609 , n55767 );
or ( n376136 , n55774 , n55775 );
not ( n55777 , n376136 );
nand ( n55778 , n608 , n610 );
nand ( n55779 , n55777 , n55778 );
nand ( n376140 , n55772 , n55779 , n608 );
nor ( n376141 , n55761 , n376140 );
and ( n55782 , n55685 , n55729 , n376141 );
not ( n376143 , n55782 );
xor ( n55784 , n55597 , n55598 );
xor ( n376145 , n55784 , n55606 );
xor ( n55786 , n55634 , n375996 );
xor ( n55787 , n55786 , n376016 );
xor ( n55788 , n376145 , n55787 );
xor ( n376149 , n375960 , n55601 );
xor ( n376150 , n376149 , n375963 );
xor ( n55791 , n613 , n55629 );
xor ( n55792 , n55791 , n55631 );
xor ( n55793 , n376150 , n55792 );
xor ( n376154 , n375998 , n376005 );
xor ( n376155 , n376154 , n376013 );
and ( n55796 , n55793 , n376155 );
and ( n55797 , n376150 , n55792 );
or ( n376158 , n55796 , n55797 );
xor ( n376159 , n55788 , n376158 );
and ( n55800 , n608 , n621 );
and ( n376161 , n611 , n618 );
xor ( n55802 , n55800 , n376161 );
and ( n376163 , n613 , n616 );
and ( n55804 , n55802 , n376163 );
and ( n55805 , n55800 , n376161 );
or ( n376166 , n55804 , n55805 );
and ( n55807 , n614 , n615 );
xor ( n376168 , n614 , n55807 );
and ( n55809 , n612 , n617 );
and ( n55810 , n376168 , n55809 );
and ( n376171 , n614 , n55807 );
or ( n55812 , n55810 , n376171 );
xor ( n376173 , n376166 , n55812 );
xor ( n376174 , n55639 , n55640 );
xor ( n376175 , n376174 , n376002 );
and ( n55816 , n376173 , n376175 );
and ( n376177 , n376166 , n55812 );
or ( n376178 , n55816 , n376177 );
xor ( n55819 , n376150 , n55792 );
xor ( n376180 , n55819 , n376155 );
xor ( n376181 , n376178 , n376180 );
xor ( n376182 , n376007 , n376008 );
xor ( n55823 , n376182 , n55650 );
and ( n376184 , n610 , n619 );
and ( n376185 , n609 , n620 );
xor ( n55826 , n376184 , n376185 );
and ( n376187 , n614 , n616 );
and ( n376188 , n613 , n617 );
xor ( n55829 , n376187 , n376188 );
and ( n55830 , n611 , n619 );
and ( n376191 , n55829 , n55830 );
and ( n376192 , n376187 , n376188 );
or ( n55833 , n376191 , n376192 );
and ( n55834 , n55826 , n55833 );
and ( n376195 , n376184 , n376185 );
or ( n376196 , n55834 , n376195 );
xor ( n55837 , n55823 , n376196 );
and ( n376198 , n610 , n620 );
and ( n55839 , n612 , n618 );
xor ( n55840 , n376198 , n55839 );
and ( n55841 , n609 , n621 );
and ( n376202 , n55840 , n55841 );
and ( n55843 , n376198 , n55839 );
or ( n376204 , n376202 , n55843 );
xor ( n55845 , n614 , n55807 );
xor ( n55846 , n55845 , n55809 );
xor ( n376207 , n376204 , n55846 );
xor ( n376208 , n55800 , n376161 );
xor ( n55849 , n376208 , n376163 );
and ( n376210 , n376207 , n55849 );
and ( n376211 , n376204 , n55846 );
or ( n55852 , n376210 , n376211 );
and ( n376213 , n55837 , n55852 );
and ( n376214 , n55823 , n376196 );
or ( n376215 , n376213 , n376214 );
and ( n376216 , n376181 , n376215 );
and ( n376217 , n376178 , n376180 );
or ( n376218 , n376216 , n376217 );
nor ( n376219 , n376159 , n376218 );
xor ( n376220 , n376145 , n55787 );
and ( n55856 , n376220 , n376158 );
and ( n376222 , n376145 , n55787 );
or ( n376223 , n55856 , n376222 );
xor ( n55859 , n375969 , n55627 );
xor ( n376225 , n55859 , n55659 );
nor ( n376226 , n376223 , n376225 );
nor ( n55862 , n376219 , n376226 );
not ( n376228 , n55862 );
xor ( n55864 , n376166 , n55812 );
xor ( n376230 , n55864 , n376175 );
xor ( n55866 , n55823 , n376196 );
xor ( n376232 , n55866 , n55852 );
xor ( n55868 , n376230 , n376232 );
xor ( n55869 , n376184 , n376185 );
xor ( n376235 , n55869 , n55833 );
and ( n376236 , n608 , n622 );
and ( n55872 , n615 , n616 );
and ( n376238 , n615 , n55872 );
xor ( n376239 , n376236 , n376238 );
and ( n55875 , n613 , n618 );
and ( n376241 , n609 , n622 );
xor ( n376242 , n55875 , n376241 );
and ( n55878 , n608 , n623 );
and ( n376244 , n376242 , n55878 );
and ( n55880 , n55875 , n376241 );
or ( n376246 , n376244 , n55880 );
and ( n376247 , n376239 , n376246 );
and ( n55883 , n376236 , n376238 );
or ( n55884 , n376247 , n55883 );
xor ( n376250 , n376235 , n55884 );
and ( n376251 , n612 , n619 );
and ( n55887 , n614 , n617 );
xor ( n376253 , n376251 , n55887 );
and ( n376254 , n611 , n620 );
and ( n55890 , n376253 , n376254 );
and ( n376256 , n376251 , n55887 );
or ( n376257 , n55890 , n376256 );
xor ( n55893 , n376198 , n55839 );
xor ( n376259 , n55893 , n55841 );
xor ( n55895 , n376257 , n376259 );
xor ( n55896 , n376187 , n376188 );
xor ( n376262 , n55896 , n55830 );
and ( n376263 , n55895 , n376262 );
and ( n55899 , n376257 , n376259 );
or ( n376265 , n376263 , n55899 );
and ( n376266 , n376250 , n376265 );
and ( n55902 , n376235 , n55884 );
or ( n376268 , n376266 , n55902 );
and ( n55904 , n55868 , n376268 );
and ( n55905 , n376230 , n376232 );
or ( n376271 , n55904 , n55905 );
xor ( n376272 , n376178 , n376180 );
xor ( n55908 , n376272 , n376215 );
or ( n376274 , n376271 , n55908 );
not ( n376275 , n376274 );
xor ( n55911 , n376230 , n376232 );
xor ( n376277 , n55911 , n376268 );
xor ( n55913 , n376204 , n55846 );
xor ( n55914 , n55913 , n55849 );
xor ( n55915 , n376235 , n55884 );
xor ( n376281 , n55915 , n376265 );
xor ( n376282 , n55914 , n376281 );
and ( n55918 , n610 , n621 );
xor ( n376284 , n615 , n55872 );
xor ( n55920 , n55918 , n376284 );
and ( n55921 , n614 , n618 );
and ( n55922 , n615 , n617 );
and ( n55923 , n55921 , n55922 );
and ( n376289 , n55920 , n55923 );
and ( n55925 , n55918 , n376284 );
or ( n55926 , n376289 , n55925 );
xor ( n55927 , n376236 , n376238 );
xor ( n376293 , n55927 , n376246 );
xor ( n376294 , n55926 , n376293 );
and ( n55930 , n612 , n620 );
and ( n376296 , n611 , n621 );
xor ( n376297 , n55930 , n376296 );
and ( n55933 , n613 , n619 );
and ( n55934 , n376297 , n55933 );
and ( n55935 , n55930 , n376296 );
or ( n55936 , n55934 , n55935 );
xor ( n55937 , n376251 , n55887 );
xor ( n55938 , n55937 , n376254 );
xor ( n55939 , n55936 , n55938 );
xor ( n55940 , n55875 , n376241 );
xor ( n55941 , n55940 , n55878 );
and ( n55942 , n55939 , n55941 );
and ( n55943 , n55936 , n55938 );
or ( n55944 , n55942 , n55943 );
and ( n376310 , n376294 , n55944 );
and ( n55946 , n55926 , n376293 );
or ( n376312 , n376310 , n55946 );
and ( n376313 , n376282 , n376312 );
and ( n55949 , n55914 , n376281 );
or ( n376315 , n376313 , n55949 );
nor ( n376316 , n376277 , n376315 );
nor ( n376317 , n376275 , n376316 );
not ( n55953 , n376317 );
xor ( n376319 , n55914 , n376281 );
xor ( n55955 , n376319 , n376312 );
xor ( n376321 , n376257 , n376259 );
xor ( n376322 , n376321 , n376262 );
and ( n55958 , n610 , n622 );
and ( n376324 , n609 , n623 );
xor ( n376325 , n55958 , n376324 );
xor ( n55961 , n55921 , n55922 );
and ( n376327 , n376325 , n55961 );
and ( n376328 , n55958 , n376324 );
or ( n55964 , n376327 , n376328 );
xor ( n376330 , n55918 , n376284 );
xor ( n376331 , n376330 , n55923 );
xor ( n55967 , n55964 , n376331 );
nand ( n55968 , n616 , n617 );
not ( n55969 , n55968 );
and ( n376335 , n614 , n619 );
and ( n376336 , n610 , n623 );
xor ( n55972 , n376335 , n376336 );
and ( n55973 , n613 , n620 );
and ( n376339 , n55972 , n55973 );
and ( n376340 , n376335 , n376336 );
or ( n55976 , n376339 , n376340 );
xor ( n55977 , n55969 , n55976 );
and ( n55978 , n615 , n618 );
and ( n55979 , n612 , n621 );
xor ( n55980 , n55978 , n55979 );
and ( n55981 , n611 , n622 );
and ( n55982 , n55980 , n55981 );
and ( n55983 , n55978 , n55979 );
or ( n55984 , n55982 , n55983 );
and ( n55985 , n55977 , n55984 );
and ( n55986 , n55969 , n55976 );
or ( n376352 , n55985 , n55986 );
and ( n55988 , n55967 , n376352 );
and ( n376354 , n55964 , n376331 );
or ( n376355 , n55988 , n376354 );
xor ( n55991 , n376322 , n376355 );
xor ( n55992 , n55926 , n376293 );
xor ( n55993 , n55992 , n55944 );
and ( n55994 , n55991 , n55993 );
and ( n55995 , n376322 , n376355 );
or ( n376361 , n55994 , n55995 );
nor ( n55997 , n55955 , n376361 );
xor ( n55998 , n376322 , n376355 );
xor ( n376364 , n55998 , n55993 );
xor ( n56000 , n55936 , n55938 );
xor ( n376366 , n56000 , n55941 );
xor ( n56002 , n55930 , n376296 );
xor ( n56003 , n56002 , n55933 );
xor ( n376369 , n55958 , n376324 );
xor ( n376370 , n376369 , n55961 );
xor ( n376371 , n56003 , n376370 );
and ( n376372 , n615 , n619 );
and ( n376373 , n616 , n618 );
and ( n376374 , n376372 , n376373 );
not ( n376375 , n616 );
not ( n376376 , n55968 );
or ( n376377 , n376375 , n376376 );
nand ( n376378 , n376377 , C1 );
xor ( n376379 , n376374 , n376378 );
and ( n376380 , n613 , n621 );
and ( n376381 , n612 , n622 );
xor ( n376382 , n376380 , n376381 );
and ( n376383 , n614 , n620 );
and ( n376384 , n376382 , n376383 );
and ( n376385 , n376380 , n376381 );
or ( n376386 , n376384 , n376385 );
and ( n376387 , n376379 , n376386 );
and ( n376388 , n376374 , n376378 );
or ( n376389 , n376387 , n376388 );
and ( n376390 , n376371 , n376389 );
and ( n376391 , n56003 , n376370 );
or ( n376392 , n376390 , n376391 );
xor ( n376393 , n376366 , n376392 );
xor ( n376394 , n55964 , n376331 );
xor ( n376395 , n376394 , n376352 );
and ( n376396 , n376393 , n376395 );
and ( n376397 , n376366 , n376392 );
or ( n376398 , n376396 , n376397 );
nor ( n376399 , n376364 , n376398 );
not ( n376400 , n376399 );
xor ( n376401 , n376366 , n376392 );
xor ( n376402 , n376401 , n376395 );
xor ( n376403 , n55969 , n55976 );
xor ( n376404 , n376403 , n55984 );
xor ( n56005 , n55978 , n55979 );
xor ( n56006 , n56005 , n55981 );
xor ( n56007 , n376335 , n376336 );
xor ( n376408 , n56007 , n55973 );
xor ( n376409 , n56006 , n376408 );
and ( n56010 , n611 , n623 );
xor ( n376411 , n376372 , n376373 );
xor ( n56012 , n56010 , n376411 );
and ( n376413 , n617 , n618 );
and ( n56014 , n617 , n376413 );
and ( n376415 , n56012 , n56014 );
and ( n56016 , n56010 , n376411 );
or ( n56017 , n376415 , n56016 );
and ( n56018 , n376409 , n56017 );
and ( n56019 , n56006 , n376408 );
or ( n56020 , n56018 , n56019 );
xor ( n56021 , n376404 , n56020 );
xor ( n56022 , n56003 , n376370 );
xor ( n56023 , n56022 , n376389 );
and ( n376424 , n56021 , n56023 );
and ( n376425 , n376404 , n56020 );
or ( n56026 , n376424 , n376425 );
or ( n376427 , n376402 , n56026 );
nand ( n56028 , n376400 , n376427 );
nor ( n56029 , n55997 , n56028 );
xor ( n376430 , n376404 , n56020 );
xor ( n376431 , n376430 , n56023 );
xor ( n56032 , n376374 , n376378 );
xor ( n376433 , n56032 , n376386 );
xor ( n376434 , n56006 , n376408 );
xor ( n56035 , n376434 , n56017 );
xor ( n376436 , n376433 , n56035 );
and ( n376437 , n615 , n620 );
and ( n56038 , n614 , n621 );
xor ( n376439 , n376437 , n56038 );
and ( n56040 , n616 , n619 );
and ( n56041 , n376439 , n56040 );
and ( n376442 , n376437 , n56038 );
or ( n376443 , n56041 , n376442 );
xor ( n56044 , n376380 , n376381 );
xor ( n376445 , n56044 , n376383 );
xor ( n376446 , n376443 , n376445 );
and ( n56047 , n613 , n622 );
and ( n376448 , n612 , n623 );
xor ( n56049 , n56047 , n376448 );
and ( n56050 , n616 , n620 );
and ( n56051 , n617 , n619 );
and ( n56052 , n56050 , n56051 );
and ( n56053 , n56049 , n56052 );
and ( n56054 , n56047 , n376448 );
or ( n56055 , n56053 , n56054 );
and ( n56056 , n376446 , n56055 );
and ( n56057 , n376443 , n376445 );
or ( n376458 , n56056 , n56057 );
and ( n56059 , n376436 , n376458 );
and ( n376460 , n376433 , n56035 );
or ( n376461 , n56059 , n376460 );
nor ( n56062 , n376431 , n376461 );
xor ( n376463 , n376433 , n56035 );
xor ( n376464 , n376463 , n376458 );
xor ( n56065 , n56010 , n376411 );
xor ( n376466 , n56065 , n56014 );
xor ( n376467 , n617 , n376413 );
and ( n56068 , n614 , n622 );
and ( n376469 , n613 , n623 );
xor ( n376470 , n56068 , n376469 );
and ( n56071 , n615 , n621 );
and ( n56072 , n376470 , n56071 );
and ( n56073 , n56068 , n376469 );
or ( n376474 , n56072 , n56073 );
xor ( n376475 , n376467 , n376474 );
xor ( n56076 , n376437 , n56038 );
xor ( n56077 , n56076 , n56040 );
and ( n56078 , n376475 , n56077 );
and ( n376479 , n376467 , n376474 );
or ( n376480 , n56078 , n376479 );
xor ( n56081 , n376466 , n376480 );
xor ( n56082 , n376443 , n376445 );
xor ( n376483 , n56082 , n56055 );
and ( n56084 , n56081 , n376483 );
and ( n376485 , n376466 , n376480 );
or ( n376486 , n56084 , n376485 );
nor ( n56087 , n376464 , n376486 );
nor ( n376488 , n56062 , n56087 );
not ( n56089 , n376488 );
xor ( n376490 , n376466 , n376480 );
xor ( n376491 , n376490 , n376483 );
xor ( n56092 , n56047 , n376448 );
xor ( n56093 , n56092 , n56052 );
xor ( n56094 , n56050 , n56051 );
and ( n56095 , n618 , n619 );
and ( n376496 , n618 , n56095 );
xor ( n56097 , n56094 , n376496 );
and ( n56098 , n616 , n621 );
and ( n376499 , n615 , n622 );
xor ( n56100 , n56098 , n376499 );
and ( n376501 , n617 , n620 );
and ( n376502 , n56100 , n376501 );
and ( n56103 , n56098 , n376499 );
or ( n56104 , n376502 , n56103 );
and ( n56105 , n56097 , n56104 );
and ( n56106 , n56094 , n376496 );
or ( n56107 , n56105 , n56106 );
xor ( n376508 , n56093 , n56107 );
xor ( n376509 , n376467 , n376474 );
xor ( n56110 , n376509 , n56077 );
and ( n376511 , n376508 , n56110 );
and ( n376512 , n56093 , n56107 );
or ( n56113 , n376511 , n376512 );
nor ( n376514 , n376491 , n56113 );
xor ( n376515 , n56093 , n56107 );
xor ( n376516 , n376515 , n56110 );
xor ( n56117 , n56068 , n376469 );
xor ( n376518 , n56117 , n56071 );
and ( n56119 , n614 , n623 );
xor ( n56120 , n618 , n56095 );
xor ( n56121 , n56119 , n56120 );
and ( n56122 , n617 , n621 );
and ( n56123 , n618 , n620 );
and ( n56124 , n56122 , n56123 );
and ( n56125 , n56121 , n56124 );
and ( n376526 , n56119 , n56120 );
or ( n376527 , n56125 , n376526 );
xor ( n56128 , n376518 , n376527 );
xor ( n376529 , n56094 , n376496 );
xor ( n376530 , n376529 , n56104 );
and ( n56131 , n56128 , n376530 );
and ( n376532 , n376518 , n376527 );
or ( n376533 , n56131 , n376532 );
nor ( n56134 , n376516 , n376533 );
nor ( n56135 , n376514 , n56134 );
not ( n56136 , n56135 );
xor ( n376537 , n376518 , n376527 );
xor ( n376538 , n376537 , n376530 );
xor ( n56139 , n56098 , n376499 );
xor ( n56140 , n56139 , n376501 );
and ( n56141 , n615 , n623 );
and ( n56142 , n616 , n622 );
xor ( n56143 , n56141 , n56142 );
and ( n376544 , n619 , n620 );
and ( n56145 , n619 , n376544 );
and ( n376546 , n56143 , n56145 );
and ( n376547 , n56141 , n56142 );
or ( n56148 , n376546 , n376547 );
xor ( n376549 , n56140 , n56148 );
xor ( n56150 , n56119 , n56120 );
xor ( n376551 , n56150 , n56124 );
and ( n56152 , n376549 , n376551 );
and ( n56153 , n56140 , n56148 );
or ( n376554 , n56152 , n56153 );
nor ( n376555 , n376538 , n376554 );
xor ( n56156 , n56140 , n56148 );
xor ( n376557 , n56156 , n376551 );
xor ( n376558 , n56122 , n56123 );
and ( n56159 , n617 , n622 );
and ( n376560 , n616 , n623 );
xor ( n376561 , n56159 , n376560 );
and ( n56162 , n618 , n621 );
and ( n376563 , n376561 , n56162 );
and ( n56164 , n56159 , n376560 );
or ( n56165 , n376563 , n56164 );
xor ( n376566 , n376558 , n56165 );
xor ( n376567 , n56141 , n56142 );
xor ( n56168 , n376567 , n56145 );
and ( n376569 , n376566 , n56168 );
and ( n376570 , n376558 , n56165 );
or ( n56171 , n376569 , n376570 );
nor ( n376572 , n376557 , n56171 );
nor ( n376573 , n376555 , n376572 );
not ( n56174 , n376573 );
xor ( n56175 , n619 , n376544 );
and ( n56176 , n618 , n622 );
and ( n376577 , n619 , n621 );
and ( n56178 , n56176 , n376577 );
xor ( n376579 , n56175 , n56178 );
xor ( n56180 , n56159 , n376560 );
xor ( n376581 , n56180 , n56162 );
and ( n56182 , n376579 , n376581 );
and ( n56183 , n56175 , n56178 );
or ( n376584 , n56182 , n56183 );
xor ( n56185 , n376558 , n56165 );
xor ( n376586 , n56185 , n56168 );
xor ( n56187 , n376584 , n376586 );
xor ( n56188 , n56175 , n56178 );
xor ( n376589 , n56188 , n376581 );
and ( n376590 , n617 , n623 );
xor ( n56191 , n56176 , n376577 );
xor ( n376592 , n376590 , n56191 );
nand ( n376593 , n620 , n621 );
not ( n56194 , n376593 );
and ( n376595 , n376592 , n56194 );
and ( n376596 , n376590 , n56191 );
or ( n376597 , n376595 , n376596 );
or ( n56198 , n376589 , n376597 );
not ( n56199 , n56198 );
xor ( n376600 , n376590 , n56191 );
xor ( n376601 , n376600 , n56194 );
and ( n56202 , n618 , n623 );
and ( n376603 , n619 , n622 );
xor ( n56204 , n56202 , n376603 );
not ( n56205 , n620 );
not ( n376606 , n376593 );
or ( n376607 , n56205 , n376606 );
nand ( n56208 , n376607 , C1 );
and ( n376609 , n56204 , n56208 );
and ( n376610 , n56202 , n376603 );
or ( n56211 , n376609 , n376610 );
or ( n376612 , n376601 , n56211 );
not ( n376613 , n376612 );
nand ( n56214 , n621 , n623 );
nand ( n376615 , n622 , n623 );
nor ( n56216 , n56214 , n376615 );
not ( n56217 , n56216 );
nand ( n376618 , n621 , n622 );
not ( n376619 , n376618 );
not ( n56220 , n621 );
nand ( n376621 , n620 , n623 );
not ( n376622 , n376621 );
or ( n56223 , n56220 , n376622 );
or ( n376624 , n376621 , n621 );
nand ( n56225 , n56223 , n376624 );
nand ( n56226 , n376619 , n56225 );
nand ( n56227 , n56217 , n56226 );
not ( n56228 , n56227 );
and ( n376629 , n619 , n623 );
not ( n376630 , n376629 );
nand ( n56231 , n620 , n622 );
not ( n376632 , n56231 );
and ( n376633 , n376630 , n376632 );
and ( n56234 , n376629 , n56231 );
nor ( n376635 , n376633 , n56234 );
nand ( n56236 , n56194 , n623 );
nand ( n56237 , n376635 , n56236 );
not ( n376638 , n56237 );
or ( n56239 , n56228 , n376638 );
or ( n376640 , n376635 , n56236 );
nand ( n376641 , n56239 , n376640 );
not ( n56242 , n376641 );
xor ( n56243 , n56202 , n376603 );
xor ( n376644 , n56243 , n56208 );
not ( n376645 , n376603 );
nor ( n56246 , n376645 , n376621 );
nor ( n376647 , n376644 , n56246 );
or ( n376648 , n56242 , n376647 );
nand ( n56249 , n376644 , n56246 );
nand ( n376650 , n376648 , n56249 );
not ( n376651 , n376650 );
or ( n56252 , n376613 , n376651 );
nand ( n376653 , n376601 , n56211 );
nand ( n376654 , n56252 , n376653 );
not ( n56255 , n376654 );
or ( n376656 , n56199 , n56255 );
nand ( n376657 , n376589 , n376597 );
nand ( n56258 , n376656 , n376657 );
and ( n56259 , n56187 , n56258 );
and ( n376660 , n376584 , n376586 );
or ( n376661 , n56259 , n376660 );
not ( n56262 , n376661 );
or ( n56263 , n56174 , n56262 );
not ( n376664 , n376555 );
nand ( n56265 , n376557 , n56171 );
not ( n376666 , n56265 );
and ( n376667 , n376664 , n376666 );
nand ( n56268 , n376538 , n376554 );
not ( n376669 , n56268 );
nor ( n56270 , n376667 , n376669 );
nand ( n56271 , n56263 , n56270 );
not ( n376672 , n56271 );
or ( n376673 , n56136 , n376672 );
not ( n56274 , n376514 );
nand ( n56275 , n376516 , n376533 );
not ( n376676 , n56275 );
and ( n376677 , n56274 , n376676 );
and ( n56278 , n376491 , n56113 );
nor ( n376679 , n376677 , n56278 );
nand ( n56280 , n376673 , n376679 );
not ( n56281 , n56280 );
or ( n376682 , n56089 , n56281 );
not ( n376683 , n56062 );
nand ( n56284 , n376464 , n376486 );
not ( n56285 , n56284 );
and ( n376686 , n376683 , n56285 );
nand ( n376687 , n376431 , n376461 );
not ( n56288 , n376687 );
nor ( n56289 , n376686 , n56288 );
nand ( n376690 , n376682 , n56289 );
nand ( n56291 , n56029 , n376690 );
nand ( n376692 , n376402 , n56026 );
or ( n56293 , n376399 , n376692 );
nand ( n56294 , n376364 , n376398 );
nand ( n376695 , n56293 , n56294 );
or ( n376696 , n55955 , n376361 );
nand ( n56297 , n376695 , n376696 );
nand ( n376698 , n55955 , n376361 );
nand ( n376699 , n56291 , n56297 , n376698 );
not ( n56300 , n376699 );
or ( n376701 , n55953 , n56300 );
not ( n376702 , n376274 );
and ( n56303 , n376277 , n376315 );
not ( n376704 , n56303 );
or ( n56305 , n376702 , n376704 );
nand ( n56306 , n376271 , n55908 );
nand ( n376707 , n56305 , n56306 );
not ( n376708 , n376707 );
nand ( n56309 , n376701 , n376708 );
not ( n376710 , n56309 );
or ( n376711 , n376228 , n376710 );
nand ( n56312 , n376159 , n376218 );
or ( n376713 , n56312 , n376226 );
nand ( n376714 , n376223 , n376225 );
nand ( n56315 , n376713 , n376714 );
not ( n376716 , n56315 );
nand ( n56317 , n376711 , n376716 );
not ( n56318 , n56317 );
or ( n56319 , n376143 , n56318 );
not ( n56320 , n55729 );
nand ( n56321 , n376022 , n55684 );
or ( n56322 , n56320 , n56321 );
nand ( n376723 , n376067 , n376049 );
or ( n376724 , n376723 , n55728 );
nand ( n376725 , n55712 , n55727 );
nand ( n376726 , n376724 , n376725 );
not ( n376727 , n376726 );
nand ( n376728 , n56322 , n376727 );
and ( n56324 , n376728 , n376141 );
nor ( n376730 , n376094 , n55746 );
and ( n376731 , n376730 , n376120 );
and ( n376732 , n376111 , n376119 );
nor ( n376733 , n376731 , n376732 );
or ( n376734 , n376733 , n376140 );
nor ( n376735 , n55766 , n55771 );
and ( n56326 , n376735 , n55779 );
nor ( n56327 , n55777 , n55778 );
nor ( n56328 , n56326 , n56327 , n609 );
not ( n56329 , n608 );
or ( n376740 , n56328 , n56329 );
nand ( n376741 , n376734 , n376740 );
nor ( n56332 , n56324 , n376741 );
nand ( n376743 , n56319 , n56332 );
buf ( n376744 , n376743 );
not ( n56335 , n580 );
nor ( n376746 , n56335 , n564 );
not ( n56337 , n581 );
nor ( n56338 , n56337 , n565 );
nor ( n376749 , n376746 , n56338 );
not ( n376750 , n566 );
nand ( n56341 , n376750 , n582 );
not ( n376752 , n56341 );
nor ( n376753 , n323556 , n567 );
nor ( n56344 , n376752 , n376753 );
and ( n376755 , n376749 , n56344 );
not ( n376756 , n562 );
nand ( n56347 , n376756 , n578 );
not ( n376758 , n563 );
nand ( n376759 , n376758 , n579 );
and ( n56350 , n56347 , n376759 );
not ( n376761 , n561 );
nand ( n56352 , n376761 , n577 );
and ( n56353 , n56350 , n56352 );
and ( n376764 , n376755 , n56353 );
not ( n56355 , n376764 );
not ( n376766 , n589 );
nand ( n56357 , n376766 , n573 );
not ( n376768 , n588 );
nand ( n376769 , n376768 , n572 );
and ( n56360 , n56357 , n376769 );
not ( n376771 , n56360 );
not ( n376772 , n573 );
nand ( n376773 , n376772 , n589 );
not ( n56364 , n376773 );
not ( n376775 , n56364 );
not ( n56366 , n574 );
nand ( n56367 , n56366 , n590 );
not ( n376778 , n575 );
nand ( n376779 , n376778 , n591 );
not ( n56370 , n376779 );
nand ( n376781 , n320740 , n574 );
nand ( n376782 , n56370 , n376781 );
nand ( n56373 , n376775 , n56367 , n376782 );
not ( n376784 , n56373 );
or ( n376785 , n376771 , n376784 );
not ( n56376 , n570 );
nand ( n376787 , n56376 , n586 );
not ( n56378 , n571 );
nand ( n56379 , n56378 , n587 );
nand ( n376790 , n376787 , n56379 );
not ( n56381 , n572 );
nand ( n376792 , n56381 , n588 );
not ( n56383 , n568 );
nand ( n376794 , n56383 , n584 );
not ( n376795 , n569 );
nand ( n56386 , n376795 , n585 );
nand ( n376797 , n376792 , n376794 , n56386 );
nor ( n376798 , n376790 , n376797 );
nand ( n56389 , n376785 , n376798 );
not ( n376800 , n571 );
nor ( n56391 , n376800 , n587 );
nand ( n56392 , n376787 , n56391 );
not ( n56393 , n56392 );
not ( n56394 , n586 );
nand ( n56395 , n56394 , n570 );
not ( n56396 , n584 );
nand ( n376807 , n56396 , n568 );
nand ( n56398 , n56395 , n376807 );
not ( n56399 , n569 );
nor ( n376810 , n56399 , n585 );
nor ( n376811 , n56398 , n376810 );
not ( n56402 , n376811 );
or ( n376813 , n56393 , n56402 );
not ( n376814 , n56386 );
not ( n56405 , n376794 );
or ( n376816 , n376814 , n56405 );
nand ( n376817 , n376816 , n376807 );
nand ( n56408 , n376813 , n376817 );
nand ( n56409 , n56389 , n56408 );
not ( n56410 , n56409 );
or ( n376821 , n56355 , n56410 );
not ( n56412 , n567 );
nor ( n56413 , n56412 , n583 );
not ( n376824 , n56413 );
not ( n56415 , n56341 );
or ( n56416 , n376824 , n56415 );
not ( n376827 , n582 );
nand ( n56418 , n376827 , n566 );
nand ( n376829 , n56416 , n56418 );
not ( n56420 , n376829 );
not ( n56421 , n376749 );
or ( n376832 , n56420 , n56421 );
not ( n376833 , n376746 );
not ( n56424 , n565 );
nor ( n376835 , n56424 , n581 );
and ( n376836 , n376833 , n376835 );
not ( n56427 , n564 );
nor ( n376838 , n56427 , n580 );
nor ( n376839 , n376836 , n376838 );
nand ( n56430 , n376832 , n376839 );
and ( n376841 , n56430 , n56353 );
not ( n56432 , n56352 );
not ( n56433 , n563 );
nor ( n56434 , n56433 , n579 );
not ( n376845 , n56434 );
not ( n56436 , n56347 );
or ( n376847 , n376845 , n56436 );
not ( n56438 , n578 );
nand ( n56439 , n56438 , n562 );
nand ( n56440 , n376847 , n56439 );
not ( n56441 , n56440 );
or ( n56442 , n56432 , n56441 );
not ( n376853 , n577 );
nand ( n56444 , n376853 , n561 );
nand ( n376855 , n56442 , n56444 );
nor ( n56446 , n376841 , n376855 );
nand ( n56447 , n376821 , n56446 );
not ( n376858 , n576 );
nor ( n376859 , n376858 , n560 );
not ( n56450 , n560 );
nor ( n376861 , n56450 , n576 );
nor ( n376862 , n376859 , n376861 );
xor ( n56453 , n56447 , n376862 );
buf ( n376864 , n56453 );
not ( n56455 , n376864 );
buf ( n376866 , n56455 );
buf ( n376867 , n376866 );
and ( n376868 , n376744 , n376867 );
buf ( n376869 , n376743 );
not ( n376870 , n376869 );
buf ( n376871 , n376870 );
buf ( n376872 , n376871 );
buf ( n376873 , n376866 );
not ( n56464 , n376873 );
buf ( n376875 , n56464 );
buf ( n376876 , n376875 );
and ( n56467 , n376872 , n376876 );
nor ( n376878 , n376868 , n56467 );
buf ( n376879 , n376878 );
buf ( n376880 , n376879 );
and ( n376881 , n376755 , n56350 );
not ( n376882 , n376881 );
not ( n56473 , n56409 );
or ( n376884 , n376882 , n56473 );
and ( n376885 , n56430 , n56350 );
nor ( n56476 , n376885 , n56440 );
nand ( n376887 , n376884 , n56476 );
nand ( n376888 , n56352 , n56444 );
xnor ( n376889 , n376887 , n376888 );
buf ( n376890 , n376889 );
and ( n376891 , n376755 , n376759 );
not ( n376892 , n376891 );
not ( n56483 , n56409 );
or ( n376894 , n376892 , n56483 );
and ( n376895 , n56430 , n376759 );
nor ( n56486 , n376895 , n56434 );
nand ( n376897 , n376894 , n56486 );
nand ( n56488 , n56347 , n56439 );
not ( n56489 , n56488 );
and ( n376900 , n376897 , n56489 );
not ( n56491 , n376897 );
and ( n376902 , n56491 , n56488 );
nor ( n376903 , n376900 , n376902 );
buf ( n376904 , n376903 );
xnor ( n56495 , n376890 , n376904 );
buf ( n376906 , n56495 );
buf ( n376907 , n376906 );
buf ( n376908 , n376889 );
not ( n376909 , n376908 );
buf ( n376910 , n376909 );
buf ( n376911 , n376910 );
buf ( n376912 , n376866 );
and ( n56503 , n376911 , n376912 );
buf ( n376914 , n376889 );
buf ( n376915 , n56453 );
and ( n56506 , n376914 , n376915 );
nor ( n376917 , n56503 , n56506 );
buf ( n376918 , n376917 );
buf ( n376919 , n376918 );
and ( n376920 , n376907 , n376919 );
buf ( n376921 , n376920 );
buf ( n376922 , n376921 );
not ( n376923 , n376922 );
buf ( n376924 , n376923 );
buf ( n376925 , n376924 );
or ( n376926 , n376880 , n376925 );
buf ( n56517 , n376906 );
buf ( n376928 , n56517 );
buf ( n376929 , n376866 );
nor ( n56520 , n376928 , n376929 );
buf ( n376931 , n56520 );
buf ( n376932 , n376931 );
not ( n376933 , n376932 );
buf ( n376934 , n376933 );
buf ( n376935 , n376934 );
nand ( n376936 , n376926 , n376935 );
buf ( n376937 , n376936 );
buf ( n376938 , n376937 );
nor ( n376939 , n56329 , n609 );
not ( n376940 , n55729 );
and ( n56531 , n376120 , n55772 );
nand ( n376942 , n56531 , n55779 );
not ( n376943 , n376107 );
nor ( n56534 , n376940 , n376942 , n376943 );
not ( n376945 , n56534 );
nand ( n376946 , n55862 , n55685 );
nor ( n56537 , n376945 , n376946 );
not ( n56538 , n56537 );
not ( n56539 , n56309 );
or ( n376950 , n56538 , n56539 );
not ( n376951 , n55685 );
not ( n56542 , n56315 );
or ( n376953 , n376951 , n56542 );
nand ( n56544 , n376953 , n56321 );
and ( n376955 , n56544 , n56534 );
and ( n376956 , n376726 , n376107 );
nor ( n56547 , n376956 , n376730 );
or ( n376958 , n56547 , n376942 );
and ( n376959 , n376732 , n55772 );
nor ( n56550 , n376959 , n376735 );
not ( n376961 , n56550 );
and ( n56552 , n376961 , n55779 );
nor ( n56553 , n56552 , n56327 );
nand ( n376964 , n376958 , n56553 );
nor ( n56555 , n376955 , n376964 );
nand ( n376966 , n376950 , n56555 );
not ( n56557 , n376966 );
and ( n376968 , n376939 , n56557 );
not ( n376969 , n376939 );
and ( n56560 , n376969 , n376966 );
or ( n376971 , n376968 , n56560 );
buf ( n376972 , n376971 );
not ( n56563 , n56352 );
nor ( n376974 , n56563 , n376859 );
and ( n56565 , n56350 , n376974 );
nand ( n56566 , n56409 , n376755 , n56565 );
and ( n56567 , n56430 , n56565 );
not ( n376978 , n376974 );
not ( n376979 , n56440 );
or ( n56570 , n376978 , n376979 );
not ( n376981 , n56444 );
not ( n376982 , n376859 );
and ( n56573 , n376981 , n376982 );
nor ( n376984 , n56573 , n376861 );
nand ( n376985 , n56570 , n376984 );
nor ( n56576 , n56567 , n376985 );
and ( n376987 , n56566 , n56576 );
buf ( n376988 , n376987 );
buf ( n56579 , n376988 );
buf ( n376990 , n56579 );
buf ( n376991 , n376990 );
and ( n56582 , n376972 , n376991 );
not ( n376993 , n376971 );
buf ( n376994 , n376993 );
buf ( n376995 , n376990 );
not ( n376996 , n376995 );
buf ( n376997 , n376996 );
buf ( n376998 , n376997 );
and ( n376999 , n376994 , n376998 );
buf ( n377000 , n56453 );
buf ( n377001 , n376987 );
xnor ( n377002 , n377000 , n377001 );
buf ( n377003 , n377002 );
buf ( n377004 , n377003 );
nor ( n377005 , n56582 , n376999 , n377004 );
buf ( n377006 , n377005 );
buf ( n377007 , n377006 );
or ( n377008 , n376938 , n377007 );
buf ( n377009 , n377008 );
buf ( n377010 , n377009 );
buf ( n377011 , n376871 );
buf ( n377012 , n376997 );
and ( n56603 , n377011 , n377012 );
buf ( n377014 , n376743 );
buf ( n377015 , n376990 );
and ( n56606 , n377014 , n377015 );
buf ( n377017 , n377003 );
nor ( n56608 , n56603 , n56606 , n377017 );
buf ( n377019 , n56608 );
buf ( n377020 , n377019 );
and ( n56611 , n377010 , n377020 );
buf ( n377022 , n377009 );
not ( n56613 , n377022 );
buf ( n377024 , n377019 );
not ( n377025 , n377024 );
and ( n377026 , n56613 , n377025 );
buf ( n377027 , n376921 );
buf ( n377028 , n376866 );
not ( n377029 , n377028 );
buf ( n377030 , n377029 );
buf ( n377031 , n377030 );
nand ( n56622 , n377027 , n377031 );
buf ( n56623 , n56622 );
buf ( n377034 , n56623 );
buf ( n377035 , n376934 );
nand ( n377036 , n377034 , n377035 );
buf ( n377037 , n377036 );
buf ( n377038 , n377037 );
nor ( n377039 , n377026 , n377038 );
buf ( n377040 , n377039 );
buf ( n377041 , n377040 );
nor ( n377042 , n56611 , n377041 );
buf ( n377043 , n377042 );
buf ( n377044 , n377043 );
not ( n377045 , n377044 );
buf ( n377046 , n377003 );
buf ( n377047 , n376997 );
nor ( n56638 , n377046 , n377047 );
buf ( n56639 , n56638 );
buf ( n56640 , n56639 );
not ( n56641 , n56640 );
buf ( n377052 , n56641 );
buf ( n377053 , n377052 );
nand ( n377054 , n377045 , n377053 );
buf ( n377055 , n377054 );
buf ( n377056 , n377055 );
nand ( n377057 , n375940 , n375956 , n377056 );
buf ( n377058 , n377057 );
buf ( n377059 , n377058 );
xor ( n377060 , n55567 , n377059 );
buf ( n377061 , n377060 );
buf ( n377062 , n377061 );
xor ( n377063 , n349135 , n349163 );
xor ( n56654 , n377063 , n349178 );
buf ( n377065 , n56654 );
buf ( n377066 , n377065 );
buf ( n377067 , n377066 );
buf ( n377068 , n377067 );
buf ( n377069 , n377068 );
not ( n377070 , n377069 );
buf ( n377071 , n377070 );
buf ( n377072 , n377071 );
not ( n56663 , n377072 );
buf ( n377074 , n359800 );
not ( n377075 , n377074 );
buf ( n377076 , n377075 );
buf ( n377077 , n377076 );
not ( n377078 , n377077 );
or ( n56669 , n56663 , n377078 );
buf ( n377080 , n359800 );
buf ( n377081 , n377068 );
nand ( n56672 , n377080 , n377081 );
buf ( n56673 , n56672 );
buf ( n377084 , n56673 );
nand ( n56675 , n56669 , n377084 );
buf ( n377086 , n56675 );
not ( n377087 , n377086 );
not ( n56678 , n359685 );
or ( n56679 , n377087 , n56678 );
and ( n56680 , n349152 , n349159 );
nor ( n377091 , n56680 , n349162 );
buf ( n377092 , n377091 );
buf ( n377093 , n377092 );
buf ( n377094 , n377093 );
buf ( n377095 , n377094 );
not ( n56686 , n377095 );
buf ( n56687 , n56686 );
buf ( n377098 , n56687 );
not ( n56689 , n377098 );
buf ( n377100 , n377076 );
not ( n377101 , n377100 );
or ( n56692 , n56689 , n377101 );
buf ( n377103 , n359800 );
buf ( n377104 , n377094 );
nand ( n56695 , n377103 , n377104 );
buf ( n377106 , n56695 );
buf ( n377107 , n377106 );
nand ( n377108 , n56692 , n377107 );
buf ( n377109 , n377108 );
nand ( n377110 , n377109 , n359804 , n39588 );
nand ( n377111 , n56679 , n377110 );
buf ( n377112 , n377111 );
xor ( n56703 , n377062 , n377112 );
or ( n377114 , n360038 , n39203 );
nand ( n56705 , n39203 , n360046 );
nand ( n377116 , n377114 , n56705 );
buf ( n56707 , n30931 );
buf ( n56708 , n56707 );
buf ( n377119 , n56708 );
buf ( n377120 , n377119 );
buf ( n56711 , n377120 );
buf ( n377122 , n56711 );
buf ( n377123 , n377122 );
buf ( n377124 , n360068 );
and ( n56715 , n377123 , n377124 );
not ( n56716 , n377123 );
buf ( n377127 , n365528 );
and ( n56718 , n56716 , n377127 );
nor ( n56719 , n56715 , n56718 );
buf ( n377130 , n56719 );
not ( n377131 , n377130 );
buf ( n377132 , n360164 );
nand ( n56723 , n377131 , n377132 );
and ( n377134 , n377116 , n56723 );
not ( n377135 , n377116 );
buf ( n377136 , n360065 );
not ( n56727 , n377136 );
buf ( n377138 , n350988 );
buf ( n377139 , n377138 );
buf ( n377140 , n377139 );
buf ( n377141 , n377140 );
buf ( n56732 , n377141 );
buf ( n377143 , n56732 );
buf ( n377144 , n377143 );
not ( n377145 , n377144 );
buf ( n377146 , n377145 );
buf ( n377147 , n377146 );
not ( n377148 , n377147 );
and ( n56739 , n56727 , n377148 );
buf ( n377150 , n363119 );
buf ( n56741 , n377143 );
not ( n377152 , n56741 );
buf ( n377153 , n377152 );
buf ( n377154 , n377153 );
and ( n56745 , n377150 , n377154 );
nor ( n377156 , n56739 , n56745 );
buf ( n377157 , n377156 );
and ( n56748 , n377135 , n377157 );
nor ( n377159 , n377134 , n56748 );
buf ( n377160 , n377159 );
xnor ( n377161 , n56703 , n377160 );
buf ( n377162 , n377161 );
buf ( n377163 , n377162 );
not ( n377164 , n377163 );
or ( n56755 , n375868 , n377164 );
buf ( n377166 , n366393 );
buf ( n377167 , n377166 );
buf ( n377168 , n377167 );
buf ( n377169 , n377168 );
not ( n377170 , n377169 );
buf ( n377171 , n377170 );
not ( n56762 , n377171 );
xor ( n377173 , n342654 , n352209 );
not ( n377174 , n377173 );
or ( n56765 , n56762 , n377174 );
buf ( n377176 , n50782 );
not ( n377177 , n377176 );
buf ( n377178 , n375951 );
nand ( n377179 , n377177 , n377178 );
buf ( n377180 , n377179 );
nand ( n377181 , n56765 , n377180 );
buf ( n377182 , n377181 );
not ( n56773 , n45553 );
not ( n56774 , n31072 );
xor ( n377185 , n365670 , n56774 );
not ( n377186 , n377185 );
or ( n56777 , n56773 , n377186 );
buf ( n377188 , n365670 );
not ( n56779 , n377188 );
buf ( n377190 , n56779 );
buf ( n377191 , n377190 );
not ( n56782 , n377191 );
buf ( n377193 , n364867 );
not ( n377194 , n377193 );
or ( n377195 , n56782 , n377194 );
buf ( n377196 , n365670 );
buf ( n377197 , n351364 );
nand ( n56788 , n377196 , n377197 );
buf ( n56789 , n56788 );
buf ( n377200 , n56789 );
nand ( n56791 , n377195 , n377200 );
buf ( n377202 , n56791 );
buf ( n56793 , n377202 );
buf ( n56794 , n45491 );
buf ( n377205 , n56794 );
nand ( n377206 , n56793 , n377205 );
buf ( n377207 , n377206 );
nand ( n56798 , n56777 , n377207 );
buf ( n377209 , n56798 );
xor ( n56800 , n377182 , n377209 );
and ( n377211 , n351229 , n342338 );
not ( n377212 , n351229 );
and ( n56803 , n377212 , n342335 );
or ( n377214 , n377211 , n56803 );
not ( n377215 , n377214 );
not ( n56806 , n48558 );
or ( n377217 , n377215 , n56806 );
and ( n377218 , n365490 , n342335 );
not ( n377219 , n365490 );
and ( n56810 , n377219 , n45592 );
nor ( n377221 , n377218 , n56810 );
not ( n377222 , n377221 );
not ( n377223 , n362383 );
not ( n56814 , n362392 );
or ( n377225 , n377223 , n56814 );
nand ( n377226 , n377225 , n362403 );
not ( n56817 , n377226 );
nand ( n377228 , n377222 , n56817 );
nand ( n377229 , n377217 , n377228 );
buf ( n377230 , n377229 );
xnor ( n377231 , n56800 , n377230 );
buf ( n377232 , n377231 );
buf ( n377233 , n377232 );
not ( n377234 , n375948 );
not ( n377235 , n377168 );
and ( n56826 , n377234 , n377235 );
nor ( n56827 , n50782 , n375937 );
nor ( n377238 , n56826 , n56827 );
or ( n377239 , n377238 , n377055 );
nand ( n377240 , n377239 , n377058 );
not ( n56831 , n377240 );
not ( n377242 , n56831 );
not ( n377243 , n377242 );
buf ( n377244 , n377052 );
not ( n56835 , n377244 );
buf ( n377246 , n377043 );
not ( n377247 , n377246 );
or ( n56838 , n56835 , n377247 );
buf ( n377249 , n377043 );
buf ( n377250 , n377052 );
or ( n377251 , n377249 , n377250 );
nand ( n377252 , n56838 , n377251 );
buf ( n377253 , n377252 );
buf ( n377254 , n377253 );
buf ( n377255 , n31231 );
buf ( n377256 , n375944 );
and ( n56847 , n377255 , n377256 );
not ( n56848 , n377255 );
buf ( n56849 , n342654 );
buf ( n377260 , n56849 );
and ( n56851 , n56848 , n377260 );
nor ( n377262 , n56847 , n56851 );
buf ( n377263 , n377262 );
or ( n56854 , n50782 , n377263 );
not ( n56855 , n375937 );
buf ( n377266 , n366425 );
not ( n377267 , n377266 );
buf ( n377268 , n377267 );
buf ( n377269 , n377268 );
not ( n377270 , n377269 );
buf ( n377271 , n377270 );
nand ( n56862 , n56855 , n377271 );
nand ( n377273 , n56854 , n56862 );
buf ( n377274 , n377273 );
xor ( n377275 , n377254 , n377274 );
buf ( n377276 , n352209 );
buf ( n377277 , n375901 );
not ( n377278 , n377277 );
buf ( n377279 , n377278 );
buf ( n377280 , n377279 );
and ( n56871 , n377276 , n377280 );
not ( n377282 , n377276 );
buf ( n377283 , n375901 );
and ( n377284 , n377282 , n377283 );
nor ( n56875 , n56871 , n377284 );
buf ( n377286 , n56875 );
buf ( n56877 , n377286 );
not ( n377288 , n56877 );
buf ( n377289 , n377288 );
buf ( n377290 , n377289 );
not ( n377291 , n377290 );
buf ( n377292 , n46463 );
not ( n377293 , n377292 );
or ( n377294 , n377291 , n377293 );
buf ( n377295 , n375901 );
not ( n56886 , n377295 );
not ( n377297 , n351290 );
buf ( n377298 , n377297 );
not ( n56889 , n377298 );
or ( n377300 , n56886 , n56889 );
not ( n377301 , n377297 );
buf ( n377302 , n377301 );
buf ( n377303 , n46474 );
nand ( n377304 , n377302 , n377303 );
buf ( n377305 , n377304 );
buf ( n377306 , n377305 );
nand ( n56897 , n377300 , n377306 );
buf ( n377308 , n56897 );
buf ( n377309 , n377308 );
buf ( n377310 , n46521 );
nand ( n377311 , n377309 , n377310 );
buf ( n377312 , n377311 );
buf ( n377313 , n377312 );
nand ( n377314 , n377294 , n377313 );
buf ( n377315 , n377314 );
buf ( n377316 , n377315 );
and ( n377317 , n377275 , n377316 );
and ( n377318 , n377254 , n377274 );
or ( n56909 , n377317 , n377318 );
buf ( n377320 , n56909 );
not ( n56911 , n377320 );
or ( n56912 , n377243 , n56911 );
not ( n56913 , n377320 );
not ( n377324 , n56913 );
not ( n56915 , n56831 );
or ( n56916 , n377324 , n56915 );
not ( n56917 , n365115 );
and ( n377328 , n30911 , n364978 );
not ( n377329 , n30911 );
and ( n56920 , n377329 , n364981 );
or ( n56921 , n377328 , n56920 );
not ( n377332 , n56921 );
or ( n56923 , n56917 , n377332 );
and ( n377334 , n364981 , n364867 );
not ( n377335 , n364981 );
and ( n377336 , n377335 , n351367 );
or ( n56927 , n377334 , n377336 );
buf ( n377338 , n56927 );
buf ( n377339 , n365033 );
nand ( n56930 , n377338 , n377339 );
buf ( n56931 , n56930 );
nand ( n377342 , n56923 , n56931 );
nand ( n377343 , n56916 , n377342 );
nand ( n56934 , n56912 , n377343 );
buf ( n377345 , n56934 );
xor ( n56936 , n377233 , n377345 );
buf ( n377347 , n352404 );
not ( n56938 , n377347 );
buf ( n377349 , n56938 );
buf ( n56940 , n377349 );
buf ( n377351 , n56940 );
buf ( n377352 , n377351 );
not ( n377353 , n377352 );
buf ( n377354 , n377353 );
not ( n56945 , n377354 );
buf ( n377356 , n366277 );
not ( n377357 , n377356 );
or ( n56948 , n56945 , n377357 );
buf ( n377359 , n362452 );
buf ( n377360 , n377352 );
nand ( n56951 , n377359 , n377360 );
buf ( n377362 , n56951 );
buf ( n377363 , n377362 );
nand ( n56954 , n56948 , n377363 );
buf ( n377365 , n56954 );
buf ( n377366 , n377365 );
not ( n56957 , n377366 );
buf ( n377368 , n40474 );
not ( n377369 , n377368 );
buf ( n377370 , n377369 );
buf ( n377371 , n377370 );
not ( n377372 , n377371 );
or ( n377373 , n56957 , n377372 );
not ( n56964 , n352368 );
not ( n377375 , n56964 );
not ( n377376 , n352364 );
not ( n56967 , n377376 );
or ( n377378 , n377375 , n56967 );
nand ( n377379 , n377378 , n352378 );
buf ( n56970 , n377379 );
buf ( n377381 , n56970 );
not ( n377382 , n377381 );
buf ( n377383 , n365468 );
not ( n377384 , n377383 );
or ( n56975 , n377382 , n377384 );
buf ( n377386 , n362452 );
buf ( n377387 , n56970 );
not ( n56978 , n377387 );
buf ( n377389 , n56978 );
buf ( n377390 , n377389 );
nand ( n377391 , n377386 , n377390 );
buf ( n377392 , n377391 );
buf ( n377393 , n377392 );
nand ( n56984 , n56975 , n377393 );
buf ( n377395 , n56984 );
buf ( n377396 , n377395 );
buf ( n377397 , n371732 );
nand ( n56988 , n377396 , n377397 );
buf ( n377399 , n56988 );
buf ( n377400 , n377399 );
nand ( n377401 , n377373 , n377400 );
buf ( n377402 , n377401 );
buf ( n377403 , n377402 );
xor ( n56994 , n56936 , n377403 );
buf ( n377405 , n56994 );
buf ( n377406 , n377405 );
nand ( n377407 , n56755 , n377406 );
buf ( n377408 , n377407 );
buf ( n377409 , n377408 );
buf ( n377410 , n55536 );
not ( n377411 , n377410 );
buf ( n377412 , n377411 );
buf ( n377413 , n377412 );
buf ( n377414 , n377162 );
not ( n57005 , n377414 );
buf ( n57006 , n57005 );
buf ( n377417 , n57006 );
nand ( n57008 , n377413 , n377417 );
buf ( n377419 , n57008 );
buf ( n377420 , n377419 );
nand ( n57011 , n377409 , n377420 );
buf ( n57012 , n57011 );
buf ( n377423 , n57012 );
buf ( n377424 , n361911 );
not ( n377425 , n377424 );
buf ( n377426 , n45336 );
not ( n57017 , n377426 );
and ( n377428 , n377425 , n57017 );
buf ( n377429 , n366329 );
buf ( n377430 , n45336 );
and ( n57021 , n377429 , n377430 );
nor ( n57022 , n377428 , n57021 );
buf ( n377433 , n57022 );
not ( n377434 , n377433 );
not ( n57025 , n377434 );
not ( n57026 , n368724 );
or ( n57027 , n57025 , n57026 );
buf ( n377438 , n351160 );
not ( n57029 , n377438 );
buf ( n377440 , n364763 );
not ( n57031 , n377440 );
or ( n57032 , n57029 , n57031 );
nand ( n377443 , n361591 , n364915 );
buf ( n377444 , n377443 );
nand ( n57035 , n57032 , n377444 );
buf ( n377446 , n57035 );
nand ( n57037 , n366339 , n377446 , n361967 , n41807 );
nand ( n57038 , n57027 , n57037 );
buf ( n377449 , n57038 );
buf ( n377450 , n364821 );
xor ( n57041 , n365422 , n40860 );
xnor ( n377452 , n57041 , n40866 );
buf ( n377453 , n377452 );
or ( n57044 , n377450 , n377453 );
buf ( n377455 , n365619 );
buf ( n377456 , n365393 );
not ( n377457 , n377456 );
buf ( n377458 , n364832 );
not ( n377459 , n377458 );
or ( n377460 , n377457 , n377459 );
buf ( n377461 , n45455 );
buf ( n377462 , n365408 );
nand ( n377463 , n377461 , n377462 );
buf ( n377464 , n377463 );
buf ( n377465 , n377464 );
nand ( n377466 , n377460 , n377465 );
buf ( n377467 , n377466 );
buf ( n377468 , n377467 );
buf ( n377469 , n362020 );
nand ( n377470 , n377455 , n377468 , n377469 );
buf ( n377471 , n377470 );
buf ( n377472 , n377471 );
nand ( n377473 , n57044 , n377472 );
buf ( n377474 , n377473 );
buf ( n377475 , n377474 );
xor ( n377476 , n377449 , n377475 );
buf ( n377477 , n368994 );
not ( n377478 , n377477 );
buf ( n377479 , n365267 );
not ( n377480 , n377479 );
or ( n57051 , n377478 , n377480 );
buf ( n377482 , n365293 );
buf ( n57053 , n48791 );
buf ( n377484 , n57053 );
nand ( n377485 , n377482 , n377484 );
buf ( n377486 , n377485 );
buf ( n377487 , n377486 );
nand ( n377488 , n57051 , n377487 );
buf ( n377489 , n377488 );
buf ( n377490 , n377489 );
not ( n377491 , n377490 );
buf ( n377492 , n361013 );
not ( n57063 , n377492 );
or ( n377494 , n377491 , n57063 );
buf ( n377495 , n365303 );
and ( n377496 , n40891 , n368665 );
not ( n57067 , n40891 );
and ( n57068 , n57067 , n368662 );
or ( n377499 , n377496 , n57068 );
buf ( n377500 , n377499 );
nand ( n377501 , n377495 , n377500 );
buf ( n377502 , n377501 );
buf ( n377503 , n377502 );
nand ( n377504 , n377494 , n377503 );
buf ( n377505 , n377504 );
buf ( n377506 , n377505 );
xor ( n377507 , n377476 , n377506 );
buf ( n377508 , n377507 );
buf ( n377509 , n377508 );
xor ( n377510 , n375893 , n375925 );
and ( n377511 , n377510 , n377059 );
and ( n57082 , n375893 , n375925 );
or ( n377513 , n377511 , n57082 );
buf ( n377514 , n377513 );
not ( n377515 , n365115 );
not ( n57086 , n364981 );
not ( n377517 , n366077 );
or ( n377518 , n57086 , n377517 );
buf ( n377519 , n42355 );
buf ( n377520 , n364978 );
nand ( n377521 , n377519 , n377520 );
buf ( n377522 , n377521 );
nand ( n377523 , n377518 , n377522 );
not ( n57093 , n377523 );
or ( n377525 , n377515 , n57093 );
or ( n377526 , n364978 , n351762 );
nand ( n57096 , n364978 , n351762 );
nand ( n377528 , n377526 , n57096 );
buf ( n377529 , n377528 );
buf ( n377530 , n365033 );
nand ( n57100 , n377529 , n377530 );
buf ( n57101 , n57100 );
nand ( n377533 , n377525 , n57101 );
xor ( n57103 , n377514 , n377533 );
and ( n57104 , n46303 , n366086 );
not ( n377536 , n46303 );
and ( n377537 , n377536 , n45908 );
or ( n57107 , n57104 , n377537 );
not ( n377539 , n57107 );
not ( n377540 , n366518 );
or ( n57110 , n377539 , n377540 );
buf ( n377542 , n365980 );
not ( n57112 , n377542 );
buf ( n377544 , n44717 );
not ( n57114 , n377544 );
or ( n57115 , n57112 , n57114 );
buf ( n377547 , n45414 );
buf ( n377548 , n365989 );
nand ( n57118 , n377547 , n377548 );
buf ( n377550 , n57118 );
buf ( n377551 , n377550 );
nand ( n57121 , n57115 , n377551 );
buf ( n377553 , n57121 );
nand ( n57123 , n369589 , n377553 );
nand ( n377555 , n57110 , n57123 );
xor ( n377556 , n57103 , n377555 );
buf ( n377557 , n377556 );
xor ( n57127 , n377509 , n377557 );
xor ( n377559 , n377233 , n377345 );
and ( n377560 , n377559 , n377403 );
and ( n57130 , n377233 , n377345 );
or ( n57131 , n377560 , n57130 );
buf ( n377563 , n57131 );
buf ( n377564 , n377563 );
xor ( n377565 , n57127 , n377564 );
buf ( n377566 , n377565 );
buf ( n377567 , n377566 );
xor ( n57137 , n377423 , n377567 );
buf ( n377569 , n23104 );
buf ( n377570 , n377569 );
buf ( n377571 , n377570 );
and ( n57141 , n342385 , n377571 );
not ( n377573 , n342385 );
buf ( n377574 , n377571 );
not ( n57144 , n377574 );
buf ( n57145 , n57144 );
and ( n57146 , n377573 , n57145 );
or ( n57147 , n57141 , n57146 );
not ( n377579 , n57147 );
buf ( n377580 , n377579 );
buf ( n377581 , n377580 );
not ( n377582 , n377581 );
buf ( n377583 , n49579 );
buf ( n377584 , n377583 );
buf ( n377585 , n377584 );
buf ( n377586 , n377585 );
not ( n377587 , n377586 );
buf ( n377588 , n366725 );
not ( n377589 , n377588 );
or ( n377590 , n377587 , n377589 );
buf ( n377591 , n366722 );
not ( n377592 , n377584 );
buf ( n377593 , n377592 );
nand ( n377594 , n377591 , n377593 );
buf ( n377595 , n377594 );
buf ( n377596 , n377595 );
nand ( n57150 , n377590 , n377596 );
buf ( n377598 , n57150 );
buf ( n377599 , n377598 );
not ( n57153 , n377599 );
or ( n57154 , n377582 , n57153 );
not ( n57155 , n377579 );
buf ( n57156 , n342385 );
buf ( n57157 , n57156 );
buf ( n57158 , n57157 );
buf ( n377606 , n57158 );
buf ( n377607 , n343039 );
and ( n57161 , n377606 , n377607 );
not ( n57162 , n377606 );
buf ( n377610 , n343039 );
not ( n377611 , n377610 );
buf ( n377612 , n377611 );
buf ( n377613 , n377612 );
and ( n57167 , n57162 , n377613 );
nor ( n377615 , n57161 , n57167 );
buf ( n377616 , n377615 );
nand ( n57170 , n57155 , n377616 );
buf ( n377618 , n57170 );
buf ( n377619 , n377618 );
not ( n57173 , n377619 );
not ( n377621 , n377585 );
not ( n377622 , n369022 );
or ( n57176 , n377621 , n377622 );
nand ( n377624 , n40251 , n377592 );
nand ( n377625 , n57176 , n377624 );
buf ( n377626 , n377625 );
nand ( n377627 , n57173 , n377626 );
buf ( n377628 , n377627 );
buf ( n377629 , n377628 );
nand ( n57183 , n57154 , n377629 );
buf ( n377631 , n57183 );
not ( n377632 , n377631 );
buf ( n377633 , n369444 );
not ( n377634 , n377633 );
buf ( n377635 , n368554 );
buf ( n377636 , n362288 );
and ( n377637 , n377635 , n377636 );
not ( n377638 , n377635 );
buf ( n377639 , n362285 );
and ( n377640 , n377638 , n377639 );
nor ( n57194 , n377637 , n377640 );
buf ( n377642 , n57194 );
buf ( n377643 , n377642 );
not ( n57197 , n377643 );
or ( n377645 , n377634 , n57197 );
buf ( n377646 , n368611 );
buf ( n377647 , n368549 );
not ( n377648 , n377647 );
buf ( n377649 , n45718 );
not ( n57203 , n377649 );
or ( n377651 , n377648 , n57203 );
buf ( n377652 , n362133 );
buf ( n377653 , n368554 );
nand ( n377654 , n377652 , n377653 );
buf ( n377655 , n377654 );
buf ( n377656 , n377655 );
nand ( n57210 , n377651 , n377656 );
buf ( n377658 , n57210 );
buf ( n377659 , n377658 );
nand ( n57213 , n377646 , n377659 );
buf ( n377661 , n57213 );
buf ( n377662 , n377661 );
nand ( n377663 , n377645 , n377662 );
buf ( n377664 , n377663 );
not ( n377665 , n377664 );
or ( n57219 , n377632 , n377665 );
not ( n377667 , n377664 );
not ( n57221 , n377667 );
buf ( n377669 , n377631 );
not ( n57223 , n377669 );
buf ( n377671 , n57223 );
not ( n377672 , n377671 );
or ( n57226 , n57221 , n377672 );
buf ( n377674 , n375878 );
not ( n57228 , n363416 );
buf ( n377676 , n57228 );
nand ( n57230 , n377674 , n377676 );
buf ( n377678 , n57230 );
not ( n57232 , n377678 );
not ( n57233 , n31194 );
buf ( n57234 , n57233 );
not ( n57235 , n57234 );
not ( n377683 , n55539 );
buf ( n377684 , n377683 );
not ( n377685 , n377684 );
or ( n377686 , n57235 , n377685 );
buf ( n377687 , n22769 );
buf ( n377688 , n351228 );
nand ( n57242 , n377687 , n377688 );
buf ( n377690 , n57242 );
buf ( n377691 , n377690 );
nand ( n377692 , n377686 , n377691 );
buf ( n377693 , n377692 );
and ( n377694 , n377693 , n363428 );
nor ( n57248 , n57232 , n377694 );
buf ( n377696 , n57248 );
not ( n57250 , n377286 );
not ( n57251 , n366708 );
and ( n377699 , n57250 , n57251 );
and ( n377700 , n375905 , n46463 );
nor ( n57254 , n377699 , n377700 );
buf ( n377702 , n57254 );
xor ( n377703 , n377696 , n377702 );
not ( n57257 , n377221 );
not ( n377705 , n362385 );
and ( n57259 , n57257 , n377705 );
not ( n57260 , n368765 );
not ( n57261 , n364915 );
and ( n377709 , n57260 , n57261 );
buf ( n377710 , n342335 );
not ( n377711 , n377710 );
buf ( n377712 , n377711 );
buf ( n377713 , n377712 );
not ( n57267 , n377713 );
buf ( n377715 , n57267 );
and ( n57269 , n377715 , n364915 );
nor ( n57270 , n377709 , n57269 );
not ( n377718 , n57270 );
nor ( n377719 , n377718 , n48502 );
nor ( n57273 , n57259 , n377719 );
buf ( n377721 , n57273 );
and ( n377722 , n377703 , n377721 );
and ( n57276 , n377696 , n377702 );
or ( n57277 , n377722 , n57276 );
buf ( n377725 , n57277 );
not ( n377726 , n45018 );
not ( n57280 , n22956 );
not ( n377728 , n57280 );
or ( n377729 , n41569 , n377728 );
nand ( n57283 , n41569 , n377728 );
nand ( n377731 , n377729 , n57283 );
not ( n377732 , n377731 );
or ( n57286 , n377726 , n377732 );
buf ( n377734 , n57280 );
not ( n377735 , n377734 );
buf ( n377736 , n361664 );
not ( n377737 , n377736 );
or ( n57291 , n377735 , n377737 );
buf ( n377739 , n372889 );
buf ( n377740 , n377728 );
nand ( n377741 , n377739 , n377740 );
buf ( n377742 , n377741 );
buf ( n377743 , n377742 );
nand ( n57297 , n57291 , n377743 );
buf ( n377745 , n57297 );
buf ( n57299 , n377745 );
buf ( n57300 , n365152 );
nand ( n57301 , n57299 , n57300 );
buf ( n57302 , n57301 );
nand ( n377750 , n57286 , n57302 );
xor ( n57304 , n377725 , n377750 );
buf ( n377752 , n351013 );
buf ( n57306 , n377752 );
buf ( n377754 , n57306 );
buf ( n377755 , n377754 );
buf ( n57309 , n377755 );
buf ( n377757 , n57309 );
buf ( n377758 , n377757 );
buf ( n377759 , n359297 );
and ( n377760 , n377758 , n377759 );
not ( n57314 , n377758 );
buf ( n377762 , n365367 );
and ( n57316 , n57314 , n377762 );
nor ( n57317 , n377760 , n57316 );
buf ( n377765 , n57317 );
buf ( n377766 , n377765 );
not ( n57320 , n377766 );
buf ( n57321 , n57320 );
buf ( n377769 , n57321 );
not ( n57323 , n377769 );
buf ( n377771 , n366989 );
not ( n57325 , n377771 );
or ( n57326 , n57323 , n57325 );
buf ( n377774 , n351027 );
not ( n57328 , n377774 );
buf ( n377776 , n57328 );
buf ( n377777 , n377776 );
buf ( n377778 , n377777 );
buf ( n377779 , n377778 );
buf ( n377780 , n377779 );
not ( n57334 , n377780 );
buf ( n377782 , n57334 );
and ( n57336 , n377782 , n355579 );
not ( n377784 , n377782 );
and ( n57338 , n377784 , n365367 );
nor ( n57339 , n57336 , n57338 );
not ( n377787 , n57339 );
nand ( n377788 , n377787 , n359312 );
buf ( n377789 , n377788 );
nand ( n377790 , n57326 , n377789 );
buf ( n377791 , n377790 );
xor ( n57345 , n57304 , n377791 );
buf ( n377793 , n57345 );
not ( n377794 , n377793 );
buf ( n377795 , n377794 );
nand ( n377796 , n57226 , n377795 );
nand ( n57350 , n57219 , n377796 );
buf ( n377798 , n57350 );
not ( n377799 , n377798 );
buf ( n377800 , n377799 );
buf ( n377801 , n377800 );
xor ( n377802 , n57137 , n377801 );
buf ( n377803 , n377802 );
buf ( n377804 , n57006 );
buf ( n377805 , n377412 );
xor ( n57359 , n377804 , n377805 );
buf ( n377807 , n377405 );
xnor ( n57361 , n57359 , n377807 );
buf ( n377809 , n57361 );
not ( n377810 , n377809 );
buf ( n377811 , n377810 );
not ( n377812 , n377811 );
xor ( n57366 , n377667 , n57345 );
and ( n57367 , n57366 , n377671 );
not ( n377815 , n57366 );
and ( n377816 , n377815 , n377631 );
nor ( n57370 , n57367 , n377816 );
not ( n57371 , n57370 );
buf ( n377819 , n57371 );
not ( n57373 , n377819 );
or ( n57374 , n377812 , n57373 );
buf ( n377822 , n57370 );
not ( n57376 , n377822 );
buf ( n377824 , n377809 );
not ( n377825 , n377824 );
or ( n57379 , n57376 , n377825 );
buf ( n377827 , n342335 );
not ( n57381 , n377827 );
buf ( n377829 , n352268 );
not ( n57383 , n377829 );
or ( n377831 , n57381 , n57383 );
buf ( n377832 , n362417 );
buf ( n377833 , n44737 );
nand ( n377834 , n377832 , n377833 );
buf ( n377835 , n377834 );
buf ( n377836 , n377835 );
nand ( n377837 , n377831 , n377836 );
buf ( n377838 , n377837 );
not ( n377839 , n377838 );
not ( n377840 , n362405 );
or ( n57394 , n377839 , n377840 );
not ( n377842 , n362385 );
nand ( n57396 , n57270 , n377842 );
nand ( n57397 , n57394 , n57396 );
buf ( n377845 , n57397 );
buf ( n377846 , n365033 );
not ( n57400 , n377846 );
buf ( n377848 , n364981 );
not ( n377849 , n377848 );
buf ( n377850 , n367575 );
not ( n377851 , n377850 );
or ( n377852 , n377849 , n377851 );
buf ( n377853 , n31072 );
buf ( n377854 , n364978 );
nand ( n377855 , n377853 , n377854 );
buf ( n377856 , n377855 );
buf ( n377857 , n377856 );
nand ( n57411 , n377852 , n377857 );
buf ( n377859 , n57411 );
buf ( n377860 , n377859 );
not ( n57414 , n377860 );
or ( n377862 , n57400 , n57414 );
buf ( n377863 , n56927 );
buf ( n377864 , n365115 );
nand ( n57418 , n377863 , n377864 );
buf ( n377866 , n57418 );
buf ( n377867 , n377866 );
nand ( n57421 , n377862 , n377867 );
buf ( n377869 , n57421 );
buf ( n377870 , n377869 );
xor ( n57424 , n377845 , n377870 );
buf ( n377872 , n365226 );
not ( n377873 , n377872 );
and ( n57427 , n342881 , n365328 );
not ( n377875 , n342881 );
and ( n57429 , n377875 , n30911 );
or ( n57430 , n57427 , n57429 );
buf ( n377878 , n57430 );
not ( n57432 , n377878 );
or ( n57433 , n377873 , n57432 );
buf ( n377881 , n45075 );
buf ( n377882 , n342881 );
not ( n57436 , n377882 );
buf ( n377884 , n48496 );
not ( n57438 , n377884 );
or ( n57439 , n57436 , n57438 );
not ( n57440 , n342881 );
nand ( n57441 , n57440 , n368700 );
buf ( n377889 , n57441 );
nand ( n57443 , n57439 , n377889 );
buf ( n377891 , n57443 );
buf ( n377892 , n377891 );
nand ( n377893 , n377881 , n377892 );
buf ( n377894 , n377893 );
buf ( n377895 , n377894 );
nand ( n57449 , n57433 , n377895 );
buf ( n377897 , n57449 );
buf ( n377898 , n377897 );
xor ( n377899 , n57424 , n377898 );
buf ( n377900 , n377899 );
buf ( n377901 , n377900 );
buf ( n377902 , n377122 );
not ( n57456 , n377902 );
buf ( n377904 , n365368 );
not ( n57458 , n377904 );
or ( n57459 , n57456 , n57458 );
buf ( n377907 , n366360 );
buf ( n57461 , n377122 );
not ( n57462 , n57461 );
buf ( n57463 , n57462 );
buf ( n377911 , n57463 );
nand ( n57465 , n377907 , n377911 );
buf ( n377913 , n57465 );
buf ( n377914 , n377913 );
nand ( n57468 , n57459 , n377914 );
buf ( n377916 , n57468 );
buf ( n377917 , n377916 );
not ( n57471 , n377917 );
buf ( n377919 , n39208 );
not ( n377920 , n377919 );
or ( n57474 , n57471 , n377920 );
buf ( n377922 , n46582 );
buf ( n377923 , n377143 );
not ( n57477 , n377923 );
buf ( n377925 , n365368 );
not ( n377926 , n377925 );
or ( n377927 , n57477 , n377926 );
not ( n57481 , n359297 );
buf ( n377929 , n57481 );
buf ( n377930 , n377153 );
nand ( n57484 , n377929 , n377930 );
buf ( n377932 , n57484 );
buf ( n377933 , n377932 );
nand ( n377934 , n377927 , n377933 );
buf ( n377935 , n377934 );
buf ( n377936 , n377935 );
nand ( n377937 , n377922 , n377936 );
buf ( n377938 , n377937 );
buf ( n377939 , n377938 );
nand ( n377940 , n57474 , n377939 );
buf ( n377941 , n377940 );
buf ( n377942 , n377941 );
xor ( n377943 , n377901 , n377942 );
buf ( n377944 , n47466 );
not ( n377945 , n377944 );
buf ( n377946 , n365052 );
buf ( n377947 , n363546 );
and ( n377948 , n377946 , n377947 );
not ( n57485 , n377946 );
buf ( n377950 , n361716 );
and ( n57487 , n57485 , n377950 );
nor ( n377952 , n377948 , n57487 );
buf ( n377953 , n377952 );
buf ( n377954 , n377953 );
not ( n57489 , n377954 );
or ( n57490 , n377945 , n57489 );
buf ( n377957 , n365041 );
not ( n57492 , n377957 );
buf ( n377959 , n41528 );
not ( n57494 , n377959 );
buf ( n377961 , n57494 );
buf ( n377962 , n377961 );
not ( n57497 , n377962 );
or ( n57498 , n57492 , n57497 );
buf ( n377965 , n41528 );
buf ( n377966 , n365052 );
nand ( n377967 , n377965 , n377966 );
buf ( n377968 , n377967 );
buf ( n377969 , n377968 );
nand ( n57504 , n57498 , n377969 );
buf ( n377971 , n57504 );
buf ( n377972 , n377971 );
buf ( n377973 , n44915 );
nand ( n377974 , n377972 , n377973 );
buf ( n377975 , n377974 );
buf ( n377976 , n377975 );
nand ( n57511 , n57490 , n377976 );
buf ( n377978 , n57511 );
buf ( n377979 , n377978 );
and ( n377980 , n377943 , n377979 );
and ( n57515 , n377901 , n377942 );
or ( n57516 , n377980 , n57515 );
buf ( n377983 , n57516 );
not ( n377984 , n377983 );
not ( n377985 , n377585 );
not ( n57520 , n366673 );
or ( n377987 , n377985 , n57520 );
buf ( n377988 , n360848 );
not ( n57523 , n377988 );
buf ( n377990 , n57523 );
buf ( n377991 , n377990 );
buf ( n377992 , n377592 );
nand ( n57527 , n377991 , n377992 );
buf ( n377994 , n57527 );
nand ( n57529 , n377987 , n377994 );
not ( n57530 , n377618 );
and ( n377997 , n57529 , n57530 );
and ( n57532 , n377625 , n377580 );
nor ( n57533 , n377997 , n57532 );
buf ( n378000 , n57533 );
not ( n57535 , n378000 );
buf ( n378002 , n57535 );
not ( n378003 , n378002 );
or ( n57538 , n377984 , n378003 );
not ( n378005 , n57533 );
buf ( n378006 , n377983 );
not ( n57541 , n378006 );
buf ( n378008 , n57541 );
not ( n378009 , n378008 );
or ( n57544 , n378005 , n378009 );
buf ( n378011 , n57430 );
buf ( n378012 , n45075 );
and ( n57547 , n378011 , n378012 );
xor ( n378014 , n342881 , n351364 );
buf ( n378015 , n378014 );
not ( n57550 , n378015 );
buf ( n378017 , n365227 );
nor ( n57552 , n57550 , n378017 );
buf ( n378019 , n57552 );
buf ( n378020 , n378019 );
nor ( n378021 , n57547 , n378020 );
buf ( n378022 , n378021 );
buf ( n378023 , n378022 );
not ( n378024 , n378023 );
buf ( n378025 , n378024 );
buf ( n378026 , n378025 );
not ( n57561 , n378026 );
buf ( n57562 , n361971 );
not ( n57563 , n57562 );
buf ( n378030 , n364763 );
buf ( n57565 , n378030 );
buf ( n378032 , n57565 );
and ( n378033 , n365408 , n378032 );
not ( n378034 , n365408 );
and ( n57569 , n378034 , n366329 );
or ( n378036 , n378033 , n57569 );
buf ( n378037 , n378036 );
not ( n57572 , n378037 );
and ( n378039 , n57563 , n57572 );
not ( n378040 , n365428 );
buf ( n378041 , n365319 );
not ( n378042 , n378041 );
buf ( n378043 , n378042 );
not ( n57578 , n378043 );
or ( n378045 , n378040 , n57578 );
buf ( n378046 , n366329 );
buf ( n57581 , n365422 );
nand ( n57582 , n378046 , n57581 );
buf ( n57583 , n57582 );
nand ( n378050 , n378045 , n57583 );
not ( n57585 , n378050 );
nor ( n378052 , n57585 , n49692 );
buf ( n378053 , n378052 );
nor ( n57588 , n378039 , n378053 );
buf ( n378055 , n57588 );
buf ( n378056 , n378055 );
not ( n378057 , n378056 );
buf ( n378058 , n378057 );
buf ( n378059 , n378058 );
not ( n57594 , n378059 );
or ( n378061 , n57561 , n57594 );
buf ( n378062 , n378022 );
not ( n57597 , n378062 );
buf ( n378064 , n378036 );
not ( n57599 , n378064 );
buf ( n378066 , n361971 );
not ( n57601 , n378066 );
and ( n378068 , n57599 , n57601 );
buf ( n57603 , n378052 );
nor ( n57604 , n378068 , n57603 );
buf ( n57605 , n57604 );
buf ( n378072 , n57605 );
not ( n378073 , n378072 );
or ( n57608 , n57597 , n378073 );
not ( n378075 , n365115 );
not ( n378076 , n377859 );
or ( n57611 , n378075 , n378076 );
and ( n378078 , n364981 , n31283 );
not ( n378079 , n364981 );
and ( n57614 , n378079 , n364808 );
or ( n378081 , n378078 , n57614 );
nand ( n57616 , n365033 , n378081 );
nand ( n57617 , n57611 , n57616 );
buf ( n378084 , n57617 );
nand ( n57619 , n57608 , n378084 );
buf ( n378086 , n57619 );
buf ( n378087 , n378086 );
nand ( n57622 , n378061 , n378087 );
buf ( n378089 , n57622 );
not ( n57624 , n378089 );
xor ( n57625 , n377254 , n377274 );
xor ( n57626 , n57625 , n377316 );
buf ( n378093 , n57626 );
buf ( n378094 , n378093 );
buf ( n378095 , n359685 );
buf ( n378096 , n29121 );
buf ( n57631 , n378096 );
buf ( n378098 , n57631 );
buf ( n378099 , n378098 );
and ( n57634 , n378095 , n378099 );
buf ( n378101 , n57634 );
buf ( n378102 , n378101 );
xor ( n378103 , n378094 , n378102 );
buf ( n378104 , n378050 );
not ( n378105 , n378104 );
buf ( n378106 , n46135 );
not ( n378107 , n378106 );
or ( n57642 , n378105 , n378107 );
not ( n57643 , n361911 );
not ( n378110 , n365989 );
or ( n378111 , n57643 , n378110 );
not ( n57646 , n364766 );
nand ( n378113 , n57646 , n365980 );
nand ( n378114 , n378111 , n378113 );
nand ( n57649 , n368724 , n378114 );
buf ( n378116 , n57649 );
nand ( n378117 , n57642 , n378116 );
buf ( n378118 , n378117 );
buf ( n378119 , n378118 );
xor ( n378120 , n378103 , n378119 );
buf ( n378121 , n378120 );
buf ( n378122 , n378121 );
not ( n378123 , n378122 );
buf ( n378124 , n378123 );
nand ( n57659 , n57624 , n378124 );
not ( n378126 , n57659 );
buf ( n378127 , n377308 );
not ( n57662 , n378127 );
buf ( n378129 , n46463 );
not ( n57664 , n378129 );
or ( n378131 , n57662 , n57664 );
not ( n57666 , n32202 );
buf ( n378133 , n342614 );
buf ( n378134 , n378133 );
buf ( n378135 , n378134 );
buf ( n378136 , n378135 );
not ( n378137 , n378136 );
buf ( n378138 , n378137 );
not ( n57673 , n378138 );
or ( n378140 , n57666 , n57673 );
not ( n378141 , n32202 );
nand ( n57676 , n375914 , n378141 );
nand ( n378143 , n378140 , n57676 );
buf ( n378144 , n378143 );
buf ( n378145 , n375896 );
nand ( n378146 , n378144 , n378145 );
buf ( n378147 , n378146 );
buf ( n378148 , n378147 );
nand ( n378149 , n378131 , n378148 );
buf ( n378150 , n378149 );
not ( n57685 , n378150 );
buf ( n378152 , n351160 );
not ( n378153 , n378152 );
not ( n57688 , n22769 );
buf ( n378155 , n57688 );
not ( n378156 , n378155 );
or ( n378157 , n378153 , n378156 );
buf ( n378158 , n46693 );
buf ( n378159 , n364915 );
nand ( n378160 , n378158 , n378159 );
buf ( n378161 , n378160 );
buf ( n378162 , n378161 );
nand ( n57697 , n378157 , n378162 );
buf ( n378164 , n57697 );
not ( n378165 , n378164 );
not ( n378166 , n363429 );
or ( n57701 , n378165 , n378166 );
buf ( n378168 , n365490 );
not ( n378169 , n378168 );
buf ( n378170 , n377683 );
not ( n378171 , n378170 );
or ( n57706 , n378169 , n378171 );
buf ( n378173 , n55539 );
buf ( n378174 , n45336 );
nand ( n57709 , n378173 , n378174 );
buf ( n378176 , n57709 );
buf ( n378177 , n378176 );
nand ( n378178 , n57706 , n378177 );
buf ( n378179 , n378178 );
buf ( n378180 , n378179 );
buf ( n57715 , n57228 );
buf ( n378182 , n57715 );
buf ( n378183 , n378182 );
buf ( n378184 , n378183 );
nand ( n378185 , n378180 , n378184 );
buf ( n378186 , n378185 );
nand ( n378187 , n57701 , n378186 );
xor ( n57722 , n57685 , n378187 );
not ( n57723 , n56531 );
nor ( n57724 , n57723 , n376943 );
not ( n378191 , n57724 );
nor ( n378192 , n378191 , n56320 );
not ( n57727 , n378192 );
not ( n378194 , n376317 );
nor ( n57729 , n378194 , n376946 );
nand ( n57730 , n376699 , n57729 );
not ( n378197 , n376946 );
nand ( n57732 , n378197 , n376707 );
nand ( n378199 , n57730 , n57732 );
not ( n57734 , n378199 );
or ( n57735 , n57727 , n57734 );
not ( n378202 , n55729 );
not ( n378203 , n56544 );
or ( n57738 , n378202 , n378203 );
nand ( n378205 , n57738 , n376727 );
and ( n378206 , n57724 , n378205 );
not ( n57741 , n376733 );
and ( n378208 , n57741 , n55772 );
nor ( n378209 , n378206 , n378208 , n376735 );
nand ( n57744 , n57735 , n378209 );
not ( n378211 , n56327 );
nand ( n57746 , n378211 , n55779 );
xnor ( n57747 , n57744 , n57746 );
buf ( n378214 , n57747 );
buf ( n378215 , n378214 );
buf ( n378216 , n376990 );
and ( n378217 , n378215 , n378216 );
buf ( n378218 , n57747 );
not ( n57753 , n378218 );
buf ( n57754 , n57753 );
buf ( n378221 , n57754 );
buf ( n378222 , n376997 );
and ( n57757 , n378221 , n378222 );
buf ( n378224 , n377003 );
nor ( n57759 , n378217 , n57757 , n378224 );
buf ( n57760 , n57759 );
not ( n378227 , n376755 );
not ( n57762 , n56409 );
or ( n57763 , n378227 , n57762 );
not ( n57764 , n56430 );
nand ( n378231 , n57763 , n57764 );
not ( n378232 , n56434 );
nand ( n57767 , n378232 , n376759 );
xnor ( n57768 , n378231 , n57767 );
buf ( n378235 , n57768 );
not ( n378236 , n376833 );
nor ( n57771 , n378236 , n376838 );
not ( n57772 , n56344 );
nor ( n57773 , n57772 , n56338 );
not ( n57774 , n57773 );
nand ( n378241 , n56408 , n56389 );
not ( n57776 , n378241 );
or ( n378243 , n57774 , n57776 );
not ( n57778 , n376829 );
not ( n57779 , n57778 );
not ( n57780 , n56338 );
and ( n57781 , n57779 , n57780 );
nor ( n57782 , n57781 , n376835 );
nand ( n57783 , n378243 , n57782 );
not ( n378250 , n57783 );
and ( n57785 , n57771 , n378250 );
not ( n57786 , n57771 );
and ( n378253 , n57786 , n57783 );
or ( n378254 , n57785 , n378253 );
not ( n57789 , n378254 );
buf ( n378256 , n57789 );
and ( n57791 , n378235 , n378256 );
not ( n378258 , n378235 );
buf ( n378259 , n378254 );
and ( n378260 , n378258 , n378259 );
nor ( n57795 , n57791 , n378260 );
buf ( n378262 , n57795 );
buf ( n57797 , n378262 );
buf ( n378264 , n376903 );
not ( n57799 , n378264 );
buf ( n57800 , n57799 );
buf ( n378267 , n57800 );
buf ( n378268 , n57768 );
not ( n378269 , n378268 );
buf ( n378270 , n378269 );
buf ( n378271 , n378270 );
and ( n57806 , n378267 , n378271 );
buf ( n378273 , n376903 );
buf ( n378274 , n57768 );
and ( n57809 , n378273 , n378274 );
nor ( n378276 , n57806 , n57809 );
buf ( n378277 , n378276 );
buf ( n378278 , n378277 );
and ( n378279 , n57797 , n378278 );
buf ( n378280 , n378279 );
buf ( n378281 , n378280 );
buf ( n378282 , n57800 );
not ( n57817 , n378282 );
buf ( n378284 , n57817 );
buf ( n378285 , n378284 );
nand ( n378286 , n378281 , n378285 );
buf ( n378287 , n378286 );
buf ( n378288 , n378287 );
buf ( n378289 , n378262 );
not ( n57824 , n378289 );
buf ( n378291 , n57824 );
buf ( n378292 , n378291 );
buf ( n378293 , n378284 );
nand ( n57828 , n378292 , n378293 );
buf ( n378295 , n57828 );
buf ( n378296 , n378295 );
and ( n378297 , n378288 , n378296 );
buf ( n378298 , n378297 );
xor ( n378299 , n57760 , n378298 );
buf ( n57834 , n376971 );
buf ( n57835 , n376866 );
and ( n57836 , n57834 , n57835 );
buf ( n378303 , n376993 );
buf ( n378304 , n376875 );
and ( n378305 , n378303 , n378304 );
nor ( n57840 , n57836 , n378305 );
buf ( n378307 , n57840 );
buf ( n378308 , n378307 );
buf ( n378309 , n376924 );
or ( n57844 , n378308 , n378309 );
buf ( n378311 , n376879 );
buf ( n378312 , n56517 );
or ( n57847 , n378311 , n378312 );
nand ( n378314 , n57844 , n57847 );
buf ( n378315 , n378314 );
and ( n57850 , n378299 , n378315 );
and ( n378317 , n57760 , n378298 );
or ( n57852 , n57850 , n378317 );
buf ( n378319 , n57852 );
buf ( n378320 , n377006 );
not ( n57855 , n378320 );
buf ( n378322 , n376937 );
not ( n378323 , n378322 );
or ( n57858 , n57855 , n378323 );
buf ( n378325 , n377009 );
nand ( n57860 , n57858 , n378325 );
buf ( n378327 , n57860 );
buf ( n378328 , n378327 );
xor ( n57863 , n378319 , n378328 );
buf ( n378330 , n376743 );
buf ( n378331 , n57800 );
and ( n57866 , n378330 , n378331 );
buf ( n378333 , n376871 );
buf ( n378334 , n378284 );
and ( n57869 , n378333 , n378334 );
nor ( n57870 , n57866 , n57869 );
buf ( n378337 , n57870 );
buf ( n378338 , n378337 );
buf ( n378339 , n378280 );
not ( n57874 , n378339 );
buf ( n378341 , n57874 );
buf ( n378342 , n378341 );
or ( n57877 , n378338 , n378342 );
buf ( n378344 , n378295 );
nand ( n57879 , n57877 , n378344 );
buf ( n378346 , n57879 );
buf ( n378347 , n378346 );
not ( n378348 , n55772 );
nor ( n57883 , n378348 , n376735 );
not ( n378350 , n57883 );
nor ( n57885 , n56320 , n55761 );
not ( n378352 , n57885 );
not ( n378353 , n56544 );
and ( n57888 , n57732 , n378353 );
and ( n57889 , n57730 , n57888 );
not ( n57890 , n57889 );
not ( n378357 , n57890 );
or ( n57892 , n378352 , n378357 );
not ( n57893 , n56547 );
and ( n57894 , n57893 , n376120 );
nor ( n57895 , n57894 , n376732 );
nand ( n57896 , n57892 , n57895 );
not ( n57897 , n57896 );
not ( n57898 , n57897 );
or ( n57899 , n378350 , n57898 );
not ( n57900 , n57883 );
nand ( n57901 , n57900 , n57896 );
nand ( n378368 , n57899 , n57901 );
buf ( n378369 , n378368 );
buf ( n378370 , n376990 );
and ( n378371 , n378369 , n378370 );
not ( n378372 , n378368 );
buf ( n378373 , n378372 );
buf ( n378374 , n376997 );
and ( n378375 , n378373 , n378374 );
buf ( n378376 , n377003 );
nor ( n57911 , n378371 , n378375 , n378376 );
buf ( n57912 , n57911 );
buf ( n57913 , n57912 );
or ( n57914 , n378347 , n57913 );
buf ( n378381 , n57914 );
xor ( n57916 , n57760 , n378298 );
xor ( n378383 , n57916 , n378315 );
and ( n57918 , n378381 , n378383 );
buf ( n378385 , n57912 );
not ( n378386 , n378385 );
buf ( n378387 , n378346 );
not ( n57922 , n378387 );
or ( n378389 , n378386 , n57922 );
buf ( n57924 , n378381 );
nand ( n57925 , n378389 , n57924 );
buf ( n57926 , n57925 );
buf ( n378393 , n378214 );
buf ( n378394 , n376866 );
and ( n57929 , n378393 , n378394 );
buf ( n378396 , n57754 );
buf ( n378397 , n376875 );
and ( n57932 , n378396 , n378397 );
nor ( n57933 , n57929 , n57932 );
buf ( n378400 , n57933 );
buf ( n378401 , n378400 );
buf ( n378402 , n376924 );
or ( n378403 , n378401 , n378402 );
buf ( n378404 , n378307 );
buf ( n378405 , n56517 );
or ( n57940 , n378404 , n378405 );
nand ( n57941 , n378403 , n57940 );
buf ( n378408 , n57941 );
xor ( n57943 , n57926 , n378408 );
buf ( n378410 , n376971 );
buf ( n378411 , n57800 );
and ( n378412 , n378410 , n378411 );
buf ( n378413 , n376993 );
buf ( n378414 , n378284 );
and ( n57949 , n378413 , n378414 );
nor ( n57950 , n378412 , n57949 );
buf ( n378417 , n57950 );
buf ( n378418 , n378417 );
buf ( n378419 , n378341 );
or ( n57954 , n378418 , n378419 );
buf ( n378421 , n378337 );
buf ( n57956 , n378291 );
not ( n57957 , n57956 );
buf ( n378424 , n57957 );
buf ( n378425 , n378424 );
or ( n378426 , n378421 , n378425 );
nand ( n57961 , n57954 , n378426 );
buf ( n378428 , n57961 );
buf ( n378429 , n378428 );
not ( n57964 , n56344 );
not ( n378431 , n378241 );
or ( n57966 , n57964 , n378431 );
nand ( n378433 , n57966 , n57778 );
nor ( n57968 , n56338 , n376835 );
xor ( n57969 , n378433 , n57968 );
not ( n57970 , n57969 );
not ( n378437 , n376753 );
not ( n57972 , n378437 );
not ( n57973 , n378241 );
or ( n57974 , n57972 , n57973 );
not ( n57975 , n56413 );
nand ( n57976 , n57974 , n57975 );
not ( n378443 , n57976 );
nand ( n57978 , n56418 , n56341 );
not ( n378445 , n57978 );
and ( n57980 , n378443 , n378445 );
and ( n378447 , n57976 , n57978 );
nor ( n57982 , n57980 , n378447 );
not ( n57983 , n57982 );
not ( n378450 , n57983 );
or ( n378451 , n57970 , n378450 );
or ( n57986 , n57969 , n57983 );
nand ( n378453 , n378451 , n57986 );
buf ( n378454 , n378453 );
buf ( n378455 , n57789 );
buf ( n378456 , n57969 );
not ( n378457 , n378456 );
buf ( n378458 , n378457 );
buf ( n378459 , n378458 );
and ( n378460 , n378455 , n378459 );
buf ( n378461 , n378254 );
buf ( n378462 , n57969 );
and ( n57997 , n378461 , n378462 );
nor ( n378464 , n378460 , n57997 );
buf ( n378465 , n378464 );
buf ( n378466 , n378465 );
and ( n378467 , n378454 , n378466 );
buf ( n378468 , n378467 );
buf ( n378469 , n378468 );
not ( n378470 , n57789 );
buf ( n378471 , n378470 );
nand ( n58006 , n378469 , n378471 );
buf ( n378473 , n58006 );
buf ( n378474 , n378473 );
not ( n58009 , n378453 );
not ( n378476 , n58009 );
buf ( n378477 , n378476 );
buf ( n378478 , n57789 );
nor ( n58013 , n378477 , n378478 );
buf ( n378480 , n58013 );
buf ( n58015 , n378480 );
not ( n378482 , n58015 );
buf ( n378483 , n378482 );
buf ( n378484 , n378483 );
and ( n378485 , n378474 , n378484 );
buf ( n378486 , n378485 );
buf ( n378487 , n378486 );
xor ( n378488 , n378429 , n378487 );
buf ( n378489 , n378368 );
buf ( n378490 , n376866 );
and ( n58025 , n378489 , n378490 );
buf ( n378492 , n378372 );
buf ( n378493 , n376875 );
and ( n378494 , n378492 , n378493 );
nor ( n58029 , n58025 , n378494 );
buf ( n58030 , n58029 );
buf ( n378497 , n58030 );
buf ( n378498 , n376924 );
or ( n378499 , n378497 , n378498 );
buf ( n378500 , n378400 );
buf ( n378501 , n56517 );
or ( n58036 , n378500 , n378501 );
nand ( n378503 , n378499 , n58036 );
buf ( n378504 , n378503 );
buf ( n378505 , n378504 );
and ( n378506 , n378488 , n378505 );
and ( n58041 , n378429 , n378487 );
or ( n378508 , n378506 , n58041 );
buf ( n378509 , n378508 );
and ( n378510 , n57943 , n378509 );
and ( n58045 , n57926 , n378408 );
or ( n58046 , n378510 , n58045 );
xor ( n378513 , n57760 , n378298 );
xor ( n378514 , n378513 , n378315 );
and ( n58049 , n58046 , n378514 );
and ( n378516 , n378381 , n58046 );
or ( n378517 , n57918 , n58049 , n378516 );
buf ( n378518 , n378517 );
xor ( n378519 , n57863 , n378518 );
buf ( n378520 , n378519 );
not ( n58055 , n46463 );
not ( n58056 , n378143 );
or ( n378523 , n58055 , n58056 );
buf ( n378524 , n375896 );
and ( n58059 , n31231 , n366659 );
not ( n378526 , n31231 );
and ( n378527 , n378526 , n378135 );
or ( n58062 , n58059 , n378527 );
buf ( n378529 , n58062 );
nand ( n378530 , n378524 , n378529 );
buf ( n378531 , n378530 );
nand ( n58066 , n378523 , n378531 );
xor ( n58067 , n378520 , n58066 );
buf ( n378534 , n365490 );
not ( n58069 , n378534 );
buf ( n378536 , n22707 );
not ( n58071 , n378536 );
or ( n378538 , n58069 , n58071 );
not ( n58073 , n375931 );
buf ( n378540 , n58073 );
buf ( n378541 , n351195 );
not ( n58076 , n378541 );
buf ( n378543 , n58076 );
buf ( n378544 , n378543 );
nand ( n58079 , n378540 , n378544 );
buf ( n378546 , n58079 );
buf ( n378547 , n378546 );
nand ( n378548 , n378538 , n378547 );
buf ( n378549 , n378548 );
buf ( n378550 , n378549 );
not ( n58085 , n378550 );
buf ( n378552 , n366396 );
not ( n378553 , n378552 );
or ( n58088 , n58085 , n378553 );
buf ( n378555 , n57233 );
not ( n58090 , n378555 );
buf ( n378557 , n55583 );
not ( n58092 , n378557 );
or ( n58093 , n58090 , n58092 );
buf ( n378560 , n58073 );
buf ( n378561 , n31194 );
nand ( n58096 , n378560 , n378561 );
buf ( n378563 , n58096 );
buf ( n378564 , n378563 );
nand ( n378565 , n58093 , n378564 );
buf ( n378566 , n378565 );
buf ( n378567 , n378566 );
buf ( n378568 , n377271 );
nand ( n58103 , n378567 , n378568 );
buf ( n378570 , n58103 );
buf ( n378571 , n378570 );
nand ( n58106 , n58088 , n378571 );
buf ( n58107 , n58106 );
and ( n378574 , n58067 , n58107 );
and ( n58109 , n378520 , n58066 );
or ( n378576 , n378574 , n58109 );
xnor ( n58111 , n57722 , n378576 );
not ( n58112 , n58111 );
not ( n58113 , n365152 );
not ( n378580 , n57280 );
not ( n58115 , n366077 );
or ( n378582 , n378580 , n58115 );
buf ( n378583 , n45916 );
buf ( n378584 , n342908 );
nand ( n378585 , n378583 , n378584 );
buf ( n378586 , n378585 );
nand ( n378587 , n378582 , n378586 );
not ( n58122 , n378587 );
or ( n58123 , n58113 , n58122 );
buf ( n58124 , n365187 );
buf ( n378591 , n22956 );
buf ( n378592 , n48496 );
and ( n378593 , n378591 , n378592 );
not ( n378594 , n378591 );
buf ( n378595 , n368700 );
and ( n378596 , n378594 , n378595 );
nor ( n58131 , n378593 , n378596 );
buf ( n378598 , n58131 );
buf ( n378599 , n378598 );
nand ( n378600 , n58124 , n378599 );
buf ( n378601 , n378600 );
nand ( n58136 , n58123 , n378601 );
not ( n378603 , n58136 );
nand ( n58138 , n58112 , n378603 );
not ( n378605 , n58138 );
buf ( n378606 , n377782 );
not ( n58141 , n378606 );
buf ( n378608 , n367600 );
not ( n378609 , n378608 );
or ( n58144 , n58141 , n378609 );
buf ( n378611 , n365293 );
buf ( n378612 , n377779 );
nand ( n378613 , n378611 , n378612 );
buf ( n378614 , n378613 );
buf ( n378615 , n378614 );
nand ( n58150 , n58144 , n378615 );
buf ( n378617 , n58150 );
not ( n58152 , n378617 );
not ( n378619 , n45376 );
not ( n378620 , n378619 );
or ( n58155 , n58152 , n378620 );
buf ( n378622 , n377353 );
not ( n58157 , n378622 );
buf ( n378624 , n45116 );
not ( n378625 , n378624 );
or ( n58160 , n58157 , n378625 );
buf ( n378627 , n365569 );
buf ( n378628 , n377352 );
nand ( n58163 , n378627 , n378628 );
buf ( n58164 , n58163 );
buf ( n58165 , n58164 );
nand ( n58166 , n58160 , n58165 );
buf ( n58167 , n58166 );
buf ( n378634 , n58167 );
not ( n58169 , n378634 );
buf ( n58170 , n58169 );
or ( n58171 , n58170 , n370050 );
nand ( n58172 , n58155 , n58171 );
not ( n58173 , n58172 );
or ( n58174 , n378605 , n58173 );
and ( n58175 , n58111 , n58136 );
not ( n378642 , n58175 );
nand ( n378643 , n58174 , n378642 );
not ( n378644 , n378643 );
or ( n58179 , n378126 , n378644 );
buf ( n378646 , n378121 );
buf ( n378647 , n378089 );
nand ( n58182 , n378646 , n378647 );
buf ( n378649 , n58182 );
nand ( n58184 , n58179 , n378649 );
nand ( n58185 , n57544 , n58184 );
nand ( n58186 , n57538 , n58185 );
buf ( n378653 , n58186 );
nand ( n378654 , n57379 , n378653 );
buf ( n378655 , n378654 );
buf ( n378656 , n378655 );
nand ( n378657 , n57374 , n378656 );
buf ( n378658 , n378657 );
and ( n58193 , n377803 , n378658 );
not ( n378660 , n377803 );
buf ( n378661 , n377810 );
not ( n58196 , n378661 );
buf ( n378663 , n57371 );
not ( n58198 , n378663 );
or ( n378665 , n58196 , n58198 );
buf ( n378666 , n378655 );
nand ( n58201 , n378665 , n378666 );
buf ( n378668 , n58201 );
not ( n378669 , n378668 );
and ( n58204 , n378660 , n378669 );
nor ( n378671 , n58193 , n58204 );
buf ( n378672 , n368611 );
not ( n58207 , n378672 );
buf ( n378674 , n377642 );
not ( n378675 , n378674 );
or ( n58210 , n58207 , n378675 );
not ( n378677 , n368549 );
not ( n58212 , n373463 );
or ( n58213 , n378677 , n58212 );
buf ( n58214 , n360885 );
buf ( n58215 , n368554 );
nand ( n58216 , n58214 , n58215 );
buf ( n58217 , n58216 );
nand ( n378684 , n58213 , n58217 );
buf ( n378685 , n378684 );
buf ( n378686 , n369444 );
nand ( n378687 , n378685 , n378686 );
buf ( n378688 , n378687 );
buf ( n378689 , n378688 );
nand ( n58224 , n58210 , n378689 );
buf ( n378691 , n58224 );
buf ( n378692 , n378691 );
not ( n58227 , n378692 );
buf ( n378694 , n58227 );
buf ( n378695 , n378694 );
not ( n378696 , n378695 );
not ( n58231 , n363416 );
not ( n378698 , n58231 );
buf ( n378699 , n31260 );
not ( n58234 , n378699 );
buf ( n378701 , n57688 );
not ( n378702 , n378701 );
or ( n58237 , n58234 , n378702 );
buf ( n378704 , n31260 );
buf ( n378705 , n377683 );
or ( n58240 , n378704 , n378705 );
buf ( n378707 , n58240 );
buf ( n378708 , n378707 );
nand ( n58243 , n58237 , n378708 );
buf ( n58244 , n58243 );
not ( n378711 , n58244 );
or ( n58246 , n378698 , n378711 );
nand ( n378713 , n375890 , n363428 );
nand ( n378714 , n58246 , n378713 );
buf ( n378715 , n378714 );
not ( n378716 , n378715 );
buf ( n378717 , n377181 );
not ( n378718 , n378717 );
buf ( n378719 , n378718 );
buf ( n378720 , n378719 );
not ( n378721 , n378720 );
and ( n378722 , n378716 , n378721 );
buf ( n378723 , n378714 );
buf ( n378724 , n378719 );
and ( n378725 , n378723 , n378724 );
nor ( n378726 , n378722 , n378725 );
buf ( n378727 , n378726 );
not ( n378728 , n378727 );
buf ( n378729 , n377214 );
not ( n378730 , n378729 );
buf ( n378731 , n368706 );
not ( n58266 , n378731 );
or ( n378733 , n378730 , n58266 );
buf ( n378734 , n365344 );
not ( n378735 , n378734 );
buf ( n378736 , n378735 );
buf ( n378737 , n378736 );
not ( n378738 , n378737 );
buf ( n378739 , n342335 );
not ( n378740 , n378739 );
or ( n58275 , n378738 , n378740 );
buf ( n378742 , n365915 );
buf ( n378743 , n49315 );
nand ( n378744 , n378742 , n378743 );
buf ( n378745 , n378744 );
buf ( n378746 , n378745 );
nand ( n378747 , n58275 , n378746 );
buf ( n378748 , n378747 );
buf ( n378749 , n378748 );
buf ( n378750 , n48490 );
nand ( n378751 , n378749 , n378750 );
buf ( n378752 , n378751 );
buf ( n378753 , n378752 );
nand ( n58288 , n378733 , n378753 );
buf ( n58289 , n58288 );
not ( n378756 , n58289 );
not ( n58291 , n378756 );
or ( n378758 , n378728 , n58291 );
or ( n378759 , n378756 , n378727 );
nand ( n58294 , n378758 , n378759 );
not ( n378761 , n45075 );
buf ( n378762 , n342881 );
not ( n58297 , n378762 );
buf ( n378764 , n366322 );
not ( n58299 , n378764 );
or ( n58300 , n58297 , n58299 );
buf ( n378767 , n361716 );
buf ( n378768 , n365202 );
nand ( n378769 , n378767 , n378768 );
buf ( n378770 , n378769 );
buf ( n378771 , n378770 );
nand ( n378772 , n58300 , n378771 );
buf ( n378773 , n378772 );
not ( n58308 , n378773 );
or ( n58309 , n378761 , n58308 );
buf ( n378776 , n365227 );
not ( n58311 , n378776 );
and ( n58312 , n362534 , n365202 );
not ( n378779 , n362534 );
and ( n58314 , n378779 , n342881 );
or ( n378781 , n58312 , n58314 );
buf ( n378782 , n378781 );
nand ( n378783 , n58311 , n378782 );
buf ( n378784 , n378783 );
nand ( n58319 , n58309 , n378784 );
and ( n378786 , n58294 , n58319 );
not ( n378787 , n58294 );
not ( n58322 , n58319 );
and ( n378789 , n378787 , n58322 );
nor ( n58324 , n378786 , n378789 );
not ( n378791 , n377395 );
not ( n58326 , n46557 );
or ( n58327 , n378791 , n58326 );
buf ( n378794 , n369374 );
not ( n378795 , n378794 );
buf ( n378796 , n365468 );
not ( n378797 , n378796 );
or ( n378798 , n378795 , n378797 );
buf ( n378799 , n360610 );
buf ( n378800 , n49178 );
nand ( n58335 , n378799 , n378800 );
buf ( n378802 , n58335 );
buf ( n378803 , n378802 );
nand ( n378804 , n378798 , n378803 );
buf ( n378805 , n378804 );
buf ( n378806 , n378805 );
buf ( n378807 , n360574 );
nand ( n58342 , n378806 , n378807 );
buf ( n378809 , n58342 );
nand ( n58344 , n58327 , n378809 );
xor ( n58345 , n58324 , n58344 );
buf ( n378812 , n58345 );
not ( n58347 , n378812 );
buf ( n378814 , n58347 );
buf ( n378815 , n378814 );
not ( n58350 , n378815 );
or ( n58351 , n378696 , n58350 );
buf ( n378818 , n58345 );
buf ( n378819 , n378691 );
nand ( n58354 , n378818 , n378819 );
buf ( n378821 , n58354 );
buf ( n378822 , n378821 );
nand ( n58357 , n58351 , n378822 );
buf ( n378824 , n58357 );
buf ( n58359 , n378824 );
not ( n58360 , n378719 );
not ( n378827 , n377229 );
or ( n378828 , n58360 , n378827 );
or ( n58363 , n378719 , n377229 );
nand ( n378830 , n58363 , n56798 );
nand ( n378831 , n378828 , n378830 );
buf ( n378832 , n39701 );
not ( n378833 , n378832 );
buf ( n378834 , n377086 );
not ( n58369 , n378834 );
or ( n378836 , n378833 , n58369 );
buf ( n378837 , n367796 );
xor ( n58372 , n349127 , n349183 );
xor ( n378839 , n58372 , n29165 );
buf ( n378840 , n378839 );
buf ( n378841 , n378840 );
buf ( n378842 , n378841 );
buf ( n378843 , n378842 );
not ( n58378 , n378843 );
buf ( n378845 , n58378 );
buf ( n58380 , n378845 );
buf ( n378847 , n58380 );
buf ( n378848 , n378847 );
not ( n58383 , n378848 );
buf ( n378850 , n45234 );
not ( n58385 , n378850 );
or ( n378852 , n58383 , n58385 );
buf ( n378853 , n366537 );
buf ( n378854 , n378847 );
not ( n58389 , n378854 );
buf ( n378856 , n58389 );
buf ( n378857 , n378856 );
nand ( n58392 , n378853 , n378857 );
buf ( n378859 , n58392 );
buf ( n378860 , n378859 );
nand ( n378861 , n378852 , n378860 );
buf ( n378862 , n378861 );
buf ( n378863 , n378862 );
nand ( n58398 , n378837 , n378863 );
buf ( n378865 , n58398 );
buf ( n378866 , n378865 );
nand ( n58401 , n378836 , n378866 );
buf ( n378868 , n58401 );
xor ( n58403 , n378831 , n378868 );
buf ( n378870 , n377157 );
not ( n378871 , n378870 );
buf ( n378872 , n378871 );
buf ( n378873 , n378872 );
not ( n378874 , n378873 );
buf ( n378875 , n40058 );
not ( n58410 , n378875 );
or ( n58411 , n378874 , n58410 );
buf ( n378878 , n377757 );
not ( n58413 , n378878 );
buf ( n378880 , n363122 );
not ( n378881 , n378880 );
or ( n58416 , n58413 , n378881 );
buf ( n378883 , n365528 );
buf ( n378884 , n377757 );
not ( n378885 , n378884 );
buf ( n378886 , n378885 );
buf ( n378887 , n378886 );
nand ( n58422 , n378883 , n378887 );
buf ( n378889 , n58422 );
buf ( n378890 , n378889 );
nand ( n58425 , n58416 , n378890 );
buf ( n58426 , n58425 );
buf ( n378893 , n58426 );
buf ( n378894 , n39949 );
nand ( n58429 , n378893 , n378894 );
buf ( n378896 , n58429 );
buf ( n378897 , n378896 );
nand ( n58432 , n58411 , n378897 );
buf ( n378899 , n58432 );
xnor ( n58434 , n58403 , n378899 );
not ( n58435 , n58434 );
buf ( n378902 , n58435 );
xor ( n378903 , n58359 , n378902 );
buf ( n378904 , n378903 );
buf ( n378905 , n378904 );
buf ( n378906 , n49609 );
not ( n378907 , n378906 );
and ( n378908 , n369769 , n40252 );
not ( n378909 , n369769 );
and ( n378910 , n378909 , n40251 );
or ( n378911 , n378908 , n378910 );
buf ( n378912 , n378911 );
not ( n378913 , n378912 );
or ( n58436 , n378907 , n378913 );
buf ( n378915 , n375864 );
buf ( n378916 , n369804 );
nand ( n58439 , n378915 , n378916 );
buf ( n378918 , n58439 );
buf ( n378919 , n378918 );
nand ( n378920 , n58436 , n378919 );
buf ( n378921 , n378920 );
buf ( n378922 , n378921 );
buf ( n378923 , n377580 );
not ( n58442 , n378923 );
buf ( n378925 , n377585 );
not ( n58444 , n378925 );
buf ( n378927 , n46902 );
not ( n58446 , n378927 );
or ( n58447 , n58444 , n58446 );
buf ( n58448 , n40199 );
buf ( n378931 , n377592 );
nand ( n378932 , n58448 , n378931 );
buf ( n378933 , n378932 );
buf ( n378934 , n378933 );
nand ( n58453 , n58447 , n378934 );
buf ( n378936 , n58453 );
buf ( n378937 , n378936 );
not ( n58456 , n378937 );
or ( n58457 , n58442 , n58456 );
buf ( n378940 , n57530 );
buf ( n378941 , n377598 );
nand ( n378942 , n378940 , n378941 );
buf ( n378943 , n378942 );
buf ( n378944 , n378943 );
nand ( n378945 , n58457 , n378944 );
buf ( n378946 , n378945 );
buf ( n378947 , n378946 );
xor ( n58462 , n378922 , n378947 );
not ( n58463 , n22707 );
buf ( n378950 , n58463 );
not ( n58465 , n378950 );
buf ( n378952 , n45125 );
not ( n378953 , n378952 );
or ( n58468 , n58465 , n378953 );
buf ( n378955 , n352192 );
not ( n378956 , n55583 );
not ( n58471 , n378956 );
buf ( n378958 , n58471 );
nand ( n58473 , n378955 , n378958 );
buf ( n378960 , n58473 );
buf ( n378961 , n378960 );
nand ( n58475 , n58468 , n378961 );
buf ( n378963 , n58475 );
buf ( n378964 , n378963 );
not ( n378965 , n378964 );
buf ( n378966 , n366428 );
not ( n58478 , n378966 );
or ( n58479 , n378965 , n58478 );
buf ( n378969 , n377173 );
buf ( n378970 , n366399 );
nand ( n58482 , n378969 , n378970 );
buf ( n378972 , n58482 );
buf ( n378973 , n378972 );
nand ( n378974 , n58479 , n378973 );
buf ( n378975 , n378974 );
not ( n58487 , n56794 );
buf ( n58488 , n350650 );
not ( n378978 , n22619 );
not ( n58490 , n30905 );
or ( n58491 , n378978 , n58490 );
or ( n378981 , n30905 , n22619 );
nand ( n58493 , n58491 , n378981 );
and ( n378983 , n58488 , n58493 );
not ( n58495 , n58488 );
not ( n58496 , n58493 );
and ( n58497 , n58495 , n58496 );
nor ( n378987 , n378983 , n58497 );
not ( n58499 , n378987 );
or ( n378989 , n58487 , n58499 );
nand ( n58501 , n45553 , n377202 );
nand ( n58502 , n378989 , n58501 );
xor ( n378992 , n378975 , n58502 );
buf ( n378993 , n46463 );
not ( n378994 , n378993 );
buf ( n378995 , n46477 );
not ( n58507 , n378995 );
buf ( n378997 , n44661 );
not ( n378998 , n378997 );
or ( n58510 , n58507 , n378998 );
buf ( n379000 , n31072 );
buf ( n379001 , n46474 );
nand ( n58513 , n379000 , n379001 );
buf ( n58514 , n58513 );
buf ( n379004 , n58514 );
nand ( n379005 , n58510 , n379004 );
buf ( n379006 , n379005 );
buf ( n379007 , n379006 );
not ( n379008 , n379007 );
or ( n58520 , n378994 , n379008 );
buf ( n379010 , n55558 );
buf ( n379011 , n46521 );
nand ( n58523 , n379010 , n379011 );
buf ( n379013 , n58523 );
buf ( n379014 , n379013 );
nand ( n58526 , n58520 , n379014 );
buf ( n379016 , n58526 );
xor ( n58528 , n378992 , n379016 );
buf ( n379018 , n58528 );
not ( n58530 , n39217 );
buf ( n379020 , n377353 );
not ( n58532 , n379020 );
buf ( n379022 , n365368 );
not ( n58534 , n379022 );
or ( n58535 , n58532 , n58534 );
buf ( n379025 , n366360 );
buf ( n379026 , n377352 );
nand ( n58538 , n379025 , n379026 );
buf ( n379028 , n58538 );
buf ( n379029 , n379028 );
nand ( n58541 , n58535 , n379029 );
buf ( n379031 , n58541 );
not ( n58543 , n379031 );
or ( n58544 , n58530 , n58543 );
not ( n58545 , n57339 );
nand ( n58546 , n58545 , n45204 );
nand ( n58547 , n58544 , n58546 );
buf ( n379037 , n58547 );
xor ( n379038 , n379018 , n379037 );
buf ( n379039 , n46397 );
not ( n379040 , n379039 );
buf ( n379041 , n41615 );
not ( n379042 , n379041 );
or ( n58554 , n379040 , n379042 );
buf ( n379044 , n41607 );
buf ( n58556 , n342909 );
nand ( n58557 , n379044 , n58556 );
buf ( n58558 , n58557 );
buf ( n379048 , n58558 );
nand ( n58560 , n58554 , n379048 );
buf ( n379050 , n58560 );
and ( n58562 , n379050 , n365152 );
and ( n379052 , n377745 , n45018 );
nor ( n379053 , n58562 , n379052 );
buf ( n379054 , n379053 );
not ( n58566 , n379054 );
buf ( n379056 , n58566 );
buf ( n379057 , n379056 );
xor ( n58569 , n379038 , n379057 );
buf ( n379059 , n58569 );
buf ( n379060 , n379059 );
xor ( n58572 , n58462 , n379060 );
buf ( n379062 , n58572 );
buf ( n379063 , n379062 );
xor ( n58575 , n378905 , n379063 );
buf ( n379065 , n58575 );
buf ( n379066 , n379065 );
xor ( n58578 , n377240 , n377320 );
xor ( n379068 , n58578 , n377342 );
buf ( n379069 , n379068 );
xor ( n379070 , n378094 , n378102 );
and ( n58582 , n379070 , n378119 );
and ( n379072 , n378094 , n378102 );
or ( n379073 , n58582 , n379072 );
buf ( n379074 , n379073 );
buf ( n379075 , n379074 );
xor ( n58587 , n379069 , n379075 );
buf ( n379077 , n364852 );
not ( n379078 , n45414 );
not ( n58590 , n368662 );
and ( n379080 , n379078 , n58590 );
buf ( n379081 , n369577 );
buf ( n379082 , n368662 );
and ( n58594 , n379081 , n379082 );
buf ( n379084 , n58594 );
nor ( n58596 , n379080 , n379084 );
buf ( n379086 , n58596 );
or ( n58598 , n379077 , n379086 );
buf ( n379088 , n365393 );
not ( n58600 , n379088 );
buf ( n379090 , n44717 );
not ( n379091 , n379090 );
or ( n58603 , n58600 , n379091 );
buf ( n379093 , n369577 );
buf ( n379094 , n365408 );
nand ( n58606 , n379093 , n379094 );
buf ( n379096 , n58606 );
buf ( n379097 , n379096 );
nand ( n58609 , n58603 , n379097 );
buf ( n58610 , n58609 );
buf ( n379100 , n58610 );
not ( n58612 , n379100 );
buf ( n58613 , n58612 );
buf ( n379103 , n58613 );
not ( n58615 , n366103 );
buf ( n379105 , n58615 );
or ( n379106 , n379103 , n379105 );
nand ( n379107 , n58598 , n379106 );
buf ( n379108 , n379107 );
not ( n379109 , n379108 );
buf ( n379110 , n378179 );
not ( n58622 , n379110 );
buf ( n379112 , n363428 );
not ( n379113 , n379112 );
or ( n58625 , n58622 , n379113 );
buf ( n379115 , n377693 );
buf ( n379116 , n57228 );
nand ( n58628 , n379115 , n379116 );
buf ( n379118 , n58628 );
buf ( n379119 , n379118 );
nand ( n58631 , n58625 , n379119 );
buf ( n58632 , n58631 );
buf ( n379122 , n58632 );
buf ( n379123 , n45553 );
not ( n379124 , n379123 );
buf ( n379125 , n377190 );
not ( n58637 , n379125 );
buf ( n379127 , n375903 );
not ( n58639 , n379127 );
or ( n58640 , n58637 , n58639 );
buf ( n58641 , n352192 );
buf ( n58642 , n365670 );
nand ( n58643 , n58641 , n58642 );
buf ( n58644 , n58643 );
buf ( n379134 , n58644 );
nand ( n58646 , n58640 , n379134 );
buf ( n379136 , n58646 );
buf ( n379137 , n379136 );
not ( n58649 , n379137 );
or ( n58650 , n379124 , n58649 );
not ( n58651 , n377190 );
not ( n58652 , n44637 );
or ( n58653 , n58651 , n58652 );
buf ( n379143 , n351317 );
buf ( n379144 , n365670 );
nand ( n58656 , n379143 , n379144 );
buf ( n379146 , n58656 );
nand ( n58658 , n58653 , n379146 );
nand ( n58659 , n58658 , n56794 );
buf ( n379149 , n58659 );
nand ( n58661 , n58650 , n379149 );
buf ( n379151 , n58661 );
buf ( n379152 , n379151 );
xor ( n379153 , n379122 , n379152 );
xor ( n58665 , n378319 , n378328 );
and ( n58666 , n58665 , n378518 );
and ( n379156 , n378319 , n378328 );
or ( n58668 , n58666 , n379156 );
buf ( n379158 , n58668 );
buf ( n379159 , n377009 );
not ( n58671 , n379159 );
buf ( n379161 , n377019 );
not ( n379162 , n379161 );
buf ( n379163 , n377037 );
not ( n379164 , n379163 );
and ( n379165 , n379162 , n379164 );
buf ( n379166 , n377019 );
buf ( n379167 , n377037 );
and ( n379168 , n379166 , n379167 );
nor ( n379169 , n379165 , n379168 );
buf ( n379170 , n379169 );
buf ( n379171 , n379170 );
not ( n379172 , n379171 );
or ( n58684 , n58671 , n379172 );
buf ( n379174 , n379170 );
buf ( n379175 , n377009 );
or ( n58687 , n379174 , n379175 );
nand ( n58688 , n58684 , n58687 );
buf ( n379178 , n58688 );
or ( n58690 , n379158 , n379178 );
not ( n58691 , n58690 );
not ( n58692 , n378566 );
not ( n58693 , n370989 );
not ( n58694 , n58693 );
or ( n58695 , n58692 , n58694 );
not ( n379185 , n377263 );
nand ( n379186 , n379185 , n377171 );
nand ( n58698 , n58695 , n379186 );
not ( n58699 , n58698 );
or ( n379189 , n58691 , n58699 );
nand ( n379190 , n379158 , n379178 );
nand ( n58702 , n379189 , n379190 );
buf ( n379192 , n58702 );
xor ( n379193 , n379153 , n379192 );
buf ( n379194 , n379193 );
not ( n58706 , n379194 );
or ( n379196 , n379109 , n58706 );
buf ( n379197 , n56794 );
not ( n379198 , n379197 );
buf ( n379199 , n379136 );
not ( n379200 , n379199 );
or ( n379201 , n379198 , n379200 );
and ( n58713 , n352209 , n365670 );
not ( n58714 , n352209 );
and ( n379204 , n58714 , n377190 );
or ( n379205 , n58713 , n379204 );
buf ( n379206 , n379205 );
buf ( n379207 , n45553 );
nand ( n379208 , n379206 , n379207 );
buf ( n379209 , n379208 );
buf ( n379210 , n379209 );
nand ( n379211 , n379201 , n379210 );
buf ( n379212 , n379211 );
xnor ( n379213 , n379158 , n379178 );
not ( n379214 , n379213 );
not ( n58726 , n58698 );
or ( n58727 , n379214 , n58726 );
or ( n379217 , n58698 , n379213 );
nand ( n379218 , n58727 , n379217 );
or ( n379219 , n379212 , n379218 );
not ( n58731 , n379219 );
not ( n379221 , n377842 );
not ( n58733 , n377838 );
or ( n379223 , n379221 , n58733 );
not ( n379224 , n365980 );
not ( n58736 , n342335 );
or ( n379226 , n379224 , n58736 );
buf ( n379227 , n342338 );
buf ( n379228 , n365989 );
nand ( n58740 , n379227 , n379228 );
buf ( n379230 , n58740 );
nand ( n58742 , n379226 , n379230 );
nand ( n58743 , n58742 , n49669 );
nand ( n58744 , n379223 , n58743 );
not ( n58745 , n58744 );
or ( n58746 , n58731 , n58745 );
nand ( n58747 , n379218 , n379212 );
nand ( n379237 , n58746 , n58747 );
not ( n379238 , n379237 );
nor ( n58750 , n379108 , n379194 );
or ( n379240 , n379238 , n58750 );
nand ( n379241 , n379196 , n379240 );
buf ( n379242 , n379241 );
and ( n58754 , n58587 , n379242 );
and ( n379244 , n379069 , n379075 );
or ( n379245 , n58754 , n379244 );
buf ( n379246 , n379245 );
buf ( n379247 , n379246 );
buf ( n379248 , n342352 );
not ( n379249 , n379248 );
buf ( n379250 , n379249 );
buf ( n379251 , n379250 );
not ( n58763 , n379251 );
buf ( n379253 , n58763 );
not ( n379254 , n379253 );
not ( n379255 , n379254 );
not ( n58767 , n342366 );
and ( n379257 , n379255 , n58767 );
and ( n379258 , n342366 , n379250 );
nor ( n58770 , n379257 , n379258 );
not ( n379260 , n58770 );
buf ( n379261 , n379260 );
buf ( n58773 , n379261 );
buf ( n379263 , n58773 );
buf ( n379264 , n379263 );
not ( n379265 , n379264 );
buf ( n379266 , n377571 );
not ( n58778 , n379266 );
buf ( n379268 , n58778 );
buf ( n58780 , n379268 );
buf ( n379270 , n58780 );
buf ( n379271 , n379270 );
buf ( n379272 , n379271 );
not ( n379273 , n379272 );
buf ( n379274 , n379273 );
and ( n379275 , n379274 , n370257 );
not ( n379276 , n379274 );
and ( n58788 , n379276 , n374422 );
or ( n379278 , n379275 , n58788 );
buf ( n379279 , n379278 );
not ( n58791 , n379279 );
or ( n58792 , n379265 , n58791 );
xor ( n379282 , n40199 , n379271 );
buf ( n379283 , n379282 );
not ( n58795 , n379283 );
buf ( n379285 , n342366 );
buf ( n379286 , n379285 );
buf ( n379287 , n379286 );
or ( n58799 , n379287 , n23104 );
buf ( n379289 , n23104 );
buf ( n379290 , n379287 );
nand ( n379291 , n379289 , n379290 );
buf ( n379292 , n379291 );
and ( n379293 , n58799 , n379292 , n58770 );
buf ( n379294 , n379293 );
not ( n379295 , n379294 );
buf ( n379296 , n379295 );
buf ( n379297 , n379296 );
not ( n58809 , n379297 );
buf ( n379299 , n58809 );
buf ( n379300 , n379299 );
nand ( n379301 , n58795 , n379300 );
buf ( n379302 , n379301 );
buf ( n379303 , n379302 );
nand ( n58815 , n58792 , n379303 );
buf ( n379305 , n58815 );
buf ( n379306 , n379305 );
xor ( n58818 , n379247 , n379306 );
buf ( n379308 , n340745 );
buf ( n379309 , n340684 );
nand ( n58821 , n379308 , n379309 );
buf ( n379311 , n58821 );
buf ( n379312 , n379311 );
buf ( n379313 , n340733 );
xnor ( n379314 , n379312 , n379313 );
buf ( n379315 , n379314 );
buf ( n379316 , n379315 );
not ( n379317 , n379316 );
buf ( n379318 , n379317 );
buf ( n379319 , n379318 );
xor ( n379320 , n340690 , n340715 );
xor ( n379321 , n379320 , n340729 );
buf ( n379322 , n379321 );
buf ( n379323 , n379322 );
not ( n58835 , n379323 );
buf ( n379325 , n58835 );
buf ( n379326 , n379325 );
nand ( n58838 , n379319 , n379326 );
buf ( n379328 , n58838 );
buf ( n379329 , n379328 );
buf ( n379330 , n379322 );
buf ( n379331 , n379315 );
nand ( n379332 , n379330 , n379331 );
buf ( n379333 , n379332 );
buf ( n379334 , n379333 );
buf ( n379335 , n20822 );
buf ( n379336 , n340711 );
and ( n379337 , n379335 , n379336 );
buf ( n379338 , n379337 );
nor ( n379339 , n340714 , n379338 );
buf ( n379340 , n379339 );
buf ( n379341 , n379325 );
and ( n58853 , n379340 , n379341 );
not ( n379343 , n379340 );
buf ( n379344 , n379322 );
and ( n58856 , n379343 , n379344 );
nor ( n58857 , n58853 , n58856 );
buf ( n379347 , n58857 );
buf ( n379348 , n379347 );
nand ( n379349 , n379329 , n379334 , n379348 );
buf ( n379350 , n379349 );
buf ( n379351 , n379350 );
not ( n379352 , n379351 );
buf ( n379353 , n379352 );
buf ( n379354 , n379353 );
buf ( n58866 , n379354 );
buf ( n58867 , n58866 );
buf ( n379357 , n58867 );
not ( n58869 , n379357 );
buf ( n379359 , n58869 );
not ( n58871 , n379359 );
buf ( n379361 , n58871 );
not ( n58873 , n379361 );
buf ( n379363 , n379318 );
buf ( n58875 , n379363 );
buf ( n379365 , n58875 );
buf ( n379366 , n379365 );
not ( n58878 , n379366 );
buf ( n379368 , n58878 );
buf ( n379369 , n379368 );
buf ( n379370 , n379369 );
buf ( n379371 , n379370 );
buf ( n379372 , n379371 );
not ( n379373 , n379372 );
buf ( n379374 , n363172 );
not ( n58886 , n379374 );
or ( n379376 , n379373 , n58886 );
buf ( n58888 , n363171 );
buf ( n379378 , n379371 );
not ( n379379 , n379378 );
buf ( n379380 , n379379 );
buf ( n379381 , n379380 );
nand ( n58893 , n58888 , n379381 );
buf ( n58894 , n58893 );
buf ( n379384 , n58894 );
nand ( n58896 , n379376 , n379384 );
buf ( n58897 , n58896 );
buf ( n379387 , n58897 );
not ( n58899 , n379387 );
or ( n379389 , n58873 , n58899 );
buf ( n379390 , n379371 );
not ( n58902 , n379390 );
buf ( n379392 , n58902 );
buf ( n379393 , n379392 );
not ( n58905 , n379393 );
buf ( n379395 , n365167 );
not ( n379396 , n379395 );
or ( n58908 , n58905 , n379396 );
buf ( n379398 , n360110 );
not ( n379399 , n379398 );
buf ( n379400 , n379371 );
nand ( n58912 , n379399 , n379400 );
buf ( n58913 , n58912 );
buf ( n379403 , n58913 );
nand ( n58915 , n58908 , n379403 );
buf ( n58916 , n58915 );
buf ( n58917 , n58916 );
buf ( n379407 , n379347 );
not ( n58919 , n379407 );
buf ( n58920 , n58919 );
buf ( n379410 , n58920 );
buf ( n58922 , n379410 );
buf ( n58923 , n58922 );
buf ( n379413 , n58923 );
nand ( n58925 , n58917 , n379413 );
buf ( n58926 , n58925 );
buf ( n58927 , n58926 );
nand ( n58928 , n379389 , n58927 );
buf ( n58929 , n58928 );
buf ( n58930 , n58929 );
and ( n58931 , n58818 , n58930 );
and ( n58932 , n379247 , n379306 );
or ( n58933 , n58931 , n58932 );
buf ( n58934 , n58933 );
buf ( n379424 , n58934 );
and ( n58936 , n379066 , n379424 );
not ( n58937 , n379066 );
buf ( n379427 , n58934 );
not ( n379428 , n379427 );
buf ( n379429 , n379428 );
buf ( n379430 , n379429 );
and ( n379431 , n58937 , n379430 );
nor ( n58943 , n58936 , n379431 );
buf ( n379433 , n58943 );
and ( n58945 , n378671 , n379433 );
not ( n379435 , n378671 );
not ( n379436 , n379433 );
and ( n58948 , n379435 , n379436 );
nor ( n379438 , n58945 , n58948 );
not ( n379439 , n379438 );
not ( n379440 , n379439 );
buf ( n379441 , n379282 );
not ( n58953 , n379441 );
buf ( n379443 , n379263 );
not ( n379444 , n379443 );
buf ( n379445 , n379444 );
buf ( n379446 , n379445 );
not ( n379447 , n379446 );
and ( n379448 , n58953 , n379447 );
and ( n379449 , n366722 , n379271 );
not ( n58961 , n366722 );
and ( n379451 , n58961 , n379274 );
or ( n379452 , n379449 , n379451 );
buf ( n379453 , n379452 );
buf ( n379454 , n379299 );
and ( n379455 , n379453 , n379454 );
nor ( n379456 , n379448 , n379455 );
buf ( n379457 , n379456 );
not ( n379458 , n379457 );
buf ( n379459 , n377130 );
buf ( n379460 , n377116 );
or ( n379461 , n379459 , n379460 );
not ( n58973 , n349202 );
buf ( n379463 , n349117 );
not ( n379464 , n379463 );
buf ( n379465 , n349211 );
nand ( n379466 , n379464 , n379465 );
buf ( n379467 , n379466 );
not ( n379468 , n379467 );
or ( n379469 , n58973 , n379468 );
not ( n58981 , n379467 );
nand ( n379471 , n58981 , n349205 );
nand ( n379472 , n379469 , n379471 );
buf ( n58984 , n379472 );
buf ( n379474 , n58984 );
not ( n379475 , n379474 );
buf ( n379476 , n360154 );
not ( n58988 , n379476 );
or ( n379478 , n379475 , n58988 );
buf ( n379479 , n360065 );
buf ( n379480 , n58984 );
not ( n379481 , n379480 );
buf ( n379482 , n379481 );
buf ( n379483 , n379482 );
nand ( n58995 , n379479 , n379483 );
buf ( n58996 , n58995 );
buf ( n379486 , n58996 );
nand ( n58998 , n379478 , n379486 );
buf ( n58999 , n58998 );
buf ( n379489 , n58999 );
buf ( n379490 , n377116 );
buf ( n379491 , n360164 );
nand ( n379492 , n379489 , n379490 , n379491 );
buf ( n379493 , n379492 );
buf ( n379494 , n379493 );
nand ( n379495 , n379461 , n379494 );
buf ( n379496 , n379495 );
buf ( n379497 , n379496 );
not ( n59009 , n377782 );
not ( n379499 , n366277 );
or ( n379500 , n59009 , n379499 );
nand ( n59012 , n366151 , n377779 );
nand ( n379502 , n379500 , n59012 );
not ( n379503 , n379502 );
not ( n59015 , n366161 );
or ( n59016 , n379503 , n59015 );
buf ( n379506 , n377365 );
buf ( n59018 , n371732 );
nand ( n59019 , n379506 , n59018 );
buf ( n59020 , n59019 );
nand ( n379510 , n59016 , n59020 );
buf ( n379511 , n379510 );
xor ( n59023 , n379497 , n379511 );
buf ( n379513 , n378098 );
not ( n379514 , n379513 );
buf ( n379515 , n379514 );
buf ( n379516 , n379515 );
buf ( n379517 , n361631 );
and ( n59029 , n379516 , n379517 );
not ( n379519 , n379516 );
buf ( n379520 , n45234 );
and ( n59032 , n379519 , n379520 );
nor ( n59033 , n59029 , n59032 );
buf ( n379523 , n59033 );
buf ( n379524 , n379523 );
not ( n379525 , n379524 );
buf ( n379526 , n39701 );
not ( n379527 , n379526 );
or ( n379528 , n379525 , n379527 );
nand ( n59040 , n367796 , n377109 );
buf ( n379530 , n59040 );
nand ( n379531 , n379528 , n379530 );
buf ( n379532 , n379531 );
buf ( n379533 , n379532 );
xnor ( n379534 , n59023 , n379533 );
buf ( n379535 , n379534 );
not ( n379536 , n379535 );
and ( n379537 , n379458 , n379536 );
xor ( n59049 , n377696 , n377702 );
xor ( n379539 , n59049 , n377721 );
buf ( n379540 , n379539 );
buf ( n379541 , n379540 );
not ( n379542 , n379541 );
buf ( n379543 , n379542 );
buf ( n379544 , n379543 );
xor ( n59056 , n362534 , n377728 );
not ( n59057 , n59056 );
not ( n59058 , n365187 );
not ( n59059 , n59058 );
and ( n59060 , n59057 , n59059 );
and ( n379550 , n377731 , n365152 );
nor ( n59062 , n59060 , n379550 );
buf ( n379552 , n59062 );
not ( n59064 , n379552 );
buf ( n379554 , n59064 );
buf ( n379555 , n379554 );
xor ( n59067 , n379544 , n379555 );
xor ( n59068 , n377845 , n377870 );
and ( n379558 , n59068 , n377898 );
and ( n379559 , n377845 , n377870 );
or ( n59071 , n379558 , n379559 );
buf ( n379561 , n59071 );
buf ( n379562 , n379561 );
xor ( n379563 , n59067 , n379562 );
buf ( n379564 , n379563 );
buf ( n379565 , n379457 );
buf ( n379566 , n379535 );
nand ( n59078 , n379565 , n379566 );
buf ( n59079 , n59078 );
and ( n379569 , n379564 , n59079 );
nor ( n59081 , n379537 , n379569 );
not ( n379571 , n59081 );
not ( n379572 , n379571 );
buf ( n379573 , n369444 );
not ( n379574 , n379573 );
buf ( n379575 , n377658 );
not ( n379576 , n379575 );
or ( n59088 , n379574 , n379576 );
buf ( n59089 , n46031 );
buf ( n379579 , n368554 );
nand ( n379580 , n59089 , n379579 );
buf ( n379581 , n379580 );
not ( n59093 , n379581 );
nand ( n379583 , n368549 , n369343 );
not ( n379584 , n379583 );
or ( n59096 , n59093 , n379584 );
nand ( n379586 , n59096 , n368611 );
buf ( n379587 , n379586 );
nand ( n59099 , n59088 , n379587 );
buf ( n379589 , n59099 );
buf ( n379590 , n379589 );
not ( n379591 , n379590 );
not ( n379592 , n375853 );
not ( n59104 , n369813 );
and ( n379594 , n379592 , n59104 );
buf ( n379595 , n369769 );
not ( n59107 , n379595 );
buf ( n379597 , n362288 );
not ( n59109 , n379597 );
or ( n59110 , n59107 , n59109 );
buf ( n379600 , n362285 );
buf ( n379601 , n369766 );
nand ( n59113 , n379600 , n379601 );
buf ( n379603 , n59113 );
buf ( n379604 , n379603 );
nand ( n59116 , n59110 , n379604 );
buf ( n379606 , n59116 );
and ( n59118 , n379606 , n369804 );
nor ( n59119 , n379594 , n59118 );
buf ( n379609 , n59119 );
not ( n59121 , n379609 );
buf ( n379611 , n59121 );
buf ( n379612 , n379611 );
not ( n59124 , n379612 );
or ( n379614 , n379591 , n59124 );
buf ( n379615 , n59119 );
not ( n59127 , n379615 );
buf ( n379617 , n379589 );
not ( n59129 , n379617 );
buf ( n59130 , n59129 );
buf ( n379620 , n59130 );
not ( n59132 , n379620 );
or ( n379622 , n59127 , n59132 );
buf ( n379623 , n369374 );
not ( n59135 , n379623 );
buf ( n379625 , n365626 );
not ( n59137 , n379625 );
or ( n59138 , n59135 , n59137 );
buf ( n379628 , n41892 );
buf ( n379629 , n49178 );
nand ( n59141 , n379628 , n379629 );
buf ( n379631 , n59141 );
buf ( n379632 , n379631 );
nand ( n59144 , n59138 , n379632 );
buf ( n59145 , n59144 );
buf ( n379635 , n59145 );
not ( n59147 , n379635 );
buf ( n379637 , n362027 );
not ( n379638 , n379637 );
or ( n59150 , n59147 , n379638 );
or ( n59151 , n370311 , n368994 );
nand ( n379641 , n368994 , n362033 );
nand ( n59153 , n59151 , n379641 );
buf ( n379643 , n59153 );
not ( n379644 , n379643 );
buf ( n379645 , n364824 );
nand ( n379646 , n379644 , n379645 );
buf ( n379647 , n379646 );
buf ( n379648 , n379647 );
nand ( n59160 , n59150 , n379648 );
buf ( n379650 , n59160 );
buf ( n379651 , n379650 );
not ( n59163 , n379651 );
buf ( n379653 , n377757 );
not ( n379654 , n379653 );
buf ( n379655 , n45270 );
not ( n379656 , n379655 );
or ( n59168 , n379654 , n379656 );
buf ( n379658 , n362452 );
buf ( n379659 , n378886 );
nand ( n379660 , n379658 , n379659 );
buf ( n379661 , n379660 );
buf ( n379662 , n379661 );
nand ( n59174 , n59168 , n379662 );
buf ( n379664 , n59174 );
buf ( n379665 , n379664 );
not ( n59177 , n379665 );
buf ( n379667 , n377370 );
not ( n59179 , n379667 );
or ( n379669 , n59177 , n59179 );
buf ( n379670 , n379502 );
buf ( n379671 , n366751 );
nand ( n379672 , n379670 , n379671 );
buf ( n379673 , n379672 );
buf ( n379674 , n379673 );
nand ( n379675 , n379669 , n379674 );
buf ( n379676 , n379675 );
buf ( n379677 , n379676 );
not ( n379678 , n379677 );
or ( n379679 , n59163 , n379678 );
buf ( n379680 , n379676 );
buf ( n379681 , n379650 );
or ( n379682 , n379680 , n379681 );
buf ( n379683 , n378856 );
not ( n59195 , n379683 );
buf ( n379685 , n370845 );
not ( n59197 , n379685 );
or ( n59198 , n59195 , n59197 );
buf ( n379688 , n365507 );
buf ( n379689 , n378847 );
nand ( n59201 , n379688 , n379689 );
buf ( n379691 , n59201 );
buf ( n379692 , n379691 );
nand ( n379693 , n59198 , n379692 );
buf ( n379694 , n379693 );
buf ( n379695 , n379694 );
not ( n379696 , n379695 );
buf ( n379697 , n40058 );
not ( n59209 , n379697 );
or ( n59210 , n379696 , n59209 );
buf ( n379700 , n365486 );
buf ( n379701 , n58999 );
nand ( n59213 , n379700 , n379701 );
buf ( n379703 , n59213 );
buf ( n379704 , n379703 );
nand ( n59216 , n59210 , n379704 );
buf ( n379706 , n59216 );
buf ( n379707 , n379706 );
nand ( n379708 , n379682 , n379707 );
buf ( n379709 , n379708 );
buf ( n379710 , n379709 );
nand ( n59222 , n379679 , n379710 );
buf ( n379712 , n59222 );
buf ( n379713 , n379712 );
nand ( n59225 , n379622 , n379713 );
buf ( n379715 , n59225 );
buf ( n379716 , n379715 );
nand ( n59228 , n379614 , n379716 );
buf ( n379718 , n59228 );
not ( n59230 , n379718 );
or ( n379720 , n379572 , n59230 );
buf ( n379721 , n379718 );
not ( n59233 , n379721 );
buf ( n379723 , n59233 );
not ( n59235 , n379723 );
not ( n59236 , n59081 );
or ( n59237 , n59235 , n59236 );
not ( n59238 , n366025 );
buf ( n379728 , n56970 );
not ( n379729 , n379728 );
buf ( n379730 , n365290 );
not ( n379731 , n379730 );
or ( n379732 , n379729 , n379731 );
buf ( n379733 , n365266 );
buf ( n379734 , n377389 );
nand ( n59246 , n379733 , n379734 );
buf ( n379736 , n59246 );
buf ( n379737 , n379736 );
nand ( n379738 , n379732 , n379737 );
buf ( n379739 , n379738 );
not ( n379740 , n379739 );
or ( n379741 , n59238 , n379740 );
buf ( n379742 , n369374 );
not ( n379743 , n379742 );
buf ( n379744 , n365290 );
not ( n379745 , n379744 );
or ( n59257 , n379743 , n379745 );
buf ( n379747 , n45091 );
buf ( n379748 , n49178 );
nand ( n59260 , n379747 , n379748 );
buf ( n379750 , n59260 );
buf ( n379751 , n379750 );
nand ( n379752 , n59257 , n379751 );
buf ( n379753 , n379752 );
nand ( n59265 , n365303 , n379753 );
nand ( n379755 , n379741 , n59265 );
not ( n59267 , n379755 );
not ( n379757 , n41882 );
not ( n59269 , n59153 );
and ( n379759 , n379757 , n59269 );
buf ( n379760 , n368665 );
not ( n59272 , n379760 );
buf ( n379762 , n364832 );
not ( n379763 , n379762 );
or ( n59275 , n59272 , n379763 );
buf ( n379765 , n362033 );
buf ( n379766 , n368662 );
nand ( n59278 , n379765 , n379766 );
buf ( n59279 , n59278 );
buf ( n379769 , n59279 );
nand ( n59281 , n59275 , n379769 );
buf ( n379771 , n59281 );
buf ( n379772 , n379771 );
not ( n379773 , n379772 );
buf ( n379774 , n364821 );
nor ( n379775 , n379773 , n379774 );
buf ( n379776 , n379775 );
nor ( n59288 , n379759 , n379776 );
buf ( n59289 , n59288 );
not ( n59290 , n59289 );
buf ( n59291 , n59290 );
not ( n379781 , n59291 );
or ( n379782 , n59267 , n379781 );
not ( n59294 , n59288 );
buf ( n379784 , n379755 );
not ( n379785 , n379784 );
buf ( n379786 , n379785 );
not ( n379787 , n379786 );
or ( n379788 , n59294 , n379787 );
buf ( n379789 , n377935 );
not ( n59301 , n379789 );
buf ( n379791 , n366989 );
not ( n59303 , n379791 );
or ( n59304 , n59301 , n59303 );
buf ( n379794 , n377765 );
not ( n59306 , n379794 );
buf ( n379796 , n359312 );
nand ( n59308 , n59306 , n379796 );
buf ( n379798 , n59308 );
buf ( n379799 , n379798 );
nand ( n59311 , n59304 , n379799 );
buf ( n379801 , n59311 );
nand ( n379802 , n379788 , n379801 );
nand ( n379803 , n379782 , n379802 );
not ( n59315 , n379543 );
not ( n379805 , n379554 );
or ( n379806 , n59315 , n379805 );
not ( n59318 , n379540 );
not ( n379808 , n59062 );
or ( n59320 , n59318 , n379808 );
nand ( n59321 , n59320 , n379561 );
nand ( n379811 , n379806 , n59321 );
xor ( n379812 , n379803 , n379811 );
not ( n59324 , n379510 );
buf ( n379814 , n379496 );
not ( n379815 , n379814 );
buf ( n379816 , n379815 );
nand ( n379817 , n59324 , n379816 );
not ( n59329 , n379817 );
not ( n59330 , n379532 );
or ( n59331 , n59329 , n59330 );
not ( n59332 , n379816 );
nand ( n59333 , n59332 , n379510 );
nand ( n59334 , n59331 , n59333 );
xor ( n59335 , n379812 , n59334 );
nand ( n59336 , n59237 , n59335 );
nand ( n59337 , n379720 , n59336 );
buf ( n379827 , n59337 );
not ( n59339 , n379827 );
buf ( n379829 , n59339 );
buf ( n379830 , n379829 );
not ( n59342 , n379830 );
buf ( n379832 , n59342 );
buf ( n379833 , n379832 );
not ( n379834 , n379833 );
buf ( n379835 , n371254 );
buf ( n379836 , n379253 );
buf ( n59348 , n379836 );
buf ( n379838 , n59348 );
buf ( n59350 , n379838 );
buf ( n379840 , n59350 );
buf ( n379841 , n379840 );
buf ( n379842 , n379841 );
and ( n379843 , n379835 , n379842 );
buf ( n379844 , n359974 );
buf ( n379845 , n379841 );
not ( n379846 , n379845 );
buf ( n379847 , n379846 );
buf ( n379848 , n379847 );
and ( n59360 , n379844 , n379848 );
nor ( n59361 , n379843 , n59360 );
buf ( n379851 , n59361 );
buf ( n379852 , n379851 );
not ( n59364 , n379852 );
buf ( n379854 , n379318 );
not ( n379855 , n379854 );
buf ( n379856 , n379855 );
buf ( n379857 , n379856 );
not ( n379858 , n379857 );
buf ( n379859 , n379858 );
buf ( n379860 , n379859 );
not ( n379861 , n379860 );
buf ( n379862 , n340648 );
buf ( n379863 , n340653 );
nand ( n379864 , n379862 , n379863 );
buf ( n379865 , n379864 );
buf ( n379866 , n379865 );
buf ( n379867 , n20858 );
not ( n379868 , n379867 );
buf ( n379869 , n379868 );
buf ( n379870 , n379869 );
and ( n379871 , n379866 , n379870 );
not ( n59383 , n379866 );
buf ( n379873 , n20858 );
and ( n59385 , n59383 , n379873 );
nor ( n59386 , n379871 , n59385 );
buf ( n379876 , n59386 );
buf ( n379877 , n379876 );
not ( n59389 , n379877 );
and ( n379879 , n379861 , n59389 );
buf ( n59391 , n379876 );
buf ( n379881 , n379859 );
and ( n379882 , n59391 , n379881 );
nor ( n379883 , n379879 , n379882 );
buf ( n379884 , n379883 );
buf ( n379885 , n379884 );
not ( n59397 , n379885 );
buf ( n379887 , n59397 );
buf ( n379888 , n379887 );
buf ( n59400 , n379888 );
buf ( n379890 , n59400 );
buf ( n379891 , n379890 );
not ( n379892 , n379891 );
buf ( n379893 , n379892 );
buf ( n379894 , n379893 );
not ( n379895 , n379894 );
and ( n59407 , n59364 , n379895 );
buf ( n379897 , n379841 );
not ( n379898 , n379897 );
buf ( n379899 , n366599 );
not ( n59411 , n379899 );
or ( n379901 , n379898 , n59411 );
buf ( n379902 , n359937 );
buf ( n379903 , n379847 );
nand ( n379904 , n379902 , n379903 );
buf ( n379905 , n379904 );
buf ( n379906 , n379905 );
nand ( n59418 , n379901 , n379906 );
buf ( n59419 , n59418 );
buf ( n59420 , n59419 );
xor ( n59421 , n342352 , n379876 );
nand ( n379911 , n59421 , n379884 );
not ( n379912 , n379911 );
not ( n59424 , n379912 );
buf ( n379914 , n59424 );
not ( n59426 , n379914 );
buf ( n379916 , n59426 );
buf ( n379917 , n379916 );
and ( n59429 , n59420 , n379917 );
nor ( n59430 , n59407 , n59429 );
buf ( n379920 , n59430 );
not ( n59432 , n379920 );
not ( n59433 , n59432 );
not ( n59434 , n58923 );
not ( n59435 , n379392 );
not ( n59436 , n40090 );
or ( n379926 , n59435 , n59436 );
nand ( n59438 , n41472 , n379371 );
nand ( n379928 , n379926 , n59438 );
not ( n59440 , n379928 );
or ( n59441 , n59434 , n59440 );
buf ( n379931 , n58916 );
buf ( n379932 , n58867 );
nand ( n59444 , n379931 , n379932 );
buf ( n379934 , n59444 );
nand ( n59446 , n59441 , n379934 );
not ( n59447 , n59446 );
not ( n59448 , n59447 );
not ( n59449 , n59448 );
or ( n379939 , n59433 , n59449 );
nand ( n59451 , n59447 , n379920 );
nand ( n59452 , n379939 , n59451 );
buf ( n379942 , n379445 );
not ( n379943 , n379942 );
buf ( n379944 , n379943 );
not ( n59456 , n379944 );
buf ( n379946 , n379274 );
not ( n379947 , n379946 );
buf ( n379948 , n362208 );
not ( n379949 , n379948 );
or ( n379950 , n379947 , n379949 );
buf ( n379951 , n44926 );
buf ( n379952 , n379271 );
nand ( n59464 , n379951 , n379952 );
buf ( n379954 , n59464 );
buf ( n379955 , n379954 );
nand ( n59467 , n379950 , n379955 );
buf ( n59468 , n59467 );
not ( n59469 , n59468 );
or ( n59470 , n59456 , n59469 );
buf ( n379960 , n379296 );
not ( n59472 , n379960 );
buf ( n379962 , n59472 );
nand ( n59474 , n379278 , n379962 );
nand ( n59475 , n59470 , n59474 );
xor ( n379965 , n59452 , n59475 );
not ( n379966 , n379965 );
buf ( n379967 , n352268 );
not ( n379968 , n379967 );
buf ( n379969 , n364763 );
not ( n59481 , n379969 );
or ( n379971 , n379968 , n59481 );
buf ( n379972 , n46303 );
not ( n59484 , n379972 );
buf ( n379974 , n366329 );
nand ( n379975 , n59484 , n379974 );
buf ( n379976 , n379975 );
buf ( n379977 , n379976 );
nand ( n59489 , n379971 , n379977 );
buf ( n379979 , n59489 );
buf ( n379980 , n379979 );
not ( n59492 , n379980 );
buf ( n379982 , n366315 );
not ( n59494 , n379982 );
or ( n59495 , n59492 , n59494 );
buf ( n59496 , n377446 );
buf ( n59497 , n41834 );
nand ( n59498 , n59496 , n59497 );
buf ( n59499 , n59498 );
buf ( n379989 , n59499 );
nand ( n59501 , n59495 , n379989 );
buf ( n379991 , n59501 );
not ( n59503 , n379991 );
not ( n59504 , n365115 );
not ( n379994 , n377528 );
or ( n379995 , n59504 , n379994 );
buf ( n379996 , n56921 );
buf ( n379997 , n365030 );
nand ( n379998 , n379996 , n379997 );
buf ( n379999 , n379998 );
nand ( n380000 , n379995 , n379999 );
not ( n59512 , n380000 );
nand ( n59513 , n59503 , n59512 );
not ( n380003 , n59513 );
buf ( n380004 , n45075 );
not ( n380005 , n380004 );
buf ( n380006 , n378781 );
not ( n59518 , n380006 );
or ( n380008 , n380005 , n59518 );
and ( n380009 , n32084 , n365202 );
not ( n59521 , n32084 );
and ( n380011 , n59521 , n342881 );
or ( n380012 , n380009 , n380011 );
buf ( n380013 , n380012 );
buf ( n380014 , n365226 );
nand ( n59526 , n380013 , n380014 );
buf ( n380016 , n59526 );
buf ( n380017 , n380016 );
nand ( n380018 , n380008 , n380017 );
buf ( n380019 , n380018 );
not ( n59531 , n380019 );
or ( n380021 , n380003 , n59531 );
buf ( n380022 , n59512 );
not ( n59534 , n380022 );
buf ( n380024 , n379979 );
not ( n380025 , n380024 );
buf ( n380026 , n366315 );
not ( n380027 , n380026 );
or ( n59539 , n380025 , n380027 );
buf ( n380029 , n59499 );
nand ( n59541 , n59539 , n380029 );
buf ( n380031 , n59541 );
buf ( n380032 , n380031 );
nand ( n59544 , n59534 , n380032 );
buf ( n380034 , n59544 );
nand ( n59546 , n380021 , n380034 );
buf ( n380036 , n58984 );
not ( n59548 , n380036 );
buf ( n380038 , n364919 );
not ( n59550 , n380038 );
or ( n380040 , n59548 , n59550 );
buf ( n380041 , n359944 );
buf ( n380042 , n379482 );
nand ( n380043 , n380041 , n380042 );
buf ( n380044 , n380043 );
buf ( n380045 , n380044 );
nand ( n380046 , n380040 , n380045 );
buf ( n380047 , n380046 );
buf ( n380048 , n380047 );
not ( n380049 , n380048 );
buf ( n380050 , n366226 );
not ( n380051 , n380050 );
or ( n380052 , n380049 , n380051 );
buf ( n380053 , n359993 );
buf ( n380054 , n377122 );
not ( n380055 , n380054 );
buf ( n380056 , n359947 );
not ( n380057 , n380056 );
or ( n380058 , n380055 , n380057 );
buf ( n380059 , n359944 );
buf ( n380060 , n57463 );
nand ( n380061 , n380059 , n380060 );
buf ( n380062 , n380061 );
buf ( n380063 , n380062 );
nand ( n380064 , n380058 , n380063 );
buf ( n380065 , n380064 );
buf ( n380066 , n380065 );
nand ( n380067 , n380053 , n380066 );
buf ( n380068 , n380067 );
buf ( n380069 , n380068 );
nand ( n380070 , n380052 , n380069 );
buf ( n380071 , n380070 );
xor ( n380072 , n59546 , n380071 );
buf ( n380073 , n379771 );
not ( n380074 , n380073 );
buf ( n380075 , n45438 );
not ( n59564 , n380075 );
or ( n380077 , n380074 , n59564 );
buf ( n380078 , n41915 );
buf ( n380079 , n377467 );
nand ( n59568 , n380078 , n380079 );
buf ( n380081 , n59568 );
buf ( n380082 , n380081 );
nand ( n59571 , n380077 , n380082 );
buf ( n380084 , n59571 );
buf ( n380085 , n380084 );
buf ( n380086 , n365428 );
not ( n380087 , n380086 );
buf ( n380088 , n44717 );
not ( n380089 , n380088 );
or ( n380090 , n380087 , n380089 );
buf ( n380091 , n45908 );
buf ( n380092 , n365422 );
nand ( n380093 , n380091 , n380092 );
buf ( n380094 , n380093 );
buf ( n380095 , n380094 );
nand ( n380096 , n380090 , n380095 );
buf ( n380097 , n380096 );
buf ( n380098 , n380097 );
not ( n59587 , n380098 );
not ( n59588 , n364848 );
buf ( n380101 , n59588 );
not ( n59590 , n380101 );
or ( n59591 , n59587 , n59590 );
nand ( n59592 , n377553 , n367590 );
buf ( n380105 , n59592 );
nand ( n380106 , n59591 , n380105 );
buf ( n380107 , n380106 );
buf ( n380108 , n380107 );
xor ( n380109 , n380085 , n380108 );
buf ( n380110 , n379753 );
not ( n380111 , n380110 );
buf ( n380112 , n366025 );
not ( n59601 , n380112 );
or ( n59602 , n380111 , n59601 );
buf ( n59603 , n40923 );
buf ( n380116 , n377489 );
nand ( n59605 , n59603 , n380116 );
buf ( n59606 , n59605 );
buf ( n380119 , n59606 );
nand ( n59608 , n59602 , n380119 );
buf ( n380121 , n59608 );
buf ( n380122 , n380121 );
and ( n380123 , n380109 , n380122 );
and ( n380124 , n380085 , n380108 );
or ( n59612 , n380123 , n380124 );
buf ( n380126 , n59612 );
xor ( n59614 , n380072 , n380126 );
xor ( n380128 , n380085 , n380108 );
xor ( n59616 , n380128 , n380122 );
buf ( n380130 , n59616 );
not ( n59618 , n380130 );
buf ( n380132 , n380000 );
buf ( n380133 , n379991 );
xor ( n59621 , n380132 , n380133 );
buf ( n380135 , n380019 );
xnor ( n380136 , n59621 , n380135 );
buf ( n380137 , n380136 );
buf ( n380138 , n380137 );
not ( n59626 , n365041 );
not ( n380140 , n361802 );
or ( n380141 , n59626 , n380140 );
not ( n59629 , n365041 );
nand ( n59630 , n59629 , n367453 );
nand ( n380144 , n380141 , n59630 );
buf ( n380145 , n380144 );
not ( n380146 , n380145 );
buf ( n380147 , n365083 );
not ( n59635 , n380147 );
and ( n380149 , n380146 , n59635 );
buf ( n380150 , n365041 );
not ( n59638 , n380150 );
buf ( n380152 , n41615 );
not ( n380153 , n380152 );
or ( n59641 , n59638 , n380153 );
buf ( n380155 , n41607 );
buf ( n380156 , n365052 );
nand ( n380157 , n380155 , n380156 );
buf ( n380158 , n380157 );
buf ( n380159 , n380158 );
nand ( n59647 , n59641 , n380159 );
buf ( n59648 , n59647 );
buf ( n59649 , n59648 );
buf ( n380163 , n47466 );
and ( n380164 , n59649 , n380163 );
nor ( n59652 , n380149 , n380164 );
buf ( n380166 , n59652 );
buf ( n380167 , n380166 );
nand ( n380168 , n380138 , n380167 );
buf ( n380169 , n380168 );
not ( n59657 , n380169 );
or ( n380171 , n59618 , n59657 );
buf ( n380172 , n380166 );
not ( n59660 , n380172 );
buf ( n59661 , n59660 );
buf ( n380175 , n59661 );
buf ( n380176 , n380137 );
not ( n380177 , n380176 );
buf ( n380178 , n380177 );
buf ( n380179 , n380178 );
nand ( n380180 , n380175 , n380179 );
buf ( n380181 , n380180 );
nand ( n59669 , n380171 , n380181 );
and ( n380183 , n59614 , n59669 );
not ( n380184 , n59614 );
not ( n59672 , n59669 );
and ( n380186 , n380184 , n59672 );
nor ( n380187 , n380183 , n380186 );
buf ( n380188 , n44915 );
not ( n380189 , n380188 );
xor ( n59677 , n365041 , n362130 );
buf ( n380191 , n59677 );
not ( n380192 , n380191 );
or ( n380193 , n380189 , n380192 );
not ( n59681 , n380144 );
nand ( n380195 , n59681 , n47466 );
buf ( n380196 , n380195 );
nand ( n380197 , n380193 , n380196 );
buf ( n380198 , n380197 );
buf ( n380199 , n380198 );
buf ( n380200 , n377159 );
not ( n380201 , n380200 );
buf ( n380202 , n377111 );
not ( n59690 , n380202 );
or ( n380204 , n380201 , n59690 );
buf ( n380205 , n377159 );
buf ( n380206 , n377111 );
or ( n380207 , n380205 , n380206 );
buf ( n380208 , n377061 );
nand ( n380209 , n380207 , n380208 );
buf ( n380210 , n380209 );
buf ( n380211 , n380210 );
nand ( n380212 , n380204 , n380211 );
buf ( n380213 , n380212 );
buf ( n380214 , n380213 );
xor ( n380215 , n380199 , n380214 );
nor ( n380216 , n377750 , n377791 );
or ( n59704 , n380216 , n377725 );
buf ( n380218 , n377791 );
buf ( n380219 , n377750 );
nand ( n59707 , n380218 , n380219 );
buf ( n380221 , n59707 );
nand ( n380222 , n59704 , n380221 );
buf ( n380223 , n380222 );
xor ( n59711 , n380215 , n380223 );
buf ( n380225 , n59711 );
and ( n380226 , n380187 , n380225 );
not ( n59714 , n380187 );
not ( n380228 , n380225 );
and ( n380229 , n59714 , n380228 );
nor ( n59717 , n380226 , n380229 );
not ( n59718 , n59717 );
not ( n59719 , n59718 );
or ( n380233 , n379966 , n59719 );
or ( n380234 , n59718 , n379965 );
nand ( n59722 , n380233 , n380234 );
buf ( n380236 , n59722 );
not ( n59724 , n380236 );
or ( n380238 , n379834 , n59724 );
buf ( n380239 , n379832 );
buf ( n380240 , n59722 );
or ( n380241 , n380239 , n380240 );
nand ( n59729 , n380238 , n380241 );
buf ( n380243 , n59729 );
buf ( n380244 , n44915 );
not ( n380245 , n380244 );
buf ( n380246 , n59648 );
not ( n59734 , n380246 );
or ( n59735 , n380245 , n59734 );
buf ( n380249 , n377971 );
buf ( n380250 , n47466 );
nand ( n59738 , n380249 , n380250 );
buf ( n380252 , n59738 );
buf ( n380253 , n380252 );
nand ( n59741 , n59735 , n380253 );
buf ( n59742 , n59741 );
not ( n59743 , n59742 );
xor ( n59744 , n379122 , n379152 );
and ( n59745 , n59744 , n379192 );
and ( n59746 , n379122 , n379152 );
or ( n59747 , n59745 , n59746 );
buf ( n380261 , n59747 );
not ( n59749 , n45075 );
not ( n59750 , n380012 );
or ( n59751 , n59749 , n59750 );
nand ( n59752 , n365226 , n377891 );
nand ( n59753 , n59751 , n59752 );
and ( n59754 , n380261 , n59753 );
not ( n59755 , n380261 );
nand ( n59756 , n380012 , n45075 );
and ( n380270 , n59756 , n59752 );
and ( n59758 , n59755 , n380270 );
nor ( n59759 , n59754 , n59758 );
buf ( n380273 , n59759 );
not ( n380274 , n366103 );
not ( n59762 , n380097 );
or ( n59763 , n380274 , n59762 );
buf ( n59764 , n361580 );
nand ( n59765 , n41482 , n58610 , n59764 );
nand ( n59766 , n59763 , n59765 );
buf ( n380280 , n59766 );
xor ( n380281 , n380273 , n380280 );
buf ( n380282 , n380281 );
not ( n59770 , n380282 );
not ( n380284 , n59770 );
or ( n59772 , n59743 , n380284 );
not ( n59773 , n59742 );
nand ( n380287 , n380282 , n59773 );
nand ( n380288 , n59772 , n380287 );
buf ( n380289 , n379786 );
not ( n380290 , n380289 );
buf ( n380291 , n59291 );
not ( n59779 , n380291 );
or ( n59780 , n380290 , n59779 );
buf ( n380294 , n379786 );
buf ( n380295 , n59291 );
or ( n59783 , n380294 , n380295 );
nand ( n59784 , n59780 , n59783 );
buf ( n380298 , n59784 );
xor ( n59786 , n379801 , n380298 );
buf ( n59787 , n59786 );
and ( n59788 , n380288 , n59787 );
not ( n59789 , n380288 );
not ( n380303 , n59787 );
and ( n59791 , n59789 , n380303 );
nor ( n59792 , n59788 , n59791 );
buf ( n59793 , n59792 );
not ( n59794 , n59793 );
buf ( n380308 , n379589 );
buf ( n380309 , n379611 );
xor ( n380310 , n380308 , n380309 );
buf ( n380311 , n379712 );
xnor ( n59799 , n380310 , n380311 );
buf ( n380313 , n59799 );
buf ( n380314 , n380313 );
not ( n59802 , n380314 );
buf ( n59803 , n59802 );
buf ( n380317 , n59803 );
not ( n59805 , n380317 );
or ( n380319 , n59794 , n59805 );
buf ( n380320 , n59792 );
not ( n59808 , n380320 );
buf ( n380322 , n59808 );
buf ( n59810 , n380322 );
not ( n59811 , n59810 );
buf ( n59812 , n380313 );
not ( n59813 , n59812 );
or ( n59814 , n59811 , n59813 );
buf ( n380328 , n49609 );
not ( n380329 , n380328 );
buf ( n380330 , n379606 );
not ( n380331 , n380330 );
or ( n380332 , n380329 , n380331 );
buf ( n380333 , n369769 );
not ( n380334 , n380333 );
buf ( n380335 , n369085 );
not ( n380336 , n380335 );
or ( n59824 , n380334 , n380336 );
buf ( n380338 , n362136 );
buf ( n380339 , n369766 );
nand ( n59827 , n380338 , n380339 );
buf ( n59828 , n59827 );
buf ( n380342 , n59828 );
nand ( n59830 , n59824 , n380342 );
buf ( n380344 , n59830 );
buf ( n59832 , n380344 );
buf ( n59833 , n369804 );
nand ( n59834 , n59832 , n59833 );
buf ( n59835 , n59834 );
buf ( n380349 , n59835 );
nand ( n59837 , n380332 , n380349 );
buf ( n380351 , n59837 );
buf ( n380352 , n380351 );
not ( n380353 , n340710 );
buf ( n380354 , n380353 );
buf ( n380355 , n380354 );
buf ( n380356 , n380355 );
buf ( n380357 , n380356 );
not ( n380358 , n380357 );
buf ( n380359 , n379339 );
not ( n380360 , n380359 );
buf ( n380361 , n380360 );
buf ( n380362 , n380361 );
buf ( n380363 , n380362 );
buf ( n380364 , n380363 );
buf ( n380365 , n380364 );
not ( n59853 , n380365 );
buf ( n380367 , n59853 );
buf ( n380368 , n380367 );
buf ( n380369 , n380368 );
not ( n380370 , n380369 );
buf ( n380371 , n40005 );
not ( n59859 , n380371 );
buf ( n59860 , n59859 );
buf ( n380374 , n59860 );
not ( n59862 , n380374 );
or ( n59863 , n380370 , n59862 );
buf ( n380377 , n365167 );
buf ( n59865 , n380368 );
not ( n59866 , n59865 );
buf ( n59867 , n59866 );
buf ( n380381 , n59867 );
nand ( n59869 , n380377 , n380381 );
buf ( n380383 , n59869 );
buf ( n380384 , n380383 );
nand ( n59872 , n59863 , n380384 );
buf ( n59873 , n59872 );
buf ( n380387 , n59873 );
not ( n59875 , n380387 );
or ( n380389 , n380358 , n59875 );
and ( n59877 , n372458 , n380368 );
not ( n59878 , n372458 );
and ( n380392 , n59878 , n59867 );
or ( n380393 , n59877 , n380392 );
buf ( n380394 , n380393 );
buf ( n380395 , n380361 );
buf ( n380396 , n380356 );
nor ( n380397 , n380395 , n380396 );
buf ( n380398 , n380397 );
buf ( n380399 , n380398 );
buf ( n380400 , n380399 );
buf ( n380401 , n380400 );
buf ( n380402 , n380401 );
buf ( n380403 , n380402 );
buf ( n380404 , n380403 );
buf ( n380405 , n380404 );
buf ( n380406 , n380405 );
buf ( n380407 , n380406 );
buf ( n380408 , n380407 );
nand ( n380409 , n380394 , n380408 );
buf ( n380410 , n380409 );
buf ( n380411 , n380410 );
nand ( n380412 , n380389 , n380411 );
buf ( n380413 , n380412 );
buf ( n380414 , n380413 );
xor ( n380415 , n380352 , n380414 );
buf ( n380416 , n369444 );
not ( n59904 , n380416 );
buf ( n380418 , n368549 );
not ( n380419 , n380418 );
buf ( n380420 , n361751 );
not ( n380421 , n380420 );
or ( n380422 , n380419 , n380421 );
not ( n59910 , n44783 );
not ( n380424 , n368549 );
nand ( n59912 , n59910 , n380424 );
buf ( n380426 , n59912 );
nand ( n59914 , n380422 , n380426 );
buf ( n380428 , n59914 );
buf ( n380429 , n380428 );
not ( n59917 , n380429 );
or ( n59918 , n59904 , n59917 );
buf ( n380432 , n368549 );
buf ( n380433 , n365757 );
and ( n380434 , n380432 , n380433 );
not ( n59922 , n380432 );
buf ( n380436 , n365760 );
and ( n59924 , n59922 , n380436 );
nor ( n380438 , n380434 , n59924 );
buf ( n380439 , n380438 );
buf ( n380440 , n380439 );
buf ( n380441 , n368608 );
nand ( n380442 , n380440 , n380441 );
buf ( n380443 , n380442 );
buf ( n380444 , n380443 );
nand ( n380445 , n59918 , n380444 );
buf ( n380446 , n380445 );
buf ( n380447 , n380446 );
not ( n380448 , n380447 );
buf ( n380449 , n378098 );
not ( n380450 , n380449 );
buf ( n380451 , n42455 );
not ( n380452 , n380451 );
or ( n59940 , n380450 , n380452 );
buf ( n59941 , n359950 );
buf ( n59942 , n379515 );
nand ( n59943 , n59941 , n59942 );
buf ( n59944 , n59943 );
buf ( n380458 , n59944 );
nand ( n59946 , n59940 , n380458 );
buf ( n380460 , n59946 );
buf ( n380461 , n380460 );
not ( n380462 , n380461 );
buf ( n380463 , n359916 );
not ( n59951 , n380463 );
or ( n380465 , n380462 , n59951 );
buf ( n59953 , n368038 );
buf ( n59954 , n377094 );
not ( n59955 , n59954 );
buf ( n380469 , n42455 );
not ( n380470 , n380469 );
or ( n59958 , n59955 , n380470 );
buf ( n380472 , n361762 );
buf ( n380473 , n56687 );
nand ( n59961 , n380472 , n380473 );
buf ( n380475 , n59961 );
buf ( n380476 , n380475 );
nand ( n380477 , n59958 , n380476 );
buf ( n380478 , n380477 );
buf ( n380479 , n380478 );
nand ( n380480 , n59953 , n380479 );
buf ( n380481 , n380480 );
buf ( n380482 , n380481 );
nand ( n59970 , n380465 , n380482 );
buf ( n59971 , n59970 );
buf ( n380485 , n59971 );
not ( n380486 , n380485 );
or ( n380487 , n380448 , n380486 );
or ( n59975 , n59971 , n380446 );
buf ( n380489 , n47466 );
not ( n380490 , n380489 );
buf ( n380491 , n365041 );
not ( n59979 , n380491 );
buf ( n380493 , n32085 );
not ( n380494 , n380493 );
or ( n380495 , n59979 , n380494 );
buf ( n380496 , n32084 );
buf ( n380497 , n369183 );
buf ( n380498 , n380497 );
nand ( n59986 , n380496 , n380498 );
buf ( n380500 , n59986 );
buf ( n380501 , n380500 );
nand ( n380502 , n380495 , n380501 );
buf ( n380503 , n380502 );
buf ( n380504 , n380503 );
not ( n59992 , n380504 );
or ( n380506 , n380490 , n59992 );
not ( n380507 , n365052 );
and ( n59995 , n362534 , n380507 );
not ( n59996 , n362534 );
and ( n380510 , n59996 , n365052 );
nor ( n380511 , n59995 , n380510 );
nand ( n380512 , n380511 , n44915 );
buf ( n380513 , n380512 );
nand ( n380514 , n380506 , n380513 );
buf ( n380515 , n380514 );
buf ( n380516 , n380515 );
buf ( n380517 , n368665 );
not ( n380518 , n380517 );
buf ( n380519 , n378032 );
not ( n60007 , n380519 );
or ( n380521 , n380518 , n60007 );
buf ( n380522 , n365319 );
buf ( n380523 , n368662 );
nand ( n380524 , n380522 , n380523 );
buf ( n380525 , n380524 );
buf ( n380526 , n380525 );
nand ( n60014 , n380521 , n380526 );
buf ( n60015 , n60014 );
buf ( n380529 , n60015 );
not ( n380530 , n380529 );
buf ( n380531 , n44591 );
not ( n380532 , n380531 );
or ( n380533 , n380530 , n380532 );
buf ( n380534 , n378036 );
not ( n60022 , n380534 );
buf ( n380536 , n41835 );
nand ( n380537 , n60022 , n380536 );
buf ( n380538 , n380537 );
buf ( n380539 , n380538 );
nand ( n60027 , n380533 , n380539 );
buf ( n380541 , n60027 );
buf ( n380542 , n380541 );
or ( n60030 , n380516 , n380542 );
xor ( n380544 , n57760 , n378298 );
xor ( n60032 , n380544 , n378315 );
xor ( n380546 , n378381 , n58046 );
xor ( n60034 , n60032 , n380546 );
buf ( n380548 , n60034 );
buf ( n380549 , n378214 );
buf ( n380550 , n57800 );
and ( n60038 , n380549 , n380550 );
buf ( n380552 , n57754 );
buf ( n380553 , n378284 );
and ( n380554 , n380552 , n380553 );
nor ( n60042 , n60038 , n380554 );
buf ( n380556 , n60042 );
buf ( n380557 , n380556 );
buf ( n380558 , n378341 );
or ( n60046 , n380557 , n380558 );
buf ( n380560 , n378417 );
buf ( n380561 , n378424 );
or ( n60049 , n380560 , n380561 );
nand ( n60050 , n60046 , n60049 );
buf ( n380564 , n60050 );
buf ( n380565 , n380564 );
buf ( n380566 , n376743 );
not ( n60054 , n57789 );
buf ( n380568 , n60054 );
not ( n380569 , n380568 );
buf ( n380570 , n380569 );
buf ( n380571 , n380570 );
and ( n60059 , n380566 , n380571 );
buf ( n380573 , n376871 );
buf ( n380574 , n60054 );
and ( n60062 , n380573 , n380574 );
nor ( n60063 , n60059 , n60062 );
buf ( n380577 , n60063 );
buf ( n380578 , n380577 );
buf ( n380579 , n378468 );
not ( n60067 , n380579 );
buf ( n380581 , n60067 );
buf ( n380582 , n380581 );
or ( n60070 , n380578 , n380582 );
buf ( n380584 , n378483 );
nand ( n380585 , n60070 , n380584 );
buf ( n380586 , n380585 );
buf ( n380587 , n380586 );
or ( n380588 , n380565 , n380587 );
buf ( n380589 , n380588 );
and ( n380590 , n55685 , n55729 , n376107 );
not ( n380591 , n380590 );
not ( n380592 , n56317 );
or ( n60080 , n380591 , n380592 );
and ( n60081 , n376728 , n376107 );
nor ( n380595 , n60081 , n376730 );
nand ( n380596 , n60080 , n380595 );
not ( n60084 , n376732 );
nand ( n380598 , n60084 , n376120 );
nor ( n60086 , n380596 , n380598 );
not ( n380600 , n60086 );
nand ( n380601 , n380596 , n380598 );
nand ( n60089 , n380600 , n380601 );
buf ( n60090 , n60089 );
buf ( n380604 , n60090 );
buf ( n380605 , n376990 );
and ( n60093 , n380604 , n380605 );
not ( n60094 , n60089 );
buf ( n380608 , n60094 );
buf ( n380609 , n376997 );
and ( n60097 , n380608 , n380609 );
buf ( n380611 , n377003 );
nor ( n60099 , n60093 , n60097 , n380611 );
buf ( n380613 , n60099 );
xor ( n60101 , n380589 , n380613 );
xor ( n60102 , n378429 , n378487 );
xor ( n380616 , n60102 , n378505 );
buf ( n380617 , n380616 );
and ( n380618 , n60101 , n380617 );
and ( n380619 , n380589 , n380613 );
or ( n60107 , n380618 , n380619 );
xor ( n380621 , n57926 , n378408 );
xor ( n380622 , n380621 , n378509 );
and ( n60110 , n60107 , n380622 );
buf ( n380624 , n60089 );
buf ( n380625 , n376866 );
and ( n380626 , n380624 , n380625 );
buf ( n380627 , n60094 );
buf ( n380628 , n376875 );
and ( n380629 , n380627 , n380628 );
nor ( n380630 , n380626 , n380629 );
buf ( n380631 , n380630 );
buf ( n380632 , n380631 );
buf ( n380633 , n376924 );
or ( n380634 , n380632 , n380633 );
buf ( n380635 , n58030 );
buf ( n380636 , n56517 );
or ( n380637 , n380635 , n380636 );
nand ( n380638 , n380634 , n380637 );
buf ( n380639 , n380638 );
buf ( n380640 , n380639 );
nor ( n380641 , n376730 , n376943 );
not ( n60129 , n55729 );
not ( n60130 , n378199 );
or ( n60131 , n60129 , n60130 );
not ( n380645 , n378205 );
nand ( n380646 , n60131 , n380645 );
not ( n380647 , n380646 );
and ( n60135 , n380641 , n380647 );
not ( n380649 , n380641 );
and ( n60137 , n380649 , n380646 );
or ( n380651 , n60135 , n60137 );
buf ( n380652 , n380651 );
buf ( n380653 , n376990 );
and ( n380654 , n380652 , n380653 );
buf ( n380655 , n380651 );
not ( n60143 , n380655 );
buf ( n380657 , n60143 );
buf ( n380658 , n380657 );
buf ( n380659 , n376997 );
and ( n60147 , n380658 , n380659 );
buf ( n380661 , n377003 );
nor ( n380662 , n380654 , n60147 , n380661 );
buf ( n380663 , n380662 );
buf ( n380664 , n380663 );
xor ( n380665 , n380640 , n380664 );
not ( n380666 , n376723 );
not ( n60154 , n55708 );
nand ( n60155 , n60154 , n57890 );
not ( n380669 , n60155 );
or ( n380670 , n380666 , n380669 );
not ( n380671 , n55728 );
nand ( n380672 , n380671 , n376725 );
nand ( n60160 , n380670 , n380672 );
not ( n380674 , n60154 );
not ( n380675 , n57890 );
or ( n60163 , n380674 , n380675 );
not ( n60164 , n376723 );
nor ( n380678 , n60164 , n380672 );
nand ( n380679 , n60163 , n380678 );
nand ( n380680 , n60160 , n380679 );
buf ( n380681 , n380680 );
buf ( n380682 , n376990 );
and ( n380683 , n380681 , n380682 );
not ( n60171 , n380680 );
buf ( n380685 , n60171 );
buf ( n380686 , n376997 );
and ( n380687 , n380685 , n380686 );
buf ( n380688 , n377003 );
nor ( n380689 , n380683 , n380687 , n380688 );
buf ( n380690 , n380689 );
buf ( n380691 , n380690 );
not ( n380692 , n57978 );
not ( n380693 , n380692 );
and ( n60181 , n57975 , n378437 );
xor ( n60182 , n60181 , n56409 );
buf ( n380696 , n60182 );
not ( n380697 , n380696 );
nand ( n380698 , n380693 , n57976 , n380697 );
not ( n60186 , n57978 );
not ( n380700 , n57976 );
nand ( n380701 , n60186 , n380700 , n380697 );
nand ( n60189 , n57976 , n380696 , n380692 );
nand ( n60190 , n380700 , n380696 , n57978 );
nand ( n380704 , n380698 , n380701 , n60189 , n60190 );
buf ( n380705 , n380696 );
not ( n60193 , n56386 );
nor ( n60194 , n376790 , n60193 );
not ( n60195 , n60194 );
not ( n380709 , n376781 );
nand ( n380710 , n376779 , n56367 );
not ( n60198 , n380710 );
or ( n60199 , n380709 , n60198 );
and ( n60200 , n376792 , n376773 );
nand ( n380714 , n60199 , n60200 );
not ( n60202 , n56357 );
and ( n60203 , n60202 , n376792 );
not ( n60204 , n376769 );
nor ( n380718 , n60203 , n60204 );
nand ( n380719 , n380714 , n380718 );
not ( n60207 , n380719 );
or ( n380721 , n60195 , n60207 );
nand ( n380722 , n56392 , n56395 );
and ( n60210 , n380722 , n56386 );
nor ( n60211 , n60210 , n376810 );
nand ( n380725 , n380721 , n60211 );
nand ( n380726 , n376794 , n376807 );
xnor ( n60214 , n380725 , n380726 );
buf ( n380728 , n60214 );
xor ( n380729 , n380705 , n380728 );
buf ( n380730 , n380729 );
buf ( n380731 , n380730 );
not ( n380732 , n380731 );
buf ( n380733 , n380732 );
nand ( n380734 , n380704 , n380733 );
not ( n380735 , n380734 );
buf ( n380736 , n380735 );
buf ( n380737 , n57983 );
nand ( n60225 , n380736 , n380737 );
buf ( n60226 , n60225 );
buf ( n60227 , n60226 );
buf ( n380741 , n380730 );
buf ( n380742 , n57983 );
nand ( n380743 , n380741 , n380742 );
buf ( n380744 , n380743 );
buf ( n380745 , n380744 );
and ( n380746 , n60227 , n380745 );
buf ( n380747 , n380746 );
buf ( n380748 , n380747 );
xor ( n60236 , n380691 , n380748 );
buf ( n380750 , n380651 );
buf ( n380751 , n376866 );
and ( n60239 , n380750 , n380751 );
buf ( n380753 , n380657 );
buf ( n380754 , n376875 );
and ( n60242 , n380753 , n380754 );
nor ( n60243 , n60239 , n60242 );
buf ( n380757 , n60243 );
buf ( n380758 , n380757 );
buf ( n380759 , n376924 );
or ( n380760 , n380758 , n380759 );
buf ( n380761 , n380631 );
buf ( n380762 , n56517 );
or ( n60250 , n380761 , n380762 );
nand ( n380764 , n380760 , n60250 );
buf ( n380765 , n380764 );
buf ( n380766 , n380765 );
and ( n60254 , n60236 , n380766 );
and ( n380768 , n380691 , n380748 );
or ( n380769 , n60254 , n380768 );
buf ( n380770 , n380769 );
buf ( n380771 , n380770 );
and ( n380772 , n380665 , n380771 );
and ( n380773 , n380640 , n380664 );
or ( n60261 , n380772 , n380773 );
buf ( n380775 , n60261 );
xor ( n60263 , n380589 , n380613 );
xor ( n380777 , n60263 , n380617 );
and ( n380778 , n380775 , n380777 );
buf ( n380779 , n378368 );
buf ( n380780 , n57800 );
and ( n380781 , n380779 , n380780 );
buf ( n380782 , n378372 );
buf ( n380783 , n378284 );
and ( n380784 , n380782 , n380783 );
nor ( n60272 , n380781 , n380784 );
buf ( n380786 , n60272 );
buf ( n380787 , n380786 );
buf ( n380788 , n378341 );
or ( n60276 , n380787 , n380788 );
buf ( n380790 , n380556 );
buf ( n380791 , n378424 );
or ( n60279 , n380790 , n380791 );
nand ( n380793 , n60276 , n60279 );
buf ( n380794 , n380793 );
buf ( n380795 , n380794 );
buf ( n380796 , n376971 );
buf ( n380797 , n380570 );
and ( n380798 , n380796 , n380797 );
buf ( n380799 , n376993 );
buf ( n380800 , n60054 );
and ( n380801 , n380799 , n380800 );
nor ( n380802 , n380798 , n380801 );
buf ( n380803 , n380802 );
buf ( n380804 , n380803 );
buf ( n380805 , n380581 );
or ( n60293 , n380804 , n380805 );
buf ( n380807 , n380577 );
buf ( n380808 , n378453 );
or ( n60296 , n380807 , n380808 );
nand ( n60297 , n60293 , n60296 );
buf ( n380811 , n60297 );
buf ( n380812 , n380811 );
xor ( n60300 , n380795 , n380812 );
buf ( n380814 , n376743 );
buf ( n380815 , n57983 );
not ( n380816 , n380815 );
buf ( n380817 , n380816 );
buf ( n380818 , n380817 );
and ( n60306 , n380814 , n380818 );
buf ( n380820 , n376871 );
buf ( n380821 , n57983 );
and ( n60309 , n380820 , n380821 );
nor ( n60310 , n60306 , n60309 );
buf ( n380824 , n60310 );
buf ( n380825 , n380824 );
buf ( n60313 , n380734 );
buf ( n380827 , n60313 );
or ( n60315 , n380825 , n380827 );
buf ( n380829 , n380744 );
nand ( n60317 , n60315 , n380829 );
buf ( n380831 , n60317 );
buf ( n380832 , n380831 );
and ( n380833 , n60154 , n376723 );
not ( n380834 , n380833 );
and ( n60322 , n57889 , n380834 );
not ( n380836 , n57889 );
and ( n60324 , n380836 , n380833 );
nor ( n380838 , n60322 , n60324 );
buf ( n380839 , n380838 );
buf ( n380840 , n376990 );
and ( n380841 , n380839 , n380840 );
buf ( n380842 , n380838 );
not ( n380843 , n380842 );
buf ( n380844 , n380843 );
buf ( n380845 , n380844 );
buf ( n380846 , n376997 );
and ( n380847 , n380845 , n380846 );
buf ( n380848 , n377003 );
nor ( n60336 , n380841 , n380847 , n380848 );
buf ( n380850 , n60336 );
buf ( n380851 , n380850 );
or ( n60339 , n380832 , n380851 );
buf ( n380853 , n60339 );
buf ( n380854 , n380853 );
and ( n380855 , n60300 , n380854 );
and ( n60343 , n380795 , n380812 );
or ( n60344 , n380855 , n60343 );
buf ( n380858 , n60344 );
buf ( n380859 , n380586 );
not ( n60347 , n380859 );
buf ( n380861 , n380564 );
not ( n380862 , n380861 );
or ( n60350 , n60347 , n380862 );
buf ( n380864 , n380589 );
nand ( n380865 , n60350 , n380864 );
buf ( n380866 , n380865 );
xor ( n60354 , n380858 , n380866 );
xor ( n60355 , n380640 , n380664 );
xor ( n380869 , n60355 , n380771 );
buf ( n380870 , n380869 );
and ( n60358 , n60354 , n380870 );
and ( n60359 , n380858 , n380866 );
or ( n380873 , n60358 , n60359 );
xor ( n60361 , n380589 , n380613 );
xor ( n380875 , n60361 , n380617 );
and ( n60363 , n380873 , n380875 );
and ( n380877 , n380775 , n380873 );
or ( n60365 , n380778 , n60363 , n380877 );
xor ( n60366 , n57926 , n378408 );
xor ( n380880 , n60366 , n378509 );
and ( n380881 , n60365 , n380880 );
and ( n60369 , n60107 , n60365 );
or ( n380883 , n60110 , n380881 , n60369 );
buf ( n380884 , n380883 );
xor ( n60372 , n380548 , n380884 );
not ( n380886 , n375920 );
not ( n380887 , n58062 );
or ( n60375 , n380886 , n380887 );
buf ( n380889 , n57233 );
not ( n380890 , n380889 );
buf ( n380891 , n366659 );
not ( n380892 , n380891 );
or ( n60380 , n380890 , n380892 );
buf ( n380894 , n31194 );
buf ( n380895 , n378135 );
nand ( n380896 , n380894 , n380895 );
buf ( n380897 , n380896 );
buf ( n380898 , n380897 );
nand ( n380899 , n60380 , n380898 );
buf ( n380900 , n380899 );
buf ( n380901 , n366707 );
nand ( n380902 , n380900 , n380901 );
nand ( n380903 , n60375 , n380902 );
buf ( n380904 , n380903 );
and ( n380905 , n60372 , n380904 );
and ( n380906 , n380548 , n380884 );
or ( n60394 , n380905 , n380906 );
buf ( n380908 , n60394 );
buf ( n380909 , n380908 );
buf ( n380910 , n56794 );
not ( n60398 , n380910 );
buf ( n380912 , n379205 );
not ( n60400 , n380912 );
or ( n380914 , n60398 , n60400 );
buf ( n380915 , n377190 );
not ( n60403 , n380915 );
buf ( n380917 , n377297 );
not ( n60405 , n380917 );
or ( n380919 , n60403 , n60405 );
buf ( n380920 , n351291 );
buf ( n380921 , n22619 );
not ( n380922 , n380921 );
buf ( n380923 , n380922 );
buf ( n380924 , n380923 );
nand ( n60412 , n380920 , n380924 );
buf ( n380926 , n60412 );
buf ( n380927 , n380926 );
nand ( n380928 , n380919 , n380927 );
buf ( n380929 , n380928 );
buf ( n380930 , n380929 );
buf ( n380931 , n45553 );
nand ( n60419 , n380930 , n380931 );
buf ( n380933 , n60419 );
buf ( n380934 , n380933 );
nand ( n380935 , n380914 , n380934 );
buf ( n380936 , n380935 );
buf ( n380937 , n380936 );
xor ( n380938 , n380909 , n380937 );
buf ( n380939 , n364901 );
not ( n380940 , n380939 );
buf ( n380941 , n42233 );
not ( n60429 , n380941 );
or ( n380943 , n380940 , n60429 );
buf ( n380944 , n46693 );
buf ( n380945 , n44737 );
nand ( n380946 , n380944 , n380945 );
buf ( n380947 , n380946 );
buf ( n380948 , n380947 );
nand ( n60436 , n380943 , n380948 );
buf ( n60437 , n60436 );
buf ( n380951 , n60437 );
not ( n60439 , n380951 );
buf ( n380953 , n363428 );
not ( n60441 , n380953 );
or ( n380955 , n60439 , n60441 );
buf ( n380956 , n378164 );
buf ( n380957 , n58231 );
nand ( n60445 , n380956 , n380957 );
buf ( n380959 , n60445 );
buf ( n380960 , n380959 );
nand ( n380961 , n380955 , n380960 );
buf ( n380962 , n380961 );
buf ( n60450 , n380962 );
not ( n60451 , n60450 );
buf ( n60452 , n60451 );
buf ( n380966 , n60452 );
xor ( n380967 , n380938 , n380966 );
buf ( n380968 , n380967 );
buf ( n380969 , n380968 );
not ( n380970 , n380969 );
buf ( n380971 , n380970 );
buf ( n380972 , n380971 );
nand ( n60460 , n60030 , n380972 );
buf ( n380974 , n60460 );
buf ( n380975 , n380541 );
buf ( n380976 , n380515 );
nand ( n380977 , n380975 , n380976 );
buf ( n380978 , n380977 );
nand ( n380979 , n380974 , n380978 );
nand ( n60467 , n59975 , n380979 );
buf ( n380981 , n60467 );
nand ( n60469 , n380487 , n380981 );
buf ( n380983 , n60469 );
buf ( n380984 , n380983 );
and ( n380985 , n380415 , n380984 );
and ( n380986 , n380352 , n380414 );
or ( n380987 , n380985 , n380986 );
buf ( n380988 , n380987 );
buf ( n380989 , n380988 );
nand ( n380990 , n59814 , n380989 );
buf ( n380991 , n380990 );
buf ( n380992 , n380991 );
nand ( n380993 , n380319 , n380992 );
buf ( n380994 , n380993 );
not ( n60482 , n380994 );
xor ( n60483 , n379718 , n59335 );
xor ( n60484 , n60483 , n379571 );
not ( n380998 , n60484 );
or ( n60486 , n60482 , n380998 );
not ( n60487 , n60484 );
not ( n60488 , n60487 );
not ( n60489 , n380994 );
not ( n60490 , n60489 );
or ( n381004 , n60488 , n60490 );
buf ( n60492 , n377809 );
not ( n60493 , n60492 );
and ( n381007 , n57371 , n58186 );
not ( n60495 , n57371 );
not ( n60496 , n58186 );
and ( n60497 , n60495 , n60496 );
nor ( n60498 , n381007 , n60497 );
and ( n60499 , n60493 , n60498 );
not ( n60500 , n60493 );
not ( n60501 , n60498 );
and ( n60502 , n60500 , n60501 );
nor ( n60503 , n60499 , n60502 );
nand ( n60504 , n381004 , n60503 );
nand ( n60505 , n60486 , n60504 );
not ( n60506 , n60505 );
nand ( n60507 , n379440 , n380243 , n60506 );
not ( n60508 , n380243 );
nand ( n60509 , n60508 , n60505 );
nor ( n60510 , n60509 , n379439 );
not ( n60511 , n60510 );
nand ( n60512 , n60505 , n380243 );
not ( n60513 , n60512 );
nand ( n60514 , n60513 , n379439 );
nor ( n60515 , n60505 , n380243 );
nand ( n60516 , n60515 , n379439 );
nand ( n381030 , n60507 , n60511 , n60514 , n60516 );
xor ( n60517 , n379535 , n379457 );
buf ( n381032 , n60517 );
buf ( n381033 , n379564 );
buf ( n381034 , n381033 );
buf ( n381035 , n381034 );
buf ( n381036 , n381035 );
xnor ( n60520 , n381032 , n381036 );
buf ( n381038 , n60520 );
buf ( n381039 , n381038 );
not ( n60523 , n381039 );
buf ( n381041 , n377983 );
buf ( n381042 , n378002 );
xor ( n60526 , n381041 , n381042 );
buf ( n381044 , n58184 );
xor ( n60528 , n60526 , n381044 );
buf ( n381046 , n60528 );
buf ( n381047 , n381046 );
not ( n381048 , n381047 );
buf ( n381049 , n381048 );
buf ( n381050 , n381049 );
not ( n381051 , n381050 );
or ( n381052 , n60523 , n381051 );
not ( n60536 , n379890 );
and ( n381054 , n379847 , n365681 );
not ( n381055 , n379847 );
and ( n60539 , n381055 , n359781 );
nor ( n381057 , n381054 , n60539 );
not ( n381058 , n381057 );
or ( n381059 , n60536 , n381058 );
not ( n60543 , n379841 );
not ( n381061 , n46902 );
or ( n60545 , n60543 , n381061 );
nand ( n381063 , n40199 , n379847 );
nand ( n60547 , n60545 , n381063 );
nand ( n60548 , n60547 , n379916 );
nand ( n381066 , n381059 , n60548 );
buf ( n60550 , n368608 );
not ( n60551 , n60550 );
buf ( n381069 , n368549 );
not ( n381070 , n381069 );
buf ( n381071 , n43377 );
not ( n381072 , n381071 );
or ( n381073 , n381070 , n381072 );
buf ( n381074 , n361716 );
buf ( n381075 , n380424 );
nand ( n381076 , n381074 , n381075 );
buf ( n381077 , n381076 );
buf ( n381078 , n381077 );
nand ( n381079 , n381073 , n381078 );
buf ( n381080 , n381079 );
buf ( n381081 , n381080 );
not ( n381082 , n381081 );
or ( n381083 , n60551 , n381082 );
buf ( n381084 , n380439 );
buf ( n381085 , n369444 );
nand ( n381086 , n381084 , n381085 );
buf ( n381087 , n381086 );
buf ( n381088 , n381087 );
nand ( n381089 , n381083 , n381088 );
buf ( n381090 , n381089 );
buf ( n381091 , n381090 );
not ( n381092 , n381091 );
buf ( n381093 , n359993 );
buf ( n381094 , n378098 );
nand ( n381095 , n381093 , n381094 );
buf ( n381096 , n381095 );
buf ( n381097 , n381096 );
nand ( n60559 , n381092 , n381097 );
buf ( n381099 , n60559 );
buf ( n381100 , n381099 );
buf ( n381101 , n378856 );
not ( n60563 , n381101 );
buf ( n381103 , n35547 );
not ( n381104 , n381103 );
or ( n60566 , n60563 , n381104 );
buf ( n381106 , n51966 );
buf ( n381107 , n378847 );
nand ( n60569 , n381106 , n381107 );
buf ( n381109 , n60569 );
buf ( n381110 , n381109 );
nand ( n381111 , n60566 , n381110 );
buf ( n381112 , n381111 );
buf ( n381113 , n381112 );
not ( n381114 , n381113 );
buf ( n381115 , n367273 );
not ( n381116 , n381115 );
or ( n60578 , n381114 , n381116 );
buf ( n60579 , n58984 );
buf ( n60580 , n355579 );
and ( n60581 , n60579 , n60580 );
not ( n60582 , n60579 );
buf ( n381122 , n365353 );
and ( n381123 , n60582 , n381122 );
nor ( n60585 , n60581 , n381123 );
buf ( n381125 , n60585 );
buf ( n381126 , n381125 );
not ( n381127 , n381126 );
buf ( n381128 , n46582 );
nand ( n60590 , n381127 , n381128 );
buf ( n381130 , n60590 );
buf ( n381131 , n381130 );
nand ( n381132 , n60578 , n381131 );
buf ( n381133 , n381132 );
buf ( n381134 , n381133 );
and ( n381135 , n381100 , n381134 );
buf ( n381136 , n381096 );
not ( n381137 , n381136 );
buf ( n381138 , n381137 );
buf ( n381139 , n381138 );
buf ( n381140 , n381090 );
and ( n60602 , n381139 , n381140 );
buf ( n381142 , n60602 );
buf ( n381143 , n381142 );
nor ( n381144 , n381135 , n381143 );
buf ( n381145 , n381144 );
buf ( n60607 , n381145 );
not ( n60608 , n60607 );
buf ( n60609 , n60608 );
buf ( n381149 , n60609 );
not ( n60611 , n381149 );
not ( n381151 , n58170 );
not ( n381152 , n370050 );
and ( n60614 , n381151 , n381152 );
and ( n381154 , n378617 , n378619 );
nor ( n381155 , n60614 , n381154 );
nand ( n60617 , n378603 , n58111 );
nor ( n381157 , n381155 , n60617 );
not ( n381158 , n381157 );
not ( n381159 , n58138 );
nand ( n381160 , n381159 , n381155 );
nand ( n60621 , n58172 , n58112 , n58136 );
nand ( n381162 , n381155 , n58175 );
nand ( n381163 , n381158 , n381160 , n60621 , n381162 );
buf ( n381164 , n381163 );
not ( n381165 , n381164 );
buf ( n381166 , n381165 );
buf ( n381167 , n381166 );
not ( n381168 , n381167 );
or ( n60627 , n60611 , n381168 );
buf ( n381170 , n381145 );
not ( n381171 , n381170 );
buf ( n381172 , n381163 );
not ( n381173 , n381172 );
or ( n60632 , n381171 , n381173 );
buf ( n381175 , n369374 );
not ( n381176 , n381175 );
buf ( n381177 , n44717 );
not ( n60636 , n381177 );
or ( n60637 , n381176 , n60636 );
buf ( n381180 , n366096 );
buf ( n381181 , n49178 );
nand ( n381182 , n381180 , n381181 );
buf ( n381183 , n381182 );
buf ( n381184 , n381183 );
nand ( n60643 , n60637 , n381184 );
buf ( n381186 , n60643 );
buf ( n381187 , n381186 );
not ( n60646 , n381187 );
buf ( n381189 , n364849 );
not ( n381190 , n381189 );
or ( n60649 , n60646 , n381190 );
buf ( n381192 , n367590 );
buf ( n381193 , n368994 );
not ( n60652 , n381193 );
buf ( n60653 , n44717 );
not ( n60654 , n60653 );
or ( n60655 , n60652 , n60654 );
buf ( n381198 , n45414 );
buf ( n381199 , n57053 );
nand ( n60658 , n381198 , n381199 );
buf ( n381201 , n60658 );
buf ( n381202 , n381201 );
nand ( n381203 , n60655 , n381202 );
buf ( n381204 , n381203 );
buf ( n381205 , n381204 );
nand ( n60664 , n381192 , n381205 );
buf ( n381207 , n60664 );
buf ( n381208 , n381207 );
nand ( n381209 , n60649 , n381208 );
buf ( n381210 , n381209 );
buf ( n381211 , n381210 );
xor ( n60670 , n57926 , n378408 );
xor ( n60671 , n60670 , n378509 );
xor ( n60672 , n60107 , n60365 );
xor ( n60673 , n60671 , n60672 );
buf ( n381216 , n60673 );
not ( n60675 , n380901 );
buf ( n381218 , n351195 );
not ( n381219 , n381218 );
buf ( n381220 , n381219 );
buf ( n381221 , n381220 );
buf ( n381222 , n378138 );
and ( n381223 , n381221 , n381222 );
not ( n60682 , n381221 );
buf ( n381225 , n378135 );
and ( n60684 , n60682 , n381225 );
nor ( n60685 , n381223 , n60684 );
buf ( n381228 , n60685 );
not ( n381229 , n381228 );
or ( n60688 , n60675 , n381229 );
buf ( n381231 , n366649 );
not ( n381232 , n381231 );
buf ( n381233 , n380900 );
nand ( n60692 , n381232 , n381233 );
buf ( n381235 , n60692 );
nand ( n60694 , n60688 , n381235 );
buf ( n381237 , n60694 );
xor ( n381238 , n381216 , n381237 );
buf ( n381239 , n364901 );
not ( n60698 , n381239 );
buf ( n381241 , n58471 );
not ( n381242 , n381241 );
or ( n381243 , n60698 , n381242 );
buf ( n381244 , n342654 );
buf ( n381245 , n364900 );
nand ( n60704 , n381244 , n381245 );
buf ( n381247 , n60704 );
buf ( n381248 , n381247 );
nand ( n60707 , n381243 , n381248 );
buf ( n381250 , n60707 );
buf ( n381251 , n381250 );
not ( n60710 , n381251 );
buf ( n381253 , n366396 );
not ( n381254 , n381253 );
or ( n60713 , n60710 , n381254 );
buf ( n381256 , n366393 );
not ( n60715 , n381256 );
buf ( n381258 , n351160 );
not ( n60717 , n381258 );
buf ( n381260 , n375944 );
not ( n381261 , n381260 );
or ( n60720 , n60717 , n381261 );
buf ( n381263 , n378956 );
buf ( n381264 , n351160 );
not ( n60723 , n381264 );
buf ( n381266 , n60723 );
buf ( n381267 , n381266 );
nand ( n60726 , n381263 , n381267 );
buf ( n381269 , n60726 );
buf ( n381270 , n381269 );
nand ( n60729 , n60720 , n381270 );
buf ( n381272 , n60729 );
buf ( n381273 , n381272 );
nand ( n60732 , n60715 , n381273 );
buf ( n381275 , n60732 );
buf ( n381276 , n381275 );
nand ( n381277 , n60713 , n381276 );
buf ( n381278 , n381277 );
buf ( n381279 , n381278 );
and ( n381280 , n381238 , n381279 );
and ( n60739 , n381216 , n381237 );
or ( n381282 , n381280 , n60739 );
buf ( n381283 , n381282 );
buf ( n381284 , n45802 );
not ( n60743 , n381284 );
not ( n381286 , n46693 );
buf ( n381287 , n381286 );
not ( n60746 , n381287 );
or ( n381289 , n60743 , n60746 );
buf ( n381290 , n55539 );
buf ( n381291 , n45802 );
not ( n60750 , n381291 );
buf ( n60751 , n60750 );
buf ( n60752 , n60751 );
nand ( n60753 , n381290 , n60752 );
buf ( n381296 , n60753 );
buf ( n381297 , n381296 );
nand ( n381298 , n381289 , n381297 );
buf ( n381299 , n381298 );
buf ( n381300 , n381299 );
not ( n60759 , n381300 );
buf ( n381302 , n363429 );
not ( n60761 , n381302 );
or ( n381304 , n60759 , n60761 );
buf ( n381305 , n363416 );
not ( n60764 , n381305 );
buf ( n381307 , n60437 );
nand ( n60766 , n60764 , n381307 );
buf ( n381309 , n60766 );
buf ( n381310 , n381309 );
nand ( n381311 , n381304 , n381310 );
buf ( n381312 , n381311 );
xor ( n381313 , n381283 , n381312 );
buf ( n381314 , n365393 );
not ( n60773 , n381314 );
buf ( n381316 , n368765 );
not ( n381317 , n381316 );
or ( n60776 , n60773 , n381317 );
buf ( n381319 , n362417 );
buf ( n381320 , n365408 );
nand ( n381321 , n381319 , n381320 );
buf ( n381322 , n381321 );
buf ( n60781 , n381322 );
nand ( n60782 , n60776 , n60781 );
buf ( n60783 , n60782 );
buf ( n381326 , n60783 );
not ( n60785 , n381326 );
buf ( n381328 , n362405 );
not ( n60787 , n381328 );
or ( n60788 , n60785 , n60787 );
not ( n381331 , n365428 );
not ( n60790 , n368765 );
or ( n381333 , n381331 , n60790 );
buf ( n381334 , n342335 );
not ( n381335 , n381334 );
buf ( n381336 , n381335 );
buf ( n381337 , n381336 );
buf ( n381338 , n365422 );
nand ( n60797 , n381337 , n381338 );
buf ( n381340 , n60797 );
nand ( n60799 , n381333 , n381340 );
nand ( n381342 , n60799 , n48558 );
buf ( n381343 , n381342 );
nand ( n381344 , n60788 , n381343 );
buf ( n381345 , n381344 );
and ( n60804 , n381313 , n381345 );
and ( n381347 , n381283 , n381312 );
or ( n381348 , n60804 , n381347 );
buf ( n381349 , n381348 );
xor ( n381350 , n381211 , n381349 );
and ( n381351 , n377353 , n365626 );
not ( n60810 , n377353 );
and ( n381353 , n60810 , n41892 );
or ( n381354 , n381351 , n381353 );
buf ( n381355 , n381354 );
not ( n60814 , n381355 );
buf ( n381357 , n364797 );
not ( n381358 , n381357 );
or ( n60817 , n60814 , n381358 );
buf ( n381360 , n41918 );
buf ( n381361 , n56970 );
not ( n60820 , n381361 );
buf ( n381363 , n364832 );
not ( n381364 , n381363 );
or ( n60823 , n60820 , n381364 );
buf ( n381366 , n41892 );
buf ( n381367 , n377389 );
nand ( n381368 , n381366 , n381367 );
buf ( n381369 , n381368 );
buf ( n381370 , n381369 );
nand ( n60829 , n60823 , n381370 );
buf ( n381372 , n60829 );
buf ( n381373 , n381372 );
nand ( n381374 , n381360 , n381373 );
buf ( n381375 , n381374 );
buf ( n381376 , n381375 );
nand ( n381377 , n60817 , n381376 );
buf ( n381378 , n381377 );
buf ( n381379 , n381378 );
and ( n60838 , n381350 , n381379 );
and ( n60839 , n381211 , n381349 );
or ( n60840 , n60838 , n60839 );
buf ( n381383 , n60840 );
buf ( n381384 , n381383 );
nand ( n381385 , n60632 , n381384 );
buf ( n381386 , n381385 );
buf ( n381387 , n381386 );
nand ( n381388 , n60627 , n381387 );
buf ( n381389 , n381388 );
xor ( n381390 , n381066 , n381389 );
not ( n381391 , n368611 );
not ( n381392 , n380428 );
or ( n381393 , n381391 , n381392 );
not ( n381394 , n379583 );
not ( n381395 , n379581 );
or ( n381396 , n381394 , n381395 );
nand ( n381397 , n381396 , n369444 );
nand ( n381398 , n381393 , n381397 );
not ( n381399 , n380936 );
buf ( n381400 , n381399 );
not ( n381401 , n381400 );
buf ( n381402 , n60452 );
not ( n381403 , n381402 );
or ( n60843 , n381401 , n381403 );
buf ( n381405 , n380908 );
nand ( n60845 , n60843 , n381405 );
buf ( n381407 , n60845 );
buf ( n60847 , n381407 );
buf ( n381409 , n380962 );
buf ( n381410 , n380936 );
nand ( n60850 , n381409 , n381410 );
buf ( n381412 , n60850 );
buf ( n60852 , n381412 );
nand ( n60853 , n60847 , n60852 );
buf ( n60854 , n60853 );
buf ( n381416 , n60854 );
buf ( n381417 , n58596 );
buf ( n381418 , n58615 );
or ( n381419 , n381417 , n381418 );
buf ( n381420 , n381204 );
buf ( n381421 , n361580 );
not ( n381422 , n381421 );
buf ( n381423 , n381422 );
buf ( n381424 , n381423 );
not ( n60864 , n381424 );
buf ( n381426 , n60864 );
buf ( n381427 , n381426 );
not ( n60867 , n366103 );
buf ( n381429 , n60867 );
nand ( n60869 , n381420 , n381427 , n381429 );
buf ( n381431 , n60869 );
buf ( n381432 , n381431 );
nand ( n60872 , n381419 , n381432 );
buf ( n381434 , n60872 );
buf ( n60874 , n381434 );
xor ( n60875 , n381416 , n60874 );
buf ( n381437 , n381372 );
not ( n381438 , n381437 );
buf ( n381439 , n45438 );
not ( n381440 , n381439 );
or ( n381441 , n381438 , n381440 );
buf ( n381442 , n365622 );
buf ( n381443 , n59145 );
nand ( n381444 , n381442 , n381443 );
buf ( n381445 , n381444 );
buf ( n381446 , n381445 );
nand ( n381447 , n381441 , n381446 );
buf ( n381448 , n381447 );
buf ( n381449 , n381448 );
and ( n381450 , n60875 , n381449 );
and ( n381451 , n381416 , n60874 );
or ( n60891 , n381450 , n381451 );
buf ( n381453 , n60891 );
xor ( n60893 , n381398 , n381453 );
not ( n60894 , n369959 );
buf ( n381456 , n377071 );
buf ( n381457 , n366243 );
and ( n60897 , n381456 , n381457 );
not ( n381459 , n381456 );
buf ( n381460 , n364919 );
and ( n60900 , n381459 , n381460 );
nor ( n60901 , n60897 , n60900 );
buf ( n381463 , n60901 );
not ( n381464 , n381463 );
and ( n60904 , n60894 , n381464 );
not ( n60905 , n380478 );
nor ( n60906 , n60905 , n363291 );
nor ( n381468 , n60904 , n60906 );
xnor ( n381469 , n60893 , n381468 );
and ( n60909 , n381390 , n381469 );
and ( n381471 , n381066 , n381389 );
or ( n60911 , n60909 , n381471 );
buf ( n381473 , n60911 );
nand ( n381474 , n381052 , n381473 );
buf ( n381475 , n381474 );
buf ( n381476 , n381475 );
buf ( n381477 , n381046 );
buf ( n381478 , n381038 );
not ( n381479 , n381478 );
buf ( n381480 , n381479 );
buf ( n381481 , n381480 );
nand ( n60921 , n381477 , n381481 );
buf ( n381483 , n60921 );
buf ( n381484 , n381483 );
nand ( n381485 , n381476 , n381484 );
buf ( n381486 , n381485 );
buf ( n381487 , n381486 );
not ( n381488 , n380404 );
not ( n60928 , n59873 );
or ( n381490 , n381488 , n60928 );
buf ( n381491 , n380368 );
not ( n381492 , n381491 );
buf ( n381493 , n40091 );
not ( n60933 , n381493 );
or ( n381495 , n381492 , n60933 );
buf ( n381496 , n40090 );
buf ( n381497 , n59867 );
nand ( n381498 , n381496 , n381497 );
buf ( n381499 , n381498 );
buf ( n381500 , n381499 );
nand ( n60940 , n381495 , n381500 );
buf ( n381502 , n60940 );
nand ( n60942 , n381502 , n380356 );
nand ( n60943 , n381490 , n60942 );
buf ( n381505 , n60943 );
not ( n60945 , n381505 );
buf ( n381507 , n379890 );
not ( n381508 , n381507 );
buf ( n60948 , n379841 );
not ( n60949 , n60948 );
buf ( n60950 , n44925 );
not ( n60951 , n60950 );
or ( n60952 , n60949 , n60951 );
buf ( n60953 , n359756 );
buf ( n60954 , n379847 );
nand ( n60955 , n60953 , n60954 );
buf ( n60956 , n60955 );
buf ( n60957 , n60956 );
nand ( n60958 , n60952 , n60957 );
buf ( n60959 , n60958 );
buf ( n381521 , n60959 );
not ( n60961 , n381521 );
or ( n381523 , n381508 , n60961 );
not ( n60963 , n379841 );
not ( n60964 , n359781 );
or ( n381526 , n60963 , n60964 );
and ( n381527 , n379847 , n365681 );
nor ( n60967 , n381527 , n59424 );
nand ( n381529 , n381526 , n60967 );
buf ( n60969 , n381529 );
nand ( n60970 , n381523 , n60969 );
buf ( n60971 , n60970 );
buf ( n381533 , n60971 );
not ( n60973 , n381533 );
or ( n381535 , n60945 , n60973 );
buf ( n381536 , n60971 );
buf ( n381537 , n60943 );
or ( n60977 , n381536 , n381537 );
buf ( n381539 , n56794 );
not ( n381540 , n381539 );
buf ( n381541 , n377185 );
not ( n60981 , n381541 );
or ( n381543 , n381540 , n60981 );
nand ( n381544 , n58658 , n45553 );
buf ( n381545 , n381544 );
nand ( n381546 , n381543 , n381545 );
buf ( n381547 , n381546 );
buf ( n381548 , n381547 );
buf ( n381549 , n359896 );
not ( n60989 , n381549 );
buf ( n60990 , n359634 );
buf ( n381552 , n60990 );
nand ( n60992 , n60989 , n381552 );
buf ( n381554 , n60992 );
buf ( n381555 , n381554 );
buf ( n381556 , n378098 );
and ( n381557 , n381555 , n381556 );
or ( n60997 , n359904 , n359634 );
nand ( n60998 , n60997 , n366534 );
buf ( n381560 , n60998 );
nor ( n381561 , n381557 , n381560 );
buf ( n381562 , n381561 );
buf ( n381563 , n381562 );
xor ( n381564 , n381548 , n381563 );
buf ( n381565 , n378114 );
not ( n381566 , n381565 );
buf ( n381567 , n44591 );
not ( n61007 , n381567 );
or ( n381569 , n381566 , n61007 );
buf ( n381570 , n379979 );
buf ( n381571 , n365311 );
nand ( n381572 , n381570 , n381571 );
buf ( n381573 , n381572 );
buf ( n381574 , n381573 );
nand ( n61014 , n381569 , n381574 );
buf ( n381576 , n61014 );
buf ( n381577 , n381576 );
xor ( n381578 , n381564 , n381577 );
buf ( n381579 , n381578 );
buf ( n381580 , n381579 );
buf ( n381581 , n366229 );
not ( n61021 , n381581 );
buf ( n381583 , n381463 );
not ( n61023 , n381583 );
and ( n61024 , n61021 , n61023 );
buf ( n381586 , n365801 );
buf ( n381587 , n359944 );
not ( n61027 , n381587 );
buf ( n381589 , n378847 );
not ( n381590 , n381589 );
and ( n61030 , n61027 , n381590 );
buf ( n381592 , n366243 );
buf ( n381593 , n378847 );
and ( n381594 , n381592 , n381593 );
nor ( n381595 , n61030 , n381594 );
buf ( n381596 , n381595 );
buf ( n381597 , n381596 );
nor ( n61037 , n381586 , n381597 );
buf ( n381599 , n61037 );
buf ( n381600 , n381599 );
nor ( n61040 , n61024 , n381600 );
buf ( n381602 , n61040 );
buf ( n381603 , n381602 );
not ( n61043 , n381603 );
buf ( n381605 , n61043 );
buf ( n381606 , n381605 );
xor ( n381607 , n381580 , n381606 );
not ( n61047 , n378576 );
buf ( n61048 , n57685 );
not ( n381610 , n61048 );
not ( n381611 , n381610 );
or ( n61051 , n61047 , n381611 );
nor ( n381613 , n378576 , n381610 );
not ( n381614 , n378187 );
or ( n61054 , n381613 , n381614 );
nand ( n381616 , n61051 , n61054 );
buf ( n61056 , n381616 );
not ( n381618 , n378587 );
not ( n61058 , n45018 );
or ( n381620 , n381618 , n61058 );
not ( n381621 , n59056 );
nand ( n61061 , n381621 , n365152 );
nand ( n381623 , n381620 , n61061 );
buf ( n61063 , n381623 );
xor ( n61064 , n61056 , n61063 );
buf ( n381626 , n58167 );
not ( n61066 , n381626 );
buf ( n381628 , n365279 );
not ( n61068 , n381628 );
or ( n381630 , n61066 , n61068 );
buf ( n381631 , n40923 );
buf ( n381632 , n379739 );
nand ( n61072 , n381631 , n381632 );
buf ( n381634 , n61072 );
buf ( n381635 , n381634 );
nand ( n381636 , n381630 , n381635 );
buf ( n381637 , n381636 );
buf ( n381638 , n381637 );
and ( n381639 , n61064 , n381638 );
and ( n61079 , n61056 , n61063 );
or ( n381641 , n381639 , n61079 );
buf ( n381642 , n381641 );
buf ( n381643 , n381642 );
xor ( n381644 , n381607 , n381643 );
buf ( n381645 , n381644 );
buf ( n381646 , n381645 );
nand ( n61086 , n60977 , n381646 );
buf ( n381648 , n61086 );
buf ( n381649 , n381648 );
nand ( n61089 , n381535 , n381649 );
buf ( n381651 , n61089 );
xor ( n381652 , n379247 , n379306 );
xor ( n61092 , n381652 , n58930 );
buf ( n381654 , n61092 );
xor ( n381655 , n381651 , n381654 );
xor ( n381656 , n379069 , n379075 );
xor ( n61096 , n381656 , n379242 );
buf ( n381658 , n61096 );
buf ( n381659 , n381658 );
not ( n61099 , n381659 );
buf ( n61100 , n61099 );
buf ( n381662 , n61100 );
not ( n61102 , n381662 );
and ( n61103 , n379371 , n365206 );
not ( n381665 , n379371 );
and ( n61105 , n381665 , n371416 );
or ( n381667 , n61103 , n61105 );
buf ( n381668 , n381667 );
buf ( n381669 , n58871 );
and ( n381670 , n381668 , n381669 );
buf ( n381671 , n58897 );
not ( n381672 , n381671 );
buf ( n381673 , n58923 );
not ( n61113 , n381673 );
buf ( n381675 , n61113 );
buf ( n381676 , n381675 );
nor ( n61116 , n381672 , n381676 );
buf ( n381678 , n61116 );
buf ( n381679 , n381678 );
nor ( n61119 , n381670 , n381679 );
buf ( n381681 , n61119 );
buf ( n381682 , n381681 );
not ( n61122 , n381682 );
or ( n381684 , n61102 , n61122 );
not ( n381685 , n381398 );
nand ( n61125 , n381685 , n381468 );
not ( n381687 , n61125 );
not ( n381688 , n381453 );
or ( n61128 , n381687 , n381688 );
not ( n381690 , n381468 );
nand ( n61130 , n381690 , n381398 );
nand ( n61131 , n61128 , n61130 );
buf ( n381693 , n61131 );
nand ( n381694 , n381684 , n381693 );
buf ( n381695 , n381694 );
buf ( n381696 , n381695 );
buf ( n381697 , n381681 );
not ( n61137 , n381697 );
buf ( n381699 , n381658 );
nand ( n381700 , n61137 , n381699 );
buf ( n381701 , n381700 );
buf ( n381702 , n381701 );
nand ( n61142 , n381696 , n381702 );
buf ( n381704 , n61142 );
xor ( n381705 , n381655 , n381704 );
buf ( n61145 , n381705 );
xor ( n61146 , n381487 , n61145 );
buf ( n381708 , n61131 );
buf ( n381709 , n381658 );
xor ( n61149 , n381708 , n381709 );
buf ( n381711 , n381681 );
xor ( n61151 , n61149 , n381711 );
buf ( n381713 , n61151 );
buf ( n381714 , n381713 );
not ( n381715 , n381714 );
buf ( n381716 , n381715 );
buf ( n381717 , n381716 );
not ( n381718 , n381717 );
buf ( n381719 , n378089 );
buf ( n381720 , n378121 );
and ( n61160 , n381719 , n381720 );
not ( n61161 , n381719 );
buf ( n61162 , n378124 );
and ( n381724 , n61161 , n61162 );
nor ( n61164 , n61160 , n381724 );
buf ( n61165 , n61164 );
buf ( n381727 , n61165 );
buf ( n381728 , n378643 );
and ( n381729 , n381727 , n381728 );
not ( n381730 , n381727 );
buf ( n381731 , n378643 );
not ( n61171 , n381731 );
buf ( n61172 , n61171 );
buf ( n381734 , n61172 );
and ( n61174 , n381730 , n381734 );
nor ( n381736 , n381729 , n61174 );
buf ( n381737 , n381736 );
buf ( n381738 , n381737 );
not ( n381739 , n381738 );
buf ( n381740 , n379371 );
not ( n61180 , n381740 );
buf ( n381742 , n44925 );
not ( n381743 , n381742 );
or ( n61183 , n61180 , n381743 );
buf ( n381745 , n359756 );
buf ( n381746 , n379380 );
nand ( n61186 , n381745 , n381746 );
buf ( n61187 , n61186 );
buf ( n61188 , n61187 );
nand ( n61189 , n61183 , n61188 );
buf ( n61190 , n61189 );
buf ( n381752 , n61190 );
not ( n61192 , n381752 );
buf ( n381754 , n61192 );
buf ( n381755 , n381754 );
not ( n381756 , n381755 );
buf ( n381757 , n379359 );
not ( n61197 , n381757 );
and ( n381759 , n381756 , n61197 );
buf ( n381760 , n381667 );
buf ( n381761 , n58923 );
and ( n381762 , n381760 , n381761 );
nor ( n61199 , n381759 , n381762 );
buf ( n381764 , n61199 );
buf ( n381765 , n381764 );
nand ( n61202 , n381739 , n381765 );
buf ( n381767 , n61202 );
buf ( n381768 , n381767 );
xor ( n61205 , n381416 , n60874 );
xor ( n61206 , n61205 , n381449 );
buf ( n381771 , n61206 );
buf ( n381772 , n381771 );
buf ( n381773 , n49609 );
not ( n61210 , n381773 );
buf ( n381775 , n380344 );
not ( n61212 , n381775 );
or ( n61213 , n61210 , n61212 );
buf ( n381778 , n369769 );
not ( n381779 , n381778 );
buf ( n381780 , n369349 );
not ( n381781 , n381780 );
or ( n61218 , n381779 , n381781 );
buf ( n381783 , n46031 );
buf ( n381784 , n369766 );
nand ( n61221 , n381783 , n381784 );
buf ( n381786 , n61221 );
buf ( n381787 , n381786 );
nand ( n381788 , n61218 , n381787 );
buf ( n381789 , n381788 );
buf ( n381790 , n381789 );
buf ( n381791 , n369804 );
nand ( n381792 , n381790 , n381791 );
buf ( n381793 , n381792 );
buf ( n381794 , n381793 );
nand ( n61231 , n61213 , n381794 );
buf ( n61232 , n61231 );
buf ( n381797 , n61232 );
xor ( n61234 , n381772 , n381797 );
xor ( n61235 , n380548 , n380884 );
xor ( n381800 , n61235 , n380904 );
buf ( n381801 , n381800 );
not ( n381802 , n381272 );
not ( n381803 , n366399 );
or ( n381804 , n381802 , n381803 );
buf ( n381805 , n378549 );
buf ( n381806 , n366425 );
nand ( n381807 , n381805 , n381806 );
buf ( n381808 , n381807 );
nand ( n381809 , n381804 , n381808 );
not ( n61246 , n381809 );
not ( n61247 , n56794 );
not ( n61248 , n380929 );
or ( n61249 , n61247 , n61248 );
buf ( n381814 , n32202 );
buf ( n381815 , n365670 );
nand ( n61252 , n381814 , n381815 );
buf ( n381817 , n61252 );
nand ( n61254 , n378141 , n22619 );
nand ( n61255 , n381817 , n61254 );
buf ( n381820 , n61255 );
buf ( n381821 , n45553 );
nand ( n381822 , n381820 , n381821 );
buf ( n381823 , n381822 );
nand ( n61260 , n61249 , n381823 );
not ( n381825 , n61260 );
not ( n61262 , n381825 );
or ( n381827 , n61246 , n61262 );
or ( n61264 , n381809 , n381825 );
nand ( n381829 , n381827 , n61264 );
xor ( n381830 , n381801 , n381829 );
not ( n61267 , n381830 );
buf ( n381832 , n364981 );
not ( n61269 , n381832 );
buf ( n381834 , n375903 );
not ( n381835 , n381834 );
or ( n381836 , n61269 , n381835 );
buf ( n381837 , n352192 );
buf ( n381838 , n364978 );
nand ( n381839 , n381837 , n381838 );
buf ( n381840 , n381839 );
buf ( n381841 , n381840 );
nand ( n61278 , n381836 , n381841 );
buf ( n381843 , n61278 );
and ( n381844 , n381843 , n365115 );
and ( n61281 , n352209 , n364978 );
not ( n381846 , n352209 );
and ( n61283 , n381846 , n364981 );
or ( n381848 , n61281 , n61283 );
and ( n381849 , n381848 , n365030 );
nor ( n61286 , n381844 , n381849 );
buf ( n381851 , n45075 );
not ( n381852 , n381851 );
xor ( n61289 , n342881 , n31072 );
buf ( n381854 , n61289 );
not ( n381855 , n381854 );
or ( n381856 , n381852 , n381855 );
buf ( n381857 , n342881 );
not ( n381858 , n381857 );
buf ( n381859 , n44638 );
not ( n61296 , n381859 );
or ( n381861 , n381858 , n61296 );
buf ( n381862 , n364808 );
buf ( n381863 , n365202 );
nand ( n381864 , n381862 , n381863 );
buf ( n381865 , n381864 );
buf ( n381866 , n381865 );
nand ( n61303 , n381861 , n381866 );
buf ( n381868 , n61303 );
buf ( n381869 , n381868 );
buf ( n381870 , n365226 );
nand ( n381871 , n381869 , n381870 );
buf ( n381872 , n381871 );
buf ( n381873 , n381872 );
nand ( n381874 , n381856 , n381873 );
buf ( n381875 , n381874 );
buf ( n381876 , n381875 );
not ( n381877 , n381876 );
buf ( n381878 , n381877 );
nand ( n61315 , n61286 , n381878 );
not ( n381880 , n61315 );
or ( n381881 , n61267 , n381880 );
buf ( n381882 , n381875 );
buf ( n381883 , n61286 );
not ( n381884 , n381883 );
buf ( n381885 , n381884 );
buf ( n381886 , n381885 );
nand ( n381887 , n381882 , n381886 );
buf ( n381888 , n381887 );
nand ( n61325 , n381881 , n381888 );
buf ( n381890 , n61325 );
buf ( n381891 , n377757 );
not ( n61328 , n381891 );
buf ( n381893 , n373924 );
not ( n61330 , n381893 );
or ( n381895 , n61328 , n61330 );
not ( n61332 , n365267 );
buf ( n381897 , n61332 );
buf ( n381898 , n378886 );
nand ( n381899 , n381897 , n381898 );
buf ( n381900 , n381899 );
buf ( n381901 , n381900 );
nand ( n381902 , n381895 , n381901 );
buf ( n381903 , n381902 );
buf ( n381904 , n381903 );
not ( n381905 , n381904 );
buf ( n381906 , n372247 );
not ( n381907 , n381906 );
or ( n61344 , n381905 , n381907 );
buf ( n381909 , n365303 );
buf ( n381910 , n378617 );
nand ( n61347 , n381909 , n381910 );
buf ( n381912 , n61347 );
buf ( n381913 , n381912 );
nand ( n61350 , n61344 , n381913 );
buf ( n61351 , n61350 );
buf ( n381916 , n61351 );
xor ( n61353 , n381890 , n381916 );
buf ( n381918 , n365030 );
not ( n381919 , n381918 );
buf ( n381920 , n381843 );
not ( n381921 , n381920 );
or ( n61358 , n381919 , n381921 );
buf ( n381923 , n378081 );
buf ( n381924 , n365115 );
nand ( n381925 , n381923 , n381924 );
buf ( n381926 , n381925 );
buf ( n381927 , n381926 );
nand ( n381928 , n61358 , n381927 );
buf ( n381929 , n381928 );
xor ( n381930 , n378520 , n58066 );
xor ( n381931 , n381930 , n58107 );
xor ( n381932 , n381929 , n381931 );
not ( n61369 , n56817 );
not ( n381934 , n60799 );
or ( n61371 , n61369 , n381934 );
nand ( n61372 , n58742 , n362386 );
nand ( n381937 , n61371 , n61372 );
xor ( n381938 , n381932 , n381937 );
buf ( n381939 , n381938 );
and ( n381940 , n61353 , n381939 );
and ( n381941 , n381890 , n381916 );
or ( n61378 , n381940 , n381941 );
buf ( n381943 , n61378 );
buf ( n381944 , n381943 );
and ( n61381 , n61234 , n381944 );
and ( n381946 , n381772 , n381797 );
or ( n61383 , n61381 , n381946 );
buf ( n381948 , n61383 );
buf ( n381949 , n381948 );
and ( n381950 , n381768 , n381949 );
buf ( n381951 , n381737 );
not ( n381952 , n381951 );
buf ( n381953 , n381764 );
nor ( n61390 , n381952 , n381953 );
buf ( n61391 , n61390 );
buf ( n381956 , n61391 );
nor ( n61393 , n381950 , n381956 );
buf ( n381958 , n61393 );
buf ( n381959 , n381958 );
not ( n381960 , n381959 );
buf ( n381961 , n381960 );
buf ( n381962 , n381961 );
not ( n381963 , n381962 );
or ( n61400 , n381718 , n381963 );
buf ( n381965 , n381713 );
not ( n61402 , n381965 );
buf ( n381967 , n381958 );
not ( n381968 , n381967 );
or ( n381969 , n61402 , n381968 );
not ( n61406 , n360610 );
not ( n381971 , n377146 );
and ( n381972 , n61406 , n381971 );
buf ( n381973 , n362452 );
not ( n381974 , n381973 );
buf ( n381975 , n377143 );
nor ( n381976 , n381974 , n381975 );
buf ( n381977 , n381976 );
nor ( n381978 , n381972 , n381977 );
buf ( n381979 , n381978 );
not ( n61416 , n381979 );
buf ( n61417 , n61416 );
buf ( n381982 , n61417 );
not ( n61419 , n381982 );
buf ( n381984 , n377370 );
not ( n381985 , n381984 );
or ( n381986 , n61419 , n381985 );
buf ( n381987 , n379664 );
buf ( n381988 , n371732 );
nand ( n61425 , n381987 , n381988 );
buf ( n381990 , n61425 );
buf ( n381991 , n381990 );
nand ( n381992 , n381986 , n381991 );
buf ( n381993 , n381992 );
buf ( n381994 , n381993 );
or ( n61431 , n381931 , n381929 );
nand ( n381996 , n61431 , n381937 );
nand ( n61433 , n381931 , n381929 );
nand ( n381998 , n381996 , n61433 );
buf ( n381999 , n381998 );
nand ( n61436 , n381994 , n381999 );
buf ( n382001 , n61436 );
buf ( n382002 , n381993 );
buf ( n382003 , n381998 );
or ( n382004 , n382002 , n382003 );
buf ( n382005 , n45015 );
not ( n382006 , n382005 );
xor ( n61443 , n57280 , n30911 );
buf ( n382008 , n61443 );
not ( n61445 , n382008 );
or ( n382010 , n382006 , n61445 );
buf ( n382011 , n378598 );
buf ( n382012 , n365152 );
nand ( n382013 , n382011 , n382012 );
buf ( n382014 , n382013 );
buf ( n382015 , n382014 );
nand ( n382016 , n382010 , n382015 );
buf ( n382017 , n382016 );
buf ( n382018 , n382017 );
buf ( n382019 , n365226 );
not ( n382020 , n382019 );
buf ( n382021 , n61289 );
not ( n382022 , n382021 );
or ( n61459 , n382020 , n382022 );
buf ( n382024 , n378014 );
buf ( n382025 , n45075 );
nand ( n61462 , n382024 , n382025 );
buf ( n382027 , n61462 );
buf ( n382028 , n382027 );
nand ( n61465 , n61459 , n382028 );
buf ( n382030 , n61465 );
buf ( n382031 , n382030 );
or ( n61468 , n382018 , n382031 );
buf ( n61469 , n61468 );
buf ( n382034 , n61469 );
buf ( n382035 , n381809 );
not ( n61472 , n382035 );
buf ( n382037 , n61260 );
not ( n61474 , n382037 );
or ( n61475 , n61472 , n61474 );
buf ( n382040 , n61260 );
buf ( n382041 , n381809 );
or ( n382042 , n382040 , n382041 );
buf ( n382043 , n381801 );
nand ( n382044 , n382042 , n382043 );
buf ( n382045 , n382044 );
buf ( n382046 , n382045 );
nand ( n382047 , n61475 , n382046 );
buf ( n382048 , n382047 );
buf ( n382049 , n382048 );
and ( n61486 , n382034 , n382049 );
buf ( n382051 , n382030 );
buf ( n61488 , n382017 );
and ( n61489 , n382051 , n61488 );
buf ( n382054 , n61489 );
buf ( n382055 , n382054 );
nor ( n61492 , n61486 , n382055 );
buf ( n382057 , n61492 );
buf ( n382058 , n382057 );
not ( n61495 , n382058 );
buf ( n382060 , n61495 );
buf ( n382061 , n382060 );
nand ( n61498 , n382004 , n382061 );
buf ( n382063 , n61498 );
nand ( n382064 , n382001 , n382063 );
and ( n61501 , n360885 , n377592 );
not ( n61502 , n360885 );
and ( n61503 , n61502 , n377585 );
nor ( n382068 , n61501 , n61503 );
not ( n382069 , n382068 );
not ( n61506 , n377618 );
and ( n61507 , n382069 , n61506 );
and ( n61508 , n57529 , n377580 );
nor ( n382073 , n61507 , n61508 );
and ( n382074 , n382064 , n382073 );
not ( n61511 , n382064 );
not ( n61512 , n382073 );
and ( n61513 , n61511 , n61512 );
nor ( n382078 , n382074 , n61513 );
buf ( n382079 , n379299 );
not ( n61516 , n382079 );
not ( n61517 , n379274 );
not ( n61518 , n367158 );
or ( n61519 , n61517 , n61518 );
buf ( n382084 , n40251 );
buf ( n382085 , n379271 );
nand ( n61520 , n382084 , n382085 );
buf ( n382087 , n61520 );
nand ( n382088 , n61519 , n382087 );
buf ( n382089 , n382088 );
not ( n382090 , n382089 );
or ( n61525 , n61516 , n382090 );
buf ( n382092 , n379452 );
buf ( n382093 , n379263 );
nand ( n382094 , n382092 , n382093 );
buf ( n382095 , n382094 );
buf ( n382096 , n382095 );
nand ( n382097 , n61525 , n382096 );
buf ( n382098 , n382097 );
and ( n382099 , n382078 , n382098 );
not ( n61534 , n382078 );
buf ( n382101 , n382098 );
not ( n382102 , n382101 );
buf ( n382103 , n382102 );
and ( n61538 , n61534 , n382103 );
nor ( n382105 , n382099 , n61538 );
buf ( n382106 , n382105 );
not ( n61541 , n382106 );
buf ( n61542 , n61541 );
not ( n382109 , n61542 );
not ( n61544 , n56687 );
not ( n382111 , n365948 );
or ( n61546 , n61544 , n382111 );
nand ( n382113 , n377094 , n360068 );
nand ( n382114 , n61546 , n382113 );
buf ( n382115 , n382114 );
not ( n382116 , n382115 );
buf ( n382117 , n45345 );
not ( n382118 , n382117 );
or ( n382119 , n382116 , n382118 );
buf ( n382120 , n377068 );
not ( n382121 , n382120 );
buf ( n382122 , n365945 );
not ( n382123 , n382122 );
or ( n382124 , n382121 , n382123 );
buf ( n382125 , n365528 );
buf ( n382126 , n377071 );
nand ( n382127 , n382125 , n382126 );
buf ( n382128 , n382127 );
buf ( n382129 , n382128 );
nand ( n382130 , n382124 , n382129 );
buf ( n382131 , n382130 );
buf ( n382132 , n382131 );
buf ( n382133 , n365954 );
nand ( n382134 , n382132 , n382133 );
buf ( n382135 , n382134 );
buf ( n382136 , n382135 );
nand ( n382137 , n382119 , n382136 );
buf ( n382138 , n382137 );
not ( n382139 , n382138 );
buf ( n382140 , n377122 );
not ( n382141 , n382140 );
buf ( n382142 , n365468 );
not ( n382143 , n382142 );
or ( n382144 , n382141 , n382143 );
buf ( n382145 , n360610 );
buf ( n382146 , n57463 );
nand ( n382147 , n382145 , n382146 );
buf ( n382148 , n382147 );
buf ( n382149 , n382148 );
nand ( n382150 , n382144 , n382149 );
buf ( n382151 , n382150 );
not ( n382152 , n382151 );
and ( n61557 , n360583 , n40473 );
not ( n61558 , n61557 );
or ( n382155 , n382152 , n61558 );
or ( n61560 , n381978 , n360571 );
nand ( n61561 , n382155 , n61560 );
not ( n61562 , n61561 );
or ( n61563 , n382139 , n61562 );
buf ( n382160 , n61561 );
not ( n61565 , n382160 );
buf ( n382162 , n61565 );
not ( n61567 , n382162 );
buf ( n382164 , n382138 );
not ( n61569 , n382164 );
buf ( n382166 , n61569 );
not ( n61571 , n382166 );
or ( n61572 , n61567 , n61571 );
xor ( n61573 , n382051 , n61488 );
buf ( n382170 , n61573 );
buf ( n382171 , n382170 );
buf ( n382172 , n382048 );
and ( n61577 , n382171 , n382172 );
not ( n61578 , n382171 );
buf ( n382175 , n382048 );
not ( n61580 , n382175 );
buf ( n382177 , n61580 );
buf ( n382178 , n382177 );
and ( n61583 , n61578 , n382178 );
nor ( n61584 , n61577 , n61583 );
buf ( n382181 , n61584 );
buf ( n382182 , n382181 );
buf ( n382183 , n382182 );
buf ( n382184 , n382183 );
nand ( n382185 , n61572 , n382184 );
nand ( n61590 , n61563 , n382185 );
buf ( n382187 , n61590 );
not ( n61592 , n379263 );
not ( n61593 , n382088 );
or ( n382190 , n61592 , n61593 );
buf ( n382191 , n379274 );
not ( n61596 , n382191 );
buf ( n382193 , n360848 );
not ( n382194 , n382193 );
or ( n61599 , n61596 , n382194 );
buf ( n382196 , n369722 );
not ( n61601 , n382196 );
buf ( n382198 , n379271 );
nand ( n61603 , n61601 , n382198 );
buf ( n382200 , n61603 );
buf ( n382201 , n382200 );
nand ( n61606 , n61599 , n382201 );
buf ( n382203 , n61606 );
buf ( n382204 , n382203 );
buf ( n382205 , n379299 );
nand ( n61610 , n382204 , n382205 );
buf ( n382207 , n61610 );
nand ( n61612 , n382190 , n382207 );
buf ( n382209 , n61612 );
xor ( n382210 , n382187 , n382209 );
not ( n61613 , n379893 );
nand ( n61614 , n61613 , n60547 );
and ( n61615 , n379841 , n366725 );
not ( n61616 , n379841 );
and ( n61617 , n61616 , n366722 );
or ( n61618 , n61615 , n61617 );
buf ( n382217 , n61618 );
buf ( n382218 , n379916 );
nand ( n382219 , n382217 , n382218 );
buf ( n382220 , n382219 );
nand ( n61623 , n61614 , n382220 );
buf ( n382222 , n61623 );
and ( n382223 , n382210 , n382222 );
and ( n61626 , n382187 , n382209 );
or ( n382225 , n382223 , n61626 );
buf ( n382226 , n382225 );
not ( n61629 , n382226 );
or ( n382228 , n382109 , n61629 );
not ( n382229 , n382105 );
buf ( n61632 , n382226 );
not ( n61633 , n61632 );
buf ( n61634 , n61633 );
not ( n382233 , n61634 );
or ( n61636 , n382229 , n382233 );
buf ( n382235 , n57530 );
not ( n382236 , n382235 );
buf ( n382237 , n377585 );
not ( n61640 , n382237 );
buf ( n382239 , n362288 );
not ( n61642 , n382239 );
or ( n61643 , n61640 , n61642 );
buf ( n382242 , n362285 );
buf ( n382243 , n377592 );
nand ( n61646 , n382242 , n382243 );
buf ( n382245 , n61646 );
buf ( n382246 , n382245 );
nand ( n61649 , n61643 , n382246 );
buf ( n382248 , n61649 );
buf ( n382249 , n382248 );
not ( n61652 , n382249 );
or ( n382251 , n382236 , n61652 );
buf ( n382252 , n382068 );
not ( n382253 , n382252 );
buf ( n382254 , n377580 );
nand ( n382255 , n382253 , n382254 );
buf ( n382256 , n382255 );
buf ( n382257 , n382256 );
nand ( n61660 , n382251 , n382257 );
buf ( n382259 , n61660 );
buf ( n382260 , n382259 );
not ( n61663 , n382260 );
buf ( n382262 , n58744 );
xor ( n382263 , n379218 , n379212 );
xor ( n61666 , n382262 , n382263 );
buf ( n382265 , n44915 );
not ( n382266 , n382265 );
buf ( n382267 , n377953 );
not ( n382268 , n382267 );
or ( n382269 , n382266 , n382268 );
buf ( n382270 , n380511 );
buf ( n382271 , n47466 );
nand ( n61674 , n382270 , n382271 );
buf ( n382273 , n61674 );
buf ( n382274 , n382273 );
nand ( n382275 , n382269 , n382274 );
buf ( n382276 , n382275 );
not ( n382277 , n382276 );
and ( n382278 , n61666 , n382277 );
not ( n61681 , n61666 );
and ( n382280 , n61681 , n382276 );
nor ( n382281 , n382278 , n382280 );
not ( n61684 , n382281 );
not ( n382283 , n381125 );
not ( n382284 , n39207 );
and ( n61687 , n382283 , n382284 );
and ( n61688 , n377916 , n39217 );
nor ( n61689 , n61687 , n61688 );
not ( n61690 , n61689 );
or ( n382289 , n61684 , n61690 );
not ( n382290 , n382281 );
not ( n61693 , n61689 );
nand ( n382292 , n382290 , n61693 );
nand ( n382293 , n382289 , n382292 );
buf ( n61696 , n382293 );
not ( n61697 , n61696 );
buf ( n61698 , n61697 );
buf ( n382297 , n61698 );
not ( n382298 , n382297 );
or ( n61701 , n61663 , n382298 );
buf ( n382300 , n61698 );
buf ( n382301 , n382259 );
or ( n61704 , n382300 , n382301 );
buf ( n382303 , n382057 );
buf ( n61706 , n381998 );
not ( n382305 , n61706 );
buf ( n382306 , n382305 );
buf ( n382307 , n382306 );
and ( n61710 , n382303 , n382307 );
not ( n382309 , n382303 );
buf ( n382310 , n381998 );
and ( n61713 , n382309 , n382310 );
nor ( n382312 , n61710 , n61713 );
buf ( n382313 , n382312 );
buf ( n382314 , n382313 );
not ( n382315 , n382314 );
buf ( n382316 , n381993 );
not ( n61719 , n382316 );
buf ( n61720 , n61719 );
buf ( n61721 , n61720 );
not ( n61722 , n61721 );
and ( n61723 , n382315 , n61722 );
buf ( n382322 , n61720 );
buf ( n382323 , n382313 );
and ( n61726 , n382322 , n382323 );
nor ( n382325 , n61723 , n61726 );
buf ( n382326 , n382325 );
buf ( n382327 , n382326 );
not ( n382328 , n382327 );
buf ( n382329 , n382328 );
buf ( n382330 , n382329 );
nand ( n61733 , n61704 , n382330 );
buf ( n382332 , n61733 );
buf ( n382333 , n382332 );
nand ( n382334 , n61701 , n382333 );
buf ( n382335 , n382334 );
nand ( n61738 , n61636 , n382335 );
nand ( n382337 , n382228 , n61738 );
buf ( n382338 , n382337 );
nand ( n61741 , n381969 , n382338 );
buf ( n382340 , n61741 );
buf ( n382341 , n382340 );
nand ( n61744 , n61400 , n382341 );
buf ( n382343 , n61744 );
buf ( n382344 , n382343 );
xor ( n61747 , n61146 , n382344 );
buf ( n382346 , n61747 );
buf ( n382347 , n382346 );
not ( n382348 , n382347 );
buf ( n382349 , n382337 );
not ( n61752 , n382349 );
buf ( n382351 , n381958 );
not ( n61754 , n382351 );
and ( n382353 , n61752 , n61754 );
buf ( n382354 , n382337 );
buf ( n382355 , n381958 );
and ( n382356 , n382354 , n382355 );
nor ( n61759 , n382353 , n382356 );
buf ( n61760 , n61759 );
buf ( n382359 , n61760 );
buf ( n382360 , n381713 );
buf ( n382361 , n382360 );
buf ( n382362 , n382361 );
buf ( n382363 , n382362 );
not ( n61766 , n382363 );
buf ( n382365 , n61766 );
buf ( n382366 , n382365 );
and ( n382367 , n382359 , n382366 );
not ( n61770 , n382359 );
buf ( n382369 , n382362 );
and ( n382370 , n61770 , n382369 );
nor ( n382371 , n382367 , n382370 );
buf ( n382372 , n382371 );
buf ( n382373 , n382372 );
not ( n61776 , n382373 );
buf ( n382375 , n61776 );
not ( n61778 , n382375 );
buf ( n382377 , n382335 );
buf ( n382378 , n382226 );
buf ( n61781 , n382378 );
buf ( n382380 , n61781 );
buf ( n382381 , n382380 );
xor ( n61784 , n382377 , n382381 );
buf ( n382383 , n61542 );
xor ( n61786 , n61784 , n382383 );
buf ( n382385 , n61786 );
buf ( n382386 , n381737 );
buf ( n382387 , n381948 );
xor ( n61790 , n382386 , n382387 );
buf ( n382389 , n381764 );
xnor ( n61792 , n61790 , n382389 );
buf ( n382391 , n61792 );
buf ( n382392 , n382391 );
not ( n61795 , n382392 );
buf ( n382394 , n61795 );
buf ( n382395 , n382394 );
xor ( n61798 , n381066 , n381389 );
xor ( n61799 , n61798 , n381469 );
buf ( n382398 , n61799 );
not ( n61801 , n382398 );
buf ( n382400 , n61801 );
buf ( n382401 , n382400 );
nand ( n382402 , n382395 , n382401 );
buf ( n382403 , n382402 );
and ( n61806 , n382385 , n382403 );
and ( n382405 , n382391 , n61799 );
nor ( n382406 , n61806 , n382405 );
buf ( n382407 , n382406 );
not ( n382408 , n382407 );
buf ( n382409 , n382408 );
not ( n61812 , n382409 );
or ( n382411 , n61778 , n61812 );
not ( n382412 , n382406 );
not ( n61815 , n382372 );
or ( n382414 , n382412 , n61815 );
xor ( n61817 , n381772 , n381797 );
xor ( n61818 , n61817 , n381944 );
buf ( n382417 , n61818 );
buf ( n382418 , n382417 );
not ( n61821 , n382418 );
buf ( n61822 , n61821 );
buf ( n382421 , n61822 );
not ( n61824 , n382421 );
and ( n382423 , n381383 , n381145 );
not ( n382424 , n381383 );
and ( n61827 , n382424 , n60609 );
or ( n61828 , n382423 , n61827 );
and ( n61829 , n61828 , n381163 );
not ( n382428 , n61828 );
and ( n382429 , n382428 , n381166 );
nor ( n61832 , n61829 , n382429 );
buf ( n382431 , n61832 );
not ( n61834 , n382431 );
or ( n382433 , n61824 , n61834 );
buf ( n382434 , n382259 );
not ( n61837 , n382434 );
buf ( n382436 , n382326 );
not ( n382437 , n382436 );
or ( n382438 , n61837 , n382437 );
buf ( n382439 , n382259 );
buf ( n382440 , n382326 );
or ( n61843 , n382439 , n382440 );
nand ( n382442 , n382438 , n61843 );
buf ( n382443 , n382442 );
buf ( n382444 , n382443 );
buf ( n382445 , n382293 );
and ( n382446 , n382444 , n382445 );
not ( n61849 , n382444 );
buf ( n382448 , n61698 );
and ( n382449 , n61849 , n382448 );
nor ( n61852 , n382446 , n382449 );
buf ( n61853 , n61852 );
not ( n382452 , n61853 );
buf ( n382453 , n382452 );
nand ( n382454 , n382433 , n382453 );
buf ( n382455 , n382454 );
buf ( n382456 , n382455 );
not ( n382457 , n61832 );
nand ( n382458 , n382457 , n382417 );
buf ( n382459 , n382458 );
nand ( n382460 , n382456 , n382459 );
buf ( n382461 , n382460 );
buf ( n382462 , n365152 );
not ( n382463 , n382462 );
buf ( n382464 , n61443 );
not ( n382465 , n382464 );
or ( n61868 , n382463 , n382465 );
buf ( n382467 , n57280 );
not ( n382468 , n382467 );
buf ( n382469 , n364855 );
not ( n382470 , n382469 );
or ( n61873 , n382468 , n382470 );
buf ( n382472 , n351367 );
buf ( n382473 , n377728 );
nand ( n61876 , n382472 , n382473 );
buf ( n382475 , n61876 );
buf ( n382476 , n382475 );
nand ( n382477 , n61873 , n382476 );
buf ( n382478 , n382477 );
buf ( n382479 , n382478 );
buf ( n382480 , n365186 );
nand ( n61883 , n382479 , n382480 );
buf ( n382482 , n61883 );
buf ( n382483 , n382482 );
nand ( n61886 , n61868 , n382483 );
buf ( n382485 , n61886 );
buf ( n382486 , n382485 );
buf ( n382487 , n56794 );
not ( n382488 , n382487 );
buf ( n382489 , n61255 );
not ( n382490 , n382489 );
or ( n61893 , n382488 , n382490 );
buf ( n382492 , n22619 );
not ( n382493 , n382492 );
buf ( n382494 , n31231 );
not ( n382495 , n382494 );
buf ( n382496 , n382495 );
buf ( n382497 , n382496 );
not ( n61900 , n382497 );
or ( n382499 , n382493 , n61900 );
buf ( n382500 , n31231 );
not ( n61903 , n342564 );
buf ( n382502 , n61903 );
nand ( n382503 , n382500 , n382502 );
buf ( n382504 , n382503 );
buf ( n382505 , n382504 );
nand ( n382506 , n382499 , n382505 );
buf ( n382507 , n382506 );
buf ( n382508 , n382507 );
buf ( n382509 , n45553 );
nand ( n61912 , n382508 , n382509 );
buf ( n382511 , n61912 );
buf ( n382512 , n382511 );
nand ( n61915 , n61893 , n382512 );
buf ( n382514 , n61915 );
xor ( n382515 , n380589 , n380613 );
xor ( n61918 , n382515 , n380617 );
xor ( n382517 , n380775 , n380873 );
xor ( n382518 , n61918 , n382517 );
not ( n61921 , n382518 );
xor ( n382520 , n380691 , n380748 );
xor ( n382521 , n382520 , n380766 );
buf ( n382522 , n382521 );
buf ( n382523 , n380680 );
buf ( n382524 , n376866 );
and ( n382525 , n382523 , n382524 );
buf ( n382526 , n60171 );
buf ( n382527 , n376875 );
and ( n382528 , n382526 , n382527 );
nor ( n382529 , n382525 , n382528 );
buf ( n382530 , n382529 );
buf ( n382531 , n382530 );
buf ( n382532 , n376924 );
or ( n61935 , n382531 , n382532 );
buf ( n382534 , n380757 );
buf ( n382535 , n56517 );
or ( n382536 , n382534 , n382535 );
nand ( n61939 , n61935 , n382536 );
buf ( n382538 , n61939 );
buf ( n382539 , n382538 );
buf ( n382540 , n378214 );
buf ( n382541 , n380570 );
and ( n382542 , n382540 , n382541 );
buf ( n382543 , n57754 );
buf ( n382544 , n60054 );
and ( n382545 , n382543 , n382544 );
nor ( n61948 , n382542 , n382545 );
buf ( n61949 , n61948 );
buf ( n382548 , n61949 );
buf ( n382549 , n380581 );
or ( n382550 , n382548 , n382549 );
buf ( n382551 , n380803 );
buf ( n382552 , n378453 );
or ( n382553 , n382551 , n382552 );
nand ( n382554 , n382550 , n382553 );
buf ( n382555 , n382554 );
buf ( n382556 , n382555 );
xor ( n382557 , n382539 , n382556 );
buf ( n382558 , n60089 );
buf ( n382559 , n57800 );
and ( n382560 , n382558 , n382559 );
buf ( n382561 , n60094 );
buf ( n382562 , n376903 );
and ( n61965 , n382561 , n382562 );
nor ( n382564 , n382560 , n61965 );
buf ( n382565 , n382564 );
buf ( n382566 , n382565 );
buf ( n382567 , n378341 );
or ( n61970 , n382566 , n382567 );
buf ( n382569 , n380786 );
buf ( n382570 , n378424 );
or ( n61973 , n382569 , n382570 );
nand ( n61974 , n61970 , n61973 );
buf ( n382573 , n61974 );
buf ( n382574 , n382573 );
and ( n61977 , n382557 , n382574 );
and ( n61978 , n382539 , n382556 );
or ( n61979 , n61977 , n61978 );
buf ( n382578 , n61979 );
xor ( n382579 , n382522 , n382578 );
xor ( n61982 , n380795 , n380812 );
xor ( n382581 , n61982 , n380854 );
buf ( n382582 , n382581 );
and ( n382583 , n382579 , n382582 );
and ( n61986 , n382522 , n382578 );
or ( n382585 , n382583 , n61986 );
xor ( n382586 , n380858 , n380866 );
xor ( n61989 , n382586 , n380870 );
and ( n382588 , n382585 , n61989 );
nand ( n382589 , n55685 , n56321 );
xnor ( n61992 , n56317 , n382589 );
buf ( n382591 , n61992 );
buf ( n382592 , n376990 );
and ( n382593 , n382591 , n382592 );
buf ( n382594 , n61992 );
not ( n61997 , n382594 );
buf ( n382596 , n61997 );
buf ( n382597 , n382596 );
buf ( n382598 , n376997 );
and ( n62001 , n382597 , n382598 );
buf ( n382600 , n377003 );
nor ( n62003 , n382593 , n62001 , n382600 );
buf ( n382602 , n62003 );
not ( n62005 , n376790 );
not ( n62006 , n62005 );
not ( n62007 , n380719 );
or ( n382606 , n62006 , n62007 );
not ( n382607 , n380722 );
nand ( n382608 , n382606 , n382607 );
nor ( n62011 , n60193 , n376810 );
xor ( n382610 , n382608 , n62011 );
buf ( n382611 , n382610 );
not ( n62014 , n56360 );
nand ( n62015 , n380710 , n376781 );
not ( n62016 , n62015 );
not ( n62017 , n62016 );
or ( n382616 , n62014 , n62017 );
and ( n62019 , n56360 , n56364 );
nand ( n382618 , n376792 , n56379 );
nor ( n62021 , n62019 , n382618 );
nand ( n62022 , n382616 , n62021 );
not ( n62023 , n56391 );
nand ( n62024 , n62022 , n62023 );
nand ( n382623 , n376787 , n56395 );
xnor ( n62026 , n62024 , n382623 );
buf ( n382625 , n62026 );
not ( n62028 , n382625 );
buf ( n382627 , n62028 );
buf ( n382628 , n382627 );
and ( n382629 , n382611 , n382628 );
not ( n382630 , n382611 );
buf ( n382631 , n62026 );
and ( n382632 , n382630 , n382631 );
nor ( n382633 , n382629 , n382632 );
buf ( n382634 , n382633 );
buf ( n382635 , n382634 );
buf ( n382636 , n60214 );
not ( n382637 , n382636 );
buf ( n382638 , n382637 );
buf ( n382639 , n382638 );
buf ( n382640 , n382610 );
not ( n62043 , n382640 );
buf ( n382642 , n62043 );
buf ( n382643 , n382642 );
and ( n62046 , n382639 , n382643 );
buf ( n382645 , n382638 );
not ( n62048 , n382645 );
buf ( n382647 , n62048 );
buf ( n382648 , n382647 );
buf ( n382649 , n382610 );
and ( n382650 , n382648 , n382649 );
nor ( n382651 , n62046 , n382650 );
buf ( n382652 , n382651 );
buf ( n382653 , n382652 );
and ( n62056 , n382635 , n382653 );
buf ( n382655 , n62056 );
buf ( n382656 , n382655 );
buf ( n382657 , n382647 );
nand ( n62060 , n382656 , n382657 );
buf ( n382659 , n62060 );
buf ( n382660 , n382659 );
buf ( n382661 , n382634 );
not ( n62064 , n382661 );
buf ( n382663 , n62064 );
buf ( n382664 , n382663 );
buf ( n382665 , n382647 );
nand ( n62068 , n382664 , n382665 );
buf ( n382667 , n62068 );
buf ( n382668 , n382667 );
and ( n382669 , n382660 , n382668 );
buf ( n382670 , n382669 );
xor ( n382671 , n382602 , n382670 );
buf ( n382672 , n378368 );
buf ( n382673 , n380570 );
and ( n382674 , n382672 , n382673 );
buf ( n382675 , n378372 );
buf ( n382676 , n60054 );
and ( n382677 , n382675 , n382676 );
nor ( n62080 , n382674 , n382677 );
buf ( n62081 , n62080 );
buf ( n382680 , n62081 );
buf ( n382681 , n380581 );
or ( n62084 , n382680 , n382681 );
buf ( n382683 , n61949 );
buf ( n382684 , n378453 );
or ( n382685 , n382683 , n382684 );
nand ( n62088 , n62084 , n382685 );
buf ( n382687 , n62088 );
and ( n382688 , n382671 , n382687 );
and ( n62091 , n382602 , n382670 );
or ( n382690 , n382688 , n62091 );
buf ( n62093 , n382690 );
buf ( n382692 , n380850 );
not ( n62095 , n382692 );
buf ( n382694 , n380831 );
not ( n62097 , n382694 );
or ( n62098 , n62095 , n62097 );
buf ( n382697 , n380853 );
nand ( n62100 , n62098 , n382697 );
buf ( n62101 , n62100 );
buf ( n382700 , n62101 );
xor ( n62103 , n62093 , n382700 );
buf ( n382702 , n380651 );
buf ( n382703 , n57800 );
and ( n62106 , n382702 , n382703 );
buf ( n382705 , n380657 );
buf ( n382706 , n376903 );
and ( n382707 , n382705 , n382706 );
nor ( n382708 , n62106 , n382707 );
buf ( n382709 , n382708 );
buf ( n382710 , n382709 );
buf ( n382711 , n378341 );
or ( n382712 , n382710 , n382711 );
buf ( n382713 , n382565 );
buf ( n382714 , n378424 );
or ( n382715 , n382713 , n382714 );
nand ( n62118 , n382712 , n382715 );
buf ( n382717 , n62118 );
buf ( n382718 , n382717 );
buf ( n382719 , n376971 );
buf ( n382720 , n380817 );
and ( n62123 , n382719 , n382720 );
buf ( n382722 , n376993 );
buf ( n382723 , n57983 );
and ( n382724 , n382722 , n382723 );
nor ( n62127 , n62123 , n382724 );
buf ( n382726 , n62127 );
buf ( n382727 , n382726 );
buf ( n382728 , n60313 );
or ( n62131 , n382727 , n382728 );
buf ( n382730 , n380824 );
buf ( n382731 , n380733 );
or ( n62134 , n382730 , n382731 );
nand ( n382733 , n62131 , n62134 );
buf ( n382734 , n382733 );
buf ( n382735 , n382734 );
xor ( n382736 , n382718 , n382735 );
buf ( n382737 , n380838 );
buf ( n382738 , n376866 );
and ( n382739 , n382737 , n382738 );
buf ( n382740 , n380844 );
buf ( n382741 , n376866 );
not ( n382742 , n382741 );
buf ( n382743 , n382742 );
buf ( n382744 , n382743 );
and ( n62147 , n382740 , n382744 );
nor ( n62148 , n382739 , n62147 );
buf ( n382747 , n62148 );
buf ( n382748 , n382747 );
buf ( n382749 , n376924 );
or ( n62152 , n382748 , n382749 );
buf ( n382751 , n382530 );
buf ( n382752 , n56517 );
or ( n382753 , n382751 , n382752 );
nand ( n382754 , n62152 , n382753 );
buf ( n382755 , n382754 );
buf ( n382756 , n382755 );
and ( n62159 , n382736 , n382756 );
and ( n62160 , n382718 , n382735 );
or ( n382759 , n62159 , n62160 );
buf ( n382760 , n382759 );
buf ( n382761 , n382760 );
and ( n382762 , n62103 , n382761 );
and ( n382763 , n62093 , n382700 );
or ( n62166 , n382762 , n382763 );
buf ( n382765 , n62166 );
xor ( n382766 , n382522 , n382578 );
xor ( n382767 , n382766 , n382582 );
and ( n62170 , n382765 , n382767 );
buf ( n382769 , n61992 );
buf ( n382770 , n376866 );
and ( n62173 , n382769 , n382770 );
buf ( n382772 , n382596 );
buf ( n382773 , n382743 );
and ( n62176 , n382772 , n382773 );
nor ( n62177 , n62173 , n62176 );
buf ( n382776 , n62177 );
buf ( n382777 , n382776 );
buf ( n382778 , n376924 );
or ( n382779 , n382777 , n382778 );
buf ( n382780 , n382747 );
buf ( n382781 , n56517 );
or ( n62184 , n382780 , n382781 );
nand ( n62185 , n382779 , n62184 );
buf ( n382784 , n62185 );
buf ( n382785 , n382784 );
not ( n382786 , n376226 );
nand ( n62189 , n382786 , n376714 );
not ( n62190 , n376219 );
not ( n382789 , n62190 );
not ( n382790 , n56309 );
or ( n62193 , n382789 , n382790 );
nand ( n382792 , n62193 , n56312 );
or ( n382793 , n62189 , n382792 );
nand ( n62196 , n382792 , n62189 );
nand ( n382795 , n382793 , n62196 );
buf ( n382796 , n382795 );
buf ( n382797 , n376990 );
and ( n382798 , n382796 , n382797 );
or ( n62201 , n62189 , n382792 );
nand ( n62202 , n62201 , n62196 );
buf ( n62203 , n62202 );
not ( n382802 , n62203 );
buf ( n382803 , n382802 );
buf ( n382804 , n382803 );
buf ( n382805 , n376997 );
and ( n62208 , n382804 , n382805 );
buf ( n382807 , n377003 );
nor ( n382808 , n382798 , n62208 , n382807 );
buf ( n382809 , n382808 );
buf ( n382810 , n382809 );
or ( n382811 , n382785 , n382810 );
buf ( n382812 , n382811 );
xor ( n382813 , n382602 , n382670 );
xor ( n62216 , n382813 , n382687 );
and ( n62217 , n382812 , n62216 );
buf ( n382816 , n378214 );
buf ( n382817 , n380817 );
and ( n62220 , n382816 , n382817 );
buf ( n382819 , n57754 );
buf ( n382820 , n57983 );
and ( n62223 , n382819 , n382820 );
nor ( n382822 , n62220 , n62223 );
buf ( n382823 , n382822 );
buf ( n382824 , n382823 );
buf ( n382825 , n60313 );
or ( n382826 , n382824 , n382825 );
buf ( n382827 , n382726 );
buf ( n382828 , n380733 );
or ( n62231 , n382827 , n382828 );
nand ( n62232 , n382826 , n62231 );
buf ( n382831 , n62232 );
buf ( n382832 , n376743 );
buf ( n382833 , n382638 );
buf ( n382834 , n382833 );
buf ( n382835 , n382834 );
buf ( n382836 , n382835 );
and ( n382837 , n382832 , n382836 );
buf ( n382838 , n376871 );
buf ( n382839 , n382835 );
not ( n62242 , n382839 );
buf ( n62243 , n62242 );
buf ( n382842 , n62243 );
and ( n62245 , n382838 , n382842 );
nor ( n382844 , n382837 , n62245 );
buf ( n382845 , n382844 );
buf ( n382846 , n382845 );
buf ( n382847 , n382655 );
not ( n62250 , n382847 );
buf ( n382849 , n62250 );
buf ( n382850 , n382849 );
or ( n62253 , n382846 , n382850 );
buf ( n382852 , n382667 );
nand ( n382853 , n62253 , n382852 );
buf ( n382854 , n382853 );
xor ( n382855 , n382831 , n382854 );
buf ( n382856 , n60089 );
buf ( n382857 , n380570 );
and ( n382858 , n382856 , n382857 );
buf ( n382859 , n60094 );
buf ( n382860 , n60054 );
and ( n382861 , n382859 , n382860 );
nor ( n62264 , n382858 , n382861 );
buf ( n382863 , n62264 );
buf ( n382864 , n382863 );
buf ( n382865 , n380581 );
or ( n62268 , n382864 , n382865 );
buf ( n382867 , n62081 );
buf ( n382868 , n378453 );
or ( n62271 , n382867 , n382868 );
nand ( n382870 , n62268 , n62271 );
buf ( n382871 , n382870 );
and ( n62274 , n382855 , n382871 );
and ( n62275 , n382831 , n382854 );
or ( n62276 , n62274 , n62275 );
xor ( n382875 , n382602 , n382670 );
xor ( n382876 , n382875 , n382687 );
and ( n62279 , n62276 , n382876 );
and ( n382878 , n382812 , n62276 );
or ( n382879 , n62217 , n62279 , n382878 );
xor ( n62282 , n382539 , n382556 );
xor ( n382881 , n62282 , n382574 );
buf ( n382882 , n382881 );
xor ( n62285 , n382879 , n382882 );
xor ( n62286 , n62093 , n382700 );
xor ( n382885 , n62286 , n382761 );
buf ( n382886 , n382885 );
and ( n62289 , n62285 , n382886 );
and ( n62290 , n382879 , n382882 );
or ( n62291 , n62289 , n62290 );
xor ( n382890 , n382522 , n382578 );
xor ( n382891 , n382890 , n382582 );
and ( n62294 , n62291 , n382891 );
and ( n62295 , n382765 , n62291 );
or ( n62296 , n62170 , n62294 , n62295 );
xor ( n382895 , n380858 , n380866 );
xor ( n382896 , n382895 , n380870 );
and ( n62299 , n62296 , n382896 );
and ( n382898 , n382585 , n62296 );
or ( n382899 , n382588 , n62299 , n382898 );
not ( n62302 , n382899 );
nand ( n382901 , n61921 , n62302 );
not ( n62304 , n382901 );
buf ( n382903 , n351160 );
not ( n382904 , n382903 );
buf ( n382905 , n366659 );
not ( n382906 , n382905 );
or ( n62309 , n382904 , n382906 );
buf ( n382908 , n378135 );
buf ( n382909 , n381266 );
nand ( n62312 , n382908 , n382909 );
buf ( n382911 , n62312 );
buf ( n382912 , n382911 );
nand ( n62314 , n62309 , n382912 );
buf ( n382914 , n62314 );
buf ( n382915 , n382914 );
not ( n62317 , n382915 );
buf ( n382917 , n375896 );
not ( n382918 , n382917 );
or ( n62319 , n62317 , n382918 );
buf ( n382920 , n381228 );
buf ( n382921 , n375920 );
nand ( n62322 , n382920 , n382921 );
buf ( n382923 , n62322 );
buf ( n382924 , n382923 );
nand ( n62325 , n62319 , n382924 );
buf ( n382926 , n62325 );
not ( n62327 , n382926 );
or ( n62328 , n62304 , n62327 );
nand ( n62329 , n382899 , n382518 );
nand ( n62330 , n62328 , n62329 );
xor ( n62331 , n382514 , n62330 );
buf ( n382932 , n365115 );
not ( n62333 , n382932 );
buf ( n382934 , n381848 );
not ( n62335 , n382934 );
or ( n62336 , n62333 , n62335 );
not ( n62337 , n22547 );
not ( n62338 , n342499 );
or ( n62339 , n62337 , n62338 );
nand ( n62340 , n62339 , n342502 );
not ( n62341 , n62340 );
not ( n62342 , n351292 );
or ( n62343 , n62341 , n62342 );
buf ( n382944 , n377301 );
not ( n62345 , n62340 );
buf ( n382946 , n62345 );
nand ( n62347 , n382944 , n382946 );
buf ( n382948 , n62347 );
nand ( n62349 , n62343 , n382948 );
buf ( n382950 , n62349 );
buf ( n382951 , n365024 );
nand ( n62352 , n382950 , n382951 );
buf ( n382953 , n62352 );
buf ( n382954 , n382953 );
nand ( n62355 , n62336 , n382954 );
buf ( n382956 , n62355 );
and ( n382957 , n62331 , n382956 );
and ( n382958 , n382514 , n62330 );
or ( n382959 , n382957 , n382958 );
buf ( n382960 , n382959 );
xor ( n382961 , n382486 , n382960 );
buf ( n382962 , n368994 );
not ( n382963 , n382962 );
buf ( n382964 , n378032 );
not ( n382965 , n382964 );
or ( n382966 , n382963 , n382965 );
buf ( n382967 , n365319 );
buf ( n382968 , n57053 );
nand ( n382969 , n382967 , n382968 );
buf ( n382970 , n382969 );
buf ( n382971 , n382970 );
nand ( n382972 , n382966 , n382971 );
buf ( n382973 , n382972 );
buf ( n382974 , n382973 );
not ( n62358 , n382974 );
buf ( n382976 , n44591 );
not ( n62360 , n382976 );
or ( n382978 , n62358 , n62360 );
buf ( n382979 , n60015 );
buf ( n382980 , n41834 );
nand ( n62364 , n382979 , n382980 );
buf ( n382982 , n62364 );
buf ( n382983 , n382982 );
nand ( n382984 , n382978 , n382983 );
buf ( n382985 , n382984 );
buf ( n382986 , n382985 );
and ( n62370 , n382961 , n382986 );
and ( n62371 , n382486 , n382960 );
or ( n382989 , n62370 , n62371 );
buf ( n382990 , n382989 );
buf ( n382991 , n382990 );
not ( n62375 , n382991 );
buf ( n382993 , n355579 );
not ( n382994 , n382993 );
buf ( n382995 , n360046 );
not ( n62379 , n382995 );
or ( n62380 , n382994 , n62379 );
buf ( n382998 , n378098 );
nand ( n382999 , n62380 , n382998 );
buf ( n383000 , n382999 );
buf ( n383001 , n383000 );
buf ( n383002 , n365528 );
buf ( n383003 , n365367 );
buf ( n383004 , n39937 );
nand ( n383005 , n383003 , n383004 );
buf ( n383006 , n383005 );
buf ( n383007 , n383006 );
and ( n62391 , n383001 , n383002 , n383007 );
buf ( n383009 , n62391 );
not ( n62393 , n383009 );
buf ( n383011 , n380497 );
buf ( n383012 , n351762 );
and ( n383013 , n383011 , n383012 );
not ( n383014 , n383011 );
buf ( n383015 , n48496 );
and ( n62399 , n383014 , n383015 );
nor ( n383017 , n383013 , n62399 );
buf ( n383018 , n383017 );
buf ( n383019 , n383018 );
not ( n383020 , n383019 );
buf ( n62404 , n44913 );
not ( n62405 , n62404 );
and ( n62406 , n383020 , n62405 );
buf ( n383024 , n380503 );
buf ( n383025 , n44915 );
and ( n62409 , n383024 , n383025 );
nor ( n62410 , n62406 , n62409 );
buf ( n383028 , n62410 );
nand ( n62412 , n62393 , n383028 );
not ( n62413 , n62412 );
buf ( n383031 , n377143 );
not ( n383032 , n383031 );
buf ( n383033 , n367600 );
not ( n62417 , n383033 );
or ( n383035 , n383032 , n62417 );
buf ( n383036 , n365569 );
buf ( n383037 , n377146 );
nand ( n383038 , n383036 , n383037 );
buf ( n383039 , n383038 );
buf ( n383040 , n383039 );
nand ( n62424 , n383035 , n383040 );
buf ( n383042 , n62424 );
buf ( n383043 , n383042 );
not ( n383044 , n383043 );
buf ( n383045 , n372247 );
not ( n62429 , n383045 );
or ( n383047 , n383044 , n62429 );
buf ( n383048 , n40923 );
buf ( n383049 , n381903 );
nand ( n383050 , n383048 , n383049 );
buf ( n383051 , n383050 );
buf ( n383052 , n383051 );
nand ( n383053 , n383047 , n383052 );
buf ( n383054 , n383053 );
not ( n383055 , n383054 );
or ( n383056 , n62413 , n383055 );
buf ( n383057 , n383028 );
not ( n383058 , n383057 );
buf ( n383059 , n383009 );
nand ( n383060 , n383058 , n383059 );
buf ( n383061 , n383060 );
nand ( n383062 , n383056 , n383061 );
buf ( n383063 , n383062 );
not ( n383064 , n383063 );
buf ( n383065 , n383064 );
buf ( n383066 , n383065 );
nand ( n383067 , n62375 , n383066 );
buf ( n383068 , n383067 );
buf ( n383069 , n383068 );
xor ( n383070 , n380968 , n380515 );
xnor ( n383071 , n383070 , n380541 );
buf ( n383072 , n383071 );
and ( n383073 , n383069 , n383072 );
buf ( n383074 , n382990 );
not ( n62456 , n383074 );
buf ( n383076 , n383065 );
nor ( n383077 , n62456 , n383076 );
buf ( n383078 , n383077 );
buf ( n383079 , n383078 );
nor ( n62461 , n383073 , n383079 );
buf ( n383081 , n62461 );
buf ( n383082 , n383081 );
not ( n383083 , n383082 );
buf ( n383084 , n383083 );
not ( n62466 , n383084 );
buf ( n383086 , n359902 );
not ( n62468 , n383086 );
buf ( n383088 , n365528 );
not ( n62470 , n383088 );
or ( n62471 , n62468 , n62470 );
buf ( n383091 , n359944 );
nand ( n62473 , n62471 , n383091 );
buf ( n383093 , n62473 );
buf ( n383094 , n383093 );
not ( n62476 , n383094 );
buf ( n383096 , n359890 );
not ( n62478 , n383096 );
buf ( n383098 , n365945 );
not ( n62480 , n383098 );
or ( n62481 , n62478 , n62480 );
buf ( n383101 , n378098 );
nand ( n62483 , n62481 , n383101 );
buf ( n383103 , n62483 );
buf ( n383104 , n383103 );
nand ( n62486 , n62476 , n383104 );
buf ( n383106 , n62486 );
not ( n62488 , n383106 );
buf ( n383108 , n382131 );
not ( n62490 , n383108 );
buf ( n383110 , n368290 );
not ( n62492 , n383110 );
or ( n62493 , n62490 , n62492 );
buf ( n383113 , n365954 );
buf ( n383114 , n379694 );
nand ( n383115 , n383113 , n383114 );
buf ( n383116 , n383115 );
buf ( n383117 , n383116 );
nand ( n383118 , n62493 , n383117 );
buf ( n383119 , n383118 );
buf ( n383120 , n383119 );
not ( n383121 , n383120 );
buf ( n383122 , n383121 );
xor ( n383123 , n62488 , n383122 );
xor ( n383124 , n57617 , n378022 );
xnor ( n383125 , n383124 , n378055 );
xnor ( n383126 , n383123 , n383125 );
buf ( n383127 , n383126 );
not ( n383128 , n383127 );
buf ( n383129 , n383128 );
not ( n383130 , n383129 );
or ( n383131 , n62466 , n383130 );
not ( n383132 , n383081 );
not ( n383133 , n383126 );
or ( n383134 , n383132 , n383133 );
xor ( n383135 , n381283 , n381312 );
xor ( n383136 , n383135 , n381345 );
buf ( n383137 , n56970 );
not ( n383138 , n383137 );
buf ( n383139 , n44717 );
not ( n383140 , n383139 );
or ( n383141 , n383138 , n383140 );
buf ( n383142 , n45414 );
buf ( n383143 , n377389 );
nand ( n383144 , n383142 , n383143 );
buf ( n383145 , n383144 );
buf ( n383146 , n383145 );
nand ( n62505 , n383141 , n383146 );
buf ( n383148 , n62505 );
buf ( n383149 , n383148 );
not ( n62508 , n383149 );
buf ( n383151 , n364849 );
not ( n62510 , n383151 );
or ( n383153 , n62508 , n62510 );
buf ( n383154 , n367590 );
buf ( n383155 , n381186 );
nand ( n383156 , n383154 , n383155 );
buf ( n383157 , n383156 );
buf ( n383158 , n383157 );
nand ( n383159 , n383153 , n383158 );
buf ( n383160 , n383159 );
or ( n383161 , n383136 , n383160 );
buf ( n383162 , n365428 );
not ( n383163 , n383162 );
buf ( n383164 , n381286 );
not ( n62523 , n383164 );
or ( n383166 , n383163 , n62523 );
buf ( n383167 , n377683 );
not ( n62526 , n383167 );
buf ( n383169 , n365422 );
nand ( n62528 , n62526 , n383169 );
buf ( n383171 , n62528 );
buf ( n383172 , n383171 );
nand ( n62531 , n383166 , n383172 );
buf ( n383174 , n62531 );
buf ( n383175 , n383174 );
not ( n62534 , n383175 );
buf ( n383177 , n363428 );
not ( n383178 , n383177 );
or ( n62537 , n62534 , n383178 );
buf ( n383180 , n381299 );
buf ( n383181 , n57228 );
nand ( n62540 , n383180 , n383181 );
buf ( n383183 , n62540 );
buf ( n383184 , n383183 );
nand ( n62543 , n62537 , n383184 );
buf ( n383186 , n62543 );
buf ( n383187 , n383186 );
xor ( n62546 , n381216 , n381237 );
xor ( n383189 , n62546 , n381279 );
buf ( n383190 , n383189 );
buf ( n383191 , n383190 );
xor ( n383192 , n383187 , n383191 );
buf ( n383193 , n382507 );
buf ( n383194 , n56794 );
and ( n383195 , n383193 , n383194 );
buf ( n383196 , n22619 );
not ( n62555 , n383196 );
buf ( n383198 , n31194 );
not ( n383199 , n383198 );
or ( n62558 , n62555 , n383199 );
buf ( n383201 , n57233 );
buf ( n383202 , n380923 );
nand ( n62561 , n383201 , n383202 );
buf ( n383204 , n62561 );
buf ( n383205 , n383204 );
nand ( n62564 , n62558 , n383205 );
buf ( n383207 , n62564 );
buf ( n383208 , n383207 );
not ( n383209 , n383208 );
buf ( n383210 , n365722 );
nor ( n383211 , n383209 , n383210 );
buf ( n383212 , n383211 );
buf ( n383213 , n383212 );
nor ( n383214 , n383195 , n383213 );
buf ( n383215 , n383214 );
buf ( n383216 , n383215 );
not ( n62575 , n383216 );
buf ( n383218 , n62575 );
buf ( n383219 , n383218 );
buf ( n383220 , n45802 );
not ( n62579 , n383220 );
buf ( n383222 , n22707 );
not ( n62581 , n383222 );
or ( n383224 , n62579 , n62581 );
buf ( n383225 , n342654 );
buf ( n383226 , n60751 );
nand ( n62585 , n383225 , n383226 );
buf ( n383228 , n62585 );
buf ( n383229 , n383228 );
nand ( n383230 , n383224 , n383229 );
buf ( n383231 , n383230 );
buf ( n62590 , n383231 );
not ( n62591 , n62590 );
buf ( n62592 , n366399 );
not ( n62593 , n62592 );
or ( n62594 , n62591 , n62593 );
buf ( n62595 , n381250 );
buf ( n383238 , n377171 );
nand ( n62597 , n62595 , n383238 );
buf ( n62598 , n62597 );
buf ( n383241 , n62598 );
nand ( n62600 , n62594 , n383241 );
buf ( n62601 , n62600 );
buf ( n383244 , n62601 );
or ( n62603 , n383219 , n383244 );
buf ( n383246 , n365108 );
not ( n383247 , n383246 );
buf ( n383248 , n62349 );
not ( n383249 , n383248 );
or ( n62608 , n383247 , n383249 );
not ( n383251 , n62340 );
not ( n62610 , n375886 );
or ( n383253 , n383251 , n62610 );
buf ( n383254 , n32202 );
buf ( n383255 , n62345 );
nand ( n383256 , n383254 , n383255 );
buf ( n383257 , n383256 );
nand ( n383258 , n383253 , n383257 );
buf ( n62617 , n383258 );
buf ( n383260 , n365024 );
nand ( n383261 , n62617 , n383260 );
buf ( n383262 , n383261 );
buf ( n62621 , n383262 );
nand ( n383264 , n62608 , n62621 );
buf ( n383265 , n383264 );
buf ( n383266 , n383265 );
nand ( n383267 , n62603 , n383266 );
buf ( n383268 , n383267 );
buf ( n383269 , n383268 );
buf ( n383270 , n62601 );
buf ( n383271 , n383218 );
nand ( n383272 , n383270 , n383271 );
buf ( n383273 , n383272 );
buf ( n383274 , n383273 );
nand ( n383275 , n383269 , n383274 );
buf ( n383276 , n383275 );
buf ( n383277 , n383276 );
and ( n62636 , n383192 , n383277 );
and ( n62637 , n383187 , n383191 );
or ( n62638 , n62636 , n62637 );
buf ( n383281 , n62638 );
nand ( n62640 , n383161 , n383281 );
buf ( n383283 , n383160 );
buf ( n383284 , n383136 );
nand ( n62643 , n383283 , n383284 );
buf ( n383286 , n62643 );
nand ( n62645 , n62640 , n383286 );
not ( n383288 , n62645 );
buf ( n383289 , n369769 );
not ( n383290 , n383289 );
buf ( n383291 , n41615 );
not ( n383292 , n383291 );
or ( n62651 , n383290 , n383292 );
buf ( n383294 , n41946 );
buf ( n383295 , n369766 );
nand ( n383296 , n383294 , n383295 );
buf ( n383297 , n383296 );
buf ( n383298 , n383297 );
nand ( n383299 , n62651 , n383298 );
buf ( n383300 , n383299 );
and ( n62659 , n383300 , n369804 );
and ( n383302 , n381789 , n49609 );
nor ( n62661 , n62659 , n383302 );
and ( n383304 , n382203 , n379263 );
not ( n62663 , n379274 );
buf ( n383306 , n360885 );
not ( n62665 , n383306 );
buf ( n383308 , n62665 );
not ( n383309 , n383308 );
or ( n62668 , n62663 , n383309 );
nand ( n383311 , n379271 , n360885 );
nand ( n383312 , n62668 , n383311 );
and ( n62671 , n383312 , n379293 );
nor ( n62672 , n383304 , n62671 );
nand ( n383315 , n62661 , n62672 );
not ( n62674 , n383315 );
or ( n62675 , n383288 , n62674 );
buf ( n383318 , n62661 );
not ( n383319 , n383318 );
buf ( n383320 , n383319 );
buf ( n383321 , n383320 );
buf ( n62680 , n62672 );
not ( n62681 , n62680 );
buf ( n383324 , n62681 );
buf ( n383325 , n383324 );
nand ( n383326 , n383321 , n383325 );
buf ( n383327 , n383326 );
nand ( n62686 , n62675 , n383327 );
nand ( n383329 , n383134 , n62686 );
nand ( n383330 , n383131 , n383329 );
buf ( n62689 , n383330 );
xor ( n62690 , n61056 , n61063 );
xor ( n383333 , n62690 , n381638 );
buf ( n383334 , n383333 );
buf ( n383335 , n383334 );
xor ( n62694 , n379194 , n379237 );
xor ( n383337 , n62694 , n379108 );
buf ( n62696 , n383337 );
xor ( n62697 , n383335 , n62696 );
buf ( n383340 , n382276 );
not ( n383341 , n383340 );
buf ( n383342 , n61693 );
not ( n383343 , n383342 );
or ( n383344 , n383341 , n383343 );
buf ( n383345 , n382277 );
not ( n383346 , n383345 );
buf ( n383347 , n61689 );
not ( n62706 , n383347 );
or ( n62707 , n383346 , n62706 );
buf ( n383350 , n61666 );
nand ( n383351 , n62707 , n383350 );
buf ( n383352 , n383351 );
buf ( n383353 , n383352 );
nand ( n383354 , n383344 , n383353 );
buf ( n383355 , n383354 );
buf ( n383356 , n383355 );
xor ( n62715 , n62697 , n383356 );
buf ( n383358 , n62715 );
buf ( n383359 , n383358 );
xor ( n62718 , n62689 , n383359 );
and ( n62719 , n383106 , n383122 );
or ( n62720 , n62719 , n383125 );
buf ( n383363 , n383119 );
buf ( n383364 , n62488 );
nand ( n62723 , n383363 , n383364 );
buf ( n383366 , n62723 );
nand ( n62725 , n62720 , n383366 );
buf ( n383368 , n62725 );
xor ( n62727 , n377901 , n377942 );
xor ( n62728 , n62727 , n377979 );
buf ( n62729 , n62728 );
buf ( n383372 , n62729 );
xor ( n62731 , n383368 , n383372 );
buf ( n383374 , n379650 );
buf ( n383375 , n379676 );
xor ( n62734 , n383374 , n383375 );
buf ( n383377 , n379706 );
xnor ( n62736 , n62734 , n383377 );
buf ( n383379 , n62736 );
buf ( n383380 , n383379 );
xnor ( n62739 , n62731 , n383380 );
buf ( n383382 , n62739 );
buf ( n383383 , n383382 );
xor ( n383384 , n62718 , n383383 );
buf ( n383385 , n383384 );
xor ( n383386 , n382461 , n383385 );
buf ( n383387 , n383126 );
buf ( n383388 , n62686 );
xor ( n62747 , n383387 , n383388 );
buf ( n383390 , n383081 );
xor ( n383391 , n62747 , n383390 );
buf ( n383392 , n383391 );
not ( n62751 , n383392 );
xor ( n383394 , n382187 , n382209 );
xor ( n383395 , n383394 , n382222 );
buf ( n383396 , n383395 );
not ( n62755 , n383396 );
or ( n383398 , n62751 , n62755 );
nor ( n383399 , n383396 , n383392 );
buf ( n383400 , n382990 );
buf ( n383401 , n383062 );
xor ( n62760 , n383400 , n383401 );
buf ( n383403 , n383071 );
xor ( n383404 , n62760 , n383403 );
buf ( n383405 , n383404 );
buf ( n383406 , n383054 );
not ( n383407 , n383406 );
buf ( n383408 , n383028 );
not ( n62767 , n383408 );
buf ( n383410 , n383009 );
not ( n383411 , n383410 );
and ( n383412 , n62767 , n383411 );
buf ( n383413 , n383028 );
buf ( n383414 , n383009 );
and ( n62773 , n383413 , n383414 );
nor ( n383416 , n383412 , n62773 );
buf ( n383417 , n383416 );
buf ( n383418 , n383417 );
not ( n62777 , n383418 );
or ( n62778 , n383407 , n62777 );
buf ( n383421 , n383417 );
buf ( n383422 , n383054 );
or ( n62781 , n383421 , n383422 );
nand ( n62782 , n62778 , n62781 );
buf ( n383425 , n62782 );
buf ( n383426 , n383425 );
buf ( n383427 , n377757 );
not ( n383428 , n383427 );
buf ( n383429 , n365626 );
not ( n62788 , n383429 );
or ( n62789 , n383428 , n62788 );
buf ( n383432 , n41892 );
buf ( n62791 , n378886 );
nand ( n62792 , n383432 , n62791 );
buf ( n62793 , n62792 );
buf ( n383436 , n62793 );
nand ( n62795 , n62789 , n383436 );
buf ( n383438 , n62795 );
buf ( n383439 , n383438 );
not ( n62798 , n383439 );
buf ( n383441 , n364797 );
not ( n383442 , n383441 );
or ( n62801 , n62798 , n383442 );
buf ( n383444 , n377782 );
not ( n383445 , n383444 );
buf ( n383446 , n365626 );
not ( n383447 , n383446 );
or ( n62806 , n383445 , n383447 );
buf ( n383449 , n45455 );
buf ( n383450 , n377779 );
nand ( n62809 , n383449 , n383450 );
buf ( n383452 , n62809 );
buf ( n383453 , n383452 );
nand ( n383454 , n62806 , n383453 );
buf ( n383455 , n383454 );
buf ( n383456 , n383455 );
buf ( n383457 , n371063 );
nand ( n383458 , n383456 , n383457 );
buf ( n383459 , n383458 );
buf ( n383460 , n383459 );
nand ( n62819 , n62801 , n383460 );
buf ( n383462 , n62819 );
buf ( n383463 , n383462 );
buf ( n383464 , n368608 );
not ( n62823 , n383464 );
buf ( n383466 , n380424 );
not ( n62825 , n383466 );
buf ( n383468 , n366078 );
not ( n383469 , n383468 );
or ( n383470 , n62825 , n383469 );
buf ( n383471 , n366077 );
buf ( n383472 , n368549 );
nand ( n383473 , n383471 , n383472 );
buf ( n383474 , n383473 );
buf ( n383475 , n383474 );
nand ( n62834 , n383470 , n383475 );
buf ( n62835 , n62834 );
buf ( n383478 , n62835 );
not ( n383479 , n383478 );
or ( n383480 , n62823 , n383479 );
buf ( n383481 , n368549 );
not ( n383482 , n383481 );
buf ( n383483 , n46126 );
not ( n62842 , n383483 );
or ( n62843 , n383482 , n62842 );
buf ( n383486 , n362534 );
buf ( n383487 , n380424 );
nand ( n383488 , n383486 , n383487 );
buf ( n383489 , n383488 );
buf ( n62848 , n383489 );
nand ( n383491 , n62843 , n62848 );
buf ( n383492 , n383491 );
buf ( n383493 , n383492 );
buf ( n383494 , n369444 );
nand ( n383495 , n383493 , n383494 );
buf ( n383496 , n383495 );
buf ( n383497 , n383496 );
nand ( n62856 , n383480 , n383497 );
buf ( n383499 , n62856 );
buf ( n383500 , n383499 );
xor ( n62859 , n383463 , n383500 );
buf ( n383502 , n365226 );
not ( n62861 , n383502 );
buf ( n383504 , n342881 );
not ( n62863 , n383504 );
buf ( n383506 , n45125 );
not ( n62865 , n383506 );
or ( n62866 , n62863 , n62865 );
buf ( n383509 , n352192 );
buf ( n383510 , n365202 );
nand ( n62869 , n383509 , n383510 );
buf ( n383512 , n62869 );
buf ( n383513 , n383512 );
nand ( n383514 , n62866 , n383513 );
buf ( n383515 , n383514 );
buf ( n383516 , n383515 );
not ( n383517 , n383516 );
or ( n62876 , n62861 , n383517 );
buf ( n383519 , n381868 );
buf ( n383520 , n45075 );
nand ( n383521 , n383519 , n383520 );
buf ( n383522 , n383521 );
buf ( n383523 , n383522 );
nand ( n383524 , n62876 , n383523 );
buf ( n383525 , n383524 );
not ( n62884 , n47466 );
buf ( n383527 , n365041 );
not ( n383528 , n383527 );
buf ( n383529 , n45152 );
not ( n383530 , n383529 );
or ( n62889 , n383528 , n383530 );
buf ( n383532 , n380497 );
buf ( n383533 , n30911 );
nand ( n62892 , n383532 , n383533 );
buf ( n383535 , n62892 );
buf ( n383536 , n383535 );
nand ( n383537 , n62889 , n383536 );
buf ( n383538 , n383537 );
not ( n62897 , n383538 );
or ( n383540 , n62884 , n62897 );
not ( n383541 , n383018 );
nand ( n62900 , n383541 , n44915 );
nand ( n62901 , n383540 , n62900 );
xor ( n383544 , n383525 , n62901 );
buf ( n383545 , n368665 );
not ( n383546 , n383545 );
buf ( n383547 , n342335 );
not ( n62906 , n383547 );
or ( n383549 , n383546 , n62906 );
buf ( n383550 , n342338 );
buf ( n383551 , n368662 );
nand ( n62910 , n383550 , n383551 );
buf ( n62911 , n62910 );
buf ( n383554 , n62911 );
nand ( n383555 , n383549 , n383554 );
buf ( n383556 , n383555 );
buf ( n383557 , n383556 );
not ( n383558 , n383557 );
buf ( n383559 , n42263 );
not ( n62918 , n383559 );
or ( n383561 , n383558 , n62918 );
buf ( n383562 , n60783 );
buf ( n383563 , n48490 );
nand ( n62922 , n383562 , n383563 );
buf ( n383565 , n62922 );
buf ( n383566 , n383565 );
nand ( n383567 , n383561 , n383566 );
buf ( n383568 , n383567 );
xor ( n383569 , n383544 , n383568 );
buf ( n383570 , n383569 );
and ( n62929 , n62859 , n383570 );
and ( n62930 , n383463 , n383500 );
or ( n383573 , n62929 , n62930 );
buf ( n383574 , n383573 );
buf ( n383575 , n383574 );
xor ( n62934 , n383426 , n383575 );
buf ( n383577 , n49609 );
not ( n383578 , n383577 );
buf ( n383579 , n369769 );
not ( n383580 , n383579 );
buf ( n383581 , n361664 );
not ( n383582 , n383581 );
or ( n383583 , n383580 , n383582 );
buf ( n383584 , n41528 );
buf ( n383585 , n369766 );
nand ( n62944 , n383584 , n383585 );
buf ( n383587 , n62944 );
buf ( n383588 , n383587 );
nand ( n62947 , n383583 , n383588 );
buf ( n383590 , n62947 );
buf ( n383591 , n383590 );
not ( n383592 , n383591 );
or ( n383593 , n383578 , n383592 );
buf ( n383594 , n369804 );
buf ( n383595 , n369769 );
not ( n383596 , n383595 );
buf ( n383597 , n51996 );
not ( n62956 , n383597 );
or ( n383599 , n383596 , n62956 );
buf ( n383600 , n361716 );
buf ( n383601 , n369766 );
nand ( n62960 , n383600 , n383601 );
buf ( n383603 , n62960 );
buf ( n383604 , n383603 );
nand ( n62963 , n383599 , n383604 );
buf ( n383606 , n62963 );
buf ( n383607 , n383606 );
nand ( n62966 , n383594 , n383607 );
buf ( n383609 , n62966 );
buf ( n383610 , n383609 );
nand ( n62969 , n383593 , n383610 );
buf ( n383612 , n62969 );
buf ( n383613 , n383612 );
not ( n383614 , n383613 );
buf ( n383615 , n383614 );
buf ( n383616 , n383615 );
not ( n383617 , n383616 );
buf ( n383618 , n377094 );
not ( n62977 , n383618 );
buf ( n383620 , n359297 );
not ( n62979 , n383620 );
or ( n383622 , n62977 , n62979 );
buf ( n383623 , n365367 );
buf ( n383624 , n56687 );
nand ( n62983 , n383623 , n383624 );
buf ( n383626 , n62983 );
buf ( n383627 , n383626 );
nand ( n383628 , n383622 , n383627 );
buf ( n383629 , n383628 );
buf ( n383630 , n383629 );
not ( n62989 , n383630 );
buf ( n383632 , n369260 );
not ( n383633 , n383632 );
or ( n62992 , n62989 , n383633 );
buf ( n383635 , n46582 );
not ( n383636 , n51966 );
not ( n62995 , n377071 );
or ( n62996 , n383636 , n62995 );
not ( n383639 , n365353 );
nand ( n383640 , n383639 , n377068 );
nand ( n62999 , n62996 , n383640 );
buf ( n383642 , n62999 );
nand ( n63001 , n383635 , n383642 );
buf ( n383644 , n63001 );
buf ( n383645 , n383644 );
nand ( n383646 , n62992 , n383645 );
buf ( n383647 , n383646 );
buf ( n383648 , n383647 );
not ( n383649 , n383648 );
buf ( n383650 , n383649 );
buf ( n383651 , n383650 );
not ( n383652 , n383651 );
or ( n383653 , n383617 , n383652 );
buf ( n383654 , n57280 );
not ( n383655 , n383654 );
buf ( n383656 , n44661 );
not ( n63015 , n383656 );
or ( n383658 , n383655 , n63015 );
buf ( n383659 , n351107 );
buf ( n383660 , n377728 );
nand ( n383661 , n383659 , n383660 );
buf ( n383662 , n383661 );
buf ( n383663 , n383662 );
nand ( n383664 , n383658 , n383663 );
buf ( n383665 , n383664 );
buf ( n383666 , n383665 );
buf ( n383667 , n365152 );
and ( n383668 , n383666 , n383667 );
buf ( n383669 , n57280 );
not ( n63028 , n383669 );
buf ( n383671 , n351318 );
not ( n383672 , n383671 );
or ( n63031 , n63028 , n383672 );
buf ( n383674 , n364808 );
buf ( n383675 , n377728 );
nand ( n63034 , n383674 , n383675 );
buf ( n383677 , n63034 );
buf ( n383678 , n383677 );
nand ( n63037 , n63031 , n383678 );
buf ( n383680 , n63037 );
buf ( n383681 , n383680 );
not ( n383682 , n383681 );
not ( n383683 , n365186 );
buf ( n383684 , n383683 );
nor ( n383685 , n383682 , n383684 );
buf ( n383686 , n383685 );
buf ( n383687 , n383686 );
nor ( n63046 , n383668 , n383687 );
buf ( n63047 , n63046 );
buf ( n383690 , n63047 );
not ( n63049 , n383690 );
buf ( n383692 , n365052 );
buf ( n383693 , n351367 );
and ( n383694 , n383692 , n383693 );
not ( n383695 , n383692 );
buf ( n383696 , n366131 );
and ( n63055 , n383695 , n383696 );
nor ( n63056 , n383694 , n63055 );
buf ( n383699 , n63056 );
not ( n383700 , n383699 );
not ( n63059 , n44913 );
and ( n63060 , n383700 , n63059 );
and ( n63061 , n383538 , n44915 );
nor ( n383704 , n63060 , n63061 );
buf ( n383705 , n383704 );
not ( n63064 , n383705 );
or ( n63065 , n63049 , n63064 );
buf ( n383708 , n383215 );
buf ( n383709 , n383265 );
xor ( n63068 , n383708 , n383709 );
buf ( n383711 , n62601 );
xnor ( n383712 , n63068 , n383711 );
buf ( n383713 , n383712 );
buf ( n383714 , n383713 );
nand ( n63073 , n63065 , n383714 );
buf ( n383716 , n63073 );
buf ( n383717 , n383716 );
buf ( n383718 , n63047 );
not ( n63077 , n383718 );
buf ( n383720 , n383704 );
not ( n63079 , n383720 );
buf ( n383722 , n63079 );
buf ( n383723 , n383722 );
nand ( n63082 , n63077 , n383723 );
buf ( n383725 , n63082 );
buf ( n383726 , n383725 );
nand ( n63085 , n383717 , n383726 );
buf ( n383728 , n63085 );
buf ( n383729 , n383728 );
nand ( n63088 , n383653 , n383729 );
buf ( n383731 , n63088 );
buf ( n383732 , n383731 );
buf ( n383733 , n383647 );
buf ( n383734 , n383612 );
nand ( n383735 , n383733 , n383734 );
buf ( n383736 , n383735 );
buf ( n383737 , n383736 );
nand ( n383738 , n383732 , n383737 );
buf ( n383739 , n383738 );
buf ( n383740 , n383739 );
and ( n383741 , n62934 , n383740 );
and ( n383742 , n383426 , n383575 );
or ( n63101 , n383741 , n383742 );
buf ( n383744 , n63101 );
xor ( n63103 , n383405 , n383744 );
not ( n383746 , n383320 );
not ( n63105 , n62672 );
or ( n63106 , n383746 , n63105 );
nand ( n63107 , n62661 , n383324 );
nand ( n383750 , n63106 , n63107 );
and ( n383751 , n383750 , n62645 );
not ( n63110 , n383750 );
not ( n383753 , n62645 );
and ( n383754 , n63110 , n383753 );
nor ( n383755 , n383751 , n383754 );
and ( n383756 , n63103 , n383755 );
and ( n63115 , n383405 , n383744 );
or ( n383758 , n383756 , n63115 );
not ( n383759 , n383758 );
or ( n63118 , n383399 , n383759 );
nand ( n383761 , n383398 , n63118 );
and ( n383762 , n383386 , n383761 );
and ( n63121 , n382461 , n383385 );
or ( n383764 , n383762 , n63121 );
nand ( n383765 , n382414 , n383764 );
nand ( n383766 , n382411 , n383765 );
buf ( n383767 , n383766 );
not ( n383768 , n383767 );
or ( n63127 , n382348 , n383768 );
or ( n383770 , n383766 , n382346 );
xor ( n63129 , n62689 , n383359 );
and ( n63130 , n63129 , n383383 );
and ( n383773 , n62689 , n383359 );
or ( n383774 , n63130 , n383773 );
buf ( n383775 , n383774 );
buf ( n383776 , n383775 );
buf ( n383777 , n383776 );
buf ( n383778 , n383777 );
buf ( n383779 , n383778 );
not ( n383780 , n383779 );
buf ( n383781 , n381480 );
not ( n63140 , n383781 );
buf ( n383783 , n381049 );
not ( n383784 , n383783 );
or ( n63143 , n63140 , n383784 );
buf ( n383786 , n381046 );
buf ( n383787 , n381038 );
nand ( n63146 , n383786 , n383787 );
buf ( n63147 , n63146 );
buf ( n383790 , n63147 );
nand ( n63149 , n63143 , n383790 );
buf ( n383792 , n63149 );
buf ( n383793 , n383792 );
buf ( n383794 , n60911 );
not ( n383795 , n383794 );
buf ( n383796 , n383795 );
buf ( n383797 , n383796 );
and ( n63156 , n383793 , n383797 );
not ( n63157 , n383793 );
buf ( n63158 , n60911 );
and ( n383801 , n63157 , n63158 );
nor ( n63160 , n63156 , n383801 );
buf ( n63161 , n63160 );
buf ( n383804 , n63161 );
not ( n63163 , n383804 );
buf ( n63164 , n63163 );
buf ( n383807 , n63164 );
not ( n63166 , n383807 );
or ( n383809 , n383780 , n63166 );
buf ( n383810 , n383778 );
not ( n383811 , n383810 );
buf ( n383812 , n383811 );
buf ( n383813 , n383812 );
not ( n383814 , n383813 );
buf ( n383815 , n63161 );
not ( n63174 , n383815 );
or ( n383817 , n383814 , n63174 );
xor ( n63176 , n380352 , n380414 );
xor ( n383819 , n63176 , n380984 );
buf ( n383820 , n383819 );
not ( n383821 , n383820 );
and ( n63180 , n380979 , n380446 );
not ( n63181 , n380979 );
not ( n383824 , n380446 );
and ( n383825 , n63181 , n383824 );
nor ( n63184 , n63180 , n383825 );
buf ( n383827 , n59971 );
not ( n383828 , n383827 );
buf ( n383829 , n383828 );
and ( n63188 , n63184 , n383829 );
not ( n63189 , n63184 );
and ( n383832 , n63189 , n59971 );
nor ( n383833 , n63188 , n383832 );
buf ( n383834 , n383833 );
xor ( n383835 , n382181 , n382162 );
buf ( n383836 , n382138 );
and ( n63195 , n383835 , n383836 );
not ( n383838 , n383835 );
and ( n383839 , n383838 , n382166 );
nor ( n63198 , n63195 , n383839 );
buf ( n383841 , n63198 );
buf ( n63200 , n377580 );
not ( n63201 , n63200 );
buf ( n63202 , n382248 );
not ( n63203 , n63202 );
or ( n63204 , n63201 , n63203 );
buf ( n383847 , n377585 );
not ( n383848 , n383847 );
buf ( n383849 , n45718 );
not ( n383850 , n383849 );
or ( n383851 , n383848 , n383850 );
buf ( n383852 , n362133 );
buf ( n383853 , n377592 );
nand ( n383854 , n383852 , n383853 );
buf ( n383855 , n383854 );
buf ( n383856 , n383855 );
nand ( n63215 , n383851 , n383856 );
buf ( n383858 , n63215 );
buf ( n63217 , n383858 );
buf ( n63218 , n57530 );
nand ( n63219 , n63217 , n63218 );
buf ( n63220 , n63219 );
buf ( n63221 , n63220 );
nand ( n63222 , n63204 , n63221 );
buf ( n63223 , n63222 );
buf ( n383866 , n63223 );
not ( n63225 , n383866 );
buf ( n383868 , n63225 );
buf ( n383869 , n383868 );
nand ( n383870 , n383841 , n383869 );
buf ( n383871 , n383870 );
buf ( n383872 , n383871 );
not ( n383873 , n381801 );
and ( n383874 , n381829 , n383873 );
not ( n63233 , n381829 );
and ( n383876 , n63233 , n381801 );
nor ( n383877 , n383874 , n383876 );
buf ( n383878 , n381885 );
not ( n383879 , n383878 );
buf ( n383880 , n381878 );
not ( n63239 , n383880 );
or ( n383882 , n383879 , n63239 );
buf ( n383883 , n381875 );
buf ( n383884 , n61286 );
nand ( n383885 , n383883 , n383884 );
buf ( n383886 , n383885 );
buf ( n383887 , n383886 );
nand ( n383888 , n383882 , n383887 );
buf ( n383889 , n383888 );
xor ( n63248 , n383877 , n383889 );
buf ( n383891 , n63248 );
not ( n383892 , n383891 );
buf ( n383893 , n383892 );
not ( n63252 , n383893 );
xor ( n383895 , n382486 , n382960 );
xor ( n383896 , n383895 , n382986 );
buf ( n383897 , n383896 );
not ( n383898 , n383897 );
or ( n63257 , n63252 , n383898 );
or ( n383900 , n383893 , n383897 );
buf ( n383901 , n365187 );
not ( n383902 , n383901 );
buf ( n383903 , n383665 );
not ( n63262 , n383903 );
or ( n383905 , n383902 , n63262 );
buf ( n383906 , n382478 );
buf ( n383907 , n365152 );
nand ( n383908 , n383906 , n383907 );
buf ( n383909 , n383908 );
buf ( n383910 , n383909 );
nand ( n383911 , n383905 , n383910 );
buf ( n383912 , n383911 );
not ( n63271 , n383912 );
buf ( n383914 , n369374 );
not ( n383915 , n383914 );
buf ( n383916 , n367248 );
not ( n63275 , n383916 );
or ( n383918 , n383915 , n63275 );
buf ( n383919 , n364744 );
buf ( n383920 , n49178 );
nand ( n383921 , n383919 , n383920 );
buf ( n383922 , n383921 );
buf ( n383923 , n383922 );
nand ( n383924 , n383918 , n383923 );
buf ( n383925 , n383924 );
buf ( n383926 , n383925 );
not ( n383927 , n383926 );
buf ( n383928 , n44591 );
not ( n63287 , n383928 );
or ( n383930 , n383927 , n63287 );
not ( n383931 , n49692 );
nand ( n63290 , n383931 , n382973 );
buf ( n383933 , n63290 );
nand ( n63292 , n383930 , n383933 );
buf ( n63293 , n63292 );
not ( n383936 , n63293 );
or ( n63295 , n63271 , n383936 );
buf ( n383938 , n383912 );
not ( n63297 , n383938 );
buf ( n383940 , n63297 );
buf ( n383941 , n383940 );
not ( n63300 , n383941 );
buf ( n383943 , n63293 );
not ( n383944 , n383943 );
buf ( n383945 , n383944 );
buf ( n383946 , n383945 );
not ( n63305 , n383946 );
or ( n63306 , n63300 , n63305 );
xor ( n383949 , n380858 , n380866 );
xor ( n383950 , n383949 , n380870 );
xor ( n63309 , n382585 , n62296 );
xor ( n63310 , n383950 , n63309 );
buf ( n383953 , n63310 );
buf ( n383954 , n56794 );
not ( n63313 , n383954 );
buf ( n383956 , n383207 );
not ( n383957 , n383956 );
or ( n63316 , n63313 , n383957 );
buf ( n383959 , n365725 );
buf ( n383960 , n22619 );
not ( n383961 , n383960 );
buf ( n383962 , n378543 );
not ( n63321 , n383962 );
or ( n383964 , n383961 , n63321 );
buf ( n383965 , n351195 );
buf ( n383966 , n380923 );
nand ( n383967 , n383965 , n383966 );
buf ( n383968 , n383967 );
buf ( n383969 , n383968 );
nand ( n383970 , n383964 , n383969 );
buf ( n383971 , n383970 );
buf ( n383972 , n383971 );
nand ( n383973 , n383959 , n383972 );
buf ( n383974 , n383973 );
buf ( n383975 , n383974 );
nand ( n383976 , n63316 , n383975 );
buf ( n383977 , n383976 );
buf ( n63336 , n383977 );
xor ( n63337 , n383953 , n63336 );
not ( n383980 , n380901 );
buf ( n383981 , n366659 );
not ( n63340 , n383981 );
buf ( n383983 , n364901 );
not ( n383984 , n383983 );
or ( n63343 , n63340 , n383984 );
buf ( n63344 , n32234 );
not ( n63345 , n63344 );
buf ( n383988 , n63345 );
not ( n383989 , n383988 );
buf ( n383990 , n342617 );
nand ( n63349 , n383989 , n383990 );
buf ( n383992 , n63349 );
buf ( n383993 , n383992 );
nand ( n383994 , n63343 , n383993 );
buf ( n383995 , n383994 );
not ( n63354 , n383995 );
or ( n63355 , n383980 , n63354 );
buf ( n383998 , n382914 );
buf ( n383999 , n375920 );
nand ( n63358 , n383998 , n383999 );
buf ( n384001 , n63358 );
nand ( n63360 , n63355 , n384001 );
buf ( n384003 , n63360 );
and ( n384004 , n63337 , n384003 );
and ( n63363 , n383953 , n63336 );
or ( n384006 , n384004 , n63363 );
buf ( n384007 , n384006 );
not ( n63366 , n384007 );
not ( n63367 , n63366 );
xor ( n63368 , n382518 , n62302 );
xnor ( n384011 , n63368 , n382926 );
not ( n63370 , n384011 );
not ( n384013 , n63370 );
and ( n384014 , n63367 , n384013 );
xor ( n63373 , n382522 , n382578 );
xor ( n63374 , n63373 , n382582 );
xor ( n384017 , n382765 , n62291 );
xor ( n63376 , n63374 , n384017 );
buf ( n384019 , n63376 );
buf ( n384020 , n382809 );
not ( n63379 , n384020 );
buf ( n384022 , n382784 );
not ( n63381 , n384022 );
or ( n63382 , n63379 , n63381 );
buf ( n384025 , n382812 );
nand ( n384026 , n63382 , n384025 );
buf ( n384027 , n384026 );
buf ( n384028 , n384027 );
buf ( n384029 , n380680 );
buf ( n384030 , n57800 );
and ( n63389 , n384029 , n384030 );
buf ( n384032 , n60171 );
buf ( n384033 , n376903 );
and ( n384034 , n384032 , n384033 );
nor ( n63393 , n63389 , n384034 );
buf ( n384036 , n63393 );
buf ( n384037 , n384036 );
buf ( n384038 , n378341 );
or ( n63397 , n384037 , n384038 );
buf ( n384040 , n382709 );
buf ( n384041 , n378424 );
or ( n63400 , n384040 , n384041 );
nand ( n63401 , n63397 , n63400 );
buf ( n384044 , n63401 );
buf ( n63403 , n384044 );
xor ( n63404 , n384028 , n63403 );
and ( n384047 , n62190 , n56312 );
xor ( n63406 , n384047 , n56309 );
buf ( n384049 , n63406 );
buf ( n384050 , n376990 );
and ( n63409 , n384049 , n384050 );
buf ( n63410 , n63406 );
not ( n384053 , n63410 );
buf ( n384054 , n384053 );
buf ( n384055 , n384054 );
buf ( n384056 , n376997 );
and ( n63415 , n384055 , n384056 );
buf ( n384058 , n377003 );
nor ( n384059 , n63409 , n63415 , n384058 );
buf ( n384060 , n384059 );
buf ( n384061 , n384060 );
and ( n63420 , n62023 , n56379 );
not ( n384063 , n63420 );
and ( n63422 , n380719 , n384063 );
not ( n384065 , n380719 );
and ( n384066 , n384065 , n63420 );
or ( n63425 , n63422 , n384066 );
buf ( n384068 , n63425 );
buf ( n384069 , n62026 );
xor ( n384070 , n384068 , n384069 );
buf ( n384071 , n384070 );
buf ( n384072 , n384071 );
buf ( n384073 , n63425 );
nand ( n384074 , n56373 , n56357 );
nand ( n384075 , n376792 , n376769 );
xnor ( n63434 , n384074 , n384075 );
buf ( n384077 , n63434 );
xor ( n63436 , n384073 , n384077 );
buf ( n384079 , n63436 );
buf ( n384080 , n384079 );
not ( n63439 , n384080 );
buf ( n384082 , n63439 );
buf ( n384083 , n384082 );
and ( n63442 , n384072 , n384083 );
buf ( n384085 , n63442 );
buf ( n384086 , n384085 );
buf ( n384087 , n62026 );
buf ( n63446 , n384087 );
buf ( n384089 , n63446 );
buf ( n384090 , n384089 );
nand ( n384091 , n384086 , n384090 );
buf ( n384092 , n384091 );
buf ( n384093 , n384092 );
buf ( n384094 , n384079 );
buf ( n384095 , n384089 );
nand ( n384096 , n384094 , n384095 );
buf ( n384097 , n384096 );
buf ( n384098 , n384097 );
and ( n63457 , n384093 , n384098 );
buf ( n384100 , n63457 );
buf ( n63459 , n384100 );
xor ( n63460 , n384061 , n63459 );
buf ( n384103 , n382795 );
buf ( n384104 , n376866 );
and ( n63463 , n384103 , n384104 );
buf ( n384106 , n382803 );
buf ( n384107 , n382743 );
and ( n63466 , n384106 , n384107 );
nor ( n384109 , n63463 , n63466 );
buf ( n384110 , n384109 );
buf ( n384111 , n384110 );
buf ( n384112 , n376924 );
or ( n63471 , n384111 , n384112 );
buf ( n384114 , n382776 );
buf ( n384115 , n56517 );
or ( n384116 , n384114 , n384115 );
nand ( n63475 , n63471 , n384116 );
buf ( n63476 , n63475 );
buf ( n384119 , n63476 );
and ( n63478 , n63460 , n384119 );
and ( n384121 , n384061 , n63459 );
or ( n63480 , n63478 , n384121 );
buf ( n384123 , n63480 );
buf ( n384124 , n384123 );
and ( n63483 , n63404 , n384124 );
and ( n384126 , n384028 , n63403 );
or ( n63485 , n63483 , n384126 );
buf ( n384128 , n63485 );
xor ( n63487 , n382718 , n382735 );
xor ( n384130 , n63487 , n382756 );
buf ( n384131 , n384130 );
xor ( n63490 , n384128 , n384131 );
xor ( n384133 , n382602 , n382670 );
xor ( n384134 , n384133 , n382687 );
xor ( n63493 , n382812 , n62276 );
xor ( n384136 , n384134 , n63493 );
and ( n63495 , n63490 , n384136 );
and ( n63496 , n384128 , n384131 );
or ( n63497 , n63495 , n63496 );
xor ( n63498 , n382879 , n382882 );
xor ( n384141 , n63498 , n382886 );
and ( n63500 , n63497 , n384141 );
buf ( n384143 , n376971 );
buf ( n384144 , n382835 );
and ( n384145 , n384143 , n384144 );
buf ( n384146 , n376993 );
buf ( n384147 , n62243 );
and ( n63506 , n384146 , n384147 );
nor ( n63507 , n384145 , n63506 );
buf ( n384150 , n63507 );
buf ( n384151 , n384150 );
buf ( n384152 , n382849 );
or ( n384153 , n384151 , n384152 );
buf ( n384154 , n382845 );
buf ( n384155 , n382663 );
not ( n63514 , n384155 );
buf ( n384157 , n63514 );
buf ( n384158 , n384157 );
or ( n384159 , n384154 , n384158 );
nand ( n63518 , n384153 , n384159 );
buf ( n63519 , n63518 );
buf ( n384162 , n63519 );
buf ( n384163 , n63406 );
buf ( n384164 , n376866 );
and ( n63523 , n384163 , n384164 );
buf ( n384166 , n384054 );
buf ( n384167 , n382743 );
and ( n384168 , n384166 , n384167 );
nor ( n63527 , n63523 , n384168 );
buf ( n384170 , n63527 );
buf ( n384171 , n384170 );
buf ( n384172 , n376924 );
or ( n63531 , n384171 , n384172 );
buf ( n384174 , n384110 );
buf ( n384175 , n56517 );
or ( n63534 , n384174 , n384175 );
nand ( n63535 , n63531 , n63534 );
buf ( n384178 , n63535 );
buf ( n384179 , n384178 );
not ( n63538 , n376316 );
not ( n384181 , n63538 );
not ( n384182 , n376699 );
or ( n63541 , n384181 , n384182 );
not ( n384184 , n56303 );
nand ( n63543 , n63541 , n384184 );
nand ( n384186 , n56306 , n376274 );
not ( n384187 , n384186 );
and ( n384188 , n63543 , n384187 );
not ( n63547 , n63543 );
and ( n384190 , n63547 , n384186 );
nor ( n63549 , n384188 , n384190 );
buf ( n384192 , n63549 );
buf ( n384193 , n376990 );
and ( n63552 , n384192 , n384193 );
and ( n384195 , n63543 , n384187 );
not ( n384196 , n63543 );
and ( n63555 , n384196 , n384186 );
nor ( n384198 , n384195 , n63555 );
not ( n384199 , n384198 );
buf ( n384200 , n384199 );
buf ( n384201 , n376997 );
and ( n384202 , n384200 , n384201 );
buf ( n384203 , n377003 );
nor ( n63562 , n63552 , n384202 , n384203 );
buf ( n384205 , n63562 );
buf ( n384206 , n384205 );
or ( n384207 , n384179 , n384206 );
buf ( n384208 , n384207 );
buf ( n384209 , n384208 );
xor ( n384210 , n384162 , n384209 );
buf ( n384211 , n378368 );
buf ( n384212 , n380817 );
and ( n384213 , n384211 , n384212 );
buf ( n384214 , n378372 );
buf ( n384215 , n57983 );
and ( n63574 , n384214 , n384215 );
nor ( n384217 , n384213 , n63574 );
buf ( n384218 , n384217 );
buf ( n384219 , n384218 );
buf ( n384220 , n60313 );
or ( n63579 , n384219 , n384220 );
buf ( n384222 , n382823 );
buf ( n384223 , n380733 );
or ( n63582 , n384222 , n384223 );
nand ( n384225 , n63579 , n63582 );
buf ( n384226 , n384225 );
buf ( n384227 , n384226 );
and ( n384228 , n384210 , n384227 );
and ( n384229 , n384162 , n384209 );
or ( n63588 , n384228 , n384229 );
buf ( n384231 , n63588 );
xor ( n384232 , n382831 , n382854 );
xor ( n384233 , n384232 , n382871 );
and ( n63592 , n384231 , n384233 );
buf ( n384235 , n380651 );
buf ( n384236 , n380570 );
and ( n63595 , n384235 , n384236 );
buf ( n384238 , n380657 );
buf ( n384239 , n60054 );
and ( n384240 , n384238 , n384239 );
nor ( n63599 , n63595 , n384240 );
buf ( n384242 , n63599 );
buf ( n384243 , n384242 );
buf ( n384244 , n380581 );
or ( n63603 , n384243 , n384244 );
buf ( n384246 , n382863 );
buf ( n384247 , n378453 );
or ( n63606 , n384246 , n384247 );
nand ( n384249 , n63603 , n63606 );
buf ( n384250 , n384249 );
buf ( n384251 , n384250 );
buf ( n384252 , n380838 );
buf ( n384253 , n57800 );
and ( n384254 , n384252 , n384253 );
buf ( n384255 , n380844 );
buf ( n384256 , n376903 );
and ( n384257 , n384255 , n384256 );
nor ( n384258 , n384254 , n384257 );
buf ( n384259 , n384258 );
buf ( n384260 , n384259 );
buf ( n384261 , n378341 );
or ( n63620 , n384260 , n384261 );
buf ( n384263 , n384036 );
buf ( n384264 , n378424 );
or ( n63623 , n384263 , n384264 );
nand ( n63624 , n63620 , n63623 );
buf ( n384267 , n63624 );
buf ( n384268 , n384267 );
xor ( n384269 , n384251 , n384268 );
xor ( n63628 , n384061 , n63459 );
xor ( n63629 , n63628 , n384119 );
buf ( n384272 , n63629 );
buf ( n384273 , n384272 );
and ( n63632 , n384269 , n384273 );
and ( n384275 , n384251 , n384268 );
or ( n384276 , n63632 , n384275 );
buf ( n384277 , n384276 );
xor ( n384278 , n382831 , n382854 );
xor ( n384279 , n384278 , n382871 );
and ( n63638 , n384277 , n384279 );
and ( n384281 , n384231 , n384277 );
or ( n384282 , n63592 , n63638 , n384281 );
xor ( n63641 , n384128 , n384131 );
xor ( n384284 , n63641 , n384136 );
and ( n63643 , n384282 , n384284 );
buf ( n384286 , n378214 );
buf ( n384287 , n382835 );
and ( n384288 , n384286 , n384287 );
buf ( n384289 , n57754 );
buf ( n384290 , n62243 );
and ( n384291 , n384289 , n384290 );
nor ( n63650 , n384288 , n384291 );
buf ( n63651 , n63650 );
buf ( n384294 , n63651 );
buf ( n384295 , n382849 );
or ( n63654 , n384294 , n384295 );
buf ( n384297 , n384150 );
buf ( n384298 , n384157 );
or ( n63657 , n384297 , n384298 );
nand ( n63658 , n63654 , n63657 );
buf ( n384301 , n63658 );
buf ( n384302 , n60089 );
buf ( n384303 , n380817 );
and ( n384304 , n384302 , n384303 );
buf ( n384305 , n60094 );
not ( n63664 , n57982 );
buf ( n384307 , n63664 );
and ( n384308 , n384305 , n384307 );
nor ( n63667 , n384304 , n384308 );
buf ( n63668 , n63667 );
buf ( n384311 , n63668 );
buf ( n384312 , n60313 );
or ( n384313 , n384311 , n384312 );
buf ( n384314 , n384218 );
buf ( n384315 , n380733 );
or ( n384316 , n384314 , n384315 );
nand ( n384317 , n384313 , n384316 );
buf ( n384318 , n384317 );
xor ( n384319 , n384301 , n384318 );
buf ( n384320 , n380680 );
buf ( n384321 , n380570 );
and ( n384322 , n384320 , n384321 );
buf ( n384323 , n60171 );
buf ( n384324 , n60054 );
and ( n63683 , n384323 , n384324 );
nor ( n384326 , n384322 , n63683 );
buf ( n384327 , n384326 );
buf ( n384328 , n384327 );
buf ( n384329 , n380581 );
or ( n63688 , n384328 , n384329 );
buf ( n384331 , n384242 );
buf ( n384332 , n378453 );
or ( n384333 , n384331 , n384332 );
nand ( n63692 , n63688 , n384333 );
buf ( n384335 , n63692 );
and ( n63694 , n384319 , n384335 );
and ( n63695 , n384301 , n384318 );
or ( n384338 , n63694 , n63695 );
buf ( n384339 , n384338 );
buf ( n384340 , n376743 );
buf ( n384341 , n384089 );
not ( n63700 , n384341 );
buf ( n384343 , n63700 );
buf ( n384344 , n384343 );
and ( n63703 , n384340 , n384344 );
buf ( n384346 , n376871 );
buf ( n384347 , n384089 );
and ( n63706 , n384346 , n384347 );
nor ( n384349 , n63703 , n63706 );
buf ( n384350 , n384349 );
buf ( n384351 , n384350 );
buf ( n384352 , n384085 );
not ( n384353 , n384352 );
buf ( n384354 , n384353 );
buf ( n384355 , n384354 );
or ( n384356 , n384351 , n384355 );
buf ( n384357 , n384097 );
nand ( n63716 , n384356 , n384357 );
buf ( n384359 , n63716 );
buf ( n384360 , n384359 );
buf ( n384361 , n61992 );
buf ( n384362 , n57800 );
and ( n63721 , n384361 , n384362 );
buf ( n63722 , n382596 );
buf ( n63723 , n376903 );
and ( n63724 , n63722 , n63723 );
nor ( n63725 , n63721 , n63724 );
buf ( n63726 , n63725 );
buf ( n384369 , n63726 );
buf ( n384370 , n378341 );
or ( n384371 , n384369 , n384370 );
buf ( n384372 , n384259 );
buf ( n384373 , n378424 );
or ( n384374 , n384372 , n384373 );
nand ( n63733 , n384371 , n384374 );
buf ( n384376 , n63733 );
buf ( n384377 , n384376 );
xor ( n384378 , n384360 , n384377 );
and ( n63737 , n63538 , n384184 );
xor ( n384380 , n63737 , n376699 );
buf ( n384381 , n384380 );
buf ( n384382 , n376990 );
and ( n384383 , n384381 , n384382 );
buf ( n384384 , n384380 );
not ( n63743 , n384384 );
buf ( n384386 , n63743 );
buf ( n384387 , n384386 );
buf ( n384388 , n376997 );
and ( n384389 , n384387 , n384388 );
buf ( n384390 , n377003 );
nor ( n384391 , n384383 , n384389 , n384390 );
buf ( n384392 , n384391 );
buf ( n384393 , n384392 );
nor ( n63752 , n60202 , n56364 );
and ( n384395 , n63752 , n62016 );
not ( n63754 , n63752 );
and ( n384397 , n63754 , n62015 );
or ( n384398 , n384395 , n384397 );
buf ( n384399 , n384398 );
not ( n384400 , n574 );
not ( n384401 , n320740 );
or ( n63760 , n384400 , n384401 );
nand ( n63761 , n63760 , n56367 );
and ( n63762 , n63761 , n56370 );
not ( n384405 , n63761 );
and ( n384406 , n384405 , n376779 );
or ( n63765 , n63762 , n384406 );
not ( n384408 , n63765 );
buf ( n384409 , n384408 );
xor ( n63768 , n384399 , n384409 );
buf ( n384411 , n63768 );
not ( n63770 , n384411 );
xor ( n63771 , n384398 , n63434 );
nand ( n384414 , n63770 , n63771 );
buf ( n384415 , n384414 );
not ( n63774 , n384415 );
buf ( n384417 , n63774 );
buf ( n63776 , n384417 );
buf ( n384419 , n63434 );
buf ( n63778 , n384419 );
buf ( n384421 , n63778 );
buf ( n384422 , n384421 );
nand ( n384423 , n63776 , n384422 );
buf ( n384424 , n384423 );
buf ( n384425 , n384424 );
buf ( n384426 , n384421 );
buf ( n384427 , n384411 );
nand ( n63786 , n384426 , n384427 );
buf ( n384429 , n63786 );
buf ( n384430 , n384429 );
and ( n384431 , n384425 , n384430 );
buf ( n384432 , n384431 );
buf ( n384433 , n384432 );
xor ( n63792 , n384393 , n384433 );
buf ( n384435 , n63549 );
buf ( n384436 , n376866 );
and ( n384437 , n384435 , n384436 );
buf ( n384438 , n384199 );
buf ( n384439 , n382743 );
and ( n384440 , n384438 , n384439 );
nor ( n63799 , n384437 , n384440 );
buf ( n63800 , n63799 );
buf ( n384443 , n63800 );
buf ( n384444 , n376924 );
or ( n384445 , n384443 , n384444 );
buf ( n384446 , n384170 );
buf ( n384447 , n56517 );
or ( n63806 , n384446 , n384447 );
nand ( n63807 , n384445 , n63806 );
buf ( n384450 , n63807 );
buf ( n384451 , n384450 );
and ( n63810 , n63792 , n384451 );
and ( n384453 , n384393 , n384433 );
or ( n384454 , n63810 , n384453 );
buf ( n384455 , n384454 );
buf ( n384456 , n384455 );
and ( n384457 , n384378 , n384456 );
and ( n63816 , n384360 , n384377 );
or ( n384459 , n384457 , n63816 );
buf ( n384460 , n384459 );
buf ( n384461 , n384460 );
xor ( n384462 , n384339 , n384461 );
xor ( n384463 , n384162 , n384209 );
xor ( n63822 , n384463 , n384227 );
buf ( n384465 , n63822 );
buf ( n384466 , n384465 );
and ( n63825 , n384462 , n384466 );
and ( n384468 , n384339 , n384461 );
or ( n384469 , n63825 , n384468 );
buf ( n384470 , n384469 );
xor ( n63829 , n384028 , n63403 );
xor ( n63830 , n63829 , n384124 );
buf ( n384473 , n63830 );
xor ( n384474 , n384470 , n384473 );
xor ( n63833 , n382831 , n382854 );
xor ( n384476 , n63833 , n382871 );
xor ( n63835 , n384231 , n384277 );
xor ( n63836 , n384476 , n63835 );
and ( n384479 , n384474 , n63836 );
and ( n384480 , n384470 , n384473 );
or ( n63839 , n384479 , n384480 );
xor ( n384482 , n384128 , n384131 );
xor ( n384483 , n384482 , n384136 );
and ( n63842 , n63839 , n384483 );
and ( n384485 , n384282 , n63839 );
or ( n63844 , n63643 , n63842 , n384485 );
xor ( n63845 , n382879 , n382882 );
xor ( n63846 , n63845 , n382886 );
and ( n384489 , n63844 , n63846 );
and ( n63848 , n63497 , n63844 );
or ( n63849 , n63500 , n384489 , n63848 );
buf ( n384492 , n63849 );
xor ( n63851 , n384019 , n384492 );
buf ( n63852 , n56794 );
not ( n63853 , n63852 );
buf ( n63854 , n383971 );
not ( n63855 , n63854 );
or ( n63856 , n63853 , n63855 );
buf ( n63857 , n365722 );
not ( n384500 , n63857 );
buf ( n384501 , n384500 );
buf ( n384502 , n384501 );
and ( n384503 , n351160 , n61903 );
not ( n63862 , n351160 );
and ( n384505 , n63862 , n22619 );
or ( n63864 , n384503 , n384505 );
buf ( n384507 , n63864 );
nand ( n63866 , n384502 , n384507 );
buf ( n384509 , n63866 );
buf ( n384510 , n384509 );
nand ( n63869 , n63856 , n384510 );
buf ( n384512 , n63869 );
buf ( n384513 , n384512 );
and ( n63872 , n63851 , n384513 );
and ( n63873 , n384019 , n384492 );
or ( n384516 , n63872 , n63873 );
buf ( n384517 , n384516 );
buf ( n384518 , n384517 );
buf ( n384519 , n365108 );
not ( n63878 , n384519 );
buf ( n384521 , n383258 );
not ( n63880 , n384521 );
or ( n63881 , n63878 , n63880 );
buf ( n384524 , n364981 );
not ( n384525 , n384524 );
buf ( n384526 , n375873 );
not ( n384527 , n384526 );
or ( n63886 , n384525 , n384527 );
buf ( n384529 , n31231 );
buf ( n384530 , n62345 );
nand ( n384531 , n384529 , n384530 );
buf ( n384532 , n384531 );
buf ( n384533 , n384532 );
nand ( n384534 , n63886 , n384533 );
buf ( n384535 , n384534 );
buf ( n384536 , n384535 );
buf ( n63895 , n365024 );
nand ( n63896 , n384536 , n63895 );
buf ( n384539 , n63896 );
buf ( n384540 , n384539 );
nand ( n384541 , n63881 , n384540 );
buf ( n384542 , n384541 );
buf ( n384543 , n384542 );
xor ( n384544 , n384518 , n384543 );
buf ( n384545 , n365428 );
not ( n384546 , n384545 );
not ( n63905 , n56849 );
buf ( n384548 , n63905 );
not ( n384549 , n384548 );
or ( n63908 , n384546 , n384549 );
buf ( n384551 , n342656 );
buf ( n384552 , n365422 );
nand ( n384553 , n384551 , n384552 );
buf ( n384554 , n384553 );
buf ( n384555 , n384554 );
nand ( n384556 , n63908 , n384555 );
buf ( n384557 , n384556 );
buf ( n384558 , n384557 );
not ( n384559 , n384558 );
buf ( n384560 , n366399 );
not ( n384561 , n384560 );
or ( n63920 , n384559 , n384561 );
buf ( n384563 , n383231 );
buf ( n384564 , n377171 );
nand ( n384565 , n384563 , n384564 );
buf ( n384566 , n384565 );
buf ( n384567 , n384566 );
nand ( n384568 , n63920 , n384567 );
buf ( n384569 , n384568 );
buf ( n384570 , n384569 );
and ( n63929 , n384544 , n384570 );
and ( n384572 , n384518 , n384543 );
or ( n63931 , n63929 , n384572 );
buf ( n384574 , n63931 );
nand ( n384575 , n63366 , n63370 );
and ( n384576 , n384574 , n384575 );
nor ( n63935 , n384014 , n384576 );
buf ( n384578 , n63935 );
not ( n384579 , n384578 );
buf ( n384580 , n384579 );
buf ( n384581 , n384580 );
nand ( n384582 , n63306 , n384581 );
buf ( n384583 , n384582 );
nand ( n384584 , n63295 , n384583 );
nand ( n63943 , n383900 , n384584 );
nand ( n63944 , n63257 , n63943 );
buf ( n384587 , n63944 );
and ( n384588 , n383872 , n384587 );
not ( n63947 , n63223 );
nor ( n384590 , n63947 , n63198 );
buf ( n63949 , n384590 );
nor ( n63950 , n384588 , n63949 );
buf ( n63951 , n63950 );
buf ( n384594 , n63951 );
xor ( n63953 , n383834 , n384594 );
buf ( n384596 , n379890 );
not ( n63955 , n384596 );
buf ( n384598 , n61618 );
not ( n63957 , n384598 );
or ( n384600 , n63955 , n63957 );
buf ( n384601 , n379847 );
buf ( n384602 , n367158 );
and ( n63961 , n384601 , n384602 );
not ( n384604 , n384601 );
buf ( n384605 , n40251 );
and ( n63964 , n384604 , n384605 );
nor ( n63965 , n63961 , n63964 );
buf ( n63966 , n63965 );
buf ( n384609 , n63966 );
buf ( n384610 , n379916 );
nand ( n63969 , n384609 , n384610 );
buf ( n384612 , n63969 );
buf ( n384613 , n384612 );
nand ( n63972 , n384600 , n384613 );
buf ( n384615 , n63972 );
xor ( n384616 , n381139 , n381140 );
buf ( n384617 , n384616 );
buf ( n384618 , n384617 );
buf ( n384619 , n381133 );
and ( n384620 , n384618 , n384619 );
not ( n384621 , n384618 );
buf ( n384622 , n381133 );
not ( n63981 , n384622 );
buf ( n63982 , n63981 );
buf ( n384625 , n63982 );
and ( n384626 , n384621 , n384625 );
nor ( n63985 , n384620 , n384626 );
buf ( n384628 , n63985 );
or ( n384629 , n384615 , n384628 );
buf ( n384630 , n384629 );
xor ( n63989 , n381890 , n381916 );
xor ( n384632 , n63989 , n381939 );
buf ( n384633 , n384632 );
buf ( n384634 , n384633 );
and ( n384635 , n384630 , n384634 );
buf ( n384636 , n384615 );
buf ( n384637 , n384628 );
and ( n384638 , n384636 , n384637 );
buf ( n384639 , n384638 );
buf ( n384640 , n384639 );
nor ( n384641 , n384635 , n384640 );
buf ( n384642 , n384641 );
buf ( n384643 , n384642 );
and ( n64002 , n63953 , n384643 );
and ( n384645 , n383834 , n384594 );
or ( n384646 , n64002 , n384645 );
buf ( n384647 , n384646 );
not ( n64006 , n384647 );
not ( n384649 , n64006 );
or ( n64008 , n383821 , n384649 );
buf ( n384651 , n383820 );
not ( n64010 , n384651 );
buf ( n384653 , n64010 );
not ( n384654 , n384653 );
not ( n384655 , n384647 );
or ( n64014 , n384654 , n384655 );
buf ( n384657 , n380407 );
not ( n64016 , n384657 );
buf ( n384659 , n380368 );
not ( n384660 , n384659 );
buf ( n384661 , n365206 );
not ( n384662 , n384661 );
or ( n384663 , n384660 , n384662 );
buf ( n384664 , n371416 );
buf ( n384665 , n380368 );
not ( n384666 , n384665 );
buf ( n384667 , n384666 );
buf ( n384668 , n384667 );
nand ( n384669 , n384664 , n384668 );
buf ( n384670 , n384669 );
buf ( n384671 , n384670 );
nand ( n64030 , n384663 , n384671 );
buf ( n384673 , n64030 );
buf ( n384674 , n384673 );
not ( n64033 , n384674 );
or ( n64034 , n64016 , n64033 );
buf ( n384677 , n380393 );
buf ( n384678 , n380356 );
nand ( n384679 , n384677 , n384678 );
buf ( n384680 , n384679 );
buf ( n384681 , n384680 );
nand ( n384682 , n64034 , n384681 );
buf ( n384683 , n384682 );
buf ( n384684 , n384683 );
buf ( n384685 , n58923 );
not ( n384686 , n384685 );
buf ( n384687 , n61190 );
not ( n64046 , n384687 );
or ( n384689 , n384686 , n64046 );
buf ( n384690 , n379371 );
not ( n384691 , n384690 );
buf ( n384692 , n364987 );
not ( n384693 , n384692 );
or ( n64052 , n384691 , n384693 );
buf ( n384695 , n359781 );
buf ( n384696 , n379380 );
nand ( n384697 , n384695 , n384696 );
buf ( n384698 , n384697 );
buf ( n384699 , n384698 );
nand ( n384700 , n64052 , n384699 );
buf ( n384701 , n384700 );
buf ( n384702 , n384701 );
buf ( n384703 , n58871 );
nand ( n64062 , n384702 , n384703 );
buf ( n384705 , n64062 );
buf ( n384706 , n384705 );
nand ( n64065 , n384689 , n384706 );
buf ( n384708 , n64065 );
buf ( n384709 , n384708 );
xor ( n64068 , n384684 , n384709 );
buf ( n384711 , n369444 );
not ( n384712 , n384711 );
buf ( n384713 , n381080 );
not ( n64072 , n384713 );
or ( n384715 , n384712 , n64072 );
buf ( n384716 , n383492 );
buf ( n384717 , n368608 );
nand ( n64076 , n384716 , n384717 );
buf ( n64077 , n64076 );
buf ( n384720 , n64077 );
nand ( n64079 , n384715 , n384720 );
buf ( n64080 , n64079 );
buf ( n384723 , n64080 );
buf ( n384724 , n383455 );
not ( n384725 , n384724 );
buf ( n384726 , n362027 );
not ( n64085 , n384726 );
or ( n384728 , n384725 , n64085 );
buf ( n384729 , n364824 );
buf ( n384730 , n381354 );
nand ( n64089 , n384729 , n384730 );
buf ( n64090 , n64089 );
buf ( n384733 , n64090 );
nand ( n384734 , n384728 , n384733 );
buf ( n384735 , n384734 );
buf ( n384736 , n384735 );
xor ( n384737 , n384723 , n384736 );
xor ( n64096 , n383525 , n62901 );
and ( n64097 , n64096 , n383568 );
and ( n384740 , n383525 , n62901 );
or ( n384741 , n64097 , n384740 );
buf ( n384742 , n384741 );
and ( n64101 , n384737 , n384742 );
and ( n64102 , n384723 , n384736 );
or ( n384745 , n64101 , n64102 );
buf ( n384746 , n384745 );
buf ( n384747 , n384746 );
xor ( n64106 , n381211 , n381349 );
xor ( n64107 , n64106 , n381379 );
buf ( n384750 , n64107 );
buf ( n384751 , n384750 );
xor ( n64110 , n384747 , n384751 );
buf ( n384753 , n62999 );
not ( n64112 , n384753 );
buf ( n384755 , n369260 );
not ( n64114 , n384755 );
or ( n384757 , n64112 , n64114 );
buf ( n384758 , n39217 );
buf ( n384759 , n381112 );
nand ( n64118 , n384758 , n384759 );
buf ( n384761 , n64118 );
buf ( n384762 , n384761 );
nand ( n64121 , n384757 , n384762 );
buf ( n384764 , n64121 );
buf ( n384765 , n384764 );
buf ( n384766 , n378098 );
not ( n64125 , n384766 );
buf ( n384768 , n39963 );
not ( n64127 , n384768 );
or ( n384770 , n64125 , n64127 );
buf ( n384771 , n365507 );
buf ( n384772 , n379515 );
nand ( n64131 , n384771 , n384772 );
buf ( n384774 , n64131 );
buf ( n384775 , n384774 );
nand ( n384776 , n384770 , n384775 );
buf ( n384777 , n384776 );
buf ( n384778 , n384777 );
not ( n384779 , n384778 );
buf ( n384780 , n40058 );
not ( n384781 , n384780 );
or ( n64140 , n384779 , n384781 );
buf ( n384783 , n39949 );
buf ( n384784 , n382114 );
nand ( n64143 , n384783 , n384784 );
buf ( n384786 , n64143 );
buf ( n384787 , n384786 );
nand ( n384788 , n64140 , n384787 );
buf ( n384789 , n384788 );
buf ( n384790 , n384789 );
xor ( n384791 , n384765 , n384790 );
buf ( n384792 , n58984 );
not ( n384793 , n384792 );
buf ( n384794 , n45270 );
not ( n64153 , n384794 );
or ( n64154 , n384793 , n64153 );
buf ( n384797 , n362452 );
buf ( n384798 , n379482 );
nand ( n384799 , n384797 , n384798 );
buf ( n384800 , n384799 );
buf ( n64159 , n384800 );
nand ( n384802 , n64154 , n64159 );
buf ( n384803 , n384802 );
buf ( n384804 , n384803 );
not ( n384805 , n384804 );
buf ( n384806 , n46557 );
not ( n64165 , n384806 );
or ( n384808 , n384805 , n64165 );
buf ( n384809 , n360577 );
buf ( n384810 , n382151 );
nand ( n384811 , n384809 , n384810 );
buf ( n384812 , n384811 );
buf ( n384813 , n384812 );
nand ( n64172 , n384808 , n384813 );
buf ( n64173 , n64172 );
buf ( n384816 , n64173 );
and ( n384817 , n384791 , n384816 );
and ( n64176 , n384765 , n384790 );
or ( n384819 , n384817 , n64176 );
buf ( n384820 , n384819 );
buf ( n384821 , n384820 );
and ( n64180 , n64110 , n384821 );
and ( n384823 , n384747 , n384751 );
or ( n384824 , n64180 , n384823 );
buf ( n384825 , n384824 );
buf ( n384826 , n384825 );
and ( n64185 , n64068 , n384826 );
and ( n384828 , n384684 , n384709 );
or ( n384829 , n64185 , n384828 );
buf ( n384830 , n384829 );
nand ( n64189 , n64014 , n384830 );
nand ( n384832 , n64008 , n64189 );
buf ( n384833 , n384832 );
nand ( n64192 , n383817 , n384833 );
buf ( n384835 , n64192 );
buf ( n384836 , n384835 );
nand ( n64195 , n383809 , n384836 );
buf ( n384838 , n64195 );
buf ( n384839 , n384838 );
nand ( n64198 , n383770 , n384839 );
buf ( n384841 , n64198 );
nand ( n384842 , n63127 , n384841 );
buf ( n384843 , n384842 );
xor ( n384844 , n381030 , n384843 );
xor ( n64203 , n381487 , n61145 );
and ( n384846 , n64203 , n382344 );
and ( n384847 , n381487 , n61145 );
or ( n64206 , n384846 , n384847 );
buf ( n384849 , n64206 );
buf ( n384850 , n384849 );
nand ( n384851 , n59770 , n59773 );
not ( n64210 , n384851 );
not ( n64211 , n59786 );
or ( n384854 , n64210 , n64211 );
nand ( n384855 , n59742 , n380282 );
nand ( n64214 , n384854 , n384855 );
buf ( n384857 , n64214 );
buf ( n384858 , n59766 );
not ( n64217 , n384858 );
buf ( n384860 , n59753 );
not ( n384861 , n384860 );
or ( n384862 , n64217 , n384861 );
buf ( n384863 , n59766 );
buf ( n384864 , n59753 );
or ( n384865 , n384863 , n384864 );
buf ( n384866 , n380261 );
nand ( n384867 , n384865 , n384866 );
buf ( n384868 , n384867 );
buf ( n384869 , n384868 );
nand ( n384870 , n384862 , n384869 );
buf ( n384871 , n384870 );
buf ( n384872 , n384871 );
xor ( n384873 , n381548 , n381563 );
and ( n384874 , n384873 , n381577 );
and ( n384875 , n381548 , n381563 );
or ( n64234 , n384874 , n384875 );
buf ( n384877 , n64234 );
buf ( n64236 , n384877 );
and ( n64237 , n384872 , n64236 );
not ( n384880 , n384872 );
not ( n384881 , n384877 );
buf ( n384882 , n384881 );
and ( n384883 , n384880 , n384882 );
nor ( n384884 , n64237 , n384883 );
buf ( n384885 , n384884 );
not ( n384886 , n384885 );
not ( n384887 , n384886 );
buf ( n384888 , n380047 );
not ( n64247 , n384888 );
buf ( n384890 , n366237 );
nor ( n64249 , n64247 , n384890 );
buf ( n384892 , n64249 );
not ( n384893 , n384892 );
not ( n384894 , n381596 );
nand ( n384895 , n384894 , n368051 );
nand ( n64254 , n384893 , n384895 );
not ( n384897 , n64254 );
not ( n384898 , n384897 );
or ( n64257 , n384887 , n384898 );
nand ( n64258 , n384885 , n64254 );
nand ( n384901 , n64257 , n64258 );
not ( n384902 , n381642 );
not ( n64261 , n381579 );
nand ( n64262 , n64261 , n381602 );
not ( n64263 , n64262 );
or ( n384906 , n384902 , n64263 );
buf ( n384907 , n381579 );
nand ( n64266 , n384907 , n381605 );
nand ( n64267 , n384906 , n64266 );
and ( n64268 , n384901 , n64267 );
not ( n384911 , n384901 );
not ( n64270 , n64267 );
and ( n64271 , n384911 , n64270 );
nor ( n64272 , n64268 , n64271 );
xnor ( n64273 , n384857 , n64272 );
buf ( n384916 , n64273 );
buf ( n384917 , n59419 );
not ( n64276 , n384917 );
buf ( n384919 , n64276 );
buf ( n384920 , n384919 );
not ( n64279 , n384920 );
buf ( n384922 , n379893 );
not ( n64281 , n384922 );
and ( n64282 , n64279 , n64281 );
buf ( n384925 , n60959 );
buf ( n384926 , n379916 );
and ( n384927 , n384925 , n384926 );
nor ( n64286 , n64282 , n384927 );
buf ( n384929 , n64286 );
buf ( n384930 , n384929 );
buf ( n64289 , n359136 );
nand ( n64290 , n64289 , n39046 , n59867 );
nand ( n384933 , n373845 , n380368 );
nand ( n384934 , n64290 , n384933 );
not ( n384935 , n384934 );
buf ( n384936 , n384935 );
not ( n384937 , n384936 );
buf ( n384938 , n380356 );
not ( n64297 , n384938 );
buf ( n384940 , n64297 );
buf ( n384941 , n384940 );
not ( n384942 , n384941 );
and ( n384943 , n384937 , n384942 );
buf ( n384944 , n381502 );
buf ( n384945 , n380404 );
and ( n64304 , n384944 , n384945 );
nor ( n384947 , n384943 , n64304 );
buf ( n384948 , n384947 );
buf ( n384949 , n384948 );
xor ( n384950 , n384930 , n384949 );
buf ( n384951 , n384950 );
buf ( n384952 , n384951 );
and ( n384953 , n380178 , n380166 );
not ( n64312 , n380178 );
and ( n64313 , n64312 , n59661 );
or ( n384956 , n384953 , n64313 );
xor ( n384957 , n384956 , n380130 );
buf ( n384958 , n384957 );
xor ( n64317 , n384952 , n384958 );
buf ( n384960 , n64317 );
buf ( n384961 , n384960 );
xor ( n64320 , n384916 , n384961 );
not ( n64321 , n62725 );
buf ( n384964 , n62729 );
not ( n384965 , n384964 );
buf ( n384966 , n384965 );
buf ( n384967 , n384966 );
buf ( n384968 , n383379 );
nand ( n384969 , n384967 , n384968 );
buf ( n384970 , n384969 );
not ( n64329 , n384970 );
or ( n64330 , n64321 , n64329 );
not ( n384973 , n383379 );
nand ( n384974 , n384973 , n62729 );
nand ( n384975 , n64330 , n384974 );
buf ( n384976 , n384975 );
xor ( n384977 , n383335 , n62696 );
and ( n384978 , n384977 , n383356 );
and ( n64337 , n383335 , n62696 );
or ( n64338 , n384978 , n64337 );
buf ( n384981 , n64338 );
buf ( n384982 , n384981 );
or ( n64341 , n384976 , n384982 );
buf ( n384984 , n61512 );
not ( n384985 , n384984 );
buf ( n384986 , n382098 );
not ( n384987 , n384986 );
or ( n384988 , n384985 , n384987 );
not ( n64347 , n382103 );
not ( n64348 , n382073 );
or ( n384991 , n64347 , n64348 );
nand ( n384992 , n384991 , n382064 );
buf ( n384993 , n384992 );
nand ( n64352 , n384988 , n384993 );
buf ( n384995 , n64352 );
buf ( n384996 , n384995 );
nand ( n64355 , n64341 , n384996 );
buf ( n384998 , n64355 );
buf ( n384999 , n384998 );
buf ( n385000 , n384975 );
buf ( n385001 , n384981 );
nand ( n64360 , n385000 , n385001 );
buf ( n385003 , n64360 );
buf ( n385004 , n385003 );
nand ( n64363 , n384999 , n385004 );
buf ( n385006 , n64363 );
buf ( n385007 , n385006 );
and ( n64366 , n64320 , n385007 );
and ( n64367 , n384916 , n384961 );
or ( n64368 , n64366 , n64367 );
buf ( n385011 , n64368 );
buf ( n385012 , n385011 );
not ( n64371 , n385012 );
buf ( n385014 , n64371 );
buf ( n385015 , n385014 );
not ( n64374 , n385015 );
buf ( n385017 , n381651 );
not ( n64376 , n385017 );
buf ( n385019 , n381654 );
not ( n64378 , n385019 );
buf ( n385021 , n64378 );
buf ( n385022 , n385021 );
nand ( n64381 , n64376 , n385022 );
buf ( n385024 , n64381 );
buf ( n385025 , n385024 );
buf ( n385026 , n381704 );
and ( n64385 , n385025 , n385026 );
buf ( n385028 , n381651 );
not ( n64387 , n385028 );
buf ( n385030 , n385021 );
nor ( n64389 , n64387 , n385030 );
buf ( n385032 , n64389 );
buf ( n385033 , n385032 );
nor ( n64392 , n64385 , n385033 );
buf ( n385035 , n64392 );
buf ( n385036 , n385035 );
not ( n64395 , n385036 );
buf ( n385038 , n64395 );
buf ( n385039 , n385038 );
not ( n385040 , n385039 );
not ( n64399 , n64270 );
not ( n64400 , n64214 );
not ( n385043 , n64400 );
or ( n385044 , n64399 , n385043 );
not ( n64403 , n64267 );
not ( n385046 , n64214 );
or ( n385047 , n64403 , n385046 );
nand ( n64406 , n385047 , n384901 );
nand ( n385049 , n385044 , n64406 );
buf ( n385050 , n385049 );
not ( n64409 , n384929 );
not ( n64410 , n384948 );
and ( n385053 , n64409 , n64410 );
buf ( n385054 , n384929 );
buf ( n385055 , n384948 );
nand ( n385056 , n385054 , n385055 );
buf ( n385057 , n385056 );
and ( n64416 , n384957 , n385057 );
nor ( n385059 , n385053 , n64416 );
buf ( n64418 , n385059 );
xor ( n64419 , n385050 , n64418 );
buf ( n385062 , n380404 );
not ( n385063 , n385062 );
buf ( n385064 , n385063 );
buf ( n385065 , n385064 );
buf ( n385066 , n384940 );
nand ( n64425 , n385065 , n385066 );
buf ( n385068 , n64425 );
nand ( n64427 , n384934 , n385068 );
buf ( n385070 , n64427 );
not ( n385071 , n384881 );
not ( n64430 , n385071 );
not ( n385073 , n64254 );
or ( n385074 , n64430 , n385073 );
or ( n64433 , n385071 , n64254 );
nand ( n385076 , n64433 , n384871 );
nand ( n64435 , n385074 , n385076 );
buf ( n385078 , n64435 );
xor ( n385079 , n385070 , n385078 );
xor ( n385080 , n379803 , n379811 );
and ( n64439 , n385080 , n59334 );
and ( n385082 , n379803 , n379811 );
or ( n64441 , n64439 , n385082 );
buf ( n385084 , n64441 );
xnor ( n64443 , n385079 , n385084 );
buf ( n64444 , n64443 );
buf ( n385087 , n64444 );
xor ( n385088 , n64419 , n385087 );
buf ( n385089 , n385088 );
buf ( n385090 , n385089 );
not ( n64449 , n385090 );
or ( n385092 , n385040 , n64449 );
buf ( n385093 , n385089 );
not ( n64452 , n385093 );
buf ( n64453 , n64452 );
buf ( n385096 , n64453 );
buf ( n385097 , n385035 );
nand ( n385098 , n385096 , n385097 );
buf ( n385099 , n385098 );
buf ( n385100 , n385099 );
nand ( n64459 , n385092 , n385100 );
buf ( n385102 , n64459 );
buf ( n385103 , n385102 );
not ( n385104 , n385103 );
or ( n64463 , n64374 , n385104 );
buf ( n385106 , n385102 );
buf ( n385107 , n385014 );
or ( n385108 , n385106 , n385107 );
nand ( n64467 , n64463 , n385108 );
buf ( n64468 , n64467 );
buf ( n385111 , n64468 );
xor ( n64470 , n384850 , n385111 );
xor ( n385113 , n384916 , n384961 );
xor ( n64472 , n385113 , n385007 );
buf ( n385115 , n64472 );
buf ( n64474 , n385115 );
buf ( n385117 , n384981 );
buf ( n385118 , n384975 );
xor ( n385119 , n385117 , n385118 );
buf ( n385120 , n384995 );
xnor ( n64479 , n385119 , n385120 );
buf ( n385122 , n64479 );
buf ( n385123 , n385122 );
not ( n64482 , n385123 );
buf ( n64483 , n64482 );
not ( n385126 , n64483 );
xor ( n64485 , n60971 , n60943 );
xor ( n385128 , n64485 , n381645 );
not ( n385129 , n385128 );
or ( n64488 , n385126 , n385129 );
buf ( n385131 , n385128 );
not ( n385132 , n385131 );
buf ( n385133 , n385132 );
not ( n385134 , n385133 );
not ( n385135 , n385122 );
or ( n64494 , n385134 , n385135 );
buf ( n385137 , n59792 );
buf ( n385138 , n59803 );
xor ( n385139 , n385137 , n385138 );
buf ( n64498 , n380988 );
xor ( n64499 , n385139 , n64498 );
buf ( n385142 , n64499 );
nand ( n64501 , n64494 , n385142 );
nand ( n385144 , n64488 , n64501 );
buf ( n64503 , n385144 );
xor ( n64504 , n64474 , n64503 );
not ( n64505 , n60503 );
or ( n385148 , n60487 , n380994 );
nand ( n64507 , n60487 , n380994 );
nand ( n385150 , n385148 , n64507 );
and ( n64509 , n64505 , n385150 );
not ( n64510 , n64505 );
and ( n64511 , n60489 , n60487 );
and ( n64512 , n64510 , n64511 );
nor ( n385155 , n64509 , n64512 );
nand ( n64514 , n60484 , n60503 , n380994 );
nand ( n385157 , n385155 , n64514 );
buf ( n385158 , n385157 );
and ( n64517 , n64504 , n385158 );
and ( n385160 , n64474 , n64503 );
or ( n64519 , n64517 , n385160 );
buf ( n385162 , n64519 );
buf ( n385163 , n385162 );
xor ( n64522 , n64470 , n385163 );
buf ( n385165 , n64522 );
xor ( n64524 , n384844 , n385165 );
buf ( n385167 , n384838 );
buf ( n385168 , n382346 );
xor ( n385169 , n385167 , n385168 );
buf ( n385170 , n383766 );
xnor ( n385171 , n385169 , n385170 );
buf ( n385172 , n385171 );
not ( n64531 , n385172 );
not ( n64532 , n64531 );
xor ( n64533 , n64474 , n64503 );
xor ( n385176 , n64533 , n385158 );
buf ( n385177 , n385176 );
not ( n385178 , n385177 );
or ( n64537 , n64532 , n385178 );
not ( n64538 , n385177 );
not ( n385181 , n64538 );
not ( n385182 , n385172 );
or ( n64541 , n385181 , n385182 );
buf ( n385184 , n385128 );
buf ( n385185 , n385142 );
xor ( n64544 , n385184 , n385185 );
buf ( n385187 , n64483 );
xnor ( n64546 , n64544 , n385187 );
buf ( n385189 , n64546 );
buf ( n385190 , n385189 );
buf ( n385191 , n383775 );
buf ( n385192 , n384832 );
xor ( n64551 , n385191 , n385192 );
buf ( n385194 , n63164 );
xnor ( n64553 , n64551 , n385194 );
buf ( n385196 , n64553 );
buf ( n385197 , n385196 );
xor ( n64556 , n385190 , n385197 );
xor ( n64557 , n382514 , n62330 );
xor ( n64558 , n64557 , n382956 );
buf ( n385201 , n64558 );
buf ( n385202 , n365393 );
not ( n64561 , n385202 );
buf ( n385204 , n342718 );
not ( n64563 , n385204 );
or ( n64564 , n64561 , n64563 );
not ( n385207 , n42233 );
nand ( n385208 , n385207 , n365408 );
buf ( n385209 , n385208 );
nand ( n385210 , n64564 , n385209 );
buf ( n385211 , n385210 );
buf ( n385212 , n385211 );
not ( n64571 , n385212 );
buf ( n385214 , n363429 );
not ( n385215 , n385214 );
or ( n385216 , n64571 , n385215 );
buf ( n385217 , n383174 );
buf ( n385218 , n57228 );
nand ( n64577 , n385217 , n385218 );
buf ( n385220 , n64577 );
buf ( n385221 , n385220 );
nand ( n64580 , n385216 , n385221 );
buf ( n385223 , n64580 );
buf ( n385224 , n385223 );
not ( n64583 , n385224 );
buf ( n385226 , n64583 );
buf ( n385227 , n385226 );
not ( n64586 , n385227 );
not ( n64587 , n377842 );
not ( n64588 , n383556 );
or ( n64589 , n64587 , n64588 );
not ( n385232 , n368994 );
not ( n64591 , n342335 );
or ( n385234 , n385232 , n64591 );
buf ( n385235 , n342338 );
buf ( n385236 , n368994 );
not ( n385237 , n385236 );
buf ( n385238 , n385237 );
buf ( n385239 , n385238 );
nand ( n64598 , n385235 , n385239 );
buf ( n385241 , n64598 );
nand ( n385242 , n385234 , n385241 );
buf ( n385243 , n362403 );
nand ( n64602 , n385242 , n385243 , n362385 );
nand ( n385245 , n64589 , n64602 );
buf ( n385246 , n385245 );
not ( n64605 , n385246 );
buf ( n64606 , n64605 );
buf ( n385249 , n64606 );
not ( n64608 , n385249 );
or ( n64609 , n64586 , n64608 );
buf ( n385252 , n45075 );
not ( n385253 , n385252 );
buf ( n385254 , n383515 );
not ( n385255 , n385254 );
or ( n385256 , n385253 , n385255 );
xor ( n385257 , n352209 , n22930 );
buf ( n385258 , n385257 );
buf ( n385259 , n365226 );
nand ( n385260 , n385258 , n385259 );
buf ( n385261 , n385260 );
buf ( n385262 , n385261 );
nand ( n385263 , n385256 , n385262 );
buf ( n385264 , n385263 );
buf ( n385265 , n385264 );
nand ( n385266 , n64609 , n385265 );
buf ( n385267 , n385266 );
buf ( n385268 , n385267 );
buf ( n385269 , n385223 );
buf ( n385270 , n385245 );
nand ( n385271 , n385269 , n385270 );
buf ( n385272 , n385271 );
buf ( n385273 , n385272 );
nand ( n385274 , n385268 , n385273 );
buf ( n385275 , n385274 );
buf ( n385276 , n385275 );
xor ( n385277 , n385201 , n385276 );
not ( n385278 , n378098 );
nor ( n385279 , n385278 , n377116 );
buf ( n385280 , n385279 );
and ( n64615 , n385277 , n385280 );
and ( n64616 , n385201 , n385276 );
or ( n385283 , n64615 , n64616 );
buf ( n385284 , n385283 );
buf ( n385285 , n385284 );
buf ( n385286 , n49609 );
not ( n64621 , n385286 );
buf ( n385288 , n383300 );
not ( n385289 , n385288 );
or ( n64624 , n64621 , n385289 );
buf ( n385291 , n383590 );
buf ( n385292 , n369804 );
nand ( n64627 , n385291 , n385292 );
buf ( n64628 , n64627 );
buf ( n385295 , n64628 );
nand ( n64630 , n64624 , n385295 );
buf ( n385297 , n64630 );
buf ( n385298 , n385297 );
xor ( n64633 , n385285 , n385298 );
buf ( n385300 , n377122 );
not ( n64635 , n385300 );
not ( n64636 , n45092 );
buf ( n385303 , n64636 );
not ( n385304 , n385303 );
or ( n64639 , n64635 , n385304 );
buf ( n385306 , n365293 );
buf ( n385307 , n57463 );
nand ( n385308 , n385306 , n385307 );
buf ( n385309 , n385308 );
buf ( n385310 , n385309 );
nand ( n64645 , n64639 , n385310 );
buf ( n385312 , n64645 );
buf ( n385313 , n385312 );
not ( n385314 , n385313 );
buf ( n385315 , n372247 );
not ( n385316 , n385315 );
or ( n385317 , n385314 , n385316 );
buf ( n385318 , n40923 );
buf ( n385319 , n383042 );
nand ( n385320 , n385318 , n385319 );
buf ( n385321 , n385320 );
buf ( n385322 , n385321 );
nand ( n385323 , n385317 , n385322 );
buf ( n385324 , n385323 );
buf ( n385325 , n385324 );
xor ( n64660 , n383187 , n383191 );
xor ( n64661 , n64660 , n383277 );
buf ( n385328 , n64661 );
buf ( n64663 , n385328 );
xor ( n64664 , n385325 , n64663 );
buf ( n385331 , n377353 );
buf ( n385332 , n361534 );
and ( n64667 , n385331 , n385332 );
not ( n385334 , n385331 );
buf ( n64669 , n369577 );
and ( n385336 , n385334 , n64669 );
nor ( n64671 , n64667 , n385336 );
buf ( n64672 , n64671 );
buf ( n385339 , n64672 );
not ( n64674 , n385339 );
buf ( n64675 , n64674 );
buf ( n385342 , n64675 );
not ( n64677 , n385342 );
buf ( n385344 , n361606 );
not ( n64679 , n385344 );
or ( n64680 , n64677 , n64679 );
buf ( n385347 , n383148 );
buf ( n385348 , n50987 );
nand ( n64683 , n385347 , n385348 );
buf ( n385350 , n64683 );
buf ( n385351 , n385350 );
nand ( n385352 , n64680 , n385351 );
buf ( n385353 , n385352 );
buf ( n385354 , n385353 );
and ( n64689 , n64664 , n385354 );
and ( n64690 , n385325 , n64663 );
or ( n385357 , n64689 , n64690 );
buf ( n385358 , n385357 );
buf ( n385359 , n385358 );
and ( n385360 , n64633 , n385359 );
and ( n385361 , n385285 , n385298 );
or ( n64696 , n385360 , n385361 );
buf ( n385363 , n64696 );
buf ( n64698 , n385363 );
buf ( n385365 , n58923 );
not ( n64700 , n385365 );
buf ( n385367 , n384701 );
not ( n64702 , n385367 );
or ( n385369 , n64700 , n64702 );
buf ( n385370 , n379371 );
not ( n385371 , n385370 );
buf ( n385372 , n42684 );
not ( n64707 , n385372 );
or ( n385374 , n385371 , n64707 );
buf ( n385375 , n40201 );
buf ( n385376 , n379380 );
nand ( n385377 , n385375 , n385376 );
buf ( n385378 , n385377 );
buf ( n385379 , n385378 );
nand ( n385380 , n385374 , n385379 );
buf ( n385381 , n385380 );
buf ( n385382 , n385381 );
buf ( n385383 , n58871 );
nand ( n385384 , n385382 , n385383 );
buf ( n385385 , n385384 );
buf ( n385386 , n385385 );
nand ( n64721 , n385369 , n385386 );
buf ( n385388 , n64721 );
buf ( n385389 , n385388 );
xor ( n385390 , n64698 , n385389 );
buf ( n385391 , n380407 );
not ( n385392 , n385391 );
and ( n64727 , n380368 , n44925 );
not ( n64728 , n380368 );
and ( n385395 , n64728 , n359756 );
or ( n385396 , n64727 , n385395 );
buf ( n385397 , n385396 );
not ( n385398 , n385397 );
or ( n385399 , n385392 , n385398 );
buf ( n385400 , n384673 );
buf ( n385401 , n380356 );
nand ( n385402 , n385400 , n385401 );
buf ( n385403 , n385402 );
buf ( n385404 , n385403 );
nand ( n385405 , n385399 , n385404 );
buf ( n385406 , n385405 );
buf ( n385407 , n385406 );
and ( n64742 , n385390 , n385407 );
and ( n385409 , n64698 , n385389 );
or ( n64744 , n64742 , n385409 );
buf ( n385411 , n64744 );
buf ( n385412 , n385411 );
xor ( n64747 , n384684 , n384709 );
xor ( n64748 , n64747 , n384826 );
buf ( n385415 , n64748 );
buf ( n385416 , n385415 );
xor ( n64751 , n385412 , n385416 );
xor ( n385418 , n384723 , n384736 );
xor ( n64753 , n385418 , n384742 );
buf ( n385420 , n64753 );
buf ( n385421 , n385420 );
and ( n385422 , n383858 , n377580 );
and ( n64757 , n377585 , n363317 );
not ( n64758 , n377585 );
and ( n385425 , n64758 , n46031 );
or ( n64760 , n64757 , n385425 );
and ( n385427 , n64760 , n57530 );
nor ( n64762 , n385422 , n385427 );
buf ( n385429 , n64762 );
not ( n64764 , n385429 );
buf ( n385431 , n64764 );
buf ( n385432 , n385431 );
or ( n64767 , n385421 , n385432 );
and ( n64768 , n383136 , n383281 );
not ( n64769 , n383136 );
buf ( n385436 , n383281 );
not ( n64771 , n385436 );
buf ( n385438 , n64771 );
and ( n64773 , n64769 , n385438 );
nor ( n64774 , n64768 , n64773 );
and ( n385441 , n64774 , n383160 );
not ( n64776 , n64774 );
buf ( n385443 , n383160 );
not ( n64778 , n385443 );
buf ( n385445 , n64778 );
and ( n385446 , n64776 , n385445 );
nor ( n385447 , n385441 , n385446 );
buf ( n64782 , n385447 );
buf ( n385449 , n64782 );
nand ( n385450 , n64767 , n385449 );
buf ( n385451 , n385450 );
buf ( n385452 , n385451 );
buf ( n385453 , n385420 );
buf ( n385454 , n385431 );
nand ( n64789 , n385453 , n385454 );
buf ( n385456 , n64789 );
buf ( n385457 , n385456 );
nand ( n64792 , n385452 , n385457 );
buf ( n385459 , n64792 );
buf ( n385460 , n385459 );
not ( n64795 , n385460 );
buf ( n385462 , n58871 );
not ( n64797 , n385462 );
buf ( n385464 , n379371 );
not ( n64799 , n385464 );
buf ( n385466 , n363391 );
not ( n64801 , n385466 );
or ( n64802 , n64799 , n64801 );
buf ( n385469 , n366719 );
buf ( n385470 , n379380 );
nand ( n385471 , n385469 , n385470 );
buf ( n385472 , n385471 );
buf ( n385473 , n385472 );
nand ( n64808 , n64802 , n385473 );
buf ( n385475 , n64808 );
buf ( n385476 , n385475 );
not ( n64811 , n385476 );
or ( n385478 , n64797 , n64811 );
buf ( n385479 , n385381 );
buf ( n385480 , n58923 );
nand ( n385481 , n385479 , n385480 );
buf ( n385482 , n385481 );
buf ( n385483 , n385482 );
nand ( n64818 , n385478 , n385483 );
buf ( n385485 , n64818 );
buf ( n385486 , n385485 );
not ( n385487 , n385486 );
buf ( n385488 , n385487 );
not ( n64823 , n385488 );
buf ( n385490 , n379890 );
not ( n385491 , n385490 );
buf ( n385492 , n63966 );
not ( n385493 , n385492 );
or ( n64828 , n385491 , n385493 );
buf ( n385495 , n379841 );
not ( n385496 , n385495 );
buf ( n385497 , n362461 );
not ( n64832 , n385497 );
or ( n385499 , n385496 , n64832 );
not ( n385500 , n366673 );
nand ( n64835 , n385500 , n379847 );
buf ( n385502 , n64835 );
nand ( n385503 , n385499 , n385502 );
buf ( n385504 , n385503 );
buf ( n385505 , n385504 );
buf ( n385506 , n379916 );
nand ( n64841 , n385505 , n385506 );
buf ( n385508 , n64841 );
buf ( n385509 , n385508 );
nand ( n64844 , n64828 , n385509 );
buf ( n385511 , n64844 );
buf ( n385512 , n385511 );
not ( n385513 , n385512 );
buf ( n385514 , n385513 );
not ( n64849 , n385514 );
and ( n385516 , n64823 , n64849 );
buf ( n64851 , n385488 );
buf ( n64852 , n385514 );
nand ( n64853 , n64851 , n64852 );
buf ( n64854 , n64853 );
xor ( n64855 , n384765 , n384790 );
xor ( n385522 , n64855 , n384816 );
buf ( n385523 , n385522 );
and ( n385524 , n64854 , n385523 );
nor ( n64859 , n385516 , n385524 );
buf ( n385526 , n64859 );
not ( n64861 , n385526 );
buf ( n385528 , n64861 );
buf ( n385529 , n385528 );
not ( n64864 , n385529 );
or ( n64865 , n64795 , n64864 );
buf ( n385532 , n385459 );
not ( n385533 , n385532 );
buf ( n385534 , n385533 );
buf ( n385535 , n385534 );
not ( n385536 , n385535 );
buf ( n385537 , n64859 );
not ( n64872 , n385537 );
or ( n385539 , n385536 , n64872 );
xor ( n385540 , n384747 , n384751 );
xor ( n64875 , n385540 , n384821 );
buf ( n385542 , n64875 );
buf ( n385543 , n385542 );
nand ( n64878 , n385539 , n385543 );
buf ( n64879 , n64878 );
buf ( n385546 , n64879 );
nand ( n64881 , n64865 , n385546 );
buf ( n385548 , n64881 );
buf ( n385549 , n385548 );
and ( n64884 , n64751 , n385549 );
and ( n64885 , n385412 , n385416 );
or ( n64886 , n64884 , n64885 );
buf ( n385553 , n64886 );
buf ( n385554 , n383820 );
buf ( n385555 , n384830 );
xor ( n64890 , n385554 , n385555 );
buf ( n385557 , n64006 );
xor ( n385558 , n64890 , n385557 );
buf ( n385559 , n385558 );
or ( n385560 , n385553 , n385559 );
buf ( n385561 , n385560 );
xor ( n64896 , n383834 , n384594 );
xor ( n64897 , n64896 , n384643 );
buf ( n385564 , n64897 );
buf ( n385565 , n385564 );
not ( n385566 , n385565 );
buf ( n385567 , n385566 );
buf ( n385568 , n385567 );
not ( n64902 , n385568 );
not ( n385570 , n61822 );
not ( n385571 , n61853 );
not ( n64905 , n385571 );
or ( n385573 , n385570 , n64905 );
buf ( n385574 , n61853 );
buf ( n385575 , n382417 );
nand ( n385576 , n385574 , n385575 );
buf ( n385577 , n385576 );
nand ( n385578 , n385573 , n385577 );
buf ( n385579 , n61832 );
and ( n64913 , n385578 , n385579 );
not ( n64914 , n385578 );
not ( n64915 , n385579 );
and ( n385583 , n64914 , n64915 );
nor ( n385584 , n64913 , n385583 );
not ( n64918 , n385584 );
buf ( n385586 , n64918 );
not ( n64920 , n385586 );
or ( n64921 , n64902 , n64920 );
buf ( n385589 , n385564 );
not ( n64923 , n385589 );
buf ( n385591 , n385584 );
not ( n64925 , n385591 );
or ( n64926 , n64923 , n64925 );
buf ( n385594 , n383868 );
not ( n385595 , n385594 );
not ( n385596 , n63198 );
buf ( n385597 , n385596 );
not ( n385598 , n385597 );
or ( n385599 , n385595 , n385598 );
buf ( n385600 , n63198 );
buf ( n385601 , n63223 );
nand ( n385602 , n385600 , n385601 );
buf ( n385603 , n385602 );
buf ( n385604 , n385603 );
nand ( n385605 , n385599 , n385604 );
buf ( n385606 , n385605 );
buf ( n385607 , n385606 );
buf ( n385608 , n63944 );
and ( n385609 , n385607 , n385608 );
not ( n385610 , n385607 );
buf ( n385611 , n63944 );
not ( n385612 , n385611 );
buf ( n385613 , n385612 );
buf ( n385614 , n385613 );
and ( n385615 , n385610 , n385614 );
nor ( n385616 , n385609 , n385615 );
buf ( n385617 , n385616 );
buf ( n385618 , n385617 );
not ( n385619 , n385618 );
xor ( n64930 , n384636 , n384637 );
buf ( n385621 , n64930 );
buf ( n385622 , n385621 );
buf ( n385623 , n384633 );
and ( n64934 , n385622 , n385623 );
not ( n385625 , n385622 );
buf ( n385626 , n384633 );
not ( n64937 , n385626 );
buf ( n385628 , n64937 );
buf ( n385629 , n385628 );
and ( n64940 , n385625 , n385629 );
nor ( n385631 , n64934 , n64940 );
buf ( n385632 , n385631 );
buf ( n64943 , n385632 );
not ( n64944 , n64943 );
or ( n64945 , n385619 , n64944 );
buf ( n385636 , n385617 );
buf ( n385637 , n385632 );
or ( n64948 , n385636 , n385637 );
buf ( n385639 , n378856 );
not ( n385640 , n385639 );
buf ( n385641 , n365468 );
not ( n385642 , n385641 );
or ( n385643 , n385640 , n385642 );
buf ( n385644 , n362452 );
buf ( n385645 , n378847 );
nand ( n64956 , n385644 , n385645 );
buf ( n385647 , n64956 );
buf ( n385648 , n385647 );
nand ( n64959 , n385643 , n385648 );
buf ( n385650 , n64959 );
buf ( n385651 , n385650 );
not ( n64962 , n385651 );
buf ( n385653 , n40475 );
not ( n64964 , n385653 );
or ( n385655 , n64962 , n64964 );
buf ( n385656 , n384803 );
buf ( n385657 , n360574 );
nand ( n385658 , n385656 , n385657 );
buf ( n385659 , n385658 );
buf ( n385660 , n385659 );
nand ( n385661 , n385655 , n385660 );
buf ( n385662 , n385661 );
buf ( n385663 , n385662 );
not ( n385664 , n385663 );
buf ( n385665 , n57530 );
not ( n64976 , n385665 );
buf ( n385667 , n377585 );
buf ( n64978 , n41607 );
and ( n64979 , n385667 , n64978 );
not ( n385670 , n385667 );
buf ( n385671 , n44783 );
and ( n385672 , n385670 , n385671 );
nor ( n385673 , n64979 , n385672 );
buf ( n385674 , n385673 );
buf ( n385675 , n385674 );
not ( n64986 , n385675 );
or ( n385677 , n64976 , n64986 );
buf ( n64988 , n64760 );
buf ( n385679 , n377580 );
nand ( n385680 , n64988 , n385679 );
buf ( n385681 , n385680 );
buf ( n385682 , n385681 );
nand ( n64993 , n385677 , n385682 );
buf ( n385684 , n64993 );
buf ( n385685 , n385684 );
not ( n64996 , n385685 );
or ( n385687 , n385664 , n64996 );
buf ( n385688 , n385684 );
buf ( n385689 , n385662 );
or ( n385690 , n385688 , n385689 );
buf ( n385691 , n45075 );
not ( n65002 , n385691 );
buf ( n385693 , n385257 );
not ( n385694 , n385693 );
or ( n65005 , n65002 , n385694 );
and ( n385696 , n22930 , n351292 );
not ( n65007 , n22930 );
and ( n385698 , n65007 , n351291 );
or ( n65009 , n385696 , n385698 );
buf ( n385700 , n65009 );
buf ( n385701 , n365226 );
nand ( n65012 , n385700 , n385701 );
buf ( n385703 , n65012 );
buf ( n385704 , n385703 );
nand ( n65015 , n65005 , n385704 );
buf ( n385706 , n65015 );
buf ( n385707 , n385706 );
xor ( n65018 , n383953 , n63336 );
xor ( n385709 , n65018 , n384003 );
buf ( n385710 , n385709 );
buf ( n385711 , n385710 );
xor ( n385712 , n385707 , n385711 );
buf ( n385713 , n368665 );
not ( n65024 , n385713 );
buf ( n385715 , n342718 );
not ( n385716 , n385715 );
or ( n65027 , n65024 , n385716 );
buf ( n385718 , n55539 );
buf ( n385719 , n368662 );
nand ( n65030 , n385718 , n385719 );
buf ( n385721 , n65030 );
buf ( n385722 , n385721 );
nand ( n65033 , n65027 , n385722 );
buf ( n65034 , n65033 );
buf ( n385725 , n65034 );
not ( n65036 , n385725 );
buf ( n385727 , n363429 );
not ( n385728 , n385727 );
or ( n385729 , n65036 , n385728 );
buf ( n385730 , n363416 );
not ( n385731 , n385730 );
buf ( n385732 , n385211 );
nand ( n65043 , n385731 , n385732 );
buf ( n65044 , n65043 );
buf ( n385735 , n65044 );
nand ( n65046 , n385729 , n385735 );
buf ( n65047 , n65046 );
buf ( n385738 , n65047 );
and ( n65049 , n385712 , n385738 );
and ( n385740 , n385707 , n385711 );
or ( n65051 , n65049 , n385740 );
buf ( n385742 , n65051 );
buf ( n385743 , n385742 );
not ( n65054 , n63366 );
not ( n65055 , n384011 );
and ( n65056 , n65054 , n65055 );
and ( n65057 , n384011 , n63366 );
nor ( n65058 , n65056 , n65057 );
xnor ( n65059 , n65058 , n384574 );
buf ( n385750 , n65059 );
xor ( n65061 , n385743 , n385750 );
buf ( n385752 , n366317 );
buf ( n385753 , n56970 );
not ( n65064 , n385753 );
buf ( n385755 , n41772 );
not ( n385756 , n385755 );
or ( n65067 , n65064 , n385756 );
buf ( n385758 , n364744 );
buf ( n385759 , n377389 );
nand ( n385760 , n385758 , n385759 );
buf ( n385761 , n385760 );
buf ( n385762 , n385761 );
nand ( n65073 , n65067 , n385762 );
buf ( n385764 , n65073 );
buf ( n385765 , n385764 );
not ( n65076 , n385765 );
buf ( n385767 , n65076 );
buf ( n385768 , n385767 );
or ( n385769 , n385752 , n385768 );
buf ( n385770 , n383925 );
not ( n385771 , n385770 );
buf ( n385772 , n385771 );
buf ( n385773 , n385772 );
buf ( n385774 , n41836 );
or ( n385775 , n385773 , n385774 );
nand ( n65086 , n385769 , n385775 );
buf ( n385777 , n65086 );
buf ( n385778 , n385777 );
and ( n65089 , n65061 , n385778 );
and ( n385780 , n385743 , n385750 );
or ( n385781 , n65089 , n385780 );
buf ( n385782 , n385781 );
buf ( n385783 , n385782 );
nand ( n385784 , n385690 , n385783 );
buf ( n385785 , n385784 );
buf ( n385786 , n385785 );
nand ( n65097 , n385687 , n385786 );
buf ( n385788 , n65097 );
buf ( n385789 , n385788 );
not ( n65100 , n385789 );
not ( n65101 , n383312 );
not ( n385792 , n65101 );
not ( n385793 , n379445 );
and ( n65104 , n385792 , n385793 );
buf ( n385795 , n379274 );
not ( n385796 , n385795 );
buf ( n385797 , n370566 );
not ( n65108 , n385797 );
or ( n65109 , n385796 , n65108 );
buf ( n385800 , n362285 );
buf ( n385801 , n379271 );
nand ( n385802 , n385800 , n385801 );
buf ( n385803 , n385802 );
buf ( n385804 , n385803 );
nand ( n385805 , n65109 , n385804 );
buf ( n385806 , n385805 );
buf ( n65117 , n379293 );
and ( n385808 , n385806 , n65117 );
nor ( n385809 , n65104 , n385808 );
buf ( n385810 , n385809 );
not ( n385811 , n385810 );
buf ( n385812 , n385811 );
buf ( n385813 , n385812 );
not ( n65124 , n385813 );
or ( n385815 , n65100 , n65124 );
buf ( n385816 , n385788 );
not ( n385817 , n385816 );
buf ( n385818 , n385817 );
buf ( n65129 , n385818 );
not ( n65130 , n65129 );
buf ( n65131 , n385809 );
not ( n65132 , n65131 );
or ( n65133 , n65130 , n65132 );
xor ( n385824 , n385201 , n385276 );
xor ( n385825 , n385824 , n385280 );
buf ( n385826 , n385825 );
buf ( n385827 , n385826 );
buf ( n385828 , n366103 );
buf ( n385829 , n64672 );
and ( n385830 , n385828 , n385829 );
not ( n65141 , n385828 );
buf ( n385832 , n377782 );
not ( n65143 , n385832 );
buf ( n385834 , n44717 );
not ( n385835 , n385834 );
or ( n65146 , n65143 , n385835 );
buf ( n385837 , n361531 );
buf ( n385838 , n377779 );
nand ( n385839 , n385837 , n385838 );
buf ( n385840 , n385839 );
buf ( n385841 , n385840 );
nand ( n385842 , n65146 , n385841 );
buf ( n385843 , n385842 );
buf ( n385844 , n385843 );
buf ( n385845 , n59764 );
nand ( n385846 , n385844 , n385845 );
buf ( n385847 , n385846 );
buf ( n385848 , n385847 );
and ( n65159 , n65141 , n385848 );
nor ( n385850 , n385830 , n65159 );
buf ( n385851 , n385850 );
buf ( n385852 , n385851 );
not ( n385853 , n385852 );
buf ( n385854 , n62835 );
buf ( n385855 , n368621 );
and ( n65166 , n385854 , n385855 );
and ( n65167 , n380424 , n351762 );
not ( n65168 , n380424 );
and ( n65169 , n65168 , n48496 );
or ( n65170 , n65167 , n65169 );
buf ( n385861 , n65170 );
not ( n65172 , n385861 );
buf ( n385863 , n368605 );
nor ( n65174 , n65172 , n385863 );
buf ( n385865 , n65174 );
buf ( n385866 , n385865 );
nor ( n385867 , n65166 , n385866 );
buf ( n385868 , n385867 );
buf ( n385869 , n385868 );
not ( n385870 , n385869 );
buf ( n385871 , n385870 );
buf ( n65182 , n385871 );
not ( n65183 , n65182 );
or ( n65184 , n385853 , n65183 );
buf ( n385875 , n385312 );
not ( n65186 , n385875 );
buf ( n385877 , n65186 );
or ( n65188 , n370050 , n385877 );
not ( n385879 , n370060 );
and ( n385880 , n379482 , n61332 );
not ( n65191 , n379482 );
and ( n385882 , n65191 , n45116 );
or ( n65193 , n385880 , n385882 );
nand ( n385884 , n385879 , n65193 );
nand ( n65195 , n65188 , n385884 );
buf ( n385886 , n65195 );
buf ( n385887 , n385851 );
not ( n65198 , n385887 );
buf ( n65199 , n65198 );
buf ( n65200 , n65199 );
buf ( n385891 , n385868 );
nand ( n385892 , n65200 , n385891 );
buf ( n385893 , n385892 );
buf ( n385894 , n385893 );
nand ( n385895 , n385886 , n385894 );
buf ( n385896 , n385895 );
buf ( n385897 , n385896 );
nand ( n385898 , n65184 , n385897 );
buf ( n385899 , n385898 );
buf ( n385900 , n385899 );
xor ( n65211 , n385827 , n385900 );
buf ( n385902 , n377143 );
not ( n65213 , n385902 );
buf ( n385904 , n44634 );
not ( n385905 , n385904 );
or ( n385906 , n65213 , n385905 );
buf ( n385907 , n41892 );
buf ( n385908 , n377146 );
nand ( n385909 , n385907 , n385908 );
buf ( n385910 , n385909 );
buf ( n385911 , n385910 );
nand ( n385912 , n385906 , n385911 );
buf ( n385913 , n385912 );
buf ( n385914 , n385913 );
not ( n65225 , n385914 );
buf ( n385916 , n366046 );
not ( n65227 , n385916 );
or ( n65228 , n65225 , n65227 );
buf ( n385919 , n371063 );
buf ( n385920 , n383438 );
nand ( n385921 , n385919 , n385920 );
buf ( n385922 , n385921 );
buf ( n385923 , n385922 );
nand ( n65234 , n65228 , n385923 );
buf ( n385925 , n65234 );
not ( n65236 , n385925 );
buf ( n385927 , n359296 );
not ( n65238 , n385927 );
buf ( n385929 , n362452 );
not ( n65240 , n385929 );
or ( n65241 , n65238 , n65240 );
buf ( n385932 , n366360 );
nand ( n385933 , n65241 , n385932 );
buf ( n385934 , n385933 );
buf ( n385935 , n385934 );
not ( n65246 , n385935 );
buf ( n385937 , n362452 );
buf ( n385938 , n359296 );
or ( n65249 , n385937 , n385938 );
buf ( n385940 , n378098 );
nand ( n65251 , n65249 , n385940 );
buf ( n385942 , n65251 );
buf ( n385943 , n385942 );
nand ( n385944 , n65246 , n385943 );
buf ( n385945 , n385944 );
buf ( n385946 , n385945 );
not ( n385947 , n385946 );
buf ( n385948 , n385947 );
not ( n385949 , n385948 );
or ( n385950 , n65236 , n385949 );
buf ( n385951 , n385925 );
buf ( n385952 , n385948 );
nor ( n65263 , n385951 , n385952 );
buf ( n385954 , n65263 );
buf ( n385955 , n366708 );
not ( n65266 , n385955 );
buf ( n385957 , n342617 );
not ( n65268 , n385957 );
buf ( n385959 , n60751 );
not ( n385960 , n385959 );
and ( n65271 , n65268 , n385960 );
buf ( n385962 , n375914 );
buf ( n385963 , n60751 );
and ( n385964 , n385962 , n385963 );
nor ( n65275 , n65271 , n385964 );
buf ( n385966 , n65275 );
buf ( n385967 , n385966 );
not ( n385968 , n385967 );
and ( n385969 , n65266 , n385968 );
not ( n65280 , n383995 );
nor ( n65281 , n65280 , n366650 );
buf ( n385972 , n65281 );
nor ( n385973 , n385969 , n385972 );
buf ( n385974 , n385973 );
buf ( n385975 , n385974 );
not ( n385976 , n385975 );
buf ( n385977 , n385976 );
buf ( n385978 , n385977 );
not ( n65289 , n385978 );
buf ( n385980 , n384535 );
not ( n385981 , n385980 );
buf ( n385982 , n365108 );
not ( n385983 , n385982 );
or ( n385984 , n385981 , n385983 );
buf ( n65295 , n364981 );
not ( n65296 , n65295 );
buf ( n65297 , n31194 );
not ( n65298 , n65297 );
or ( n65299 , n65296 , n65298 );
buf ( n385990 , n57233 );
buf ( n385991 , n62345 );
nand ( n65302 , n385990 , n385991 );
buf ( n385993 , n65302 );
buf ( n385994 , n385993 );
nand ( n65305 , n65299 , n385994 );
buf ( n385996 , n65305 );
buf ( n385997 , n385996 );
buf ( n385998 , n365024 );
nand ( n65309 , n385997 , n385998 );
buf ( n386000 , n65309 );
buf ( n386001 , n386000 );
nand ( n386002 , n385984 , n386001 );
buf ( n386003 , n386002 );
buf ( n386004 , n386003 );
not ( n386005 , n386004 );
or ( n386006 , n65289 , n386005 );
buf ( n386007 , n386003 );
buf ( n386008 , n385977 );
or ( n386009 , n386007 , n386008 );
xor ( n65320 , n384019 , n384492 );
xor ( n65321 , n65320 , n384513 );
buf ( n386012 , n65321 );
buf ( n386013 , n386012 );
nand ( n65324 , n386009 , n386013 );
buf ( n386015 , n65324 );
buf ( n386016 , n386015 );
nand ( n65327 , n386006 , n386016 );
buf ( n386018 , n65327 );
buf ( n386019 , n386018 );
not ( n386020 , n50782 );
xor ( n65331 , n58073 , n365408 );
not ( n65332 , n65331 );
and ( n65333 , n386020 , n65332 );
not ( n386024 , n384557 );
buf ( n386025 , n366428 );
not ( n65336 , n386025 );
buf ( n386027 , n65336 );
nor ( n386028 , n386024 , n386027 );
nor ( n386029 , n65333 , n386028 );
buf ( n386030 , n386029 );
not ( n386031 , n386030 );
buf ( n386032 , n386031 );
not ( n65343 , n386032 );
buf ( n386034 , n45075 );
not ( n386035 , n386034 );
buf ( n386036 , n65009 );
not ( n386037 , n386036 );
or ( n386038 , n386035 , n386037 );
buf ( n65349 , n342877 );
not ( n386040 , n65349 );
not ( n65351 , n386040 );
not ( n386042 , n65351 );
not ( n386043 , n32202 );
not ( n65354 , n386043 );
or ( n386045 , n386042 , n65354 );
or ( n65356 , n386043 , n65351 );
nand ( n386047 , n386045 , n65356 );
buf ( n386048 , n386047 );
buf ( n386049 , n365226 );
nand ( n65360 , n386048 , n386049 );
buf ( n386051 , n65360 );
buf ( n386052 , n386051 );
nand ( n65363 , n386038 , n386052 );
buf ( n386054 , n65363 );
not ( n65365 , n386054 );
or ( n65366 , n65343 , n65365 );
buf ( n386057 , n386054 );
not ( n386058 , n386057 );
buf ( n386059 , n386058 );
not ( n386060 , n386059 );
not ( n386061 , n386029 );
or ( n386062 , n386060 , n386061 );
xor ( n386063 , n382879 , n382882 );
xor ( n386064 , n386063 , n382886 );
xor ( n386065 , n63497 , n63844 );
xor ( n386066 , n386064 , n386065 );
buf ( n386067 , n386066 );
and ( n386068 , n352268 , n61903 );
not ( n386069 , n352268 );
and ( n386070 , n386069 , n22619 );
or ( n386071 , n386068 , n386070 );
buf ( n386072 , n386071 );
not ( n386073 , n386072 );
buf ( n386074 , n384501 );
not ( n386075 , n386074 );
or ( n386076 , n386073 , n386075 );
buf ( n386077 , n63864 );
buf ( n386078 , n56794 );
nand ( n386079 , n386077 , n386078 );
buf ( n386080 , n386079 );
buf ( n386081 , n386080 );
nand ( n386082 , n386076 , n386081 );
buf ( n386083 , n386082 );
buf ( n386084 , n386083 );
xor ( n386085 , n386067 , n386084 );
buf ( n386086 , n365108 );
not ( n386087 , n386086 );
buf ( n386088 , n385996 );
not ( n386089 , n386088 );
or ( n386090 , n386087 , n386089 );
not ( n386091 , n44853 );
buf ( n386092 , n386091 );
buf ( n386093 , n364975 );
buf ( n386094 , n386093 );
not ( n386095 , n386094 );
buf ( n386096 , n381220 );
not ( n65372 , n386096 );
or ( n386098 , n386095 , n65372 );
buf ( n386099 , n351195 );
buf ( n386100 , n364975 );
not ( n386101 , n386100 );
buf ( n386102 , n386101 );
buf ( n386103 , n386102 );
nand ( n386104 , n386099 , n386103 );
buf ( n386105 , n386104 );
buf ( n386106 , n386105 );
nand ( n65382 , n386098 , n386106 );
buf ( n386108 , n65382 );
buf ( n386109 , n386108 );
nand ( n65385 , n386092 , n386109 );
buf ( n386111 , n65385 );
buf ( n386112 , n386111 );
nand ( n386113 , n386090 , n386112 );
buf ( n386114 , n386113 );
buf ( n386115 , n386114 );
and ( n386116 , n386085 , n386115 );
and ( n65392 , n386067 , n386084 );
or ( n386118 , n386116 , n65392 );
buf ( n386119 , n386118 );
nand ( n386120 , n386062 , n386119 );
nand ( n65396 , n65366 , n386120 );
buf ( n386122 , n65396 );
xor ( n386123 , n386019 , n386122 );
buf ( n386124 , n369374 );
buf ( n386125 , n342335 );
and ( n386126 , n386124 , n386125 );
not ( n386127 , n386124 );
buf ( n386128 , n362417 );
and ( n386129 , n386127 , n386128 );
nor ( n386130 , n386126 , n386129 );
buf ( n386131 , n386130 );
buf ( n386132 , n386131 );
not ( n386133 , n386132 );
buf ( n386134 , n386133 );
buf ( n386135 , n386134 );
not ( n386136 , n386135 );
buf ( n386137 , n368706 );
not ( n65413 , n386137 );
or ( n386139 , n386136 , n65413 );
nand ( n65415 , n362386 , n385242 );
buf ( n386141 , n65415 );
nand ( n65417 , n386139 , n386141 );
buf ( n386143 , n65417 );
buf ( n386144 , n386143 );
and ( n65420 , n386123 , n386144 );
and ( n386146 , n386019 , n386122 );
or ( n386147 , n65420 , n386146 );
buf ( n386148 , n386147 );
buf ( n386149 , n386148 );
not ( n386150 , n386149 );
buf ( n386151 , n386150 );
or ( n386152 , n385954 , n386151 );
nand ( n65428 , n385950 , n386152 );
buf ( n386154 , n65428 );
and ( n65430 , n65211 , n386154 );
and ( n386156 , n385827 , n385900 );
or ( n65432 , n65430 , n386156 );
buf ( n386158 , n65432 );
buf ( n386159 , n386158 );
nand ( n65435 , n65133 , n386159 );
buf ( n386161 , n65435 );
buf ( n386162 , n386161 );
nand ( n386163 , n385815 , n386162 );
buf ( n386164 , n386163 );
buf ( n386165 , n386164 );
nand ( n386166 , n64948 , n386165 );
buf ( n386167 , n386166 );
buf ( n386168 , n386167 );
nand ( n386169 , n64945 , n386168 );
buf ( n386170 , n386169 );
buf ( n386171 , n386170 );
nand ( n65441 , n64926 , n386171 );
buf ( n386173 , n65441 );
buf ( n386174 , n386173 );
nand ( n65444 , n64921 , n386174 );
buf ( n386176 , n65444 );
buf ( n386177 , n386176 );
and ( n386178 , n385561 , n386177 );
buf ( n386179 , n385559 );
buf ( n386180 , n385553 );
and ( n386181 , n386179 , n386180 );
buf ( n386182 , n386181 );
buf ( n386183 , n386182 );
nor ( n386184 , n386178 , n386183 );
buf ( n386185 , n386184 );
buf ( n386186 , n386185 );
and ( n386187 , n64556 , n386186 );
and ( n386188 , n385190 , n385197 );
or ( n386189 , n386187 , n386188 );
buf ( n386190 , n386189 );
buf ( n386191 , n386190 );
not ( n386192 , n386191 );
buf ( n386193 , n386192 );
nand ( n386194 , n64541 , n386193 );
nand ( n386195 , n64537 , n386194 );
and ( n386196 , n64524 , n386195 );
not ( n65466 , n58923 );
buf ( n386198 , n379371 );
not ( n65468 , n386198 );
buf ( n386200 , n363439 );
not ( n386201 , n386200 );
or ( n386202 , n65468 , n386201 );
nand ( n65472 , n64289 , n39046 , n379380 );
buf ( n386204 , n65472 );
nand ( n386205 , n386202 , n386204 );
buf ( n386206 , n386205 );
not ( n386207 , n386206 );
or ( n386208 , n65466 , n386207 );
nand ( n65478 , n379928 , n58871 );
nand ( n386210 , n386208 , n65478 );
buf ( n386211 , n379299 );
not ( n65481 , n386211 );
buf ( n386213 , n59468 );
not ( n386214 , n386213 );
or ( n65484 , n65481 , n386214 );
buf ( n386216 , n379274 );
not ( n386217 , n386216 );
buf ( n386218 , n365206 );
not ( n386219 , n386218 );
or ( n386220 , n386217 , n386219 );
buf ( n386221 , n39830 );
buf ( n386222 , n379271 );
nand ( n386223 , n386221 , n386222 );
buf ( n386224 , n386223 );
buf ( n386225 , n386224 );
nand ( n65495 , n386220 , n386225 );
buf ( n386227 , n65495 );
buf ( n386228 , n386227 );
buf ( n386229 , n379944 );
nand ( n386230 , n386228 , n386229 );
buf ( n386231 , n386230 );
buf ( n386232 , n386231 );
nand ( n386233 , n65484 , n386232 );
buf ( n386234 , n386233 );
xor ( n386235 , n386210 , n386234 );
xor ( n386236 , n380199 , n380214 );
and ( n65506 , n386236 , n380223 );
and ( n386238 , n380199 , n380214 );
or ( n65508 , n65506 , n386238 );
buf ( n386240 , n65508 );
xnor ( n65510 , n386235 , n386240 );
not ( n386242 , n377566 );
not ( n65512 , n57350 );
or ( n386244 , n386242 , n65512 );
buf ( n386245 , n377566 );
not ( n65515 , n386245 );
buf ( n386247 , n65515 );
not ( n65517 , n386247 );
not ( n386249 , n377800 );
or ( n386250 , n65517 , n386249 );
nand ( n65520 , n386250 , n57012 );
nand ( n65521 , n386244 , n65520 );
xor ( n65522 , n65510 , n65521 );
xor ( n65523 , n377449 , n377475 );
and ( n65524 , n65523 , n377506 );
and ( n65525 , n377449 , n377475 );
or ( n65526 , n65524 , n65525 );
buf ( n386258 , n65526 );
xor ( n65528 , n377514 , n377533 );
and ( n65529 , n65528 , n377555 );
and ( n386261 , n377514 , n377533 );
or ( n65531 , n65529 , n386261 );
xor ( n386263 , n386258 , n65531 );
buf ( n386264 , n378714 );
buf ( n386265 , n377181 );
or ( n65535 , n386264 , n386265 );
buf ( n386267 , n65535 );
buf ( n386268 , n386267 );
not ( n65538 , n386268 );
buf ( n386270 , n58289 );
not ( n65540 , n386270 );
or ( n386272 , n65538 , n65540 );
buf ( n65542 , n378714 );
buf ( n386274 , n377181 );
nand ( n386275 , n65542 , n386274 );
buf ( n386276 , n386275 );
buf ( n386277 , n386276 );
nand ( n386278 , n386272 , n386277 );
buf ( n386279 , n386278 );
and ( n386280 , n365393 , n64636 );
not ( n386281 , n365393 );
and ( n65551 , n386281 , n365266 );
or ( n65552 , n386280 , n65551 );
not ( n65553 , n65552 );
not ( n386285 , n40923 );
or ( n386286 , n65553 , n386285 );
nand ( n65556 , n365279 , n377499 );
nand ( n386288 , n386286 , n65556 );
xor ( n386289 , n386279 , n386288 );
buf ( n386290 , n58426 );
not ( n386291 , n386290 );
buf ( n386292 , n45345 );
not ( n386293 , n386292 );
or ( n386294 , n386291 , n386293 );
buf ( n386295 , n377782 );
not ( n386296 , n386295 );
buf ( n386297 , n363122 );
not ( n386298 , n386297 );
or ( n386299 , n386296 , n386298 );
buf ( n386300 , n365528 );
buf ( n386301 , n377779 );
nand ( n386302 , n386300 , n386301 );
buf ( n386303 , n386302 );
buf ( n386304 , n386303 );
nand ( n386305 , n386299 , n386304 );
buf ( n386306 , n386305 );
buf ( n386307 , n386306 );
buf ( n386308 , n365486 );
nand ( n386309 , n386307 , n386308 );
buf ( n65557 , n386309 );
buf ( n386311 , n65557 );
nand ( n386312 , n386294 , n386311 );
buf ( n386313 , n386312 );
xor ( n386314 , n386289 , n386313 );
xnor ( n386315 , n386263 , n386314 );
not ( n386316 , n386315 );
xor ( n65559 , n377509 , n377557 );
and ( n386318 , n65559 , n377564 );
and ( n386319 , n377509 , n377557 );
or ( n65562 , n386318 , n386319 );
buf ( n386321 , n65562 );
not ( n65564 , n386321 );
buf ( n65565 , n45018 );
buf ( n386324 , n65565 );
not ( n386325 , n386324 );
buf ( n386326 , n379050 );
not ( n386327 , n386326 );
or ( n386328 , n386325 , n386327 );
buf ( n386329 , n46397 );
not ( n65572 , n386329 );
buf ( n386331 , n363317 );
not ( n65574 , n386331 );
or ( n65575 , n65572 , n65574 );
buf ( n386334 , n342909 );
buf ( n386335 , n367459 );
nand ( n65578 , n386334 , n386335 );
buf ( n386337 , n65578 );
buf ( n386338 , n386337 );
nand ( n386339 , n65575 , n386338 );
buf ( n386340 , n386339 );
buf ( n386341 , n386340 );
buf ( n386342 , n365152 );
nand ( n386343 , n386341 , n386342 );
buf ( n386344 , n386343 );
buf ( n386345 , n386344 );
nand ( n386346 , n386328 , n386345 );
buf ( n386347 , n386346 );
not ( n65590 , n386347 );
buf ( n386349 , n58244 );
not ( n386350 , n386349 );
buf ( n386351 , n363429 );
not ( n65594 , n386351 );
or ( n386353 , n386350 , n65594 );
not ( n386354 , n57688 );
buf ( n386355 , n386354 );
not ( n386356 , n386355 );
buf ( n386357 , n352209 );
not ( n386358 , n386357 );
buf ( n386359 , n386358 );
buf ( n386360 , n386359 );
not ( n386361 , n386360 );
or ( n386362 , n386356 , n386361 );
buf ( n386363 , n46693 );
not ( n386364 , n386363 );
buf ( n386365 , n352209 );
nand ( n386366 , n386364 , n386365 );
buf ( n386367 , n386366 );
buf ( n386368 , n386367 );
nand ( n386369 , n386362 , n386368 );
buf ( n386370 , n386369 );
buf ( n386371 , n386370 );
buf ( n386372 , n378183 );
nand ( n386373 , n386371 , n386372 );
buf ( n386374 , n386373 );
buf ( n386375 , n386374 );
nand ( n386376 , n386353 , n386375 );
buf ( n386377 , n386376 );
buf ( n386378 , n386377 );
not ( n386379 , n386378 );
buf ( n386380 , n386379 );
buf ( n386381 , n386380 );
not ( n386382 , n56794 );
buf ( n386383 , n22619 );
not ( n65613 , n386383 );
buf ( n386385 , n366187 );
not ( n386386 , n386385 );
or ( n386387 , n65613 , n386386 );
buf ( n386388 , n366187 );
not ( n386389 , n386388 );
buf ( n386390 , n386389 );
buf ( n386391 , n386390 );
buf ( n386392 , n365670 );
nand ( n65619 , n386391 , n386392 );
buf ( n386394 , n65619 );
buf ( n65621 , n386394 );
nand ( n65622 , n386387 , n65621 );
buf ( n65623 , n65622 );
not ( n386398 , n65623 );
or ( n65625 , n386382 , n386398 );
nand ( n386400 , n45553 , n378987 );
nand ( n386401 , n65625 , n386400 );
buf ( n386402 , n386401 );
xor ( n386403 , n386381 , n386402 );
buf ( n386404 , n366317 );
buf ( n386405 , n377433 );
or ( n65632 , n386404 , n386405 );
buf ( n386407 , n31197 );
not ( n386408 , n386407 );
buf ( n386409 , n41772 );
not ( n386410 , n386409 );
or ( n386411 , n386408 , n386410 );
buf ( n386412 , n366329 );
buf ( n386413 , n351229 );
nand ( n386414 , n386412 , n386413 );
buf ( n386415 , n386414 );
buf ( n386416 , n386415 );
nand ( n65643 , n386411 , n386416 );
buf ( n386418 , n65643 );
buf ( n386419 , n386418 );
not ( n65646 , n386419 );
buf ( n386421 , n65646 );
buf ( n386422 , n386421 );
buf ( n386423 , n49692 );
or ( n65650 , n386422 , n386423 );
nand ( n386425 , n65632 , n65650 );
buf ( n386426 , n386425 );
buf ( n386427 , n386426 );
xor ( n65654 , n386403 , n386427 );
buf ( n386429 , n65654 );
buf ( n386430 , n386429 );
not ( n65657 , n386430 );
buf ( n65658 , n65657 );
not ( n65659 , n65658 );
or ( n386434 , n65590 , n65659 );
buf ( n386435 , n386347 );
not ( n65662 , n386435 );
buf ( n386437 , n386429 );
nand ( n386438 , n65662 , n386437 );
buf ( n386439 , n386438 );
nand ( n65666 , n386434 , n386439 );
buf ( n386441 , n380065 );
not ( n65668 , n386441 );
buf ( n386443 , n359913 );
not ( n65670 , n386443 );
buf ( n386445 , n65670 );
buf ( n386446 , n386445 );
not ( n386447 , n386446 );
or ( n65674 , n65668 , n386447 );
buf ( n386449 , n368038 );
buf ( n386450 , n377143 );
not ( n65677 , n386450 );
buf ( n386452 , n42455 );
not ( n386453 , n386452 );
or ( n65680 , n65677 , n386453 );
buf ( n386455 , n364922 );
buf ( n386456 , n377153 );
nand ( n65683 , n386455 , n386456 );
buf ( n386458 , n65683 );
buf ( n386459 , n386458 );
nand ( n65686 , n65680 , n386459 );
buf ( n386461 , n65686 );
buf ( n386462 , n386461 );
nand ( n386463 , n386449 , n386462 );
buf ( n386464 , n386463 );
buf ( n386465 , n386464 );
nand ( n386466 , n65674 , n386465 );
buf ( n386467 , n386466 );
and ( n65694 , n65666 , n386467 );
not ( n386469 , n65666 );
not ( n386470 , n386467 );
and ( n65697 , n386469 , n386470 );
nor ( n386472 , n65694 , n65697 );
not ( n386473 , n386472 );
or ( n386474 , n65564 , n386473 );
not ( n65701 , n386472 );
not ( n386476 , n386321 );
nand ( n386477 , n65701 , n386476 );
nand ( n65704 , n386474 , n386477 );
not ( n386479 , n65704 );
not ( n386480 , n386479 );
or ( n65707 , n386316 , n386480 );
not ( n386482 , n386315 );
nand ( n65709 , n65704 , n386482 );
nand ( n65710 , n65707 , n65709 );
xnor ( n65711 , n65522 , n65710 );
buf ( n386486 , n378669 );
not ( n65713 , n386486 );
buf ( n386488 , n377803 );
not ( n65715 , n386488 );
or ( n65716 , n65713 , n65715 );
buf ( n386491 , n379433 );
nand ( n65718 , n65716 , n386491 );
buf ( n386493 , n65718 );
buf ( n386494 , n386493 );
not ( n65721 , n377803 );
nand ( n386496 , n65721 , n378668 );
buf ( n386497 , n386496 );
nand ( n65724 , n386494 , n386497 );
buf ( n386499 , n65724 );
xor ( n65726 , n65711 , n386499 );
not ( n386501 , n378814 );
nand ( n65728 , n378694 , n58434 );
not ( n65729 , n65728 );
or ( n386504 , n386501 , n65729 );
nand ( n386505 , n58435 , n378691 );
nand ( n386506 , n386504 , n386505 );
buf ( n386507 , n386506 );
buf ( n386508 , n369444 );
not ( n386509 , n386508 );
buf ( n386510 , n368549 );
not ( n386511 , n386510 );
buf ( n386512 , n360848 );
not ( n386513 , n386512 );
or ( n386514 , n386511 , n386513 );
buf ( n386515 , n362458 );
buf ( n386516 , n368554 );
nand ( n386517 , n386515 , n386516 );
buf ( n386518 , n386517 );
buf ( n386519 , n386518 );
nand ( n386520 , n386514 , n386519 );
buf ( n386521 , n386520 );
buf ( n386522 , n386521 );
not ( n386523 , n386522 );
or ( n386524 , n386509 , n386523 );
nand ( n386525 , n378684 , n368611 );
buf ( n386526 , n386525 );
nand ( n386527 , n386524 , n386526 );
buf ( n386528 , n386527 );
buf ( n386529 , n386528 );
not ( n386530 , n58322 );
not ( n386531 , n58344 );
not ( n65738 , n386531 );
or ( n65739 , n386530 , n65738 );
buf ( n386534 , n58294 );
not ( n386535 , n386534 );
buf ( n386536 , n386535 );
nand ( n65743 , n65739 , n386536 );
nand ( n65744 , n58344 , n58319 );
nand ( n65745 , n65743 , n65744 );
buf ( n386540 , n65745 );
xor ( n386541 , n386529 , n386540 );
buf ( n386542 , n378868 );
not ( n386543 , n386542 );
buf ( n386544 , n378899 );
not ( n386545 , n386544 );
or ( n386546 , n386543 , n386545 );
buf ( n386547 , n378899 );
buf ( n386548 , n378868 );
or ( n386549 , n386547 , n386548 );
buf ( n386550 , n378831 );
nand ( n65757 , n386549 , n386550 );
buf ( n386552 , n65757 );
buf ( n386553 , n386552 );
nand ( n65760 , n386546 , n386553 );
buf ( n386555 , n65760 );
buf ( n386556 , n386555 );
xor ( n386557 , n386541 , n386556 );
buf ( n386558 , n386557 );
buf ( n386559 , n386558 );
xor ( n386560 , n386507 , n386559 );
buf ( n386561 , n386560 );
buf ( n386562 , n386561 );
xor ( n65769 , n378922 , n378947 );
and ( n65770 , n65769 , n379060 );
and ( n386565 , n378922 , n378947 );
or ( n65772 , n65770 , n386565 );
buf ( n386567 , n65772 );
buf ( n386568 , n386567 );
not ( n386569 , n386568 );
buf ( n386570 , n386569 );
buf ( n386571 , n386570 );
and ( n386572 , n386562 , n386571 );
not ( n386573 , n386562 );
buf ( n386574 , n386567 );
and ( n386575 , n386573 , n386574 );
nor ( n386576 , n386572 , n386575 );
buf ( n386577 , n386576 );
buf ( n386578 , n378904 );
not ( n386579 , n386578 );
buf ( n65773 , n379062 );
not ( n65774 , n65773 );
buf ( n386582 , n65774 );
buf ( n386583 , n386582 );
nand ( n386584 , n386579 , n386583 );
buf ( n386585 , n386584 );
buf ( n386586 , n386585 );
buf ( n386587 , n58934 );
and ( n65781 , n386586 , n386587 );
and ( n386589 , n378905 , n379063 );
buf ( n386590 , n386589 );
buf ( n386591 , n386590 );
nor ( n386592 , n65781 , n386591 );
buf ( n386593 , n386592 );
xor ( n65783 , n386577 , n386593 );
buf ( n386595 , n44915 );
not ( n65785 , n386595 );
buf ( n386597 , n365041 );
not ( n65787 , n386597 );
buf ( n386599 , n370566 );
not ( n65789 , n386599 );
or ( n65790 , n65787 , n65789 );
buf ( n386602 , n362285 );
buf ( n386603 , n365052 );
nand ( n65793 , n386602 , n386603 );
buf ( n386605 , n65793 );
buf ( n386606 , n386605 );
nand ( n65796 , n65790 , n386606 );
buf ( n386608 , n65796 );
buf ( n386609 , n386608 );
not ( n65799 , n386609 );
or ( n65800 , n65785 , n65799 );
buf ( n386612 , n59677 );
buf ( n386613 , n47466 );
nand ( n65803 , n386612 , n386613 );
buf ( n386615 , n65803 );
buf ( n386616 , n386615 );
nand ( n65806 , n65800 , n386616 );
buf ( n386618 , n65806 );
buf ( n386619 , n386618 );
buf ( n386620 , n379056 );
not ( n65810 , n386620 );
buf ( n386622 , n58547 );
not ( n65812 , n386622 );
or ( n65813 , n65810 , n65812 );
buf ( n386625 , n379053 );
not ( n65815 , n386625 );
buf ( n386627 , n58547 );
not ( n386628 , n386627 );
buf ( n386629 , n386628 );
buf ( n386630 , n386629 );
not ( n65820 , n386630 );
or ( n386632 , n65815 , n65820 );
buf ( n386633 , n58528 );
buf ( n65823 , n386633 );
buf ( n386635 , n65823 );
buf ( n386636 , n386635 );
nand ( n65826 , n386632 , n386636 );
buf ( n386638 , n65826 );
buf ( n386639 , n386638 );
nand ( n386640 , n65813 , n386639 );
buf ( n386641 , n386640 );
buf ( n386642 , n386641 );
xor ( n386643 , n386619 , n386642 );
buf ( n386644 , n49609 );
not ( n65834 , n386644 );
buf ( n386646 , n369769 );
not ( n65836 , n386646 );
buf ( n386648 , n47193 );
not ( n386649 , n386648 );
or ( n65839 , n65836 , n386649 );
buf ( n386651 , n369766 );
buf ( n386652 , n40275 );
nand ( n65842 , n386651 , n386652 );
buf ( n386654 , n65842 );
buf ( n386655 , n386654 );
nand ( n65844 , n65839 , n386655 );
buf ( n386657 , n65844 );
buf ( n386658 , n386657 );
not ( n65847 , n386658 );
or ( n65848 , n65834 , n65847 );
buf ( n386661 , n378911 );
buf ( n386662 , n369804 );
nand ( n386663 , n386661 , n386662 );
buf ( n386664 , n386663 );
buf ( n386665 , n386664 );
nand ( n386666 , n65848 , n386665 );
buf ( n386667 , n386666 );
buf ( n386668 , n386667 );
xor ( n386669 , n386643 , n386668 );
buf ( n386670 , n386669 );
buf ( n386671 , n377452 );
not ( n386672 , n386671 );
buf ( n386673 , n386672 );
buf ( n386674 , n386673 );
not ( n386675 , n386674 );
buf ( n386676 , n41882 );
not ( n386677 , n386676 );
buf ( n386678 , n386677 );
buf ( n386679 , n386678 );
not ( n65865 , n386679 );
or ( n65866 , n386675 , n65865 );
not ( n65867 , n365980 );
not ( n65868 , n361009 );
or ( n65869 , n65867 , n65868 );
buf ( n386685 , n362033 );
buf ( n386686 , n365989 );
nand ( n65872 , n386685 , n386686 );
buf ( n386688 , n65872 );
nand ( n65874 , n65869 , n386688 );
nand ( n65875 , n365622 , n65874 );
buf ( n386691 , n65875 );
nand ( n65877 , n65866 , n386691 );
buf ( n386693 , n65877 );
buf ( n65879 , n386693 );
buf ( n386695 , n365115 );
not ( n65881 , n386695 );
buf ( n386697 , n364981 );
not ( n65883 , n386697 );
buf ( n386699 , n362534 );
not ( n386700 , n386699 );
buf ( n386701 , n386700 );
buf ( n386702 , n386701 );
not ( n65888 , n386702 );
or ( n65889 , n65883 , n65888 );
buf ( n65890 , n362537 );
not ( n386706 , n65890 );
buf ( n386707 , n386706 );
buf ( n386708 , n386707 );
buf ( n386709 , n364978 );
nand ( n65895 , n386708 , n386709 );
buf ( n386711 , n65895 );
buf ( n386712 , n386711 );
nand ( n65898 , n65889 , n386712 );
buf ( n386714 , n65898 );
buf ( n386715 , n386714 );
not ( n65901 , n386715 );
or ( n65902 , n65881 , n65901 );
nand ( n65903 , n365033 , n377523 );
buf ( n386719 , n65903 );
nand ( n65905 , n65902 , n386719 );
buf ( n386721 , n65905 );
buf ( n386722 , n386721 );
xor ( n65908 , n65879 , n386722 );
buf ( n386724 , n57107 );
not ( n386725 , n386724 );
buf ( n386726 , n361606 );
not ( n65912 , n386726 );
or ( n65913 , n386725 , n65912 );
buf ( n386729 , n351160 );
not ( n65915 , n386729 );
buf ( n386731 , n361534 );
not ( n386732 , n386731 );
or ( n386733 , n65915 , n386732 );
buf ( n386734 , n361531 );
buf ( n386735 , n364915 );
nand ( n65921 , n386734 , n386735 );
buf ( n386737 , n65921 );
buf ( n386738 , n386737 );
nand ( n65924 , n386733 , n386738 );
buf ( n386740 , n65924 );
buf ( n386741 , n386740 );
buf ( n386742 , n367590 );
nand ( n65928 , n386741 , n386742 );
buf ( n386744 , n65928 );
buf ( n386745 , n386744 );
nand ( n65931 , n65913 , n386745 );
buf ( n386747 , n65931 );
buf ( n386748 , n386747 );
xor ( n65934 , n65908 , n386748 );
buf ( n386750 , n65934 );
not ( n65936 , n379016 );
or ( n386752 , n378975 , n58502 );
not ( n65938 , n386752 );
or ( n65939 , n65936 , n65938 );
nand ( n386755 , n58502 , n378975 );
nand ( n65941 , n65939 , n386755 );
not ( n386757 , n65941 );
not ( n386758 , n386757 );
not ( n65944 , n45075 );
nand ( n65945 , n361664 , n342881 );
nand ( n386761 , n365757 , n365202 );
nand ( n386762 , n65945 , n386761 );
not ( n65948 , n386762 );
or ( n386764 , n65944 , n65948 );
nand ( n65950 , n378773 , n365226 );
nand ( n65951 , n386764 , n65950 );
not ( n386767 , n65951 );
not ( n65953 , n386767 );
or ( n386769 , n386758 , n65953 );
nand ( n386770 , n65941 , n65951 );
nand ( n65956 , n386769 , n386770 );
not ( n65957 , n378805 );
not ( n386773 , n377370 );
or ( n65959 , n65957 , n386773 );
buf ( n386775 , n368994 );
not ( n65961 , n386775 );
buf ( n386777 , n45270 );
not ( n386778 , n386777 );
or ( n386779 , n65961 , n386778 );
buf ( n386780 , n362452 );
buf ( n386781 , n57053 );
nand ( n65967 , n386780 , n386781 );
buf ( n65968 , n65967 );
buf ( n386784 , n65968 );
nand ( n65970 , n386779 , n386784 );
buf ( n386786 , n65970 );
buf ( n65972 , n386786 );
buf ( n386788 , n366751 );
nand ( n65974 , n65972 , n386788 );
buf ( n386790 , n65974 );
nand ( n65976 , n65959 , n386790 );
and ( n65977 , n65956 , n65976 );
not ( n386793 , n65956 );
not ( n386794 , n65976 );
and ( n65980 , n386793 , n386794 );
nor ( n386796 , n65977 , n65980 );
not ( n65982 , n386796 );
xor ( n386798 , n386750 , n65982 );
buf ( n386799 , n377271 );
not ( n65985 , n386799 );
buf ( n386801 , n342656 );
not ( n386802 , n386801 );
buf ( n386803 , n44637 );
not ( n65989 , n386803 );
or ( n65990 , n386802 , n65989 );
buf ( n386806 , n364808 );
buf ( n386807 , n58073 );
not ( n65993 , n386807 );
buf ( n386809 , n65993 );
nand ( n386810 , n386806 , n386809 );
buf ( n386811 , n386810 );
buf ( n386812 , n386811 );
nand ( n65998 , n65990 , n386812 );
buf ( n386814 , n65998 );
buf ( n386815 , n386814 );
not ( n66001 , n386815 );
or ( n66002 , n65985 , n66001 );
buf ( n386818 , n378963 );
buf ( n386819 , n366399 );
nand ( n386820 , n386818 , n386819 );
buf ( n386821 , n386820 );
buf ( n386822 , n386821 );
nand ( n66008 , n66002 , n386822 );
buf ( n386824 , n66008 );
not ( n66010 , n378748 );
not ( n66011 , n362405 );
or ( n66012 , n66010 , n66011 );
not ( n66013 , n362385 );
buf ( n386829 , n365440 );
not ( n386830 , n386829 );
buf ( n386831 , n342335 );
not ( n66017 , n386831 );
or ( n386833 , n386830 , n66017 );
buf ( n386834 , n362417 );
buf ( n386835 , n32202 );
not ( n66021 , n386835 );
buf ( n386837 , n66021 );
buf ( n386838 , n386837 );
nand ( n66024 , n386834 , n386838 );
buf ( n386840 , n66024 );
buf ( n386841 , n386840 );
nand ( n386842 , n386833 , n386841 );
buf ( n386843 , n386842 );
nand ( n66029 , n66013 , n386843 );
nand ( n66030 , n66012 , n66029 );
xor ( n66031 , n386824 , n66030 );
buf ( n386847 , n46521 );
not ( n386848 , n386847 );
buf ( n386849 , n379006 );
not ( n66035 , n386849 );
or ( n386851 , n386848 , n66035 );
buf ( n386852 , n46477 );
not ( n66038 , n386852 );
buf ( n386854 , n364855 );
not ( n66040 , n386854 );
or ( n386856 , n66038 , n66040 );
buf ( n386857 , n351367 );
buf ( n386858 , n46474 );
nand ( n66044 , n386857 , n386858 );
buf ( n66045 , n66044 );
buf ( n386861 , n66045 );
nand ( n66047 , n386856 , n386861 );
buf ( n386863 , n66047 );
buf ( n386864 , n386863 );
buf ( n386865 , n46463 );
nand ( n386866 , n386864 , n386865 );
buf ( n386867 , n386866 );
buf ( n386868 , n386867 );
nand ( n66054 , n386851 , n386868 );
buf ( n386870 , n66054 );
not ( n66056 , n386870 );
xor ( n386872 , n66031 , n66056 );
not ( n386873 , n379031 );
not ( n66059 , n367273 );
or ( n386875 , n386873 , n66059 );
and ( n386876 , n56970 , n35547 );
not ( n66062 , n56970 );
and ( n66063 , n66062 , n35548 );
nor ( n66064 , n386876 , n66063 );
buf ( n386880 , n66064 );
not ( n66066 , n386880 );
buf ( n66067 , n46582 );
nand ( n66068 , n66066 , n66067 );
buf ( n386884 , n66068 );
nand ( n66070 , n386875 , n386884 );
xor ( n386886 , n386872 , n66070 );
not ( n66072 , n378862 );
not ( n386888 , n359809 );
or ( n66074 , n66072 , n386888 );
not ( n66075 , n42373 );
not ( n66076 , n379482 );
not ( n386892 , n366534 );
or ( n66078 , n66076 , n386892 );
nand ( n386894 , n361631 , n58984 );
nand ( n66080 , n66078 , n386894 );
nand ( n66081 , n66075 , n66080 );
nand ( n386897 , n66074 , n66081 );
xor ( n66083 , n386886 , n386897 );
xor ( n386899 , n386798 , n66083 );
xor ( n386900 , n386670 , n386899 );
buf ( n386901 , n379851 );
not ( n386902 , n386901 );
buf ( n386903 , n59424 );
not ( n66089 , n386903 );
and ( n66090 , n386902 , n66089 );
buf ( n386906 , n379841 );
not ( n66092 , n386906 );
buf ( n386908 , n363866 );
not ( n66094 , n386908 );
or ( n66095 , n66092 , n66094 );
buf ( n386911 , n59860 );
not ( n66097 , n386911 );
buf ( n386913 , n379847 );
nand ( n66099 , n66097 , n386913 );
buf ( n386915 , n66099 );
buf ( n386916 , n386915 );
nand ( n66102 , n66095 , n386916 );
buf ( n386918 , n66102 );
buf ( n386919 , n386918 );
buf ( n386920 , n379890 );
and ( n386921 , n386919 , n386920 );
nor ( n66107 , n66090 , n386921 );
buf ( n386923 , n66107 );
buf ( n386924 , n386923 );
not ( n66110 , n386924 );
buf ( n386926 , n66110 );
not ( n386927 , n386926 );
not ( n66113 , n386927 );
xor ( n66114 , n59546 , n380071 );
and ( n66115 , n66114 , n380126 );
and ( n386931 , n59546 , n380071 );
or ( n66117 , n66115 , n386931 );
buf ( n386933 , n377580 );
not ( n386934 , n386933 );
buf ( n386935 , n377585 );
not ( n386936 , n386935 );
buf ( n386937 , n364987 );
not ( n66123 , n386937 );
or ( n66124 , n386936 , n66123 );
buf ( n386940 , n359778 );
buf ( n386941 , n377592 );
buf ( n386942 , n386941 );
buf ( n386943 , n386942 );
buf ( n386944 , n386943 );
nand ( n66130 , n386940 , n386944 );
buf ( n386946 , n66130 );
buf ( n386947 , n386946 );
nand ( n386948 , n66124 , n386947 );
buf ( n386949 , n386948 );
buf ( n386950 , n386949 );
not ( n66136 , n386950 );
or ( n66137 , n386934 , n66136 );
buf ( n386953 , n378936 );
buf ( n386954 , n57530 );
nand ( n66140 , n386953 , n386954 );
buf ( n386956 , n66140 );
buf ( n386957 , n386956 );
nand ( n66143 , n66137 , n386957 );
buf ( n386959 , n66143 );
and ( n66145 , n66117 , n386959 );
not ( n386961 , n66117 );
not ( n386962 , n386959 );
and ( n386963 , n386961 , n386962 );
nor ( n66149 , n66145 , n386963 );
not ( n386965 , n66149 );
not ( n386966 , n386965 );
or ( n66152 , n66113 , n386966 );
nand ( n66153 , n66149 , n386926 );
nand ( n386969 , n66152 , n66153 );
not ( n66155 , n386969 );
and ( n386971 , n386900 , n66155 );
not ( n66157 , n386900 );
and ( n66158 , n66157 , n386969 );
nor ( n386974 , n386971 , n66158 );
xor ( n386975 , n65783 , n386974 );
not ( n66161 , n386975 );
and ( n386977 , n65726 , n66161 );
not ( n386978 , n65726 );
buf ( n66164 , n386975 );
and ( n386980 , n386978 , n66164 );
nor ( n66166 , n386977 , n386980 );
not ( n66167 , n385038 );
not ( n66168 , n64453 );
or ( n66169 , n66167 , n66168 );
not ( n386985 , n385035 );
not ( n66171 , n385089 );
or ( n66172 , n386985 , n66171 );
nand ( n66173 , n66172 , n385011 );
nand ( n386989 , n66169 , n66173 );
buf ( n66175 , n386989 );
not ( n386991 , n59337 );
not ( n66177 , n379965 );
not ( n386993 , n66177 );
or ( n66179 , n386991 , n386993 );
not ( n66180 , n379965 );
not ( n386996 , n379829 );
or ( n386997 , n66180 , n386996 );
not ( n66183 , n59718 );
nand ( n386999 , n386997 , n66183 );
nand ( n387000 , n66179 , n386999 );
not ( n66186 , n387000 );
xor ( n387002 , n385050 , n64418 );
and ( n387003 , n387002 , n385087 );
and ( n66189 , n385050 , n64418 );
or ( n387005 , n387003 , n66189 );
buf ( n387006 , n387005 );
and ( n66192 , n66186 , n387006 );
not ( n387008 , n66186 );
not ( n387009 , n387006 );
and ( n66195 , n387008 , n387009 );
nor ( n387011 , n66192 , n66195 );
buf ( n387012 , n387011 );
not ( n66198 , n59475 );
not ( n387014 , n59446 );
nand ( n387015 , n387014 , n379920 );
not ( n387016 , n387015 );
or ( n66202 , n66198 , n387016 );
nand ( n387018 , n59432 , n59446 );
nand ( n66204 , n66202 , n387018 );
buf ( n387020 , n66204 );
not ( n66206 , n387020 );
buf ( n387022 , n66206 );
not ( n387023 , n387022 );
buf ( n387024 , n64427 );
not ( n387025 , n387024 );
buf ( n387026 , n64441 );
not ( n387027 , n387026 );
or ( n387028 , n387025 , n387027 );
buf ( n387029 , n64441 );
buf ( n387030 , n64427 );
or ( n387031 , n387029 , n387030 );
buf ( n387032 , n64435 );
nand ( n66218 , n387031 , n387032 );
buf ( n387034 , n66218 );
buf ( n387035 , n387034 );
nand ( n66221 , n387028 , n387035 );
buf ( n66222 , n66221 );
not ( n387038 , n66222 );
nor ( n66224 , n387023 , n387038 );
buf ( n387040 , n66204 );
not ( n387041 , n387040 );
not ( n66227 , n387038 );
or ( n387043 , n387041 , n66227 );
not ( n66229 , n59614 );
not ( n387045 , n66229 );
not ( n66231 , n59672 );
and ( n66232 , n387045 , n66231 );
nand ( n387048 , n66229 , n59672 );
and ( n387049 , n380225 , n387048 );
nor ( n66235 , n66232 , n387049 );
nand ( n387051 , n387043 , n66235 );
or ( n387052 , n66224 , n387051 );
not ( n66238 , n66222 );
not ( n387054 , n387023 );
or ( n387055 , n66238 , n387054 );
not ( n66241 , n387040 );
and ( n387057 , n66241 , n387038 );
nor ( n66243 , n387057 , n66235 );
nand ( n66244 , n387055 , n66243 );
nand ( n387060 , n387052 , n66244 );
buf ( n387061 , n387060 );
not ( n66247 , n387061 );
buf ( n66248 , n66247 );
buf ( n387064 , n66248 );
and ( n66250 , n387012 , n387064 );
not ( n387066 , n387012 );
buf ( n66252 , n387060 );
and ( n387068 , n387066 , n66252 );
nor ( n66254 , n66250 , n387068 );
buf ( n387070 , n66254 );
buf ( n387071 , n387070 );
xor ( n66257 , n66175 , n387071 );
or ( n387073 , n60515 , n379438 );
nand ( n387074 , n387073 , n60512 );
buf ( n387075 , n387074 );
xor ( n387076 , n66257 , n387075 );
buf ( n387077 , n387076 );
xor ( n66263 , n66166 , n387077 );
xor ( n387079 , n384850 , n385111 );
and ( n387080 , n387079 , n385163 );
and ( n66266 , n384850 , n385111 );
or ( n387082 , n387080 , n66266 );
buf ( n387083 , n387082 );
xor ( n66269 , n66263 , n387083 );
not ( n66270 , n66269 );
xor ( n387086 , n381030 , n384843 );
and ( n66272 , n387086 , n385165 );
and ( n387088 , n381030 , n384843 );
or ( n387089 , n66272 , n387088 );
buf ( n387090 , n387089 );
not ( n387091 , n387090 );
buf ( n387092 , n387091 );
nand ( n387093 , n66270 , n387092 );
xor ( n387094 , n386577 , n386593 );
and ( n387095 , n387094 , n386974 );
and ( n66281 , n386577 , n386593 );
or ( n387097 , n387095 , n66281 );
buf ( n387098 , n379299 );
not ( n387099 , n387098 );
buf ( n387100 , n386227 );
not ( n66286 , n387100 );
or ( n387102 , n387099 , n66286 );
buf ( n387103 , n379274 );
not ( n66289 , n387103 );
buf ( n387105 , n372458 );
not ( n387106 , n387105 );
or ( n66292 , n66289 , n387106 );
buf ( n387108 , n39867 );
buf ( n387109 , n379271 );
nand ( n387110 , n387108 , n387109 );
buf ( n387111 , n387110 );
buf ( n387112 , n387111 );
nand ( n387113 , n66292 , n387112 );
buf ( n387114 , n387113 );
buf ( n387115 , n387114 );
buf ( n387116 , n379944 );
nand ( n66302 , n387115 , n387116 );
buf ( n387118 , n66302 );
buf ( n387119 , n387118 );
nand ( n387120 , n387102 , n387119 );
buf ( n387121 , n387120 );
buf ( n387122 , n377580 );
not ( n66308 , n387122 );
and ( n66309 , n377585 , n44925 );
not ( n387125 , n377585 );
and ( n387126 , n387125 , n359756 );
or ( n66312 , n66309 , n387126 );
buf ( n387128 , n66312 );
not ( n66314 , n387128 );
or ( n387130 , n66308 , n66314 );
buf ( n387131 , n386949 );
buf ( n387132 , n57530 );
nand ( n387133 , n387131 , n387132 );
buf ( n387134 , n387133 );
buf ( n387135 , n387134 );
nand ( n66321 , n387130 , n387135 );
buf ( n387137 , n66321 );
buf ( n66323 , n387137 );
not ( n387139 , n66323 );
buf ( n387140 , n387139 );
xor ( n387141 , n387121 , n387140 );
buf ( n387142 , n386461 );
not ( n66328 , n387142 );
buf ( n387144 , n359916 );
not ( n387145 , n387144 );
or ( n387146 , n66328 , n387145 );
buf ( n387147 , n367440 );
buf ( n387148 , n377757 );
not ( n387149 , n387148 );
buf ( n387150 , n364909 );
not ( n387151 , n387150 );
or ( n387152 , n387149 , n387151 );
buf ( n387153 , n44743 );
buf ( n387154 , n378886 );
nand ( n66340 , n387153 , n387154 );
buf ( n387156 , n66340 );
buf ( n387157 , n387156 );
nand ( n66343 , n387152 , n387157 );
buf ( n387159 , n66343 );
buf ( n387160 , n387159 );
nand ( n66346 , n387147 , n387160 );
buf ( n387162 , n66346 );
buf ( n387163 , n387162 );
nand ( n66349 , n387146 , n387163 );
buf ( n387165 , n66349 );
buf ( n387166 , n386418 );
not ( n387167 , n387166 );
buf ( n387168 , n46135 );
not ( n387169 , n387168 );
or ( n66355 , n387167 , n387169 );
buf ( n387171 , n378736 );
not ( n387172 , n387171 );
buf ( n387173 , n361597 );
not ( n66359 , n387173 );
or ( n387175 , n387172 , n66359 );
buf ( n387176 , n366329 );
buf ( n387177 , n49315 );
nand ( n387178 , n387176 , n387177 );
buf ( n387179 , n387178 );
buf ( n387180 , n387179 );
nand ( n387181 , n387175 , n387180 );
buf ( n387182 , n387181 );
buf ( n387183 , n387182 );
buf ( n387184 , n368724 );
nand ( n387185 , n387183 , n387184 );
buf ( n387186 , n387185 );
buf ( n387187 , n387186 );
nand ( n387188 , n66355 , n387187 );
buf ( n387189 , n387188 );
buf ( n387190 , n386814 );
not ( n387191 , n387190 );
buf ( n387192 , n387191 );
buf ( n387193 , n387192 );
not ( n66379 , n387193 );
buf ( n387195 , n50782 );
not ( n66381 , n387195 );
and ( n387197 , n66379 , n66381 );
buf ( n387198 , n56849 );
not ( n66384 , n387198 );
buf ( n387200 , n44661 );
not ( n66386 , n387200 );
or ( n387202 , n66384 , n66386 );
buf ( n387203 , n58471 );
buf ( n387204 , n31072 );
nand ( n66390 , n387203 , n387204 );
buf ( n387206 , n66390 );
buf ( n387207 , n387206 );
nand ( n66393 , n387202 , n387207 );
buf ( n387209 , n66393 );
buf ( n387210 , n387209 );
buf ( n387211 , n366428 );
and ( n66397 , n387210 , n387211 );
nor ( n387213 , n387197 , n66397 );
buf ( n387214 , n387213 );
buf ( n387215 , n387214 );
buf ( n387216 , n386380 );
and ( n66402 , n387215 , n387216 );
not ( n66403 , n387215 );
buf ( n387219 , n386377 );
and ( n66405 , n66403 , n387219 );
or ( n387221 , n66402 , n66405 );
buf ( n387222 , n387221 );
not ( n66408 , n387222 );
xor ( n387224 , n387189 , n66408 );
not ( n387225 , n387224 );
and ( n66411 , n387165 , n387225 );
not ( n387227 , n387165 );
and ( n387228 , n387227 , n387224 );
or ( n66414 , n66411 , n387228 );
xor ( n387230 , n65879 , n386722 );
and ( n387231 , n387230 , n386748 );
and ( n66417 , n65879 , n386722 );
or ( n387233 , n387231 , n66417 );
buf ( n387234 , n387233 );
xor ( n66420 , n66414 , n387234 );
xor ( n66421 , n387141 , n66420 );
buf ( n387237 , n66421 );
not ( n66423 , n387237 );
buf ( n387239 , n66423 );
buf ( n387240 , n379890 );
not ( n387241 , n387240 );
not ( n387242 , n379841 );
not ( n66428 , n41472 );
or ( n66429 , n387242 , n66428 );
buf ( n66430 , n40899 );
buf ( n66431 , n379847 );
nand ( n66432 , n66430 , n66431 );
buf ( n66433 , n66432 );
nand ( n387249 , n66429 , n66433 );
buf ( n387250 , n387249 );
not ( n387251 , n387250 );
or ( n387252 , n387241 , n387251 );
buf ( n387253 , n379916 );
buf ( n66439 , n386918 );
nand ( n66440 , n387253 , n66439 );
buf ( n66441 , n66440 );
buf ( n387257 , n66441 );
nand ( n387258 , n387252 , n387257 );
buf ( n387259 , n387258 );
buf ( n387260 , n387259 );
buf ( n387261 , n66083 );
not ( n387262 , n387261 );
not ( n387263 , n386750 );
nand ( n66449 , n387263 , n386796 );
buf ( n387265 , n66449 );
nand ( n387266 , n387262 , n387265 );
buf ( n387267 , n387266 );
buf ( n387268 , n387267 );
nand ( n66454 , n65982 , n386750 );
buf ( n387270 , n66454 );
nand ( n66456 , n387268 , n387270 );
buf ( n387272 , n66456 );
buf ( n387273 , n387272 );
xor ( n66459 , n387260 , n387273 );
buf ( n387275 , n386258 );
not ( n387276 , n387275 );
buf ( n387277 , n386314 );
not ( n66463 , n387277 );
or ( n387279 , n387276 , n66463 );
buf ( n387280 , n386258 );
buf ( n387281 , n386314 );
or ( n387282 , n387280 , n387281 );
buf ( n387283 , n65531 );
nand ( n66469 , n387282 , n387283 );
buf ( n66470 , n66469 );
buf ( n387286 , n66470 );
nand ( n66472 , n387279 , n387286 );
buf ( n66473 , n66472 );
buf ( n387289 , n66473 );
xor ( n66475 , n66459 , n387289 );
buf ( n387291 , n66475 );
xor ( n387292 , n387239 , n387291 );
or ( n66478 , n386506 , n386558 );
and ( n387294 , n66478 , n386567 );
and ( n387295 , n386507 , n386559 );
buf ( n387296 , n387295 );
nor ( n387297 , n387294 , n387296 );
buf ( n387298 , n387297 );
buf ( n66484 , n387298 );
buf ( n387300 , n66484 );
and ( n387301 , n387292 , n387300 );
not ( n387302 , n387292 );
not ( n66488 , n387300 );
and ( n387304 , n387302 , n66488 );
nor ( n387305 , n387301 , n387304 );
xor ( n387306 , n387097 , n387305 );
not ( n387307 , n387060 );
not ( n66493 , n66186 );
and ( n387309 , n387307 , n66493 );
not ( n387310 , n387000 );
nand ( n66496 , n387310 , n387060 );
buf ( n387312 , n387006 );
not ( n387313 , n387312 );
buf ( n387314 , n387313 );
and ( n387315 , n66496 , n387314 );
nor ( n66501 , n387309 , n387315 );
xor ( n387317 , n387306 , n66501 );
xor ( n387318 , n66175 , n387071 );
and ( n66504 , n387318 , n387075 );
and ( n66505 , n66175 , n387071 );
or ( n387321 , n66504 , n66505 );
buf ( n387322 , n387321 );
buf ( n387323 , n387322 );
not ( n66509 , n387323 );
buf ( n387325 , n66509 );
xor ( n66511 , n387317 , n387325 );
not ( n387327 , n45075 );
buf ( n387328 , n342881 );
not ( n387329 , n387328 );
buf ( n387330 , n44783 );
not ( n66516 , n387330 );
or ( n387332 , n387329 , n66516 );
buf ( n387333 , n41607 );
buf ( n387334 , n365202 );
nand ( n66520 , n387333 , n387334 );
buf ( n66521 , n66520 );
buf ( n387337 , n66521 );
nand ( n387338 , n387332 , n387337 );
buf ( n387339 , n387338 );
not ( n387340 , n387339 );
or ( n387341 , n387327 , n387340 );
not ( n66527 , n65945 );
not ( n66528 , n386761 );
or ( n387344 , n66527 , n66528 );
nand ( n66530 , n387344 , n365226 );
nand ( n66531 , n387341 , n66530 );
buf ( n387347 , n365152 );
not ( n387348 , n387347 );
buf ( n387349 , n46397 );
not ( n66535 , n387349 );
buf ( n387351 , n45718 );
not ( n387352 , n387351 );
or ( n66538 , n66535 , n387352 );
buf ( n387354 , n362133 );
buf ( n387355 , n342909 );
buf ( n387356 , n387355 );
nand ( n387357 , n387354 , n387356 );
buf ( n387358 , n387357 );
buf ( n387359 , n387358 );
nand ( n66545 , n66538 , n387359 );
buf ( n66546 , n66545 );
buf ( n387362 , n66546 );
not ( n387363 , n387362 );
or ( n66549 , n387348 , n387363 );
buf ( n387365 , n386340 );
buf ( n387366 , n365189 );
nand ( n66552 , n387365 , n387366 );
buf ( n387368 , n66552 );
buf ( n387369 , n387368 );
nand ( n387370 , n66549 , n387369 );
buf ( n387371 , n387370 );
xor ( n387372 , n66531 , n387371 );
not ( n66558 , n56794 );
not ( n387374 , n22619 );
not ( n387375 , n366077 );
or ( n66561 , n387374 , n387375 );
buf ( n387377 , n32084 );
buf ( n387378 , n365670 );
nand ( n387379 , n387377 , n387378 );
buf ( n387380 , n387379 );
nand ( n66566 , n66561 , n387380 );
not ( n387382 , n66566 );
or ( n387383 , n66558 , n387382 );
buf ( n387384 , n65623 );
buf ( n387385 , n45553 );
nand ( n387386 , n387384 , n387385 );
buf ( n387387 , n387386 );
nand ( n66573 , n387383 , n387387 );
buf ( n387389 , n66573 );
not ( n387390 , n65874 );
not ( n66576 , n45438 );
or ( n387392 , n387390 , n66576 );
buf ( n387393 , n44737 );
buf ( n387394 , n45455 );
and ( n387395 , n387393 , n387394 );
not ( n387396 , n387393 );
buf ( n387397 , n365626 );
and ( n66583 , n387396 , n387397 );
nor ( n387399 , n387395 , n66583 );
buf ( n387400 , n387399 );
buf ( n387401 , n387400 );
not ( n66587 , n387401 );
buf ( n387403 , n365622 );
nand ( n387404 , n66587 , n387403 );
buf ( n387405 , n387404 );
nand ( n66591 , n387392 , n387405 );
buf ( n387407 , n66591 );
xor ( n387408 , n387389 , n387407 );
buf ( n387409 , n386740 );
not ( n66595 , n387409 );
buf ( n387411 , n364849 );
not ( n66597 , n387411 );
or ( n66598 , n66595 , n66597 );
buf ( n387414 , n365490 );
not ( n66600 , n387414 );
buf ( n387416 , n41386 );
not ( n387417 , n387416 );
or ( n66603 , n66600 , n387417 );
buf ( n387419 , n41386 );
not ( n387420 , n387419 );
buf ( n387421 , n387420 );
buf ( n387422 , n387421 );
buf ( n387423 , n45336 );
nand ( n66609 , n387422 , n387423 );
buf ( n66610 , n66609 );
buf ( n66611 , n66610 );
nand ( n387427 , n66603 , n66611 );
buf ( n387428 , n387427 );
buf ( n387429 , n387428 );
buf ( n387430 , n367590 );
nand ( n387431 , n387429 , n387430 );
buf ( n387432 , n387431 );
buf ( n387433 , n387432 );
nand ( n66619 , n66598 , n387433 );
buf ( n387435 , n66619 );
buf ( n387436 , n387435 );
xor ( n66622 , n387408 , n387436 );
buf ( n387438 , n66622 );
xnor ( n387439 , n387372 , n387438 );
buf ( n387440 , n387439 );
xor ( n66626 , n386619 , n386642 );
and ( n387442 , n66626 , n386668 );
and ( n387443 , n386619 , n386642 );
or ( n66629 , n387442 , n387443 );
buf ( n387445 , n66629 );
buf ( n387446 , n387445 );
xor ( n66632 , n387440 , n387446 );
xor ( n66633 , n386279 , n386288 );
and ( n387449 , n66633 , n386313 );
and ( n387450 , n386279 , n386288 );
or ( n66636 , n387449 , n387450 );
not ( n66637 , n386767 );
not ( n387453 , n386794 );
or ( n387454 , n66637 , n387453 );
nand ( n66640 , n387454 , n65941 );
nand ( n66641 , n65976 , n65951 );
nand ( n66642 , n66640 , n66641 );
xor ( n387458 , n66636 , n66642 );
nor ( n387459 , n386897 , n66070 );
or ( n66645 , n387459 , n386872 );
nand ( n66646 , n386897 , n66070 );
nand ( n66647 , n66645 , n66646 );
xor ( n387463 , n387458 , n66647 );
buf ( n387464 , n387463 );
xnor ( n66650 , n66632 , n387464 );
buf ( n387466 , n66650 );
buf ( n387467 , n387466 );
buf ( n387468 , n386670 );
not ( n66654 , n387468 );
buf ( n387470 , n66654 );
nand ( n387471 , n386969 , n387470 );
buf ( n387472 , n386899 );
not ( n66658 , n387472 );
buf ( n387474 , n66658 );
and ( n66660 , n387471 , n387474 );
nor ( n66661 , n386969 , n387470 );
nor ( n66662 , n66660 , n66661 );
buf ( n387478 , n66662 );
not ( n66664 , n387478 );
buf ( n387480 , n66664 );
buf ( n387481 , n387480 );
xor ( n66667 , n387467 , n387481 );
not ( n66668 , n386923 );
not ( n66669 , n386962 );
or ( n66670 , n66668 , n66669 );
nand ( n66671 , n66670 , n66117 );
not ( n66672 , n386962 );
nand ( n66673 , n386926 , n66672 );
nand ( n66674 , n66671 , n66673 );
buf ( n387490 , n47466 );
not ( n66676 , n387490 );
buf ( n387492 , n386608 );
not ( n66678 , n387492 );
or ( n66679 , n66676 , n66678 );
buf ( n387495 , n365041 );
not ( n66681 , n387495 );
buf ( n387497 , n368474 );
not ( n66683 , n387497 );
or ( n66684 , n66681 , n66683 );
buf ( n387500 , n360885 );
buf ( n387501 , n365052 );
nand ( n66687 , n387500 , n387501 );
buf ( n387503 , n66687 );
buf ( n387504 , n387503 );
nand ( n66690 , n66684 , n387504 );
buf ( n387506 , n66690 );
buf ( n387507 , n387506 );
buf ( n387508 , n44915 );
nand ( n387509 , n387507 , n387508 );
buf ( n387510 , n387509 );
buf ( n387511 , n387510 );
nand ( n387512 , n66679 , n387511 );
buf ( n387513 , n387512 );
buf ( n387514 , n387513 );
buf ( n387515 , n369804 );
not ( n387516 , n387515 );
buf ( n387517 , n386657 );
not ( n387518 , n387517 );
or ( n387519 , n387516 , n387518 );
buf ( n387520 , n369769 );
not ( n387521 , n387520 );
buf ( n387522 , n46902 );
not ( n66708 , n387522 );
or ( n66709 , n387521 , n66708 );
buf ( n387525 , n40199 );
buf ( n387526 , n369766 );
nand ( n387527 , n387525 , n387526 );
buf ( n387528 , n387527 );
buf ( n66714 , n387528 );
nand ( n387530 , n66709 , n66714 );
buf ( n387531 , n387530 );
buf ( n387532 , n387531 );
buf ( n387533 , n49609 );
nand ( n387534 , n387532 , n387533 );
buf ( n387535 , n387534 );
buf ( n387536 , n387535 );
nand ( n387537 , n387519 , n387536 );
buf ( n387538 , n387537 );
buf ( n387539 , n387538 );
xor ( n66725 , n387514 , n387539 );
buf ( n387541 , n66725 );
buf ( n387542 , n369444 );
buf ( n387543 , n387542 );
not ( n66729 , n387543 );
buf ( n387545 , n368549 );
not ( n387546 , n387545 );
buf ( n387547 , n40252 );
not ( n66733 , n387547 );
or ( n387549 , n387546 , n66733 );
buf ( n387550 , n54491 );
buf ( n387551 , n368554 );
nand ( n66737 , n387550 , n387551 );
buf ( n66738 , n66737 );
buf ( n387554 , n66738 );
nand ( n66740 , n387549 , n387554 );
buf ( n387556 , n66740 );
buf ( n387557 , n387556 );
not ( n387558 , n387557 );
or ( n66744 , n66729 , n387558 );
buf ( n387560 , n386521 );
buf ( n387561 , n368611 );
nand ( n66747 , n387560 , n387561 );
buf ( n387563 , n66747 );
buf ( n387564 , n387563 );
nand ( n387565 , n66744 , n387564 );
buf ( n387566 , n387565 );
buf ( n387567 , n387566 );
not ( n387568 , n387567 );
buf ( n387569 , n387568 );
and ( n387570 , n387541 , n387569 );
not ( n387571 , n387541 );
buf ( n66757 , n387566 );
and ( n66758 , n387571 , n66757 );
nor ( n66759 , n387570 , n66758 );
xor ( n387575 , n66674 , n66759 );
not ( n66761 , n66080 );
not ( n387577 , n359809 );
or ( n387578 , n66761 , n387577 );
buf ( n387579 , n362521 );
buf ( n387580 , n377122 );
not ( n387581 , n387580 );
buf ( n387582 , n366537 );
not ( n66768 , n387582 );
or ( n387584 , n387581 , n66768 );
buf ( n387585 , n39621 );
buf ( n387586 , n57463 );
nand ( n66772 , n387585 , n387586 );
buf ( n387588 , n66772 );
buf ( n387589 , n387588 );
nand ( n66775 , n387584 , n387589 );
buf ( n387591 , n66775 );
buf ( n387592 , n387591 );
nand ( n387593 , n387579 , n387592 );
buf ( n387594 , n387593 );
nand ( n387595 , n387578 , n387594 );
not ( n66781 , n387595 );
not ( n387597 , n66781 );
not ( n387598 , n65552 );
not ( n66784 , n361013 );
or ( n66785 , n387598 , n66784 );
not ( n387601 , n365428 );
not ( n387602 , n365290 );
or ( n387603 , n387601 , n387602 );
buf ( n387604 , n365266 );
buf ( n387605 , n365422 );
nand ( n387606 , n387604 , n387605 );
buf ( n387607 , n387606 );
nand ( n66793 , n387603 , n387607 );
nand ( n387609 , n66793 , n365303 );
nand ( n387610 , n66785 , n387609 );
not ( n66796 , n387610 );
not ( n387612 , n365033 );
not ( n66798 , n386714 );
or ( n387614 , n387612 , n66798 );
not ( n387615 , n364981 );
not ( n66801 , n366322 );
or ( n387617 , n387615 , n66801 );
buf ( n387618 , n361716 );
buf ( n387619 , n364978 );
nand ( n66805 , n387618 , n387619 );
buf ( n66806 , n66805 );
nand ( n387622 , n387617 , n66806 );
nand ( n66808 , n387622 , n365115 );
nand ( n387624 , n387614 , n66808 );
not ( n387625 , n387624 );
and ( n66811 , n66796 , n387625 );
not ( n66812 , n66796 );
and ( n387628 , n66812 , n387624 );
nor ( n387629 , n66811 , n387628 );
not ( n66815 , n387629 );
or ( n66816 , n387597 , n66815 );
or ( n387632 , n387629 , n66781 );
nand ( n387633 , n66816 , n387632 );
buf ( n387634 , n387633 );
not ( n66820 , n386824 );
not ( n66821 , n66030 );
or ( n387637 , n66820 , n66821 );
or ( n66823 , n66030 , n386824 );
nand ( n66824 , n66823 , n386870 );
nand ( n66825 , n387637 , n66824 );
buf ( n387641 , n386306 );
not ( n66827 , n387641 );
buf ( n387643 , n40058 );
not ( n66829 , n387643 );
or ( n66830 , n66827 , n66829 );
not ( n66831 , n365495 );
not ( n66832 , n377352 );
or ( n66833 , n66831 , n66832 );
nand ( n66834 , n365945 , n377353 );
nand ( n66835 , n66833 , n66834 );
nand ( n387651 , n365486 , n66835 );
buf ( n387652 , n387651 );
nand ( n66838 , n66830 , n387652 );
buf ( n387654 , n66838 );
xor ( n387655 , n66825 , n387654 );
xor ( n387656 , n386381 , n386402 );
and ( n387657 , n387656 , n386427 );
and ( n66843 , n386381 , n386402 );
or ( n387659 , n387657 , n66843 );
buf ( n387660 , n387659 );
xor ( n66846 , n387655 , n387660 );
buf ( n387662 , n66846 );
xor ( n387663 , n387634 , n387662 );
buf ( n387664 , n43261 );
not ( n387665 , n387664 );
buf ( n387666 , n55539 );
not ( n387667 , n387666 );
buf ( n387668 , n32160 );
not ( n66854 , n387668 );
or ( n66855 , n387667 , n66854 );
buf ( n387671 , n352192 );
buf ( n387672 , n381286 );
nand ( n387673 , n387671 , n387672 );
buf ( n387674 , n387673 );
buf ( n387675 , n387674 );
nand ( n387676 , n66855 , n387675 );
buf ( n387677 , n387676 );
buf ( n387678 , n387677 );
not ( n66864 , n387678 );
or ( n387680 , n387665 , n66864 );
buf ( n387681 , n363429 );
buf ( n387682 , n386370 );
nand ( n66868 , n387681 , n387682 );
buf ( n387684 , n66868 );
buf ( n387685 , n387684 );
nand ( n66871 , n387680 , n387685 );
buf ( n387687 , n66871 );
not ( n387688 , n46463 );
not ( n387689 , n46477 );
not ( n387690 , n365328 );
or ( n66876 , n387689 , n387690 );
buf ( n387692 , n375901 );
not ( n387693 , n387692 );
buf ( n387694 , n30911 );
nand ( n66880 , n387693 , n387694 );
buf ( n66881 , n66880 );
nand ( n387697 , n66876 , n66881 );
not ( n387698 , n387697 );
or ( n66884 , n387688 , n387698 );
buf ( n387700 , n386863 );
buf ( n387701 , n46521 );
nand ( n66887 , n387700 , n387701 );
buf ( n387703 , n66887 );
nand ( n387704 , n66884 , n387703 );
xor ( n66890 , n387687 , n387704 );
not ( n66891 , n386843 );
not ( n387707 , n368706 );
or ( n66893 , n66891 , n387707 );
not ( n66894 , n377297 );
buf ( n387710 , n66894 );
buf ( n387711 , n342335 );
and ( n66897 , n387710 , n387711 );
not ( n66898 , n387710 );
buf ( n387714 , n365915 );
and ( n66900 , n66898 , n387714 );
nor ( n66901 , n66897 , n66900 );
buf ( n387717 , n66901 );
not ( n66903 , n387717 );
nand ( n387719 , n66903 , n362386 );
nand ( n66905 , n66893 , n387719 );
xor ( n66906 , n66890 , n66905 );
buf ( n387722 , n66906 );
buf ( n387723 , n386786 );
not ( n66909 , n387723 );
buf ( n387725 , n46113 );
not ( n66911 , n387725 );
or ( n66912 , n66909 , n66911 );
not ( n66913 , n368665 );
not ( n66914 , n365468 );
or ( n66915 , n66913 , n66914 );
buf ( n387731 , n362452 );
buf ( n387732 , n368662 );
nand ( n66918 , n387731 , n387732 );
buf ( n387734 , n66918 );
nand ( n387735 , n66915 , n387734 );
buf ( n387736 , n387735 );
buf ( n387737 , n366757 );
nand ( n66923 , n387736 , n387737 );
buf ( n387739 , n66923 );
buf ( n387740 , n387739 );
nand ( n66926 , n66912 , n387740 );
buf ( n387742 , n66926 );
buf ( n387743 , n387742 );
xor ( n387744 , n387722 , n387743 );
buf ( n387745 , n367273 );
not ( n387746 , n387745 );
buf ( n387747 , n387746 );
buf ( n387748 , n387747 );
buf ( n387749 , n66064 );
or ( n387750 , n387748 , n387749 );
buf ( n66936 , n39218 );
and ( n66937 , n365367 , n49178 );
not ( n387753 , n365367 );
and ( n387754 , n387753 , n369374 );
nor ( n66940 , n66937 , n387754 );
buf ( n387756 , n66940 );
or ( n66942 , n66936 , n387756 );
nand ( n66943 , n387750 , n66942 );
buf ( n387759 , n66943 );
buf ( n387760 , n387759 );
xor ( n66946 , n387744 , n387760 );
buf ( n66947 , n66946 );
buf ( n387763 , n66947 );
xor ( n66949 , n387663 , n387763 );
buf ( n387765 , n66949 );
buf ( n387766 , n387765 );
not ( n387767 , n387766 );
buf ( n387768 , n387767 );
and ( n387769 , n387575 , n387768 );
not ( n66955 , n387575 );
and ( n387771 , n66955 , n387765 );
nor ( n66957 , n387769 , n387771 );
buf ( n387773 , n66957 );
xor ( n387774 , n66667 , n387773 );
buf ( n387775 , n387774 );
buf ( n387776 , n387775 );
not ( n387777 , n387776 );
not ( n387778 , n66204 );
buf ( n387779 , n66235 );
not ( n387780 , n387779 );
buf ( n387781 , n387780 );
not ( n66967 , n387781 );
or ( n387783 , n387778 , n66967 );
not ( n66969 , n66235 );
not ( n66970 , n387022 );
or ( n66971 , n66969 , n66970 );
nand ( n66972 , n66971 , n66222 );
nand ( n66973 , n387783 , n66972 );
buf ( n387789 , n66973 );
buf ( n387790 , n65710 );
not ( n66976 , n387790 );
not ( n66977 , n65510 );
buf ( n387793 , n66977 );
not ( n387794 , n387793 );
or ( n66980 , n66976 , n387794 );
or ( n387796 , n65710 , n66977 );
nand ( n387797 , n387796 , n65521 );
buf ( n387798 , n387797 );
nand ( n66984 , n66980 , n387798 );
buf ( n387800 , n66984 );
buf ( n387801 , n387800 );
xor ( n387802 , n387789 , n387801 );
buf ( n387803 , n386210 );
buf ( n387804 , n386234 );
nand ( n387805 , n387803 , n387804 );
buf ( n387806 , n387805 );
or ( n387807 , n386234 , n386210 );
nand ( n387808 , n387807 , n386240 );
nand ( n66994 , n387806 , n387808 );
not ( n66995 , n66994 );
not ( n387811 , n386482 );
not ( n66997 , n386472 );
or ( n387813 , n387811 , n66997 );
not ( n66999 , n386315 );
not ( n387815 , n65701 );
or ( n67001 , n66999 , n387815 );
nand ( n67002 , n67001 , n386321 );
nand ( n387818 , n387813 , n67002 );
xor ( n387819 , n66995 , n387818 );
xor ( n67005 , n386529 , n386540 );
and ( n387821 , n67005 , n386556 );
and ( n387822 , n386529 , n386540 );
or ( n67008 , n387821 , n387822 );
buf ( n387824 , n67008 );
buf ( n387825 , n386206 );
not ( n67011 , n387825 );
buf ( n387827 , n58867 );
buf ( n387828 , n58923 );
nor ( n67014 , n387827 , n387828 );
buf ( n387830 , n67014 );
buf ( n67016 , n387830 );
nor ( n67017 , n67011 , n67016 );
buf ( n67018 , n67017 );
not ( n387834 , n67018 );
not ( n67020 , n386467 );
not ( n387836 , n386347 );
or ( n387837 , n67020 , n387836 );
buf ( n387838 , n386467 );
buf ( n387839 , n386347 );
nor ( n67025 , n387838 , n387839 );
buf ( n387841 , n67025 );
or ( n387842 , n387841 , n65658 );
nand ( n67028 , n387837 , n387842 );
not ( n67029 , n67028 );
and ( n67030 , n387834 , n67029 );
not ( n387846 , n387834 );
and ( n67032 , n387846 , n67028 );
nor ( n67033 , n67030 , n67032 );
xor ( n67034 , n387824 , n67033 );
xor ( n387850 , n387819 , n67034 );
buf ( n387851 , n387850 );
xor ( n67037 , n387802 , n387851 );
buf ( n387853 , n67037 );
not ( n67039 , n387853 );
buf ( n387855 , n67039 );
not ( n67041 , n387855 );
or ( n387857 , n387777 , n67041 );
buf ( n387858 , n387775 );
not ( n387859 , n387858 );
buf ( n387860 , n387853 );
nand ( n67046 , n387859 , n387860 );
buf ( n387862 , n67046 );
buf ( n387863 , n387862 );
nand ( n67049 , n387857 , n387863 );
buf ( n387865 , n67049 );
buf ( n387866 , n387865 );
buf ( n387867 , n65711 );
not ( n387868 , n387867 );
buf ( n387869 , n387868 );
buf ( n387870 , n387869 );
not ( n387871 , n387870 );
buf ( n387872 , n386975 );
not ( n67058 , n387872 );
or ( n387874 , n387871 , n67058 );
buf ( n387875 , n386499 );
nand ( n387876 , n387874 , n387875 );
buf ( n387877 , n387876 );
not ( n387878 , n387869 );
nand ( n67064 , n66161 , n387878 );
nand ( n387880 , n387877 , n67064 );
buf ( n387881 , n387880 );
not ( n67067 , n387881 );
buf ( n67068 , n67067 );
buf ( n387884 , n67068 );
and ( n67070 , n387866 , n387884 );
not ( n67071 , n387866 );
buf ( n387887 , n387877 );
buf ( n387888 , n67064 );
nand ( n67074 , n387887 , n387888 );
buf ( n67075 , n67074 );
buf ( n67076 , n67075 );
and ( n67077 , n67071 , n67076 );
nor ( n387893 , n67070 , n67077 );
buf ( n387894 , n387893 );
xor ( n67080 , n66511 , n387894 );
buf ( n387896 , n387077 );
not ( n387897 , n387896 );
buf ( n387898 , n387897 );
not ( n387899 , n387898 );
buf ( n67085 , n66166 );
not ( n67086 , n67085 );
buf ( n387902 , n67086 );
not ( n387903 , n387902 );
and ( n387904 , n387899 , n387903 );
buf ( n67090 , n387083 );
buf ( n387906 , n387898 );
buf ( n67092 , n387902 );
nand ( n67093 , n387906 , n67092 );
buf ( n67094 , n67093 );
and ( n67095 , n67090 , n67094 );
nor ( n67096 , n387904 , n67095 );
nand ( n67097 , n67080 , n67096 );
nand ( n67098 , n386196 , n387093 , n67097 );
buf ( n387914 , n66269 );
buf ( n387915 , n387089 );
nand ( n67101 , n387914 , n387915 );
buf ( n387917 , n67101 );
not ( n67103 , n387917 );
nand ( n387919 , n67103 , n67097 );
not ( n387920 , n67096 );
not ( n67106 , n67080 );
and ( n387922 , n387920 , n67106 );
xor ( n67108 , n387097 , n387305 );
and ( n67109 , n67108 , n66501 );
and ( n67110 , n387097 , n387305 );
or ( n67111 , n67109 , n67110 );
buf ( n387927 , n67111 );
not ( n67113 , n67039 );
buf ( n387929 , n67113 );
not ( n67115 , n387929 );
buf ( n387931 , n387775 );
not ( n67117 , n387931 );
or ( n387933 , n67115 , n67117 );
buf ( n387934 , n387880 );
buf ( n387935 , n387775 );
not ( n387936 , n387935 );
buf ( n387937 , n67039 );
nand ( n387938 , n387936 , n387937 );
buf ( n387939 , n387938 );
buf ( n387940 , n387939 );
nand ( n387941 , n387934 , n387940 );
buf ( n387942 , n387941 );
buf ( n387943 , n387942 );
nand ( n387944 , n387933 , n387943 );
buf ( n387945 , n387944 );
buf ( n387946 , n387945 );
not ( n387947 , n387946 );
buf ( n387948 , n387947 );
buf ( n387949 , n387948 );
xor ( n387950 , n387927 , n387949 );
not ( n67118 , n387114 );
not ( n67119 , n65117 );
or ( n387953 , n67118 , n67119 );
buf ( n387954 , n365167 );
not ( n387955 , n387954 );
buf ( n387956 , n379271 );
not ( n387957 , n387956 );
and ( n67125 , n387955 , n387957 );
buf ( n387959 , n41406 );
buf ( n387960 , n379271 );
and ( n387961 , n387959 , n387960 );
nor ( n67129 , n67125 , n387961 );
buf ( n67130 , n67129 );
not ( n387964 , n67130 );
nand ( n67132 , n387964 , n379263 );
nand ( n387966 , n387953 , n67132 );
not ( n387967 , n387966 );
or ( n67135 , n66531 , n387371 );
nand ( n387969 , n67135 , n387438 );
buf ( n387970 , n387371 );
buf ( n387971 , n66531 );
nand ( n387972 , n387970 , n387971 );
buf ( n387973 , n387972 );
nand ( n67141 , n387969 , n387973 );
not ( n387975 , n67141 );
or ( n387976 , n387967 , n387975 );
or ( n67144 , n67141 , n387966 );
nand ( n387978 , n387976 , n67144 );
not ( n387979 , n57530 );
not ( n387980 , n66312 );
or ( n67148 , n387979 , n387980 );
buf ( n387982 , n377585 );
not ( n67150 , n387982 );
buf ( n387984 , n366600 );
not ( n67152 , n387984 );
or ( n387986 , n67150 , n67152 );
buf ( n387987 , n39830 );
buf ( n387988 , n386943 );
nand ( n387989 , n387987 , n387988 );
buf ( n387990 , n387989 );
buf ( n387991 , n387990 );
nand ( n387992 , n387986 , n387991 );
buf ( n387993 , n387992 );
buf ( n387994 , n387993 );
buf ( n387995 , n377580 );
nand ( n67163 , n387994 , n387995 );
buf ( n387997 , n67163 );
nand ( n67165 , n67148 , n387997 );
buf ( n67166 , n67165 );
and ( n67167 , n387978 , n67166 );
not ( n388001 , n387978 );
not ( n388002 , n67165 );
and ( n67170 , n388001 , n388002 );
nor ( n388004 , n67167 , n67170 );
xor ( n67172 , n387260 , n387273 );
and ( n67173 , n67172 , n387289 );
and ( n67174 , n387260 , n387273 );
or ( n388008 , n67173 , n67174 );
buf ( n388009 , n388008 );
xor ( n67177 , n388004 , n388009 );
not ( n67178 , n66757 );
not ( n388012 , n387541 );
and ( n388013 , n67178 , n388012 );
not ( n67181 , n387569 );
and ( n67182 , n67181 , n387541 );
nor ( n67183 , n388013 , n67182 );
buf ( n388017 , n67183 );
buf ( n388018 , n66674 );
or ( n67186 , n388017 , n388018 );
buf ( n388020 , n387765 );
nand ( n67188 , n67186 , n388020 );
buf ( n388022 , n67188 );
buf ( n388023 , n388022 );
not ( n388024 , n66673 );
not ( n67192 , n66671 );
or ( n67193 , n388024 , n67192 );
nand ( n388027 , n67193 , n67183 );
buf ( n67195 , n388027 );
nand ( n67196 , n388023 , n67195 );
buf ( n67197 , n67196 );
xor ( n388031 , n67177 , n67197 );
buf ( n388032 , n388031 );
not ( n388033 , n388032 );
buf ( n388034 , n388033 );
not ( n67202 , n388034 );
not ( n67203 , n387466 );
not ( n388037 , n387480 );
or ( n67205 , n67203 , n388037 );
not ( n388039 , n66662 );
buf ( n388040 , n387466 );
not ( n67208 , n388040 );
buf ( n388042 , n67208 );
not ( n388043 , n388042 );
or ( n67211 , n388039 , n388043 );
nand ( n388045 , n67211 , n66957 );
nand ( n388046 , n67205 , n388045 );
not ( n67214 , n388046 );
not ( n388048 , n67214 );
or ( n388049 , n67202 , n388048 );
buf ( n388050 , n388046 );
buf ( n388051 , n388031 );
nand ( n388052 , n388050 , n388051 );
buf ( n388053 , n388052 );
nand ( n67221 , n388049 , n388053 );
buf ( n388055 , n387463 );
not ( n388056 , n388055 );
buf ( n388057 , n388056 );
not ( n67225 , n388057 );
buf ( n388059 , n387439 );
buf ( n388060 , n388059 );
buf ( n388061 , n388060 );
not ( n67229 , n388061 );
and ( n388063 , n67225 , n67229 );
buf ( n388064 , n388057 );
buf ( n388065 , n388061 );
nand ( n67233 , n388064 , n388065 );
buf ( n388067 , n67233 );
and ( n388068 , n388067 , n387445 );
nor ( n67236 , n388063 , n388068 );
and ( n388070 , n351160 , n362033 );
not ( n67237 , n351160 );
and ( n67238 , n67237 , n364832 );
nor ( n67239 , n388070 , n67238 );
not ( n388074 , n67239 );
not ( n67241 , n41915 );
or ( n388076 , n388074 , n67241 );
not ( n67243 , n387400 );
nand ( n67244 , n67243 , n386678 );
nand ( n388079 , n388076 , n67244 );
buf ( n388080 , n46336 );
and ( n67247 , n351229 , n41386 );
not ( n388082 , n351229 );
and ( n388083 , n388082 , n387421 );
or ( n67250 , n67247 , n388083 );
buf ( n388085 , n67250 );
and ( n388086 , n388080 , n388085 );
not ( n388087 , n388080 );
buf ( n388088 , n387428 );
buf ( n388089 , n59764 );
nand ( n388090 , n388088 , n388089 );
buf ( n388091 , n388090 );
buf ( n388092 , n388091 );
and ( n388093 , n388087 , n388092 );
nor ( n67260 , n388086 , n388093 );
buf ( n388095 , n67260 );
xor ( n388096 , n388079 , n388095 );
buf ( n388097 , n45553 );
not ( n67264 , n388097 );
buf ( n388099 , n66566 );
not ( n67266 , n388099 );
or ( n67267 , n67264 , n67266 );
xnor ( n388102 , n362534 , n365670 );
buf ( n388103 , n388102 );
buf ( n388104 , n56794 );
nand ( n388105 , n388103 , n388104 );
buf ( n388106 , n388105 );
buf ( n388107 , n388106 );
nand ( n67274 , n67267 , n388107 );
buf ( n388109 , n67274 );
xor ( n67276 , n388096 , n388109 );
not ( n67277 , n44915 );
buf ( n388112 , n365041 );
not ( n67279 , n388112 );
buf ( n388114 , n369722 );
not ( n388115 , n388114 );
or ( n67282 , n67279 , n388115 );
buf ( n388117 , n362458 );
buf ( n388118 , n365052 );
nand ( n388119 , n388117 , n388118 );
buf ( n388120 , n388119 );
buf ( n388121 , n388120 );
nand ( n67288 , n67282 , n388121 );
buf ( n388123 , n67288 );
not ( n388124 , n388123 );
or ( n388125 , n67277 , n388124 );
buf ( n388126 , n387506 );
buf ( n388127 , n47466 );
nand ( n388128 , n388126 , n388127 );
buf ( n388129 , n388128 );
nand ( n67296 , n388125 , n388129 );
not ( n67297 , n67296 );
xor ( n388132 , n67276 , n67297 );
or ( n388133 , n387742 , n387759 );
nand ( n67300 , n388133 , n66906 );
buf ( n388135 , n387742 );
buf ( n388136 , n387759 );
nand ( n67303 , n388135 , n388136 );
buf ( n67304 , n67303 );
nand ( n388139 , n67300 , n67304 );
xor ( n67306 , n388132 , n388139 );
buf ( n388141 , n67306 );
buf ( n67308 , n387513 );
not ( n67309 , n67308 );
buf ( n388144 , n387538 );
not ( n67311 , n388144 );
or ( n67312 , n67309 , n67311 );
buf ( n388147 , n387538 );
buf ( n388148 , n387513 );
or ( n388149 , n388147 , n388148 );
buf ( n388150 , n387566 );
nand ( n67317 , n388149 , n388150 );
buf ( n388152 , n67317 );
buf ( n388153 , n388152 );
nand ( n67320 , n67312 , n388153 );
buf ( n67321 , n67320 );
buf ( n388156 , n67321 );
xor ( n67323 , n388141 , n388156 );
xor ( n388158 , n387634 , n387662 );
and ( n388159 , n388158 , n387763 );
and ( n67326 , n387634 , n387662 );
or ( n388161 , n388159 , n67326 );
buf ( n388162 , n388161 );
buf ( n388163 , n388162 );
xor ( n67330 , n67323 , n388163 );
buf ( n388165 , n67330 );
xor ( n67332 , n67236 , n388165 );
not ( n388167 , n387624 );
not ( n67334 , n387610 );
or ( n67335 , n388167 , n67334 );
not ( n388170 , n66796 );
not ( n67337 , n387625 );
or ( n388172 , n388170 , n67337 );
nand ( n67339 , n388172 , n387595 );
nand ( n67340 , n67335 , n67339 );
buf ( n67341 , n387591 );
not ( n67342 , n67341 );
buf ( n67343 , n39701 );
not ( n67344 , n67343 );
or ( n67345 , n67342 , n67344 );
buf ( n67346 , n367796 );
buf ( n388181 , n377143 );
not ( n67348 , n388181 );
buf ( n388183 , n366537 );
not ( n388184 , n388183 );
or ( n67351 , n67348 , n388184 );
buf ( n388186 , n366534 );
buf ( n388187 , n377146 );
nand ( n67354 , n388186 , n388187 );
buf ( n388189 , n67354 );
buf ( n388190 , n388189 );
nand ( n388191 , n67351 , n388190 );
buf ( n388192 , n388191 );
buf ( n388193 , n388192 );
nand ( n388194 , n67346 , n388193 );
buf ( n388195 , n388194 );
buf ( n388196 , n388195 );
nand ( n67363 , n67345 , n388196 );
buf ( n388198 , n67363 );
not ( n67365 , n368290 );
not ( n388200 , n66835 );
or ( n67367 , n67365 , n388200 );
buf ( n388202 , n56970 );
not ( n67369 , n388202 );
buf ( n388204 , n370845 );
not ( n388205 , n388204 );
or ( n388206 , n67369 , n388205 );
buf ( n388207 , n365507 );
buf ( n388208 , n377389 );
nand ( n388209 , n388207 , n388208 );
buf ( n388210 , n388209 );
buf ( n388211 , n388210 );
nand ( n67378 , n388206 , n388211 );
buf ( n388213 , n67378 );
buf ( n388214 , n388213 );
buf ( n388215 , n365954 );
nand ( n67382 , n388214 , n388215 );
buf ( n67383 , n67382 );
nand ( n67384 , n67367 , n67383 );
xor ( n67385 , n388198 , n67384 );
buf ( n388220 , n366986 );
not ( n67387 , n388220 );
buf ( n388222 , n66940 );
not ( n67389 , n388222 );
and ( n388224 , n67387 , n67389 );
buf ( n388225 , n46188 );
buf ( n388226 , n57053 );
buf ( n388227 , n365367 );
and ( n388228 , n388226 , n388227 );
not ( n67395 , n388226 );
buf ( n388230 , n355579 );
and ( n388231 , n67395 , n388230 );
nor ( n67398 , n388228 , n388231 );
buf ( n67399 , n67398 );
buf ( n388234 , n67399 );
nor ( n67401 , n388225 , n388234 );
buf ( n388236 , n67401 );
buf ( n388237 , n388236 );
nor ( n67404 , n388224 , n388237 );
buf ( n388239 , n67404 );
and ( n67406 , n67385 , n388239 );
not ( n388241 , n67385 );
buf ( n388242 , n388239 );
not ( n67409 , n388242 );
buf ( n388244 , n67409 );
and ( n388245 , n388241 , n388244 );
nor ( n67412 , n67406 , n388245 );
not ( n388247 , n67412 );
xor ( n388248 , n67340 , n388247 );
buf ( n388249 , n368549 );
not ( n388250 , n388249 );
buf ( n67417 , n363391 );
not ( n67418 , n67417 );
or ( n67419 , n388250 , n67418 );
buf ( n67420 , n368554 );
buf ( n67421 , n363388 );
nand ( n67422 , n67420 , n67421 );
buf ( n67423 , n67422 );
buf ( n67424 , n67423 );
nand ( n67425 , n67419 , n67424 );
buf ( n67426 , n67425 );
buf ( n67427 , n67426 );
not ( n67428 , n67427 );
buf ( n388263 , n67428 );
not ( n67430 , n388263 );
not ( n67431 , n368624 );
and ( n67432 , n67430 , n67431 );
and ( n67433 , n387556 , n368611 );
nor ( n388268 , n67432 , n67433 );
not ( n67435 , n388268 );
xnor ( n388270 , n388248 , n67435 );
buf ( n388271 , n388270 );
not ( n67438 , n388271 );
buf ( n388273 , n67438 );
buf ( n388274 , n388273 );
not ( n67441 , n388274 );
not ( n67442 , n365152 );
not ( n388277 , n362285 );
not ( n67444 , n342909 );
or ( n67445 , n388277 , n67444 );
nand ( n388280 , n362288 , n46397 );
nand ( n388281 , n67445 , n388280 );
not ( n67448 , n388281 );
or ( n67449 , n67442 , n67448 );
buf ( n388284 , n66546 );
buf ( n67451 , n65565 );
buf ( n67452 , n67451 );
nand ( n67453 , n388284 , n67452 );
buf ( n67454 , n67453 );
nand ( n388289 , n67449 , n67454 );
buf ( n388290 , n388289 );
xor ( n388291 , n66825 , n387654 );
and ( n388292 , n388291 , n387660 );
and ( n67459 , n66825 , n387654 );
or ( n67460 , n388292 , n67459 );
buf ( n388295 , n67460 );
xor ( n388296 , n388290 , n388295 );
xor ( n67463 , n387687 , n387704 );
and ( n388298 , n67463 , n66905 );
and ( n67465 , n387687 , n387704 );
or ( n67466 , n388298 , n67465 );
not ( n388301 , n366751 );
not ( n388302 , n365393 );
not ( n67469 , n365468 );
or ( n388304 , n388302 , n67469 );
buf ( n388305 , n360610 );
buf ( n388306 , n365408 );
nand ( n388307 , n388305 , n388306 );
buf ( n388308 , n388307 );
nand ( n67475 , n388304 , n388308 );
not ( n388310 , n67475 );
or ( n67477 , n388301 , n388310 );
nand ( n67478 , n387735 , n46557 );
nand ( n67479 , n67477 , n67478 );
xor ( n67480 , n67466 , n67479 );
nand ( n388315 , n387622 , n365033 );
buf ( n388316 , n364978 );
not ( n388317 , n388316 );
buf ( n388318 , n41528 );
not ( n388319 , n388318 );
or ( n67486 , n388317 , n388319 );
buf ( n388321 , n372889 );
buf ( n388322 , n364978 );
or ( n67489 , n388321 , n388322 );
buf ( n388324 , n67489 );
buf ( n388325 , n388324 );
nand ( n67492 , n67486 , n388325 );
buf ( n67493 , n67492 );
buf ( n388328 , n67493 );
buf ( n388329 , n365115 );
nand ( n388330 , n388328 , n388329 );
buf ( n388331 , n388330 );
nand ( n67498 , n388315 , n388331 );
xor ( n67499 , n67480 , n67498 );
buf ( n388334 , n67499 );
xor ( n388335 , n388296 , n388334 );
buf ( n388336 , n388335 );
buf ( n388337 , n388336 );
not ( n388338 , n388337 );
buf ( n388339 , n388338 );
buf ( n388340 , n388339 );
not ( n67507 , n388340 );
or ( n388342 , n67441 , n67507 );
nand ( n67509 , n388336 , n388270 );
buf ( n388344 , n67509 );
nand ( n67511 , n388342 , n388344 );
buf ( n388346 , n67511 );
buf ( n388347 , n388346 );
buf ( n388348 , n67028 );
not ( n67515 , n388348 );
buf ( n388350 , n67018 );
nand ( n388351 , n67515 , n388350 );
buf ( n388352 , n388351 );
buf ( n388353 , n388352 );
not ( n388354 , n388353 );
buf ( n388355 , n387824 );
not ( n67522 , n388355 );
or ( n388357 , n388354 , n67522 );
buf ( n388358 , n67018 );
not ( n388359 , n388358 );
buf ( n67526 , n67028 );
nand ( n67527 , n388359 , n67526 );
buf ( n67528 , n67527 );
buf ( n67529 , n67528 );
nand ( n67530 , n388357 , n67529 );
buf ( n67531 , n67530 );
buf ( n67532 , n67531 );
not ( n388367 , n67532 );
buf ( n388368 , n388367 );
buf ( n388369 , n388368 );
and ( n67536 , n388347 , n388369 );
not ( n388371 , n388347 );
buf ( n388372 , n67531 );
and ( n67539 , n388371 , n388372 );
nor ( n388374 , n67536 , n67539 );
buf ( n388375 , n388374 );
xor ( n67542 , n67332 , n388375 );
not ( n388377 , n67542 );
not ( n388378 , n388377 );
and ( n67545 , n67221 , n388378 );
not ( n67546 , n67221 );
and ( n67547 , n67546 , n388377 );
nor ( n388382 , n67545 , n67547 );
not ( n388383 , n388382 );
not ( n67550 , n66994 );
nand ( n67551 , n67550 , n67034 );
not ( n67552 , n67551 );
not ( n388387 , n387818 );
or ( n388388 , n67552 , n388387 );
buf ( n388389 , n67034 );
not ( n388390 , n388389 );
buf ( n388391 , n66994 );
nand ( n388392 , n388390 , n388391 );
buf ( n388393 , n388392 );
nand ( n67560 , n388388 , n388393 );
buf ( n388395 , n67560 );
not ( n388396 , n387297 );
not ( n67563 , n388396 );
not ( n388398 , n387239 );
or ( n67565 , n67563 , n388398 );
not ( n67566 , n66421 );
not ( n388401 , n387297 );
or ( n67568 , n67566 , n388401 );
nand ( n388403 , n67568 , n387291 );
nand ( n67570 , n67565 , n388403 );
buf ( n388405 , n67570 );
xor ( n388406 , n388395 , n388405 );
buf ( n388407 , n387159 );
not ( n388408 , n388407 );
buf ( n388409 , n386445 );
not ( n67576 , n388409 );
or ( n388411 , n388408 , n67576 );
buf ( n388412 , n368038 );
buf ( n388413 , n377782 );
not ( n388414 , n388413 );
buf ( n388415 , n364909 );
not ( n388416 , n388415 );
or ( n388417 , n388414 , n388416 );
buf ( n388418 , n361762 );
buf ( n388419 , n377779 );
nand ( n388420 , n388418 , n388419 );
buf ( n388421 , n388420 );
buf ( n388422 , n388421 );
nand ( n388423 , n388417 , n388422 );
buf ( n388424 , n388423 );
buf ( n388425 , n388424 );
nand ( n388426 , n388412 , n388425 );
buf ( n388427 , n388426 );
buf ( n388428 , n388427 );
nand ( n67581 , n388411 , n388428 );
buf ( n388430 , n67581 );
buf ( n388431 , n388430 );
not ( n67584 , n363429 );
not ( n67585 , n387677 );
or ( n67586 , n67584 , n67585 );
buf ( n388435 , n55539 );
not ( n67588 , n388435 );
buf ( n388437 , n44637 );
not ( n67590 , n388437 );
or ( n388439 , n67588 , n67590 );
buf ( n388440 , n364808 );
buf ( n388441 , n381286 );
nand ( n388442 , n388440 , n388441 );
buf ( n388443 , n388442 );
buf ( n388444 , n388443 );
nand ( n388445 , n388439 , n388444 );
buf ( n388446 , n388445 );
buf ( n388447 , n388446 );
buf ( n388448 , n378183 );
nand ( n388449 , n388447 , n388448 );
buf ( n388450 , n388449 );
nand ( n67603 , n67586 , n388450 );
not ( n388452 , n67603 );
buf ( n388453 , n365440 );
not ( n67606 , n388453 );
buf ( n388455 , n364763 );
not ( n67608 , n388455 );
or ( n67609 , n67606 , n67608 );
buf ( n388458 , n366329 );
buf ( n388459 , n386837 );
nand ( n67612 , n388458 , n388459 );
buf ( n388461 , n67612 );
buf ( n388462 , n388461 );
nand ( n388463 , n67609 , n388462 );
buf ( n388464 , n388463 );
buf ( n388465 , n388464 );
buf ( n388466 , n365311 );
nand ( n67619 , n388465 , n388466 );
buf ( n388468 , n67619 );
nand ( n388469 , n387182 , n366315 );
nand ( n67622 , n388468 , n388469 );
xor ( n388471 , n388452 , n67622 );
not ( n67624 , n366025 );
not ( n67625 , n66793 );
or ( n67626 , n67624 , n67625 );
buf ( n388475 , n365303 );
buf ( n388476 , n365980 );
not ( n388477 , n388476 );
buf ( n388478 , n365290 );
not ( n67631 , n388478 );
or ( n388480 , n388477 , n67631 );
buf ( n388481 , n45091 );
buf ( n388482 , n365989 );
nand ( n67635 , n388481 , n388482 );
buf ( n388484 , n67635 );
buf ( n388485 , n388484 );
nand ( n67638 , n388480 , n388485 );
buf ( n388487 , n67638 );
buf ( n388488 , n388487 );
nand ( n67641 , n388475 , n388488 );
buf ( n388490 , n67641 );
nand ( n67643 , n67626 , n388490 );
xor ( n67644 , n388471 , n67643 );
buf ( n388493 , n67644 );
xor ( n67646 , n388431 , n388493 );
xor ( n388495 , n387389 , n387407 );
and ( n388496 , n388495 , n387436 );
and ( n67649 , n387389 , n387407 );
or ( n67650 , n388496 , n67649 );
buf ( n388499 , n67650 );
buf ( n388500 , n388499 );
xor ( n388501 , n67646 , n388500 );
buf ( n388502 , n388501 );
buf ( n388503 , n388502 );
not ( n67656 , n388503 );
not ( n67657 , n379912 );
not ( n67658 , n387249 );
or ( n67659 , n67657 , n67658 );
not ( n388508 , n379893 );
buf ( n388509 , n379841 );
not ( n67662 , n388509 );
buf ( n388511 , n363439 );
not ( n388512 , n388511 );
or ( n67665 , n67662 , n388512 );
buf ( n388514 , n48344 );
buf ( n388515 , n379847 );
nand ( n67668 , n388514 , n388515 );
buf ( n67669 , n67668 );
buf ( n388518 , n67669 );
nand ( n67671 , n67665 , n388518 );
buf ( n388520 , n67671 );
nand ( n388521 , n388508 , n388520 );
nand ( n67674 , n67659 , n388521 );
not ( n67675 , n67674 );
buf ( n388524 , n67675 );
not ( n67677 , n388524 );
or ( n388526 , n67656 , n67677 );
buf ( n388527 , n67675 );
buf ( n388528 , n388502 );
or ( n388529 , n388527 , n388528 );
nand ( n388530 , n388526 , n388529 );
buf ( n388531 , n388530 );
xor ( n388532 , n66636 , n66642 );
and ( n388533 , n388532 , n66647 );
and ( n67686 , n66636 , n66642 );
or ( n388535 , n388533 , n67686 );
xor ( n388536 , n388531 , n388535 );
not ( n67689 , n387121 );
nand ( n388538 , n67689 , n387140 );
not ( n67691 , n388538 );
not ( n67692 , n66420 );
or ( n388541 , n67691 , n67692 );
buf ( n388542 , n387137 );
buf ( n388543 , n387121 );
nand ( n388544 , n388542 , n388543 );
buf ( n388545 , n388544 );
nand ( n67698 , n388541 , n388545 );
buf ( n388547 , n67698 );
not ( n67700 , n366399 );
not ( n67701 , n387209 );
or ( n67702 , n67700 , n67701 );
buf ( n388551 , n342656 );
not ( n67704 , n388551 );
buf ( n388553 , n364855 );
not ( n67706 , n388553 );
or ( n388555 , n67704 , n67706 );
buf ( n388556 , n351367 );
buf ( n388557 , n58471 );
nand ( n388558 , n388556 , n388557 );
buf ( n388559 , n388558 );
buf ( n388560 , n388559 );
nand ( n388561 , n388555 , n388560 );
buf ( n388562 , n388561 );
nand ( n388563 , n366428 , n388562 );
nand ( n67716 , n67702 , n388563 );
not ( n67717 , n67716 );
buf ( n388566 , n46521 );
not ( n67719 , n388566 );
buf ( n388568 , n387697 );
not ( n67721 , n388568 );
or ( n67722 , n67719 , n67721 );
nand ( n67723 , n46477 , n364771 );
not ( n67724 , n67723 );
buf ( n67725 , n368700 );
buf ( n388574 , n375901 );
not ( n67727 , n388574 );
buf ( n388576 , n67727 );
buf ( n388577 , n388576 );
nand ( n388578 , n67725 , n388577 );
buf ( n388579 , n388578 );
not ( n67732 , n388579 );
or ( n388581 , n67724 , n67732 );
nand ( n388582 , n388581 , n46463 );
buf ( n388583 , n388582 );
nand ( n388584 , n67722 , n388583 );
buf ( n388585 , n388584 );
not ( n388586 , n388585 );
xor ( n388587 , n67717 , n388586 );
buf ( n388588 , n368777 );
buf ( n388589 , n387717 );
or ( n388590 , n388588 , n388589 );
buf ( n388591 , n45592 );
not ( n388592 , n388591 );
buf ( n388593 , n386359 );
not ( n67746 , n388593 );
and ( n67747 , n388592 , n67746 );
buf ( n388596 , n377712 );
buf ( n388597 , n365259 );
and ( n67750 , n388596 , n388597 );
nor ( n67751 , n67747 , n67750 );
buf ( n388600 , n67751 );
buf ( n388601 , n388600 );
not ( n67754 , n377842 );
buf ( n388603 , n67754 );
or ( n67756 , n388601 , n388603 );
nand ( n388605 , n388590 , n67756 );
buf ( n388606 , n388605 );
not ( n388607 , n388606 );
xor ( n67759 , n388587 , n388607 );
buf ( n388609 , n387214 );
buf ( n388610 , n386380 );
nand ( n67762 , n388609 , n388610 );
buf ( n388612 , n67762 );
not ( n67764 , n388612 );
not ( n67765 , n387189 );
or ( n67766 , n67764 , n67765 );
or ( n67767 , n387214 , n386380 );
nand ( n67768 , n67766 , n67767 );
not ( n67769 , n67768 );
xor ( n67770 , n67759 , n67769 );
not ( n67771 , n45075 );
buf ( n388621 , n363317 );
buf ( n388622 , n45060 );
and ( n67774 , n388621 , n388622 );
buf ( n388624 , n367459 );
buf ( n388625 , n365202 );
and ( n67777 , n388624 , n388625 );
nor ( n67778 , n67774 , n67777 );
buf ( n388628 , n67778 );
not ( n67780 , n388628 );
not ( n67781 , n67780 );
or ( n67782 , n67771 , n67781 );
nand ( n67783 , n387339 , n365226 );
nand ( n67784 , n67782 , n67783 );
not ( n67785 , n67784 );
xor ( n67786 , n67770 , n67785 );
not ( n67787 , n67786 );
not ( n388637 , n67787 );
not ( n388638 , n49609 );
not ( n388639 , n359778 );
not ( n388640 , n369766 );
or ( n67792 , n388639 , n388640 );
nand ( n388642 , n364987 , n369769 );
nand ( n67794 , n67792 , n388642 );
not ( n388644 , n67794 );
or ( n388645 , n388638 , n388644 );
buf ( n388646 , n387531 );
buf ( n388647 , n369804 );
nand ( n67799 , n388646 , n388647 );
buf ( n388649 , n67799 );
nand ( n388650 , n388645 , n388649 );
not ( n67802 , n388650 );
not ( n67803 , n67802 );
or ( n67804 , n388637 , n67803 );
buf ( n388654 , n67786 );
buf ( n388655 , n388650 );
nand ( n388656 , n388654 , n388655 );
buf ( n388657 , n388656 );
nand ( n388658 , n67804 , n388657 );
not ( n388659 , n387165 );
nand ( n388660 , n388659 , n387225 );
not ( n388661 , n388660 );
not ( n388662 , n387234 );
or ( n388663 , n388661 , n388662 );
not ( n388664 , n387225 );
nand ( n388665 , n388664 , n387165 );
nand ( n388666 , n388663 , n388665 );
not ( n388667 , n388666 );
and ( n388668 , n388658 , n388667 );
not ( n388669 , n388658 );
and ( n388670 , n388669 , n388666 );
nor ( n388671 , n388668 , n388670 );
buf ( n388672 , n388671 );
not ( n388673 , n388672 );
buf ( n388674 , n388673 );
buf ( n388675 , n388674 );
and ( n388676 , n388547 , n388675 );
not ( n388677 , n388547 );
buf ( n388678 , n388671 );
and ( n388679 , n388677 , n388678 );
nor ( n388680 , n388676 , n388679 );
buf ( n388681 , n388680 );
xor ( n67808 , n388536 , n388681 );
buf ( n388683 , n67808 );
xor ( n388684 , n388406 , n388683 );
buf ( n388685 , n388684 );
buf ( n388686 , n388685 );
xor ( n67810 , n387789 , n387801 );
and ( n388688 , n67810 , n387851 );
and ( n388689 , n387789 , n387801 );
or ( n388690 , n388688 , n388689 );
buf ( n388691 , n388690 );
buf ( n388692 , n388691 );
and ( n388693 , n388686 , n388692 );
not ( n388694 , n388686 );
buf ( n388695 , n388691 );
not ( n388696 , n388695 );
buf ( n388697 , n388696 );
buf ( n388698 , n388697 );
and ( n388699 , n388694 , n388698 );
nor ( n388700 , n388693 , n388699 );
buf ( n388701 , n388700 );
not ( n388702 , n388701 );
and ( n388703 , n388383 , n388702 );
not ( n388704 , n388383 );
and ( n388705 , n388704 , n388701 );
nor ( n388706 , n388703 , n388705 );
buf ( n388707 , n388706 );
xor ( n388708 , n387950 , n388707 );
buf ( n388709 , n388708 );
not ( n67814 , n388709 );
xor ( n388711 , n387317 , n387325 );
and ( n67816 , n388711 , n387894 );
and ( n388713 , n387317 , n387325 );
or ( n67818 , n67816 , n388713 );
not ( n388715 , n67818 );
and ( n67820 , n67814 , n388715 );
nor ( n388717 , n387922 , n67820 );
nand ( n67822 , n67098 , n387919 , n388717 );
not ( n67823 , n67822 );
buf ( n388720 , n67130 );
not ( n388721 , n388720 );
buf ( n388722 , n379296 );
not ( n388723 , n388722 );
and ( n388724 , n388721 , n388723 );
not ( n67829 , n379274 );
not ( n388726 , n41472 );
or ( n388727 , n67829 , n388726 );
buf ( n388728 , n40090 );
buf ( n388729 , n379271 );
nand ( n388730 , n388728 , n388729 );
buf ( n388731 , n388730 );
nand ( n67836 , n388727 , n388731 );
buf ( n388733 , n67836 );
buf ( n388734 , n379263 );
and ( n67839 , n388733 , n388734 );
nor ( n388736 , n388724 , n67839 );
buf ( n388737 , n388736 );
not ( n67842 , n388737 );
not ( n388739 , n57530 );
not ( n67843 , n387993 );
or ( n388741 , n388739 , n67843 );
not ( n67845 , n377585 );
not ( n67846 , n372458 );
or ( n388744 , n67845 , n67846 );
nand ( n67848 , n386943 , n39867 );
nand ( n67849 , n388744 , n67848 );
nand ( n67850 , n67849 , n377580 );
nand ( n388748 , n388741 , n67850 );
not ( n67852 , n388748 );
or ( n67853 , n67842 , n67852 );
not ( n67854 , n388748 );
buf ( n388752 , n67854 );
buf ( n388753 , n388737 );
not ( n67857 , n388753 );
buf ( n388755 , n67857 );
buf ( n388756 , n388755 );
nand ( n67860 , n388752 , n388756 );
buf ( n388758 , n67860 );
nand ( n67862 , n67853 , n388758 );
buf ( n388760 , n388139 );
not ( n67864 , n388760 );
buf ( n388762 , n67276 );
not ( n67866 , n388762 );
buf ( n388764 , n67297 );
nand ( n67868 , n67866 , n388764 );
buf ( n388766 , n67868 );
buf ( n388767 , n388766 );
not ( n67871 , n388767 );
or ( n67872 , n67864 , n67871 );
buf ( n67873 , n67296 );
buf ( n67874 , n67276 );
nand ( n67875 , n67873 , n67874 );
buf ( n67876 , n67875 );
buf ( n388774 , n67876 );
nand ( n67878 , n67872 , n388774 );
buf ( n388776 , n67878 );
buf ( n67880 , n388776 );
not ( n388778 , n67880 );
buf ( n388779 , n388778 );
and ( n388780 , n67862 , n388779 );
not ( n67884 , n67862 );
not ( n388782 , n388779 );
and ( n67886 , n67884 , n388782 );
nor ( n67887 , n388780 , n67886 );
not ( n67888 , n67643 );
nand ( n67889 , n388468 , n388469 , n67603 );
not ( n388787 , n67889 );
or ( n67891 , n67888 , n388787 );
buf ( n388789 , n67622 );
buf ( n388790 , n388452 );
nand ( n67894 , n388789 , n388790 );
buf ( n388792 , n67894 );
nand ( n67896 , n67891 , n388792 );
buf ( n388794 , n43261 );
not ( n67898 , n388794 );
buf ( n388796 , n369497 );
not ( n388797 , n388796 );
buf ( n388798 , n31073 );
not ( n67902 , n388798 );
or ( n388800 , n388797 , n67902 );
buf ( n388801 , n31072 );
buf ( n388802 , n342718 );
nand ( n67906 , n388801 , n388802 );
buf ( n67907 , n67906 );
buf ( n388805 , n67907 );
nand ( n67909 , n388800 , n388805 );
buf ( n388807 , n67909 );
buf ( n388808 , n388807 );
not ( n67912 , n388808 );
or ( n388810 , n67898 , n67912 );
buf ( n388811 , n388446 );
buf ( n67915 , n363429 );
nand ( n67916 , n388811 , n67915 );
buf ( n67917 , n67916 );
buf ( n67918 , n67917 );
nand ( n67919 , n388810 , n67918 );
buf ( n67920 , n67919 );
buf ( n388818 , n342656 );
not ( n388819 , n388818 );
buf ( n388820 , n365328 );
not ( n67924 , n388820 );
or ( n388822 , n388819 , n67924 );
buf ( n388823 , n58463 );
not ( n67927 , n388823 );
buf ( n388825 , n30911 );
nand ( n388826 , n67927 , n388825 );
buf ( n388827 , n388826 );
buf ( n388828 , n388827 );
nand ( n67932 , n388822 , n388828 );
buf ( n388830 , n67932 );
not ( n67934 , n388830 );
not ( n388832 , n377271 );
or ( n388833 , n67934 , n388832 );
buf ( n67937 , n388562 );
buf ( n67938 , n366399 );
nand ( n67939 , n67937 , n67938 );
buf ( n388837 , n67939 );
nand ( n67941 , n388833 , n388837 );
xor ( n388839 , n67920 , n67941 );
not ( n388840 , n368706 );
not ( n67944 , n388600 );
not ( n67945 , n67944 );
or ( n67946 , n388840 , n67945 );
buf ( n388844 , n377712 );
not ( n388845 , n388844 );
buf ( n388846 , n45125 );
not ( n67950 , n388846 );
or ( n388848 , n388845 , n67950 );
buf ( n388849 , n342335 );
buf ( n388850 , n352192 );
nand ( n388851 , n388849 , n388850 );
buf ( n388852 , n388851 );
buf ( n388853 , n388852 );
nand ( n388854 , n388848 , n388853 );
buf ( n388855 , n388854 );
nand ( n388856 , n388855 , n48558 );
nand ( n388857 , n67946 , n388856 );
not ( n388858 , n388857 );
xor ( n388859 , n388839 , n388858 );
xor ( n388860 , n67896 , n388859 );
not ( n388861 , n388095 );
not ( n388862 , n388079 );
not ( n388863 , n388862 );
not ( n388864 , n388863 );
or ( n388865 , n388861 , n388864 );
buf ( n388866 , n388095 );
not ( n388867 , n388866 );
buf ( n388868 , n388867 );
buf ( n388869 , n388868 );
not ( n67954 , n388869 );
buf ( n388871 , n388862 );
not ( n67956 , n388871 );
or ( n67957 , n67954 , n67956 );
buf ( n388874 , n388109 );
nand ( n388875 , n67957 , n388874 );
buf ( n388876 , n388875 );
nand ( n67961 , n388865 , n388876 );
xnor ( n388878 , n388860 , n67961 );
buf ( n388879 , n388878 );
buf ( n67964 , n388424 );
not ( n67965 , n67964 );
buf ( n67966 , n386445 );
not ( n67967 , n67966 );
or ( n67968 , n67965 , n67967 );
or ( n388885 , n359947 , n377353 );
nand ( n388886 , n377353 , n359904 );
nand ( n67971 , n388885 , n388886 );
nand ( n388888 , n67971 , n359993 );
buf ( n67973 , n388888 );
nand ( n67974 , n67968 , n67973 );
buf ( n67975 , n67974 );
buf ( n388892 , n67975 );
buf ( n388893 , n365115 );
not ( n388894 , n388893 );
buf ( n388895 , n44819 );
not ( n67980 , n388895 );
buf ( n388897 , n41615 );
not ( n388898 , n388897 );
or ( n67983 , n67980 , n388898 );
buf ( n388900 , n41607 );
buf ( n388901 , n364994 );
nand ( n67986 , n388900 , n388901 );
buf ( n67987 , n67986 );
buf ( n388904 , n67987 );
nand ( n388905 , n67983 , n388904 );
buf ( n388906 , n388905 );
buf ( n67991 , n388906 );
not ( n67992 , n67991 );
or ( n67993 , n388894 , n67992 );
buf ( n67994 , n365033 );
buf ( n67995 , n67493 );
nand ( n67996 , n67994 , n67995 );
buf ( n67997 , n67996 );
buf ( n67998 , n67997 );
nand ( n67999 , n67993 , n67998 );
buf ( n68000 , n67999 );
buf ( n388917 , n68000 );
xor ( n68002 , n388892 , n388917 );
buf ( n388919 , n67603 );
buf ( n388920 , n388464 );
not ( n68005 , n388920 );
buf ( n388922 , n68005 );
not ( n388923 , n388922 );
not ( n68008 , n361971 );
and ( n388925 , n388923 , n68008 );
buf ( n388926 , n31260 );
not ( n68011 , n388926 );
buf ( n388928 , n364783 );
not ( n388929 , n388928 );
or ( n68014 , n68011 , n388929 );
buf ( n388931 , n361911 );
buf ( n388932 , n351292 );
nand ( n68017 , n388931 , n388932 );
buf ( n388934 , n68017 );
buf ( n388935 , n388934 );
nand ( n68020 , n68014 , n388935 );
buf ( n68021 , n68020 );
buf ( n388938 , n68021 );
buf ( n388939 , n41834 );
and ( n388940 , n388938 , n388939 );
buf ( n388941 , n388940 );
nor ( n68026 , n388925 , n388941 );
buf ( n388943 , n68026 );
xor ( n388944 , n388919 , n388943 );
not ( n388945 , n67239 );
not ( n68030 , n386678 );
or ( n388947 , n388945 , n68030 );
buf ( n388948 , n371063 );
buf ( n388949 , n365490 );
not ( n388950 , n388949 );
buf ( n388951 , n44634 );
not ( n388952 , n388951 );
or ( n68037 , n388950 , n388952 );
buf ( n388954 , n41892 );
buf ( n388955 , n45336 );
nand ( n388956 , n388954 , n388955 );
buf ( n388957 , n388956 );
buf ( n388958 , n388957 );
nand ( n388959 , n68037 , n388958 );
buf ( n388960 , n388959 );
buf ( n388961 , n388960 );
nand ( n388962 , n388948 , n388961 );
buf ( n388963 , n388962 );
nand ( n68048 , n388947 , n388963 );
buf ( n388965 , n68048 );
xnor ( n68050 , n388944 , n388965 );
buf ( n388967 , n68050 );
buf ( n388968 , n388967 );
xor ( n68053 , n68002 , n388968 );
buf ( n388970 , n68053 );
buf ( n388971 , n388970 );
xor ( n68056 , n388879 , n388971 );
buf ( n388973 , n49609 );
not ( n68058 , n388973 );
buf ( n388975 , n369769 );
not ( n68060 , n388975 );
buf ( n388977 , n40999 );
not ( n68062 , n388977 );
or ( n68063 , n68060 , n68062 );
buf ( n388980 , n359756 );
buf ( n388981 , n369766 );
nand ( n68066 , n388980 , n388981 );
buf ( n388983 , n68066 );
buf ( n388984 , n388983 );
nand ( n68069 , n68063 , n388984 );
buf ( n388986 , n68069 );
buf ( n388987 , n388986 );
not ( n68072 , n388987 );
or ( n388989 , n68058 , n68072 );
buf ( n388990 , n67794 );
buf ( n388991 , n369804 );
nand ( n388992 , n388990 , n388991 );
buf ( n388993 , n388992 );
buf ( n388994 , n388993 );
nand ( n388995 , n388989 , n388994 );
buf ( n388996 , n388995 );
buf ( n388997 , n388996 );
xnor ( n388998 , n68056 , n388997 );
buf ( n388999 , n388998 );
buf ( n389000 , n388999 );
not ( n68085 , n389000 );
buf ( n389002 , n68085 );
and ( n389003 , n67887 , n389002 );
not ( n389004 , n67887 );
and ( n68089 , n389004 , n388999 );
or ( n389006 , n389003 , n68089 );
buf ( n389007 , n389006 );
buf ( n389008 , n67321 );
not ( n389009 , n389008 );
buf ( n389010 , n389009 );
buf ( n389011 , n389010 );
not ( n68096 , n389011 );
buf ( n389013 , n67306 );
not ( n389014 , n389013 );
or ( n389015 , n68096 , n389014 );
buf ( n389016 , n388162 );
nand ( n389017 , n389015 , n389016 );
buf ( n389018 , n389017 );
buf ( n389019 , n389018 );
buf ( n389020 , n67306 );
not ( n389021 , n389020 );
buf ( n389022 , n67321 );
nand ( n389023 , n389021 , n389022 );
buf ( n389024 , n389023 );
buf ( n389025 , n389024 );
nand ( n389026 , n389019 , n389025 );
buf ( n389027 , n389026 );
buf ( n389028 , n389027 );
buf ( n389029 , n389028 );
buf ( n389030 , n389029 );
buf ( n389031 , n389030 );
xnor ( n389032 , n389007 , n389031 );
buf ( n389033 , n389032 );
buf ( n389034 , n389033 );
xor ( n389035 , n67236 , n388165 );
and ( n68120 , n389035 , n388375 );
and ( n68121 , n67236 , n388165 );
or ( n68122 , n68120 , n68121 );
buf ( n389039 , n68122 );
xor ( n68124 , n389034 , n389039 );
buf ( n389041 , n388273 );
not ( n68126 , n389041 );
buf ( n389043 , n388336 );
not ( n68128 , n389043 );
or ( n389045 , n68126 , n68128 );
buf ( n389046 , n388270 );
not ( n68131 , n389046 );
buf ( n389048 , n388339 );
not ( n68133 , n389048 );
or ( n389050 , n68131 , n68133 );
buf ( n389051 , n67531 );
nand ( n389052 , n389050 , n389051 );
buf ( n389053 , n389052 );
buf ( n389054 , n389053 );
nand ( n389055 , n389045 , n389054 );
buf ( n389056 , n389055 );
xor ( n68141 , n388290 , n388295 );
and ( n389058 , n68141 , n388334 );
and ( n68143 , n388290 , n388295 );
or ( n68144 , n389058 , n68143 );
buf ( n389061 , n68144 );
buf ( n389062 , n46303 );
not ( n68147 , n389062 );
buf ( n389064 , n365267 );
not ( n68149 , n389064 );
or ( n68150 , n68147 , n68149 );
buf ( n389067 , n365290 );
not ( n68152 , n389067 );
buf ( n389069 , n44737 );
nand ( n389070 , n68152 , n389069 );
buf ( n389071 , n389070 );
buf ( n389072 , n389071 );
nand ( n68157 , n68150 , n389072 );
buf ( n389074 , n68157 );
buf ( n389075 , n389074 );
buf ( n389076 , n40923 );
nand ( n68161 , n389075 , n389076 );
buf ( n389078 , n68161 );
nand ( n68163 , n388487 , n366025 );
nand ( n389080 , n389078 , n68163 );
not ( n389081 , n389080 );
not ( n68166 , n389081 );
buf ( n389083 , n366683 );
not ( n389084 , n389083 );
buf ( n389085 , n42355 );
not ( n389086 , n389085 );
or ( n389087 , n389084 , n389086 );
buf ( n389088 , n45916 );
not ( n68173 , n389088 );
buf ( n389090 , n46477 );
nand ( n389091 , n68173 , n389090 );
buf ( n389092 , n389091 );
buf ( n389093 , n389092 );
nand ( n389094 , n389087 , n389093 );
buf ( n389095 , n389094 );
buf ( n389096 , n389095 );
buf ( n389097 , n46463 );
and ( n389098 , n389096 , n389097 );
nand ( n389099 , n388579 , n67723 );
buf ( n389100 , n389099 );
buf ( n68185 , n46521 );
and ( n68186 , n389100 , n68185 );
buf ( n389103 , n68186 );
buf ( n389104 , n389103 );
nor ( n68189 , n389098 , n389104 );
buf ( n389106 , n68189 );
buf ( n389107 , n389106 );
not ( n389108 , n389107 );
buf ( n389109 , n389108 );
not ( n389110 , n389109 );
or ( n389111 , n68166 , n389110 );
buf ( n389112 , n389106 );
buf ( n389113 , n389080 );
nand ( n389114 , n389112 , n389113 );
buf ( n389115 , n389114 );
nand ( n68200 , n389111 , n389115 );
not ( n68201 , n366103 );
buf ( n389118 , n45177 );
not ( n389119 , n389118 );
buf ( n389120 , n366086 );
not ( n68205 , n389120 );
or ( n68206 , n389119 , n68205 );
nand ( n68207 , n45414 , n365344 );
buf ( n389124 , n68207 );
nand ( n68209 , n68206 , n389124 );
buf ( n389126 , n68209 );
not ( n68211 , n389126 );
not ( n68212 , n68211 );
or ( n68213 , n68201 , n68212 );
or ( n68214 , n67250 , n381423 );
nand ( n68215 , n68214 , n60867 );
nand ( n68216 , n68213 , n68215 );
not ( n68217 , n68216 );
and ( n389134 , n68200 , n68217 );
not ( n68219 , n68200 );
and ( n389136 , n68219 , n68216 );
nor ( n389137 , n389134 , n389136 );
buf ( n389138 , n389137 );
not ( n68223 , n45075 );
buf ( n389140 , n45060 );
not ( n389141 , n389140 );
buf ( n389142 , n362145 );
not ( n68227 , n389142 );
or ( n389144 , n389141 , n68227 );
buf ( n389145 , n362133 );
buf ( n389146 , n45065 );
nand ( n68231 , n389145 , n389146 );
buf ( n389148 , n68231 );
buf ( n389149 , n389148 );
nand ( n68234 , n389144 , n389149 );
buf ( n68235 , n68234 );
not ( n389152 , n68235 );
or ( n389153 , n68223 , n389152 );
buf ( n389154 , n388628 );
not ( n389155 , n389154 );
buf ( n389156 , n365226 );
nand ( n68241 , n389155 , n389156 );
buf ( n389158 , n68241 );
nand ( n389159 , n389153 , n389158 );
buf ( n389160 , n389159 );
and ( n389161 , n389138 , n389160 );
not ( n68246 , n389138 );
not ( n389163 , n389159 );
buf ( n389164 , n389163 );
and ( n68249 , n68246 , n389164 );
nor ( n389166 , n389161 , n68249 );
buf ( n389167 , n389166 );
buf ( n389168 , n389167 );
buf ( n389169 , n67384 );
buf ( n389170 , n388244 );
nand ( n68255 , n389169 , n389170 );
buf ( n389172 , n68255 );
buf ( n389173 , n67384 );
not ( n389174 , n389173 );
buf ( n389175 , n389174 );
buf ( n389176 , n389175 );
not ( n68261 , n389176 );
buf ( n389178 , n388239 );
not ( n389179 , n389178 );
or ( n68264 , n68261 , n389179 );
buf ( n389181 , n388198 );
nand ( n389182 , n68264 , n389181 );
buf ( n389183 , n389182 );
nand ( n68268 , n389172 , n389183 );
buf ( n389185 , n68268 );
and ( n389186 , n389168 , n389185 );
not ( n389187 , n389168 );
buf ( n389188 , n68268 );
not ( n68273 , n389188 );
buf ( n389190 , n68273 );
buf ( n389191 , n389190 );
and ( n68276 , n389187 , n389191 );
nor ( n68277 , n389186 , n68276 );
buf ( n389194 , n68277 );
xor ( n68279 , n389061 , n389194 );
not ( n68280 , n388268 );
not ( n68281 , n68280 );
not ( n68282 , n67340 );
or ( n68283 , n68281 , n68282 );
buf ( n389200 , n67340 );
not ( n68285 , n389200 );
buf ( n389202 , n68285 );
not ( n68287 , n389202 );
not ( n389204 , n388268 );
or ( n389205 , n68287 , n389204 );
nand ( n68290 , n389205 , n388247 );
nand ( n68291 , n68283 , n68290 );
buf ( n389208 , n68291 );
xor ( n389209 , n68279 , n389208 );
xor ( n68294 , n389056 , n389209 );
buf ( n389211 , n68294 );
xor ( n389212 , n67466 , n67479 );
and ( n68297 , n389212 , n67498 );
and ( n389214 , n67466 , n67479 );
or ( n389215 , n68297 , n389214 );
buf ( n389216 , n368611 );
not ( n68301 , n389216 );
buf ( n389218 , n67426 );
not ( n389219 , n389218 );
or ( n389220 , n68301 , n389219 );
buf ( n389221 , n368549 );
not ( n389222 , n389221 );
buf ( n389223 , n45523 );
not ( n68308 , n389223 );
or ( n68309 , n389222 , n68308 );
buf ( n389226 , n40199 );
buf ( n389227 , n368554 );
nand ( n389228 , n389226 , n389227 );
buf ( n389229 , n389228 );
buf ( n389230 , n389229 );
nand ( n389231 , n68309 , n389230 );
buf ( n389232 , n389231 );
buf ( n389233 , n389232 );
buf ( n389234 , n369444 );
nand ( n389235 , n389233 , n389234 );
buf ( n389236 , n389235 );
buf ( n389237 , n389236 );
nand ( n68322 , n389220 , n389237 );
buf ( n389239 , n68322 );
xor ( n389240 , n389215 , n389239 );
buf ( n389241 , n388192 );
not ( n68326 , n389241 );
buf ( n389243 , n363038 );
not ( n389244 , n389243 );
or ( n68329 , n68326 , n389244 );
buf ( n389246 , n362521 );
buf ( n389247 , n378886 );
not ( n68332 , n389247 );
buf ( n389249 , n366534 );
not ( n389250 , n389249 );
or ( n68335 , n68332 , n389250 );
buf ( n389252 , n45231 );
buf ( n389253 , n377757 );
nand ( n389254 , n389252 , n389253 );
buf ( n389255 , n389254 );
buf ( n389256 , n389255 );
nand ( n389257 , n68335 , n389256 );
buf ( n389258 , n389257 );
buf ( n389259 , n389258 );
nand ( n68344 , n389246 , n389259 );
buf ( n68345 , n68344 );
buf ( n389262 , n68345 );
nand ( n389263 , n68329 , n389262 );
buf ( n389264 , n389263 );
not ( n68349 , n389264 );
buf ( n389266 , n388213 );
not ( n389267 , n389266 );
buf ( n389268 , n40058 );
not ( n68353 , n389268 );
or ( n389270 , n389267 , n68353 );
buf ( n389271 , n369374 );
not ( n389272 , n389271 );
buf ( n389273 , n370845 );
not ( n389274 , n389273 );
or ( n389275 , n389272 , n389274 );
buf ( n389276 , n363119 );
buf ( n389277 , n49178 );
nand ( n389278 , n389276 , n389277 );
buf ( n389279 , n389278 );
buf ( n389280 , n389279 );
nand ( n389281 , n389275 , n389280 );
buf ( n389282 , n389281 );
buf ( n68367 , n389282 );
buf ( n389284 , n39949 );
nand ( n389285 , n68367 , n389284 );
buf ( n389286 , n389285 );
buf ( n389287 , n389286 );
nand ( n68372 , n389270 , n389287 );
buf ( n389289 , n68372 );
not ( n389290 , n389289 );
xor ( n68375 , n67717 , n388586 );
and ( n389292 , n68375 , n388607 );
and ( n389293 , n67717 , n388586 );
or ( n68378 , n389292 , n389293 );
nand ( n68379 , n68349 , n389290 , n68378 );
not ( n389296 , n68349 );
nor ( n389297 , n389289 , n68378 );
nand ( n68382 , n389296 , n389297 );
not ( n389299 , n68349 );
nand ( n389300 , n389299 , n389289 , n68378 );
not ( n389301 , n68378 );
nand ( n68386 , n389289 , n68349 , n389301 );
nand ( n68387 , n68379 , n68382 , n389300 , n68386 );
and ( n389304 , n389240 , n68387 );
not ( n389305 , n389240 );
not ( n68390 , n68387 );
and ( n68391 , n389305 , n68390 );
nor ( n68392 , n389304 , n68391 );
not ( n389309 , n68392 );
buf ( n389310 , n67451 );
not ( n68395 , n389310 );
buf ( n389312 , n388281 );
not ( n68397 , n389312 );
or ( n389314 , n68395 , n68397 );
buf ( n389315 , n46397 );
not ( n68400 , n389315 );
buf ( n389317 , n373463 );
not ( n68402 , n389317 );
or ( n389319 , n68400 , n68402 );
buf ( n389320 , n360885 );
buf ( n389321 , n342909 );
nand ( n68406 , n389320 , n389321 );
buf ( n389323 , n68406 );
buf ( n389324 , n389323 );
nand ( n68409 , n389319 , n389324 );
buf ( n389326 , n68409 );
buf ( n389327 , n389326 );
buf ( n389328 , n365152 );
nand ( n68413 , n389327 , n389328 );
buf ( n389330 , n68413 );
buf ( n389331 , n389330 );
nand ( n68416 , n389314 , n389331 );
buf ( n389333 , n68416 );
buf ( n389334 , n388123 );
not ( n68419 , n389334 );
buf ( n389336 , n68419 );
buf ( n389337 , n389336 );
not ( n389338 , n389337 );
buf ( n389339 , n44913 );
not ( n68424 , n389339 );
and ( n389341 , n389338 , n68424 );
and ( n389342 , n40251 , n365052 );
not ( n68427 , n40251 );
and ( n389344 , n68427 , n365041 );
or ( n389345 , n389342 , n389344 );
buf ( n389346 , n389345 );
buf ( n389347 , n44915 );
and ( n389348 , n389346 , n389347 );
nor ( n389349 , n389341 , n389348 );
buf ( n389350 , n389349 );
xor ( n389351 , n389333 , n389350 );
buf ( n389352 , n365676 );
not ( n68437 , n389352 );
buf ( n389354 , n43377 );
not ( n68439 , n389354 );
or ( n68440 , n68437 , n68439 );
buf ( n389357 , n361716 );
buf ( n389358 , n365673 );
nand ( n389359 , n389357 , n389358 );
buf ( n389360 , n389359 );
buf ( n389361 , n389360 );
nand ( n68446 , n68440 , n389361 );
buf ( n389363 , n68446 );
buf ( n389364 , n389363 );
buf ( n389365 , n45492 );
and ( n68450 , n389364 , n389365 );
buf ( n389367 , n388102 );
not ( n389368 , n389367 );
buf ( n389369 , n366732 );
nor ( n68454 , n389368 , n389369 );
buf ( n389371 , n68454 );
buf ( n389372 , n389371 );
nor ( n68457 , n68450 , n389372 );
buf ( n389374 , n68457 );
not ( n389375 , n389374 );
buf ( n389376 , n67399 );
not ( n68461 , n389376 );
buf ( n389378 , n68461 );
not ( n68463 , n389378 );
not ( n389380 , n369260 );
or ( n68465 , n68463 , n389380 );
not ( n68466 , n368665 );
not ( n389383 , n359297 );
or ( n389384 , n68466 , n389383 );
nand ( n389385 , n51966 , n368662 );
nand ( n389386 , n389384 , n389385 );
nand ( n68471 , n389386 , n359312 );
nand ( n389388 , n68465 , n68471 );
not ( n389389 , n389388 );
or ( n68474 , n389375 , n389389 );
not ( n68475 , n389388 );
not ( n389392 , n389374 );
nand ( n389393 , n68475 , n389392 );
nand ( n389394 , n68474 , n389393 );
not ( n68479 , n389394 );
not ( n389396 , n371732 );
not ( n389397 , n366151 );
not ( n68482 , n365422 );
or ( n68483 , n389397 , n68482 );
nand ( n389400 , n365428 , n366277 );
nand ( n389401 , n68483 , n389400 );
not ( n68486 , n389401 );
or ( n389403 , n389396 , n68486 );
nand ( n68488 , n46113 , n67475 );
nand ( n389405 , n389403 , n68488 );
not ( n68490 , n389405 );
and ( n68491 , n68479 , n68490 );
and ( n389408 , n389394 , n389405 );
nor ( n389409 , n68491 , n389408 );
xor ( n68494 , n389351 , n389409 );
not ( n389411 , n68494 );
not ( n389412 , n389411 );
not ( n68497 , n67787 );
not ( n68498 , n388650 );
or ( n389415 , n68497 , n68498 );
not ( n389416 , n67802 );
not ( n389417 , n67786 );
or ( n68502 , n389416 , n389417 );
nand ( n68503 , n68502 , n388666 );
nand ( n389420 , n389415 , n68503 );
not ( n389421 , n389420 );
not ( n68506 , n389421 );
or ( n68507 , n389412 , n68506 );
nand ( n68508 , n68494 , n389420 );
nand ( n389425 , n68507 , n68508 );
not ( n389426 , n389425 );
or ( n68511 , n389309 , n389426 );
not ( n68512 , n389411 );
not ( n68513 , n389421 );
or ( n389430 , n68512 , n68513 );
nand ( n389431 , n389430 , n68508 );
buf ( n68516 , n68392 );
or ( n68517 , n389431 , n68516 );
nand ( n68518 , n68511 , n68517 );
buf ( n389435 , n68518 );
buf ( n389436 , n389435 );
not ( n68521 , n389436 );
buf ( n389438 , n68521 );
buf ( n389439 , n389438 );
and ( n389440 , n389211 , n389439 );
not ( n389441 , n389211 );
buf ( n389442 , n389435 );
and ( n68527 , n389441 , n389442 );
nor ( n389444 , n389440 , n68527 );
buf ( n389445 , n389444 );
buf ( n389446 , n389445 );
xor ( n68531 , n68124 , n389446 );
buf ( n389448 , n68531 );
not ( n68533 , n388046 );
not ( n68534 , n68533 );
not ( n389451 , n67542 );
or ( n68536 , n68534 , n389451 );
nand ( n68537 , n68536 , n388034 );
not ( n68538 , n68533 );
nand ( n68539 , n68538 , n388377 );
nand ( n68540 , n68537 , n68539 );
not ( n68541 , n68540 );
not ( n68542 , n67698 );
nand ( n68543 , n68542 , n388671 );
not ( n389460 , n68543 );
not ( n68545 , n388536 );
or ( n68546 , n389460 , n68545 );
buf ( n389463 , n67698 );
buf ( n389464 , n388674 );
nand ( n68549 , n389463 , n389464 );
buf ( n389466 , n68549 );
nand ( n68551 , n68546 , n389466 );
not ( n389468 , n68551 );
xor ( n68553 , n388431 , n388493 );
and ( n68554 , n68553 , n388500 );
and ( n68555 , n388431 , n388493 );
or ( n389472 , n68554 , n68555 );
buf ( n389473 , n389472 );
buf ( n389474 , n389473 );
not ( n68559 , n389474 );
buf ( n389476 , n68559 );
not ( n68561 , n67759 );
not ( n68562 , n67785 );
or ( n68563 , n68561 , n68562 );
nand ( n68564 , n68563 , n67768 );
not ( n68565 , n67759 );
not ( n68566 , n67785 );
nand ( n68567 , n68565 , n68566 );
nand ( n68568 , n68564 , n68567 );
not ( n68569 , n379893 );
not ( n68570 , n59424 );
or ( n68571 , n68569 , n68570 );
nand ( n68572 , n68571 , n388520 );
and ( n68573 , n68568 , n68572 );
not ( n68574 , n68568 );
not ( n389491 , n379893 );
not ( n68576 , n59424 );
or ( n68577 , n389491 , n68576 );
nand ( n68578 , n68577 , n388520 );
not ( n68579 , n68578 );
and ( n68580 , n68574 , n68579 );
nor ( n68581 , n68573 , n68580 );
or ( n68582 , n389476 , n68581 );
nand ( n68583 , n68581 , n389476 );
nand ( n68584 , n68582 , n68583 );
buf ( n389501 , n68584 );
not ( n68586 , n67165 );
not ( n68587 , n67141 );
or ( n68588 , n68586 , n68587 );
or ( n68589 , n67165 , n67141 );
nand ( n68590 , n68589 , n387966 );
nand ( n68591 , n68588 , n68590 );
buf ( n389508 , n68591 );
xor ( n68593 , n389501 , n389508 );
buf ( n389510 , n388502 );
not ( n389511 , n389510 );
buf ( n389512 , n389511 );
buf ( n389513 , n389512 );
not ( n68598 , n389513 );
buf ( n389515 , n67675 );
not ( n389516 , n389515 );
or ( n389517 , n68598 , n389516 );
buf ( n389518 , n388535 );
nand ( n389519 , n389517 , n389518 );
buf ( n389520 , n389519 );
buf ( n389521 , n389520 );
buf ( n389522 , n67675 );
not ( n389523 , n389522 );
buf ( n68608 , n388502 );
nand ( n68609 , n389523 , n68608 );
buf ( n68610 , n68609 );
buf ( n389527 , n68610 );
nand ( n68612 , n389521 , n389527 );
buf ( n68613 , n68612 );
buf ( n389530 , n68613 );
xor ( n68615 , n68593 , n389530 );
buf ( n389532 , n68615 );
not ( n68617 , n389532 );
not ( n68618 , n68617 );
or ( n68619 , n389468 , n68618 );
not ( n68620 , n68551 );
nand ( n389537 , n68620 , n389532 );
nand ( n68622 , n68619 , n389537 );
buf ( n389539 , n388004 );
not ( n68624 , n389539 );
buf ( n389541 , n68624 );
not ( n389542 , n389541 );
not ( n389543 , n388009 );
not ( n68628 , n389543 );
not ( n68629 , n68628 );
or ( n389546 , n389542 , n68629 );
buf ( n389547 , n388004 );
not ( n68632 , n389547 );
buf ( n389549 , n389543 );
not ( n389550 , n389549 );
or ( n389551 , n68632 , n389550 );
buf ( n389552 , n67197 );
nand ( n68637 , n389551 , n389552 );
buf ( n389554 , n68637 );
nand ( n68639 , n389546 , n389554 );
and ( n68640 , n68622 , n68639 );
not ( n389557 , n68622 );
not ( n68642 , n68639 );
and ( n68643 , n389557 , n68642 );
nor ( n68644 , n68640 , n68643 );
xor ( n68645 , n388395 , n388405 );
and ( n68646 , n68645 , n388683 );
and ( n68647 , n388395 , n388405 );
or ( n68648 , n68646 , n68647 );
buf ( n389565 , n68648 );
and ( n68650 , n68644 , n389565 );
not ( n389567 , n68644 );
buf ( n389568 , n389565 );
not ( n68653 , n389568 );
buf ( n389570 , n68653 );
and ( n68655 , n389567 , n389570 );
nor ( n389572 , n68650 , n68655 );
xor ( n389573 , n68541 , n389572 );
xor ( n68658 , n389448 , n389573 );
nand ( n389575 , n388685 , n388691 );
not ( n389576 , n389575 );
not ( n389577 , n388382 );
or ( n68662 , n389576 , n389577 );
or ( n389579 , n388691 , n388685 );
nand ( n68664 , n68662 , n389579 );
xor ( n68665 , n68658 , n68664 );
buf ( n68666 , n68665 );
not ( n389583 , n68666 );
buf ( n389584 , n389583 );
buf ( n389585 , n389584 );
xor ( n389586 , n387927 , n387949 );
and ( n68671 , n389586 , n388707 );
and ( n389588 , n387927 , n387949 );
or ( n389589 , n68671 , n389588 );
buf ( n389590 , n389589 );
buf ( n389591 , n389590 );
not ( n68676 , n389591 );
buf ( n389593 , n68676 );
buf ( n389594 , n389593 );
nand ( n389595 , n389585 , n389594 );
buf ( n389596 , n389595 );
not ( n389597 , n389596 );
xor ( n389598 , n389034 , n389039 );
and ( n68683 , n389598 , n389446 );
and ( n389600 , n389034 , n389039 );
or ( n389601 , n68683 , n389600 );
buf ( n389602 , n389601 );
buf ( n389603 , n389602 );
not ( n68688 , n68540 );
buf ( n389605 , n389570 );
not ( n68690 , n68644 );
buf ( n389607 , n68690 );
nand ( n68692 , n389605 , n389607 );
buf ( n389609 , n68692 );
not ( n389610 , n389609 );
or ( n389611 , n68688 , n389610 );
buf ( n389612 , n68690 );
buf ( n389613 , n389570 );
or ( n389614 , n389612 , n389613 );
buf ( n389615 , n389614 );
nand ( n389616 , n389611 , n389615 );
buf ( n389617 , n389616 );
not ( n68702 , n389617 );
buf ( n389619 , n68702 );
buf ( n389620 , n389619 );
xor ( n68705 , n389603 , n389620 );
buf ( n389622 , n68291 );
buf ( n389623 , n389194 );
or ( n68708 , n389622 , n389623 );
buf ( n389625 , n389061 );
nand ( n389626 , n68708 , n389625 );
buf ( n389627 , n389626 );
buf ( n389628 , n389627 );
buf ( n389629 , n68291 );
buf ( n389630 , n389194 );
nand ( n389631 , n389629 , n389630 );
buf ( n389632 , n389631 );
buf ( n68717 , n389632 );
nand ( n68718 , n389628 , n68717 );
buf ( n68719 , n68718 );
not ( n389636 , n68719 );
buf ( n389637 , n379299 );
not ( n389638 , n389637 );
buf ( n389639 , n67836 );
not ( n68724 , n389639 );
or ( n68725 , n389638 , n68724 );
not ( n68726 , n379271 );
not ( n389643 , n48344 );
or ( n68728 , n68726 , n389643 );
or ( n68729 , n48344 , n379271 );
nand ( n389646 , n68728 , n68729 );
nand ( n389647 , n389646 , n379263 );
buf ( n389648 , n389647 );
nand ( n389649 , n68725 , n389648 );
buf ( n389650 , n389649 );
buf ( n389651 , n389650 );
buf ( n389652 , n369804 );
not ( n68737 , n389652 );
buf ( n389654 , n388986 );
not ( n68739 , n389654 );
or ( n68740 , n68737 , n68739 );
buf ( n389657 , n369769 );
not ( n389658 , n389657 );
buf ( n389659 , n366600 );
not ( n68744 , n389659 );
or ( n389661 , n389658 , n68744 );
buf ( n389662 , n369766 );
buf ( n389663 , n39830 );
nand ( n389664 , n389662 , n389663 );
buf ( n68745 , n389664 );
buf ( n389666 , n68745 );
nand ( n389667 , n389661 , n389666 );
buf ( n389668 , n389667 );
buf ( n389669 , n389668 );
buf ( n389670 , n49609 );
nand ( n68750 , n389669 , n389670 );
buf ( n389672 , n68750 );
buf ( n389673 , n389672 );
nand ( n389674 , n68740 , n389673 );
buf ( n389675 , n389674 );
buf ( n389676 , n389675 );
xor ( n389677 , n389651 , n389676 );
buf ( n389678 , n389137 );
not ( n68758 , n389678 );
buf ( n389680 , n389159 );
not ( n389681 , n389680 );
or ( n389682 , n68758 , n389681 );
not ( n68762 , n389183 );
not ( n389684 , n389172 );
or ( n68764 , n68762 , n389684 );
not ( n68765 , n389137 );
nand ( n68766 , n68765 , n389163 );
nand ( n68767 , n68764 , n68766 );
buf ( n389689 , n68767 );
nand ( n68769 , n389682 , n389689 );
buf ( n389691 , n68769 );
buf ( n389692 , n389691 );
xor ( n68772 , n389677 , n389692 );
buf ( n389694 , n68772 );
buf ( n389695 , n389694 );
buf ( n389696 , n45075 );
not ( n389697 , n389696 );
buf ( n68777 , n342881 );
not ( n68778 , n68777 );
buf ( n68779 , n362288 );
not ( n68780 , n68779 );
or ( n68781 , n68778 , n68780 );
buf ( n68782 , n362285 );
buf ( n68783 , n45065 );
nand ( n68784 , n68782 , n68783 );
buf ( n68785 , n68784 );
buf ( n68786 , n68785 );
nand ( n68787 , n68781 , n68786 );
buf ( n68788 , n68787 );
buf ( n389710 , n68788 );
not ( n389711 , n389710 );
or ( n68791 , n389697 , n389711 );
buf ( n389713 , n68235 );
buf ( n389714 , n45058 );
nand ( n68794 , n389713 , n389714 );
buf ( n389716 , n68794 );
buf ( n389717 , n389716 );
nand ( n68797 , n68791 , n389717 );
buf ( n389719 , n68797 );
buf ( n389720 , n389719 );
xor ( n68800 , n388892 , n388917 );
and ( n68801 , n68800 , n388968 );
and ( n68802 , n388892 , n388917 );
or ( n389724 , n68801 , n68802 );
buf ( n389725 , n389724 );
buf ( n389726 , n389725 );
xor ( n389727 , n389720 , n389726 );
buf ( n389728 , n377580 );
not ( n68808 , n389728 );
xor ( n389730 , n377585 , n41406 );
buf ( n389731 , n389730 );
not ( n68811 , n389731 );
or ( n389733 , n68808 , n68811 );
nand ( n68813 , n67849 , n57530 );
buf ( n389735 , n68813 );
nand ( n68815 , n389733 , n389735 );
buf ( n389737 , n68815 );
buf ( n389738 , n389737 );
xor ( n389739 , n389727 , n389738 );
buf ( n389740 , n389739 );
buf ( n389741 , n389740 );
and ( n389742 , n389695 , n389741 );
not ( n389743 , n389695 );
not ( n68823 , n389740 );
buf ( n389745 , n68823 );
and ( n389746 , n389743 , n389745 );
nor ( n68826 , n389742 , n389746 );
buf ( n68827 , n68826 );
not ( n389749 , n68827 );
not ( n389750 , n389749 );
or ( n68830 , n389636 , n389750 );
not ( n389752 , n68719 );
nand ( n68832 , n389752 , n68827 );
nand ( n68833 , n68830 , n68832 );
not ( n68834 , n389056 );
not ( n68835 , n389209 );
or ( n68836 , n68834 , n68835 );
or ( n68837 , n389209 , n389056 );
nand ( n68838 , n68837 , n68518 );
nand ( n68839 , n68836 , n68838 );
xor ( n68840 , n68833 , n68839 );
xor ( n68841 , n389501 , n389508 );
and ( n68842 , n68841 , n389530 );
and ( n68843 , n389501 , n389508 );
or ( n68844 , n68842 , n68843 );
buf ( n389766 , n68844 );
buf ( n389767 , n389766 );
not ( n389768 , n389767 );
buf ( n389769 , n389768 );
buf ( n389770 , n389769 );
not ( n389771 , n389770 );
not ( n389772 , n68494 );
not ( n68852 , n68392 );
and ( n389774 , n389772 , n68852 );
nand ( n389775 , n68494 , n68392 );
and ( n68855 , n389775 , n389420 );
nor ( n389777 , n389774 , n68855 );
buf ( n389778 , n389777 );
buf ( n389779 , n388855 );
not ( n389780 , n389779 );
buf ( n389781 , n42263 );
not ( n68861 , n389781 );
or ( n389783 , n389780 , n68861 );
and ( n68863 , n351318 , n365915 );
not ( n68864 , n351318 );
and ( n68865 , n68864 , n377715 );
or ( n68866 , n68863 , n68865 );
buf ( n389788 , n68866 );
buf ( n389789 , n48490 );
nand ( n68869 , n389788 , n389789 );
buf ( n389791 , n68869 );
buf ( n389792 , n389791 );
nand ( n68872 , n389783 , n389792 );
buf ( n389794 , n68872 );
buf ( n389795 , n46521 );
not ( n68875 , n389795 );
buf ( n389797 , n389095 );
not ( n389798 , n389797 );
or ( n68878 , n68875 , n389798 );
buf ( n389800 , n46477 );
not ( n68880 , n389800 );
buf ( n389802 , n368976 );
not ( n68882 , n389802 );
or ( n389804 , n68880 , n68882 );
buf ( n389805 , n362537 );
not ( n68885 , n389805 );
buf ( n389807 , n68885 );
buf ( n389808 , n389807 );
buf ( n389809 , n366683 );
nand ( n389810 , n389808 , n389809 );
buf ( n389811 , n389810 );
buf ( n389812 , n389811 );
nand ( n389813 , n389804 , n389812 );
buf ( n389814 , n389813 );
buf ( n389815 , n389814 );
buf ( n389816 , n366654 );
nand ( n68896 , n389815 , n389816 );
buf ( n389818 , n68896 );
buf ( n389819 , n389818 );
nand ( n389820 , n68878 , n389819 );
buf ( n389821 , n389820 );
xor ( n389822 , n389794 , n389821 );
buf ( n389823 , n389074 );
not ( n68903 , n389823 );
buf ( n389825 , n365279 );
not ( n389826 , n389825 );
or ( n68906 , n68903 , n389826 );
buf ( n389828 , n40923 );
buf ( n389829 , n351160 );
not ( n68909 , n389829 );
buf ( n389831 , n372882 );
not ( n68911 , n389831 );
or ( n68912 , n68909 , n68911 );
buf ( n389834 , n365569 );
buf ( n389835 , n364915 );
nand ( n389836 , n389834 , n389835 );
buf ( n389837 , n389836 );
buf ( n389838 , n389837 );
nand ( n68918 , n68912 , n389838 );
buf ( n389840 , n68918 );
buf ( n389841 , n389840 );
nand ( n68921 , n389828 , n389841 );
buf ( n389843 , n68921 );
buf ( n389844 , n389843 );
nand ( n68924 , n68906 , n389844 );
buf ( n389846 , n68924 );
xnor ( n68926 , n389822 , n389846 );
not ( n68927 , n389405 );
not ( n68928 , n68927 );
not ( n68929 , n68475 );
or ( n68930 , n68928 , n68929 );
nand ( n389852 , n68930 , n389392 );
nand ( n389853 , n389405 , n389388 );
nand ( n68933 , n389852 , n389853 );
xor ( n389855 , n68926 , n68933 );
buf ( n389856 , n389264 );
not ( n68936 , n389856 );
buf ( n389858 , n389289 );
not ( n68938 , n389858 );
or ( n68939 , n68936 , n68938 );
not ( n68940 , n68349 );
not ( n68941 , n389290 );
or ( n68942 , n68940 , n68941 );
nand ( n68943 , n68942 , n389301 );
buf ( n389865 , n68943 );
nand ( n68945 , n68939 , n389865 );
buf ( n389867 , n68945 );
xor ( n68947 , n389855 , n389867 );
buf ( n389869 , n365152 );
not ( n68949 , n389869 );
not ( n68950 , n342909 );
not ( n68951 , n362458 );
or ( n68952 , n68950 , n68951 );
not ( n68953 , n387355 );
nand ( n68954 , n68953 , n360848 );
nand ( n389876 , n68952 , n68954 );
buf ( n389877 , n389876 );
not ( n389878 , n389877 );
or ( n68958 , n68949 , n389878 );
buf ( n389880 , n389326 );
buf ( n389881 , n365189 );
nand ( n389882 , n389880 , n389881 );
buf ( n389883 , n389882 );
buf ( n389884 , n389883 );
nand ( n389885 , n68958 , n389884 );
buf ( n389886 , n389885 );
buf ( n389887 , n389886 );
buf ( n389888 , n363291 );
buf ( n389889 , n67971 );
not ( n68969 , n389889 );
buf ( n389891 , n68969 );
buf ( n389892 , n389891 );
or ( n68972 , n389888 , n389892 );
buf ( n389894 , n365801 );
buf ( n389895 , n56970 );
not ( n68975 , n389895 );
buf ( n389897 , n41623 );
not ( n68977 , n389897 );
or ( n389899 , n68975 , n68977 );
buf ( n389900 , n361762 );
buf ( n389901 , n377389 );
nand ( n68981 , n389900 , n389901 );
buf ( n389903 , n68981 );
buf ( n389904 , n389903 );
nand ( n68984 , n389899 , n389904 );
buf ( n68985 , n68984 );
buf ( n389907 , n68985 );
not ( n68987 , n389907 );
buf ( n389909 , n68987 );
buf ( n389910 , n389909 );
or ( n68990 , n389894 , n389910 );
nand ( n389912 , n68972 , n68990 );
buf ( n389913 , n389912 );
buf ( n389914 , n389913 );
xor ( n68994 , n389887 , n389914 );
buf ( n389916 , n388960 );
not ( n389917 , n389916 );
buf ( n389918 , n364797 );
not ( n68998 , n389918 );
or ( n389920 , n389917 , n68998 );
not ( n389921 , n364832 );
not ( n69001 , n31197 );
or ( n389923 , n389921 , n69001 );
nand ( n69003 , n41892 , n351229 );
nand ( n389925 , n389923 , n69003 );
nand ( n69005 , n365622 , n389925 );
buf ( n389927 , n69005 );
nand ( n389928 , n389920 , n389927 );
buf ( n389929 , n389928 );
buf ( n389930 , n389929 );
not ( n389931 , n59588 );
not ( n69011 , n389126 );
or ( n69012 , n389931 , n69011 );
buf ( n389934 , n365440 );
not ( n389935 , n389934 );
buf ( n389936 , n366086 );
not ( n389937 , n389936 );
or ( n389938 , n389935 , n389937 );
buf ( n389939 , n366096 );
buf ( n389940 , n365452 );
nand ( n389941 , n389939 , n389940 );
buf ( n389942 , n389941 );
buf ( n389943 , n389942 );
nand ( n389944 , n389938 , n389943 );
buf ( n389945 , n389944 );
buf ( n389946 , n389945 );
buf ( n69026 , n366518 );
nand ( n69027 , n389946 , n69026 );
buf ( n389949 , n69027 );
nand ( n389950 , n69012 , n389949 );
buf ( n389951 , n389950 );
xor ( n69031 , n389930 , n389951 );
buf ( n389953 , n389386 );
not ( n389954 , n389953 );
buf ( n389955 , n369260 );
not ( n389956 , n389955 );
or ( n69036 , n389954 , n389956 );
buf ( n389958 , n46582 );
not ( n389959 , n365408 );
not ( n69039 , n365367 );
or ( n389961 , n389959 , n69039 );
nand ( n69041 , n373150 , n365393 );
nand ( n389963 , n389961 , n69041 );
buf ( n389964 , n389963 );
nand ( n69044 , n389958 , n389964 );
buf ( n69045 , n69044 );
buf ( n389967 , n69045 );
nand ( n69047 , n69036 , n389967 );
buf ( n69048 , n69047 );
buf ( n389970 , n69048 );
xor ( n69050 , n69031 , n389970 );
buf ( n389972 , n69050 );
buf ( n389973 , n389972 );
xor ( n69053 , n68994 , n389973 );
buf ( n389975 , n69053 );
buf ( n389976 , n389333 );
not ( n69056 , n389976 );
buf ( n389978 , n69056 );
not ( n69058 , n389978 );
not ( n69059 , n389350 );
or ( n389981 , n69058 , n69059 );
nand ( n389982 , n389981 , n389409 );
buf ( n389983 , n389982 );
buf ( n389984 , n389350 );
not ( n69064 , n389984 );
buf ( n389986 , n389333 );
nand ( n69066 , n69064 , n389986 );
buf ( n389988 , n69066 );
buf ( n389989 , n389988 );
nand ( n69069 , n389983 , n389989 );
buf ( n389991 , n69069 );
and ( n69071 , n389975 , n389991 );
not ( n389993 , n389975 );
not ( n69073 , n389991 );
and ( n389995 , n389993 , n69073 );
nor ( n389996 , n69071 , n389995 );
xor ( n69076 , n68947 , n389996 );
not ( n389998 , n69076 );
buf ( n389999 , n389998 );
and ( n390000 , n389778 , n389999 );
not ( n69080 , n389778 );
buf ( n390002 , n69076 );
and ( n390003 , n69080 , n390002 );
nor ( n390004 , n390000 , n390003 );
buf ( n390005 , n390004 );
buf ( n390006 , n390005 );
not ( n390007 , n390006 );
or ( n69087 , n389771 , n390007 );
buf ( n390009 , n390005 );
buf ( n390010 , n389769 );
or ( n69090 , n390009 , n390010 );
nand ( n69091 , n69087 , n69090 );
buf ( n390013 , n69091 );
xor ( n69093 , n68840 , n390013 );
not ( n390015 , n68620 );
not ( n390016 , n68617 );
or ( n69096 , n390015 , n390016 );
nand ( n390018 , n69096 , n68639 );
not ( n69098 , n390018 );
and ( n69099 , n389532 , n68551 );
nor ( n390021 , n69098 , n69099 );
buf ( n390022 , n390021 );
not ( n390023 , n390022 );
not ( n69103 , n68568 );
nand ( n69104 , n69103 , n68579 );
not ( n390026 , n69104 );
not ( n390027 , n389473 );
or ( n69107 , n390026 , n390027 );
nand ( n390029 , n68568 , n68578 );
nand ( n390030 , n69107 , n390029 );
buf ( n390031 , n390030 );
buf ( n390032 , n389215 );
buf ( n69112 , n390032 );
not ( n69113 , n69112 );
buf ( n69114 , n389239 );
not ( n69115 , n69114 );
or ( n69116 , n69113 , n69115 );
buf ( n390038 , n390032 );
buf ( n390039 , n389239 );
or ( n69119 , n390038 , n390039 );
buf ( n390041 , n68390 );
nand ( n390042 , n69119 , n390041 );
buf ( n390043 , n390042 );
buf ( n390044 , n390043 );
nand ( n69124 , n69116 , n390044 );
buf ( n390046 , n69124 );
buf ( n390047 , n390046 );
xor ( n390048 , n390031 , n390047 );
not ( n390049 , n47466 );
not ( n69129 , n389345 );
or ( n390051 , n390049 , n69129 );
not ( n69131 , n365052 );
not ( n69132 , n366719 );
or ( n390054 , n69131 , n69132 );
nand ( n390055 , n366725 , n365041 );
nand ( n69135 , n390054 , n390055 );
nand ( n390057 , n69135 , n44915 );
nand ( n390058 , n390051 , n390057 );
buf ( n390059 , n389258 );
not ( n390060 , n390059 );
buf ( n390061 , n39701 );
not ( n69141 , n390061 );
or ( n69142 , n390060 , n69141 );
buf ( n390064 , n367796 );
buf ( n390065 , n377779 );
not ( n69145 , n390065 );
buf ( n390067 , n39621 );
not ( n390068 , n390067 );
or ( n69148 , n69145 , n390068 );
buf ( n390070 , n45231 );
buf ( n390071 , n377782 );
nand ( n69151 , n390070 , n390071 );
buf ( n390073 , n69151 );
buf ( n390074 , n390073 );
nand ( n69154 , n69148 , n390074 );
buf ( n390076 , n69154 );
buf ( n390077 , n390076 );
nand ( n390078 , n390064 , n390077 );
buf ( n390079 , n390078 );
buf ( n390080 , n390079 );
nand ( n390081 , n69142 , n390080 );
buf ( n390082 , n390081 );
buf ( n390083 , n390082 );
not ( n69163 , n67941 );
not ( n69164 , n388857 );
or ( n69165 , n69163 , n69164 );
not ( n69166 , n67941 );
not ( n69167 , n69166 );
not ( n390089 , n388858 );
or ( n69169 , n69167 , n390089 );
nand ( n390091 , n69169 , n67920 );
nand ( n69171 , n69165 , n390091 );
buf ( n390093 , n69171 );
xor ( n69173 , n390083 , n390093 );
buf ( n390095 , n389401 );
not ( n69175 , n390095 );
buf ( n390097 , n46113 );
not ( n69177 , n390097 );
or ( n69178 , n69175 , n69177 );
buf ( n390100 , n365980 );
buf ( n390101 , n366277 );
and ( n390102 , n390100 , n390101 );
not ( n69182 , n390100 );
buf ( n390104 , n362452 );
and ( n390105 , n69182 , n390104 );
nor ( n390106 , n390102 , n390105 );
buf ( n390107 , n390106 );
buf ( n390108 , n390107 );
not ( n390109 , n390108 );
buf ( n390110 , n360574 );
nand ( n69190 , n390109 , n390110 );
buf ( n390112 , n69190 );
buf ( n390113 , n390112 );
nand ( n69193 , n69178 , n390113 );
buf ( n69194 , n69193 );
buf ( n390116 , n69194 );
xor ( n69196 , n69173 , n390116 );
buf ( n390118 , n69196 );
and ( n69198 , n390058 , n390118 );
not ( n390120 , n390058 );
not ( n69200 , n390118 );
and ( n390122 , n390120 , n69200 );
nor ( n390123 , n69198 , n390122 );
not ( n69203 , n45345 );
not ( n390125 , n389282 );
or ( n390126 , n69203 , n390125 );
buf ( n390127 , n368994 );
not ( n390128 , n390127 );
buf ( n390129 , n363116 );
not ( n69209 , n390129 );
or ( n69210 , n390128 , n69209 );
buf ( n390132 , n370845 );
not ( n390133 , n390132 );
buf ( n390134 , n57053 );
nand ( n69214 , n390133 , n390134 );
buf ( n69215 , n69214 );
buf ( n69216 , n69215 );
nand ( n69217 , n69210 , n69216 );
buf ( n69218 , n69217 );
buf ( n390140 , n69218 );
buf ( n390141 , n39946 );
nand ( n390142 , n390140 , n390141 );
buf ( n390143 , n390142 );
nand ( n390144 , n390126 , n390143 );
not ( n69224 , n45492 );
not ( n390146 , n365676 );
not ( n69226 , n365760 );
or ( n390148 , n390146 , n69226 );
buf ( n390149 , n41528 );
buf ( n390150 , n365673 );
nand ( n390151 , n390149 , n390150 );
buf ( n390152 , n390151 );
nand ( n69232 , n390148 , n390152 );
not ( n390154 , n69232 );
or ( n390155 , n69224 , n390154 );
nand ( n69235 , n389363 , n45553 );
nand ( n390157 , n390155 , n69235 );
and ( n390158 , n390144 , n390157 );
not ( n69238 , n390144 );
buf ( n390160 , n45553 );
not ( n390161 , n390160 );
buf ( n390162 , n389363 );
not ( n390163 , n390162 );
or ( n390164 , n390161 , n390163 );
nand ( n69244 , n69232 , n45492 );
buf ( n390166 , n69244 );
nand ( n69246 , n390164 , n390166 );
buf ( n390168 , n69246 );
buf ( n390169 , n390168 );
not ( n69249 , n390169 );
buf ( n390171 , n69249 );
and ( n69251 , n69238 , n390171 );
or ( n390173 , n390158 , n69251 );
buf ( n390174 , n46135 );
not ( n69254 , n390174 );
buf ( n390176 , n68021 );
not ( n390177 , n390176 );
or ( n69257 , n69254 , n390177 );
buf ( n390179 , n365319 );
not ( n69259 , n390179 );
buf ( n390181 , n352212 );
nor ( n69261 , n69259 , n390181 );
buf ( n390183 , n69261 );
not ( n69263 , n378032 );
nor ( n69264 , n69263 , n365259 );
nor ( n390186 , n390183 , n69264 );
buf ( n390187 , n390186 );
buf ( n390188 , n365312 );
or ( n69268 , n390187 , n390188 );
nand ( n390190 , n69257 , n69268 );
buf ( n390191 , n390190 );
not ( n390192 , n366428 );
not ( n69272 , n386807 );
not ( n69273 , n366187 );
or ( n390195 , n69272 , n69273 );
buf ( n69275 , n351762 );
buf ( n390197 , n65993 );
nand ( n390198 , n69275 , n390197 );
buf ( n390199 , n390198 );
nand ( n390200 , n390195 , n390199 );
not ( n69280 , n390200 );
or ( n69281 , n390192 , n69280 );
buf ( n390203 , n388830 );
buf ( n390204 , n366399 );
nand ( n390205 , n390203 , n390204 );
buf ( n390206 , n390205 );
nand ( n69286 , n69281 , n390206 );
buf ( n390208 , n366131 );
buf ( n390209 , n22769 );
and ( n69289 , n390208 , n390209 );
buf ( n390211 , n42233 );
buf ( n390212 , n351367 );
and ( n69292 , n390211 , n390212 );
nor ( n69293 , n69289 , n69292 );
buf ( n69294 , n69293 );
buf ( n390216 , n69294 );
not ( n390217 , n390216 );
buf ( n390218 , n58231 );
not ( n69298 , n390218 );
buf ( n390220 , n69298 );
buf ( n390221 , n390220 );
not ( n69301 , n390221 );
and ( n69302 , n390217 , n69301 );
buf ( n390224 , n388807 );
buf ( n390225 , n363429 );
and ( n390226 , n390224 , n390225 );
nor ( n69306 , n69302 , n390226 );
buf ( n390228 , n69306 );
not ( n390229 , n390228 );
and ( n69309 , n69286 , n390229 );
not ( n69310 , n69286 );
and ( n390232 , n69310 , n390228 );
nor ( n390233 , n69309 , n390232 );
xor ( n69313 , n390191 , n390233 );
xor ( n69314 , n390173 , n69313 );
not ( n390236 , n69314 );
and ( n69316 , n390123 , n390236 );
not ( n390238 , n390123 );
and ( n390239 , n390238 , n69314 );
nor ( n390240 , n69316 , n390239 );
buf ( n390241 , n390240 );
xor ( n390242 , n390048 , n390241 );
buf ( n390243 , n390242 );
buf ( n390244 , n388999 );
not ( n390245 , n390244 );
buf ( n390246 , n67887 );
not ( n390247 , n390246 );
or ( n390248 , n390245 , n390247 );
buf ( n390249 , n389027 );
nand ( n390250 , n390248 , n390249 );
buf ( n390251 , n390250 );
buf ( n69331 , n390251 );
buf ( n390253 , n67887 );
not ( n69333 , n390253 );
buf ( n390255 , n389002 );
nand ( n390256 , n69333 , n390255 );
buf ( n390257 , n390256 );
buf ( n390258 , n390257 );
nand ( n390259 , n69331 , n390258 );
buf ( n390260 , n390259 );
xor ( n69340 , n390243 , n390260 );
buf ( n390262 , n388755 );
not ( n390263 , n390262 );
buf ( n390264 , n388748 );
not ( n69344 , n390264 );
or ( n69345 , n390263 , n69344 );
buf ( n390267 , n388737 );
not ( n390268 , n390267 );
buf ( n390269 , n67854 );
not ( n69349 , n390269 );
or ( n390271 , n390268 , n69349 );
buf ( n390272 , n388776 );
nand ( n69352 , n390271 , n390272 );
buf ( n390274 , n69352 );
buf ( n390275 , n390274 );
nand ( n390276 , n69345 , n390275 );
buf ( n390277 , n390276 );
buf ( n390278 , n390277 );
not ( n390279 , n67961 );
buf ( n69359 , n67896 );
not ( n390281 , n69359 );
or ( n390282 , n390279 , n390281 );
buf ( n390283 , n67961 );
buf ( n390284 , n69359 );
or ( n69364 , n390283 , n390284 );
buf ( n390286 , n388859 );
not ( n390287 , n390286 );
buf ( n390288 , n390287 );
buf ( n390289 , n390288 );
nand ( n69366 , n69364 , n390289 );
buf ( n390291 , n69366 );
nand ( n69368 , n390282 , n390291 );
not ( n390293 , n387542 );
buf ( n390294 , n368549 );
not ( n390295 , n390294 );
buf ( n390296 , n364987 );
not ( n390297 , n390296 );
or ( n390298 , n390295 , n390297 );
buf ( n390299 , n359778 );
buf ( n390300 , n368554 );
nand ( n390301 , n390299 , n390300 );
buf ( n390302 , n390301 );
buf ( n390303 , n390302 );
nand ( n390304 , n390298 , n390303 );
buf ( n390305 , n390304 );
not ( n390306 , n390305 );
or ( n390307 , n390293 , n390306 );
buf ( n390308 , n368614 );
not ( n390309 , n390308 );
buf ( n390310 , n389232 );
nand ( n390311 , n390309 , n390310 );
buf ( n390312 , n390311 );
nand ( n390313 , n390307 , n390312 );
not ( n390314 , n390313 );
and ( n390315 , n69368 , n390314 );
not ( n390316 , n69368 );
and ( n390317 , n390316 , n390313 );
nor ( n390318 , n390315 , n390317 );
buf ( n390319 , n67603 );
not ( n69373 , n390319 );
buf ( n390321 , n68026 );
not ( n69375 , n390321 );
buf ( n390323 , n69375 );
buf ( n390324 , n390323 );
not ( n69378 , n390324 );
or ( n390326 , n69373 , n69378 );
not ( n390327 , n388452 );
not ( n69381 , n68026 );
or ( n390329 , n390327 , n69381 );
nand ( n390330 , n390329 , n68048 );
buf ( n390331 , n390330 );
nand ( n390332 , n390326 , n390331 );
buf ( n390333 , n390332 );
buf ( n390334 , n390333 );
buf ( n390335 , n365033 );
not ( n69389 , n390335 );
buf ( n390337 , n388906 );
not ( n390338 , n390337 );
or ( n390339 , n69389 , n390338 );
buf ( n390340 , n44819 );
not ( n390341 , n390340 );
buf ( n390342 , n367459 );
not ( n69396 , n390342 );
buf ( n69397 , n69396 );
buf ( n390345 , n69397 );
not ( n390346 , n390345 );
or ( n69400 , n390341 , n390346 );
buf ( n390348 , n361802 );
buf ( n390349 , n364978 );
nand ( n69403 , n390348 , n390349 );
buf ( n390351 , n69403 );
buf ( n390352 , n390351 );
nand ( n69406 , n69400 , n390352 );
buf ( n390354 , n69406 );
buf ( n69408 , n390354 );
buf ( n69409 , n365115 );
nand ( n69410 , n69408 , n69409 );
buf ( n69411 , n69410 );
buf ( n69412 , n69411 );
nand ( n69413 , n390339 , n69412 );
buf ( n69414 , n69413 );
buf ( n69415 , n69414 );
xor ( n69416 , n390334 , n69415 );
not ( n390364 , n389081 );
not ( n69418 , n68216 );
and ( n390366 , n390364 , n69418 );
buf ( n390367 , n389081 );
buf ( n390368 , n68216 );
nand ( n390369 , n390367 , n390368 );
buf ( n390370 , n390369 );
and ( n390371 , n390370 , n389109 );
nor ( n390372 , n390366 , n390371 );
buf ( n390373 , n390372 );
xor ( n390374 , n69416 , n390373 );
buf ( n390375 , n390374 );
not ( n390376 , n390375 );
and ( n69430 , n390318 , n390376 );
not ( n390378 , n390318 );
and ( n390379 , n390378 , n390375 );
nor ( n69433 , n69430 , n390379 );
not ( n390381 , n69433 );
buf ( n390382 , n390381 );
xor ( n69436 , n390278 , n390382 );
buf ( n390384 , n388970 );
buf ( n390385 , n388996 );
or ( n69439 , n390384 , n390385 );
buf ( n390387 , n388878 );
buf ( n390388 , n390387 );
nand ( n390389 , n69439 , n390388 );
buf ( n390390 , n390389 );
buf ( n390391 , n390390 );
buf ( n390392 , n388996 );
buf ( n390393 , n388970 );
nand ( n69447 , n390392 , n390393 );
buf ( n390395 , n69447 );
buf ( n390396 , n390395 );
nand ( n69450 , n390391 , n390396 );
buf ( n390398 , n69450 );
buf ( n390399 , n390398 );
xor ( n69453 , n69436 , n390399 );
buf ( n390401 , n69453 );
xor ( n69455 , n69340 , n390401 );
buf ( n390403 , n69455 );
not ( n69457 , n390403 );
and ( n69458 , n390023 , n69457 );
buf ( n390406 , n69455 );
buf ( n390407 , n390021 );
and ( n69461 , n390406 , n390407 );
nor ( n69462 , n69458 , n69461 );
buf ( n390410 , n69462 );
xor ( n69464 , n69093 , n390410 );
buf ( n390412 , n69464 );
xor ( n390413 , n68705 , n390412 );
buf ( n390414 , n390413 );
buf ( n390415 , n390414 );
not ( n390416 , n390415 );
buf ( n390417 , n390416 );
buf ( n69471 , n390417 );
xor ( n69472 , n389448 , n389573 );
and ( n390420 , n69472 , n68664 );
and ( n390421 , n389448 , n389573 );
or ( n69475 , n390420 , n390421 );
buf ( n390423 , n69475 );
not ( n69477 , n390423 );
buf ( n390425 , n69477 );
buf ( n390426 , n390425 );
nand ( n69480 , n69471 , n390426 );
buf ( n390428 , n69480 );
not ( n69482 , n390428 );
or ( n69483 , n389597 , n69482 );
nand ( n69484 , n390414 , n69475 );
buf ( n69485 , n69484 );
nand ( n69486 , n69483 , n69485 );
xor ( n69487 , n389887 , n389914 );
and ( n69488 , n69487 , n389973 );
and ( n69489 , n389887 , n389914 );
or ( n390437 , n69488 , n69489 );
buf ( n390438 , n390437 );
buf ( n390439 , n389668 );
buf ( n390440 , n369804 );
and ( n69494 , n390439 , n390440 );
nor ( n390442 , n369769 , n369813 );
not ( n390443 , n390442 );
not ( n69497 , n363171 );
or ( n390445 , n390443 , n69497 );
nor ( n390446 , n369766 , n369813 );
nand ( n69500 , n41907 , n390446 );
nand ( n390448 , n390445 , n69500 );
buf ( n390449 , n390448 );
nor ( n390450 , n69494 , n390449 );
buf ( n390451 , n390450 );
not ( n390452 , n390451 );
not ( n69506 , n387542 );
not ( n69507 , n359756 );
not ( n69508 , n368554 );
or ( n69509 , n69507 , n69508 );
buf ( n69510 , n368549 );
nand ( n390458 , n362208 , n69510 );
nand ( n390459 , n69509 , n390458 );
not ( n390460 , n390459 );
or ( n69514 , n69506 , n390460 );
not ( n390462 , n368614 );
nand ( n390463 , n390462 , n390305 );
nand ( n69517 , n69514 , n390463 );
not ( n390465 , n69517 );
or ( n390466 , n390452 , n390465 );
buf ( n390467 , n390451 );
not ( n390468 , n390467 );
buf ( n390469 , n390468 );
not ( n69523 , n69517 );
nand ( n390471 , n390469 , n69523 );
nand ( n390472 , n390466 , n390471 );
xor ( n69526 , n390438 , n390472 );
buf ( n390474 , n69526 );
buf ( n390475 , n390372 );
not ( n69529 , n390475 );
not ( n69530 , n69414 );
buf ( n390478 , n69530 );
not ( n390479 , n390478 );
or ( n390480 , n69529 , n390479 );
buf ( n390481 , n390333 );
nand ( n390482 , n390480 , n390481 );
buf ( n390483 , n390482 );
buf ( n390484 , n390483 );
buf ( n390485 , n390372 );
not ( n69538 , n390485 );
buf ( n390487 , n69414 );
nand ( n69540 , n69538 , n390487 );
buf ( n390489 , n69540 );
buf ( n390490 , n390489 );
nand ( n69543 , n390484 , n390490 );
buf ( n69544 , n69543 );
buf ( n390493 , n69544 );
not ( n69546 , n57530 );
not ( n69547 , n389730 );
or ( n390496 , n69546 , n69547 );
not ( n390497 , n377585 );
not ( n69550 , n362179 );
or ( n390499 , n390497 , n69550 );
buf ( n390500 , n40899 );
buf ( n390501 , n386943 );
nand ( n390502 , n390500 , n390501 );
buf ( n390503 , n390502 );
nand ( n390504 , n390499 , n390503 );
nand ( n390505 , n390504 , n377580 );
nand ( n69558 , n390496 , n390505 );
buf ( n390507 , n69558 );
xor ( n390508 , n390493 , n390507 );
not ( n69561 , n68985 );
not ( n390510 , n386445 );
or ( n69563 , n69561 , n390510 );
buf ( n69564 , n369374 );
not ( n69565 , n69564 );
buf ( n69566 , n359904 );
not ( n69567 , n69566 );
or ( n69568 , n69565 , n69567 );
buf ( n390517 , n366243 );
buf ( n390518 , n49178 );
nand ( n69571 , n390517 , n390518 );
buf ( n390520 , n69571 );
buf ( n390521 , n390520 );
nand ( n390522 , n69568 , n390521 );
buf ( n390523 , n390522 );
nand ( n69576 , n390523 , n368038 );
nand ( n390525 , n69563 , n69576 );
buf ( n390526 , n390525 );
not ( n69579 , n390526 );
not ( n390528 , n45492 );
not ( n390529 , n41607 );
not ( n390530 , n365673 );
or ( n390531 , n390529 , n390530 );
nand ( n69584 , n44783 , n365676 );
nand ( n390533 , n390531 , n69584 );
not ( n69586 , n390533 );
or ( n390535 , n390528 , n69586 );
buf ( n390536 , n45553 );
buf ( n390537 , n69232 );
nand ( n390538 , n390536 , n390537 );
buf ( n390539 , n390538 );
nand ( n390540 , n390535 , n390539 );
buf ( n390541 , n390540 );
not ( n69594 , n390541 );
buf ( n390543 , n69594 );
buf ( n390544 , n390543 );
not ( n69597 , n390544 );
or ( n390546 , n69579 , n69597 );
not ( n390547 , n390525 );
nand ( n69600 , n390547 , n390540 );
buf ( n390549 , n69600 );
nand ( n390550 , n390546 , n390549 );
buf ( n390551 , n390550 );
buf ( n390552 , n390551 );
buf ( n390553 , n389794 );
not ( n390554 , n390553 );
buf ( n390555 , n390554 );
or ( n69608 , n389846 , n390555 );
nand ( n390557 , n69608 , n389821 );
buf ( n390558 , n389846 );
buf ( n390559 , n390555 );
nand ( n390560 , n390558 , n390559 );
buf ( n390561 , n390560 );
nand ( n69614 , n390557 , n390561 );
buf ( n390563 , n69614 );
xor ( n69616 , n390552 , n390563 );
buf ( n390565 , n69616 );
buf ( n390566 , n390565 );
xor ( n69619 , n390508 , n390566 );
buf ( n390568 , n69619 );
buf ( n390569 , n390568 );
xor ( n69622 , n390474 , n390569 );
buf ( n390571 , n69622 );
not ( n390572 , n390571 );
not ( n69625 , n68947 );
not ( n69626 , n389975 );
nand ( n69627 , n69626 , n69073 );
not ( n69628 , n69627 );
or ( n69629 , n69625 , n69628 );
not ( n69630 , n69073 );
nand ( n390579 , n69630 , n389975 );
nand ( n69632 , n69629 , n390579 );
or ( n390581 , n390572 , n69632 );
not ( n69634 , n69632 );
or ( n69635 , n390571 , n69634 );
nand ( n69636 , n390581 , n69635 );
buf ( n390585 , n69636 );
buf ( n390586 , n389777 );
not ( n390587 , n390586 );
not ( n69640 , n69076 );
buf ( n69641 , n69640 );
not ( n69642 , n69641 );
or ( n69643 , n390587 , n69642 );
buf ( n390592 , n389766 );
nand ( n390593 , n69643 , n390592 );
buf ( n390594 , n390593 );
buf ( n390595 , n390594 );
buf ( n390596 , n389777 );
not ( n69649 , n390596 );
buf ( n390598 , n69076 );
nand ( n69651 , n69649 , n390598 );
buf ( n390600 , n69651 );
buf ( n390601 , n390600 );
nand ( n69654 , n390595 , n390601 );
buf ( n390603 , n69654 );
buf ( n390604 , n390603 );
xor ( n390605 , n390585 , n390604 );
buf ( n390606 , n390605 );
not ( n69659 , n390606 );
not ( n390608 , n69659 );
xor ( n69661 , n390031 , n390047 );
and ( n390610 , n69661 , n390241 );
and ( n69663 , n390031 , n390047 );
or ( n69664 , n390610 , n69663 );
buf ( n390613 , n69664 );
buf ( n390614 , n390613 );
not ( n69667 , n390058 );
not ( n390616 , n69667 );
not ( n390617 , n69200 );
or ( n69670 , n390616 , n390617 );
not ( n390619 , n390058 );
not ( n390620 , n390118 );
or ( n69673 , n390619 , n390620 );
nand ( n390622 , n69673 , n69314 );
nand ( n69675 , n69670 , n390622 );
not ( n69676 , n69675 );
xor ( n390625 , n68926 , n68933 );
and ( n390626 , n390625 , n389867 );
and ( n69679 , n68926 , n68933 );
or ( n390628 , n390626 , n69679 );
not ( n390629 , n390628 );
buf ( n390630 , n40474 );
not ( n390631 , n390630 );
buf ( n390632 , n390107 );
not ( n390633 , n390632 );
and ( n69686 , n390631 , n390633 );
buf ( n390635 , n366754 );
buf ( n390636 , n46303 );
buf ( n390637 , n365468 );
and ( n390638 , n390636 , n390637 );
not ( n390639 , n390636 );
buf ( n390640 , n362452 );
and ( n390641 , n390639 , n390640 );
nor ( n390642 , n390638 , n390641 );
buf ( n390643 , n390642 );
buf ( n390644 , n390643 );
nor ( n390645 , n390635 , n390644 );
buf ( n390646 , n390645 );
buf ( n390647 , n390646 );
nor ( n69700 , n69686 , n390647 );
buf ( n390649 , n69700 );
buf ( n390650 , n390649 );
not ( n390651 , n390650 );
not ( n69704 , n366654 );
not ( n390653 , n43377 );
not ( n390654 , n46477 );
or ( n69707 , n390653 , n390654 );
buf ( n390656 , n41569 );
buf ( n390657 , n366683 );
nand ( n69710 , n390656 , n390657 );
buf ( n390659 , n69710 );
nand ( n390660 , n69707 , n390659 );
not ( n69713 , n390660 );
or ( n390662 , n69704 , n69713 );
buf ( n390663 , n389814 );
buf ( n390664 , n46521 );
nand ( n390665 , n390663 , n390664 );
buf ( n390666 , n390665 );
nand ( n69719 , n390662 , n390666 );
buf ( n390668 , n69719 );
not ( n390669 , n390668 );
or ( n69722 , n390651 , n390669 );
buf ( n390671 , n390649 );
buf ( n390672 , n69719 );
or ( n69725 , n390671 , n390672 );
nand ( n390674 , n69722 , n69725 );
buf ( n390675 , n390674 );
not ( n69728 , n390675 );
buf ( n390677 , n40058 );
not ( n69730 , n390677 );
buf ( n390679 , n69218 );
not ( n390680 , n390679 );
or ( n390681 , n69730 , n390680 );
not ( n69734 , n368662 );
not ( n390683 , n365948 );
or ( n390684 , n69734 , n390683 );
nand ( n69737 , n368665 , n363116 );
nand ( n390686 , n390684 , n69737 );
buf ( n390687 , n390686 );
buf ( n390688 , n39949 );
nand ( n390689 , n390687 , n390688 );
buf ( n390690 , n390689 );
buf ( n390691 , n390690 );
nand ( n69744 , n390681 , n390691 );
buf ( n390693 , n69744 );
buf ( n390694 , n390693 );
not ( n69747 , n390694 );
buf ( n390696 , n69747 );
not ( n390697 , n390696 );
not ( n69750 , n390697 );
or ( n390699 , n69728 , n69750 );
not ( n390700 , n390675 );
nand ( n69753 , n390700 , n390696 );
nand ( n390702 , n390699 , n69753 );
not ( n69755 , n390702 );
not ( n390704 , n69755 );
buf ( n390705 , n389794 );
buf ( n390706 , n389945 );
not ( n390707 , n390706 );
buf ( n390708 , n369589 );
not ( n390709 , n390708 );
or ( n390710 , n390707 , n390709 );
buf ( n390711 , n45300 );
not ( n69764 , n390711 );
buf ( n390713 , n366086 );
not ( n69766 , n390713 );
or ( n69767 , n69764 , n69766 );
buf ( n390716 , n369577 );
buf ( n390717 , n365474 );
nand ( n69770 , n390716 , n390717 );
buf ( n390719 , n69770 );
buf ( n390720 , n390719 );
nand ( n69773 , n69767 , n390720 );
buf ( n390722 , n69773 );
buf ( n69775 , n390722 );
buf ( n390724 , n366518 );
nand ( n69777 , n69775 , n390724 );
buf ( n390726 , n69777 );
buf ( n390727 , n390726 );
nand ( n390728 , n390710 , n390727 );
buf ( n390729 , n390728 );
buf ( n390730 , n390729 );
xor ( n69783 , n390705 , n390730 );
not ( n69784 , n389925 );
not ( n390733 , n362027 );
or ( n390734 , n69784 , n390733 );
buf ( n390735 , n364824 );
buf ( n390736 , n45177 );
not ( n390737 , n390736 );
buf ( n390738 , n365626 );
not ( n390739 , n390738 );
or ( n390740 , n390737 , n390739 );
buf ( n390741 , n362033 );
buf ( n390742 , n365357 );
nand ( n69795 , n390741 , n390742 );
buf ( n390744 , n69795 );
buf ( n390745 , n390744 );
nand ( n390746 , n390740 , n390745 );
buf ( n390747 , n390746 );
buf ( n390748 , n390747 );
nand ( n69801 , n390735 , n390748 );
buf ( n390750 , n69801 );
nand ( n69803 , n390734 , n390750 );
buf ( n390752 , n69803 );
xnor ( n390753 , n69783 , n390752 );
buf ( n390754 , n390753 );
not ( n69807 , n390754 );
not ( n390756 , n365115 );
buf ( n390757 , n44819 );
not ( n69810 , n390757 );
buf ( n390759 , n362145 );
not ( n390760 , n390759 );
or ( n69813 , n69810 , n390760 );
buf ( n390762 , n362136 );
buf ( n390763 , n364994 );
nand ( n69816 , n390762 , n390763 );
buf ( n390765 , n69816 );
buf ( n390766 , n390765 );
nand ( n69819 , n69813 , n390766 );
buf ( n69820 , n69819 );
not ( n390769 , n69820 );
or ( n69822 , n390756 , n390769 );
buf ( n390771 , n390354 );
buf ( n390772 , n365033 );
nand ( n69825 , n390771 , n390772 );
buf ( n390774 , n69825 );
nand ( n69827 , n69822 , n390774 );
not ( n390776 , n69827 );
not ( n390777 , n390776 );
or ( n69830 , n69807 , n390777 );
buf ( n390779 , n390754 );
not ( n390780 , n390779 );
buf ( n390781 , n390780 );
nand ( n390782 , n390781 , n69827 );
nand ( n69835 , n69830 , n390782 );
and ( n390784 , n390704 , n69835 );
not ( n390785 , n390704 );
not ( n69838 , n69835 );
and ( n390787 , n390785 , n69838 );
nor ( n69840 , n390784 , n390787 );
nand ( n69841 , n390629 , n69840 );
not ( n390790 , n390704 );
not ( n390791 , n390790 );
not ( n69844 , n69838 );
or ( n390793 , n390791 , n69844 );
nand ( n69846 , n390704 , n69835 );
nand ( n69847 , n390793 , n69846 );
nand ( n390796 , n69847 , n390628 );
nand ( n390797 , n69841 , n390796 );
not ( n69850 , n390797 );
or ( n390799 , n69676 , n69850 );
not ( n390800 , n69675 );
nand ( n69853 , n390796 , n69841 , n390800 );
nand ( n390802 , n390799 , n69853 );
buf ( n390803 , n390802 );
xor ( n69856 , n390614 , n390803 );
xor ( n390805 , n389930 , n389951 );
and ( n69858 , n390805 , n389970 );
and ( n69859 , n389930 , n389951 );
or ( n390808 , n69858 , n69859 );
buf ( n390809 , n390808 );
buf ( n390810 , n390809 );
xor ( n390811 , n390083 , n390093 );
and ( n390812 , n390811 , n390116 );
and ( n69865 , n390083 , n390093 );
or ( n390814 , n390812 , n69865 );
buf ( n390815 , n390814 );
buf ( n390816 , n390815 );
xor ( n390817 , n390810 , n390816 );
buf ( n390818 , n389840 );
not ( n390819 , n390818 );
buf ( n390820 , n372247 );
not ( n69873 , n390820 );
or ( n390822 , n390819 , n69873 );
buf ( n390823 , n40923 );
buf ( n390824 , n365490 );
not ( n390825 , n390824 );
buf ( n390826 , n365290 );
not ( n69879 , n390826 );
or ( n390828 , n390825 , n69879 );
buf ( n390829 , n45092 );
buf ( n390830 , n45336 );
nand ( n390831 , n390829 , n390830 );
buf ( n390832 , n390831 );
buf ( n390833 , n390832 );
nand ( n390834 , n390828 , n390833 );
buf ( n390835 , n390834 );
buf ( n390836 , n390835 );
nand ( n390837 , n390823 , n390836 );
buf ( n390838 , n390837 );
buf ( n390839 , n390838 );
nand ( n390840 , n390822 , n390839 );
buf ( n390841 , n390840 );
not ( n69894 , n390200 );
not ( n69895 , n69894 );
not ( n69896 , n50782 );
and ( n390845 , n69895 , n69896 );
buf ( n390846 , n56849 );
not ( n69899 , n390846 );
buf ( n390848 , n45915 );
not ( n390849 , n390848 );
or ( n69902 , n69899 , n390849 );
buf ( n390851 , n45916 );
buf ( n390852 , n63905 );
nand ( n390853 , n390851 , n390852 );
buf ( n390854 , n390853 );
buf ( n390855 , n390854 );
nand ( n69908 , n69902 , n390855 );
buf ( n390857 , n69908 );
and ( n390858 , n390857 , n366428 );
nor ( n69911 , n390845 , n390858 );
xor ( n69912 , n390841 , n69911 );
buf ( n390861 , n69912 );
not ( n69914 , n390861 );
not ( n69915 , n389963 );
not ( n69916 , n39208 );
or ( n390865 , n69915 , n69916 );
not ( n69918 , n365428 );
not ( n69919 , n366356 );
or ( n69920 , n69918 , n69919 );
buf ( n390869 , n366360 );
buf ( n390870 , n365422 );
nand ( n69923 , n390869 , n390870 );
buf ( n390872 , n69923 );
nand ( n69925 , n69920 , n390872 );
nand ( n69926 , n69925 , n46582 );
nand ( n69927 , n390865 , n69926 );
buf ( n390876 , n69927 );
not ( n69929 , n390876 );
and ( n69930 , n69914 , n69929 );
buf ( n390879 , n69927 );
buf ( n390880 , n69912 );
and ( n69933 , n390879 , n390880 );
nor ( n69934 , n69930 , n69933 );
buf ( n390883 , n69934 );
buf ( n390884 , n390883 );
xnor ( n69937 , n390817 , n390884 );
buf ( n390886 , n69937 );
buf ( n390887 , n390886 );
not ( n69940 , n47466 );
not ( n69941 , n69135 );
or ( n69942 , n69940 , n69941 );
buf ( n390891 , n365052 );
buf ( n390892 , n40199 );
and ( n69945 , n390891 , n390892 );
not ( n69946 , n390891 );
buf ( n390895 , n45523 );
and ( n69948 , n69946 , n390895 );
nor ( n69949 , n69945 , n69948 );
buf ( n390898 , n69949 );
buf ( n390899 , n390898 );
not ( n69952 , n390899 );
buf ( n390901 , n44915 );
nand ( n390902 , n69952 , n390901 );
buf ( n390903 , n390902 );
nand ( n69956 , n69942 , n390903 );
buf ( n390905 , n69956 );
buf ( n390906 , n45058 );
not ( n390907 , n390906 );
buf ( n390908 , n68788 );
not ( n69961 , n390908 );
or ( n69962 , n390907 , n69961 );
buf ( n390911 , n360885 );
not ( n390912 , n390911 );
buf ( n390913 , n365202 );
not ( n69966 , n390913 );
and ( n69967 , n390912 , n69966 );
buf ( n69968 , n383308 );
not ( n390917 , n69968 );
buf ( n390918 , n390917 );
buf ( n390919 , n390918 );
buf ( n390920 , n45065 );
and ( n69973 , n390919 , n390920 );
nor ( n390922 , n69967 , n69973 );
buf ( n390923 , n390922 );
buf ( n390924 , n390923 );
not ( n69977 , n390924 );
buf ( n390926 , n45075 );
nand ( n390927 , n69977 , n390926 );
buf ( n390928 , n390927 );
buf ( n390929 , n390928 );
nand ( n69982 , n69962 , n390929 );
buf ( n390931 , n69982 );
buf ( n390932 , n390931 );
xor ( n69985 , n390905 , n390932 );
buf ( n390934 , n365152 );
not ( n69987 , n390934 );
buf ( n390936 , n46397 );
not ( n69989 , n390936 );
not ( n69990 , n40251 );
buf ( n390939 , n69990 );
not ( n390940 , n390939 );
or ( n390941 , n69989 , n390940 );
buf ( n390942 , n360379 );
buf ( n390943 , n342909 );
nand ( n390944 , n390942 , n390943 );
buf ( n390945 , n390944 );
buf ( n390946 , n390945 );
nand ( n390947 , n390941 , n390946 );
buf ( n390948 , n390947 );
buf ( n390949 , n390948 );
not ( n390950 , n390949 );
or ( n390951 , n69987 , n390950 );
buf ( n390952 , n389876 );
buf ( n390953 , n390952 );
buf ( n390954 , n67451 );
buf ( n390955 , n390954 );
nand ( n390956 , n390953 , n390955 );
buf ( n390957 , n390956 );
buf ( n390958 , n390957 );
nand ( n390959 , n390951 , n390958 );
buf ( n390960 , n390959 );
buf ( n390961 , n390960 );
xor ( n390962 , n69985 , n390961 );
buf ( n390963 , n390962 );
buf ( n390964 , n390963 );
xor ( n390965 , n390887 , n390964 );
xor ( n390966 , n389720 , n389726 );
and ( n390967 , n390966 , n389738 );
and ( n390968 , n389720 , n389726 );
or ( n390969 , n390967 , n390968 );
buf ( n390970 , n390969 );
buf ( n390971 , n390970 );
xor ( n390972 , n390965 , n390971 );
buf ( n390973 , n390972 );
buf ( n390974 , n390973 );
xor ( n390975 , n69856 , n390974 );
buf ( n390976 , n390975 );
not ( n390977 , n390976 );
or ( n390978 , n390608 , n390977 );
not ( n390979 , n390976 );
nand ( n69997 , n390979 , n390606 );
nand ( n390981 , n390978 , n69997 );
not ( n69999 , n390981 );
xor ( n70000 , n390243 , n390260 );
and ( n390984 , n70000 , n390401 );
and ( n390985 , n390243 , n390260 );
or ( n70003 , n390984 , n390985 );
not ( n70004 , n390277 );
not ( n390988 , n390381 );
or ( n70006 , n70004 , n390988 );
not ( n70007 , n390277 );
not ( n390991 , n70007 );
not ( n70009 , n69433 );
or ( n390993 , n390991 , n70009 );
nand ( n70011 , n390993 , n390398 );
nand ( n70012 , n70006 , n70011 );
buf ( n390996 , n70012 );
buf ( n390997 , n389740 );
not ( n70015 , n390997 );
buf ( n390999 , n389694 );
not ( n391000 , n390999 );
or ( n391001 , n70015 , n391000 );
buf ( n391002 , n389740 );
buf ( n391003 , n389694 );
or ( n391004 , n391002 , n391003 );
buf ( n391005 , n68719 );
nand ( n391006 , n391004 , n391005 );
buf ( n391007 , n391006 );
buf ( n391008 , n391007 );
nand ( n391009 , n391001 , n391008 );
buf ( n391010 , n391009 );
buf ( n391011 , n391010 );
xor ( n391012 , n390996 , n391011 );
not ( n70030 , n390168 );
not ( n391014 , n390144 );
or ( n391015 , n70030 , n391014 );
not ( n70033 , n390144 );
not ( n70034 , n70033 );
not ( n391018 , n390171 );
or ( n70036 , n70034 , n391018 );
nand ( n70037 , n70036 , n69313 );
nand ( n391021 , n391015 , n70037 );
buf ( n391022 , n391021 );
buf ( n391023 , n379445 );
not ( n70041 , n391023 );
buf ( n391025 , n379296 );
not ( n70043 , n391025 );
or ( n391027 , n70041 , n70043 );
buf ( n391028 , n389646 );
nand ( n391029 , n391027 , n391028 );
buf ( n391030 , n391029 );
buf ( n391031 , n391030 );
nor ( n70049 , n391022 , n391031 );
buf ( n391033 , n70049 );
buf ( n391034 , n391033 );
not ( n70052 , n391034 );
buf ( n391036 , n391030 );
buf ( n391037 , n391021 );
nand ( n391038 , n391036 , n391037 );
buf ( n391039 , n391038 );
buf ( n391040 , n391039 );
nand ( n70058 , n70052 , n391040 );
buf ( n391042 , n70058 );
not ( n391043 , n69286 );
not ( n391044 , n390229 );
or ( n70062 , n391043 , n391044 );
buf ( n391046 , n390228 );
not ( n391047 , n391046 );
not ( n70065 , n69286 );
buf ( n391049 , n70065 );
not ( n391050 , n391049 );
or ( n70068 , n391047 , n391050 );
buf ( n391052 , n390191 );
nand ( n70070 , n70068 , n391052 );
buf ( n391054 , n70070 );
nand ( n391055 , n70062 , n391054 );
buf ( n391056 , n390076 );
not ( n70074 , n391056 );
buf ( n391058 , n363038 );
not ( n391059 , n391058 );
or ( n70077 , n70074 , n391059 );
buf ( n391061 , n362521 );
buf ( n391062 , n377353 );
not ( n70080 , n391062 );
buf ( n391064 , n45231 );
not ( n70082 , n391064 );
or ( n70083 , n70080 , n70082 );
buf ( n391067 , n45234 );
buf ( n391068 , n377352 );
nand ( n70086 , n391067 , n391068 );
buf ( n391070 , n70086 );
buf ( n391071 , n391070 );
nand ( n70089 , n70083 , n391071 );
buf ( n391073 , n70089 );
buf ( n391074 , n391073 );
nand ( n70092 , n391061 , n391074 );
buf ( n391076 , n70092 );
buf ( n391077 , n391076 );
nand ( n70095 , n70077 , n391077 );
buf ( n391079 , n70095 );
buf ( n391080 , n391079 );
not ( n391081 , n391080 );
buf ( n391082 , n391081 );
xor ( n391083 , n391055 , n391082 );
buf ( n391084 , n48490 );
not ( n391085 , n391084 );
buf ( n391086 , n362423 );
not ( n391087 , n391086 );
buf ( n391088 , n367575 );
not ( n391089 , n391088 );
or ( n70107 , n391087 , n391089 );
buf ( n391091 , n364827 );
buf ( n70109 , n377715 );
nand ( n70110 , n391091 , n70109 );
buf ( n70111 , n70110 );
buf ( n391095 , n70111 );
nand ( n70113 , n70107 , n391095 );
buf ( n391097 , n70113 );
buf ( n391098 , n391097 );
not ( n391099 , n391098 );
or ( n70116 , n391085 , n391099 );
buf ( n391101 , n368706 );
buf ( n391102 , n68866 );
nand ( n391103 , n391101 , n391102 );
buf ( n391104 , n391103 );
buf ( n391105 , n391104 );
nand ( n70121 , n70116 , n391105 );
buf ( n391107 , n70121 );
buf ( n391108 , n391107 );
buf ( n391109 , n43261 );
not ( n70125 , n391109 );
buf ( n391111 , n370021 );
not ( n391112 , n391111 );
or ( n391113 , n70125 , n391112 );
buf ( n391114 , n69294 );
not ( n391115 , n391114 );
buf ( n391116 , n363429 );
nand ( n391117 , n391115 , n391116 );
buf ( n391118 , n391117 );
buf ( n391119 , n391118 );
nand ( n391120 , n391113 , n391119 );
buf ( n391121 , n391120 );
buf ( n391122 , n391121 );
xor ( n391123 , n391108 , n391122 );
buf ( n391124 , n366317 );
buf ( n391125 , n390186 );
or ( n391126 , n391124 , n391125 );
buf ( n391127 , n365312 );
not ( n391128 , n361911 );
not ( n391129 , n352194 );
and ( n391130 , n391128 , n391129 );
buf ( n391131 , n365319 );
not ( n391132 , n391131 );
not ( n391133 , n45125 );
buf ( n391134 , n391133 );
nor ( n391135 , n391132 , n391134 );
buf ( n391136 , n391135 );
nor ( n391137 , n391130 , n391136 );
buf ( n391138 , n391137 );
or ( n70131 , n391127 , n391138 );
nand ( n70132 , n391126 , n70131 );
buf ( n391141 , n70132 );
buf ( n391142 , n391141 );
xor ( n70135 , n391123 , n391142 );
buf ( n391144 , n70135 );
xor ( n70137 , n391083 , n391144 );
buf ( n391146 , n70137 );
not ( n391147 , n391146 );
buf ( n391148 , n391147 );
and ( n391149 , n391042 , n391148 );
not ( n70142 , n391042 );
and ( n391151 , n70142 , n70137 );
nor ( n70144 , n391149 , n391151 );
buf ( n391153 , n70144 );
not ( n391154 , n390375 );
not ( n391155 , n390313 );
not ( n70148 , n391155 );
and ( n391157 , n391154 , n70148 );
nand ( n391158 , n390375 , n391155 );
buf ( n70151 , n69368 );
and ( n391160 , n391158 , n70151 );
nor ( n391161 , n391157 , n391160 );
not ( n70154 , n391161 );
buf ( n391163 , n70154 );
xor ( n70156 , n391153 , n391163 );
buf ( n391165 , n389650 );
buf ( n391166 , n389675 );
or ( n391167 , n391165 , n391166 );
buf ( n391168 , n391167 );
not ( n391169 , n391168 );
buf ( n391170 , n389691 );
buf ( n70163 , n391170 );
buf ( n70164 , n70163 );
not ( n391173 , n70164 );
or ( n70166 , n391169 , n391173 );
buf ( n391175 , n389675 );
buf ( n391176 , n389650 );
and ( n70169 , n391175 , n391176 );
buf ( n391178 , n70169 );
not ( n70171 , n391178 );
nand ( n391180 , n70166 , n70171 );
buf ( n391181 , n391180 );
xor ( n391182 , n70156 , n391181 );
buf ( n391183 , n391182 );
buf ( n391184 , n391183 );
xnor ( n70177 , n391012 , n391184 );
buf ( n391186 , n70177 );
not ( n391187 , n391186 );
and ( n70180 , n70003 , n391187 );
not ( n70181 , n70003 );
and ( n391190 , n70181 , n391186 );
nor ( n70183 , n70180 , n391190 );
not ( n391192 , n70183 );
xor ( n70185 , n68833 , n68839 );
and ( n70186 , n70185 , n390013 );
and ( n391195 , n68833 , n68839 );
or ( n70188 , n70186 , n391195 );
not ( n391197 , n70188 );
or ( n70190 , n391192 , n391197 );
buf ( n391199 , n70183 );
not ( n391200 , n391199 );
buf ( n391201 , n391200 );
buf ( n391202 , n391201 );
buf ( n391203 , n70188 );
not ( n391204 , n391203 );
buf ( n391205 , n391204 );
buf ( n391206 , n391205 );
nand ( n391207 , n391202 , n391206 );
buf ( n391208 , n391207 );
nand ( n70201 , n70190 , n391208 );
not ( n391210 , n70201 );
or ( n391211 , n69999 , n391210 );
not ( n70204 , n390981 );
not ( n391213 , n70204 );
not ( n391214 , n70201 );
not ( n70207 , n391214 );
or ( n391216 , n391213 , n70207 );
buf ( n391217 , n69455 );
not ( n391218 , n391217 );
not ( n70211 , n69093 );
or ( n391220 , n391218 , n70211 );
buf ( n70213 , n69455 );
or ( n391222 , n69093 , n70213 );
buf ( n391223 , n390021 );
not ( n70216 , n391223 );
buf ( n70217 , n70216 );
nand ( n391226 , n391222 , n70217 );
nand ( n391227 , n391220 , n391226 );
nand ( n391228 , n391216 , n391227 );
nand ( n70221 , n391211 , n391228 );
buf ( n391230 , n70221 );
not ( n70223 , n391230 );
not ( n391232 , n390898 );
not ( n391233 , n44913 );
and ( n70226 , n391232 , n391233 );
not ( n70227 , n365041 );
not ( n70228 , n364987 );
or ( n70229 , n70227 , n70228 );
buf ( n391238 , n359778 );
buf ( n391239 , n365052 );
nand ( n70232 , n391238 , n391239 );
buf ( n391241 , n70232 );
nand ( n391242 , n70229 , n391241 );
and ( n391243 , n391242 , n44915 );
nor ( n70236 , n70226 , n391243 );
buf ( n391245 , n70236 );
not ( n70238 , n391245 );
buf ( n391247 , n70238 );
buf ( n391248 , n390525 );
not ( n70241 , n391248 );
buf ( n391250 , n70241 );
buf ( n391251 , n391250 );
not ( n391252 , n391251 );
buf ( n391253 , n390543 );
not ( n70246 , n391253 );
or ( n391255 , n391252 , n70246 );
buf ( n391256 , n69614 );
nand ( n70249 , n391255 , n391256 );
buf ( n391258 , n70249 );
buf ( n391259 , n391258 );
buf ( n391260 , n390540 );
buf ( n391261 , n390525 );
nand ( n70254 , n391260 , n391261 );
buf ( n391263 , n70254 );
buf ( n391264 , n391263 );
and ( n70257 , n391259 , n391264 );
buf ( n391266 , n70257 );
xor ( n391267 , n391247 , n391266 );
xor ( n70260 , n391108 , n391122 );
and ( n391269 , n70260 , n391142 );
and ( n391270 , n391108 , n391122 );
or ( n70263 , n391269 , n391270 );
buf ( n391272 , n70263 );
not ( n70265 , n391272 );
not ( n391274 , n390523 );
not ( n70267 , n359916 );
or ( n391276 , n391274 , n70267 );
and ( n70269 , n368994 , n364919 );
not ( n70270 , n368994 );
and ( n391279 , n70270 , n44743 );
nor ( n391280 , n70269 , n391279 );
not ( n70273 , n391280 );
nand ( n391282 , n70273 , n371846 );
nand ( n70275 , n391276 , n391282 );
not ( n70276 , n70275 );
not ( n70277 , n70276 );
or ( n70278 , n70265 , n70277 );
not ( n70279 , n391272 );
nand ( n70280 , n70279 , n70275 );
nand ( n70281 , n70278 , n70280 );
not ( n70282 , n48490 );
not ( n70283 , n369881 );
or ( n70284 , n70282 , n70283 );
nand ( n391293 , n49669 , n391097 );
nand ( n70286 , n70284 , n391293 );
not ( n70287 , n49689 );
not ( n70288 , n70287 );
not ( n70289 , n41835 );
or ( n391298 , n70288 , n70289 );
not ( n391299 , n391137 );
nand ( n70292 , n391299 , n46135 );
nand ( n391301 , n391298 , n70292 );
xor ( n391302 , n70286 , n391301 );
buf ( n391303 , n365622 );
buf ( n391304 , n365440 );
not ( n391305 , n391304 );
buf ( n391306 , n44634 );
not ( n391307 , n391306 );
or ( n70300 , n391305 , n391307 );
buf ( n391309 , n45455 );
buf ( n391310 , n365452 );
nand ( n70303 , n391309 , n391310 );
buf ( n391312 , n70303 );
buf ( n391313 , n391312 );
nand ( n391314 , n70300 , n391313 );
buf ( n391315 , n391314 );
buf ( n391316 , n391315 );
nand ( n70309 , n391303 , n391316 );
buf ( n391318 , n70309 );
nand ( n391319 , n390747 , n362027 );
and ( n70312 , n391318 , n391319 );
xnor ( n70313 , n391302 , n70312 );
and ( n391322 , n70281 , n70313 );
not ( n391323 , n70281 );
not ( n70316 , n70313 );
and ( n391325 , n391323 , n70316 );
nor ( n391326 , n391322 , n391325 );
xnor ( n391327 , n391267 , n391326 );
buf ( n391328 , n391327 );
buf ( n391329 , n57530 );
not ( n391330 , n391329 );
buf ( n391331 , n390504 );
not ( n70324 , n391331 );
or ( n391333 , n391330 , n70324 );
not ( n391334 , n377585 );
not ( n70327 , n40083 );
not ( n70328 , n39039 );
or ( n70329 , n70327 , n70328 );
nand ( n70330 , n70329 , n53517 );
not ( n70331 , n70330 );
or ( n70332 , n391334 , n70331 );
or ( n70333 , n70330 , n377585 );
nand ( n391342 , n70332 , n70333 );
nand ( n70335 , n391342 , n377580 );
buf ( n391344 , n70335 );
nand ( n391345 , n391333 , n391344 );
buf ( n391346 , n391345 );
buf ( n391347 , n391346 );
buf ( n391348 , n387542 );
not ( n391349 , n391348 );
and ( n70342 , n368549 , n359939 );
not ( n70343 , n368549 );
and ( n391352 , n70343 , n371416 );
or ( n391353 , n70342 , n391352 );
buf ( n391354 , n391353 );
not ( n70347 , n391354 );
or ( n70348 , n391349 , n70347 );
nand ( n391357 , n390459 , n368611 );
buf ( n391358 , n391357 );
nand ( n391359 , n70348 , n391358 );
buf ( n391360 , n391359 );
buf ( n391361 , n391360 );
xor ( n70354 , n391347 , n391361 );
buf ( n391363 , n390809 );
not ( n391364 , n391363 );
buf ( n391365 , n391364 );
buf ( n391366 , n391365 );
not ( n391367 , n391366 );
buf ( n391368 , n390883 );
not ( n391369 , n391368 );
or ( n70362 , n391367 , n391369 );
buf ( n391371 , n390815 );
nand ( n70364 , n70362 , n391371 );
buf ( n391373 , n70364 );
buf ( n391374 , n391373 );
buf ( n391375 , n390883 );
buf ( n391376 , n391365 );
or ( n70369 , n391375 , n391376 );
buf ( n391378 , n70369 );
buf ( n391379 , n391378 );
nand ( n70372 , n391374 , n391379 );
buf ( n70373 , n70372 );
buf ( n391382 , n70373 );
xor ( n391383 , n70354 , n391382 );
buf ( n391384 , n391383 );
buf ( n391385 , n391384 );
xor ( n391386 , n391328 , n391385 );
buf ( n391387 , n390800 );
not ( n70380 , n391387 );
buf ( n391389 , n69840 );
not ( n391390 , n391389 );
or ( n70383 , n70380 , n391390 );
not ( n70384 , n69847 );
not ( n70385 , n69675 );
or ( n391394 , n70384 , n70385 );
buf ( n391395 , n390628 );
nand ( n70388 , n391394 , n391395 );
buf ( n391397 , n70388 );
nand ( n391398 , n70383 , n391397 );
buf ( n391399 , n391398 );
buf ( n391400 , n391399 );
xor ( n391401 , n391386 , n391400 );
buf ( n391402 , n391401 );
buf ( n391403 , n391402 );
xor ( n391404 , n390614 , n390803 );
and ( n70397 , n391404 , n390974 );
and ( n70398 , n390614 , n390803 );
or ( n70399 , n70397 , n70398 );
buf ( n391408 , n70399 );
buf ( n391409 , n391408 );
xor ( n70402 , n391403 , n391409 );
not ( n70403 , n69755 );
buf ( n391412 , n69827 );
not ( n391413 , n391412 );
or ( n70406 , n70403 , n391413 );
not ( n70407 , n390776 );
not ( n391416 , n390702 );
or ( n391417 , n70407 , n391416 );
nand ( n70410 , n391417 , n390781 );
nand ( n70411 , n70406 , n70410 );
not ( n70412 , n70411 );
not ( n391421 , n70412 );
not ( n70414 , n45553 );
not ( n70415 , n390533 );
or ( n70416 , n70414 , n70415 );
buf ( n391425 , n365676 );
not ( n70418 , n391425 );
buf ( n391427 , n369343 );
not ( n70420 , n391427 );
or ( n391429 , n70418 , n70420 );
buf ( n391430 , n369352 );
buf ( n391431 , n365673 );
nand ( n70424 , n391430 , n391431 );
buf ( n391433 , n70424 );
buf ( n391434 , n391433 );
nand ( n70427 , n391429 , n391434 );
buf ( n391436 , n70427 );
buf ( n391437 , n391436 );
buf ( n391438 , n45492 );
nand ( n70431 , n391437 , n391438 );
buf ( n391440 , n70431 );
nand ( n391441 , n70416 , n391440 );
buf ( n391442 , n391441 );
buf ( n391443 , n390555 );
not ( n391444 , n391443 );
buf ( n391445 , n391444 );
buf ( n391446 , n391445 );
not ( n70439 , n391446 );
buf ( n391448 , n390729 );
buf ( n70441 , n391448 );
buf ( n391450 , n70441 );
buf ( n391451 , n391450 );
not ( n70444 , n391451 );
or ( n391453 , n70439 , n70444 );
buf ( n391454 , n391450 );
buf ( n391455 , n391445 );
or ( n391456 , n391454 , n391455 );
buf ( n391457 , n69803 );
nand ( n70450 , n391456 , n391457 );
buf ( n391459 , n70450 );
buf ( n391460 , n391459 );
nand ( n391461 , n391453 , n391460 );
buf ( n391462 , n391461 );
buf ( n391463 , n391462 );
xor ( n391464 , n391442 , n391463 );
buf ( n391465 , n49828 );
buf ( n391466 , n390835 );
not ( n70459 , n391466 );
buf ( n391468 , n372247 );
not ( n391469 , n391468 );
or ( n391470 , n70459 , n391469 );
buf ( n391471 , n370059 );
not ( n70464 , n391471 );
buf ( n391473 , n365303 );
nand ( n391474 , n70464 , n391473 );
buf ( n391475 , n391474 );
buf ( n391476 , n391475 );
nand ( n391477 , n391470 , n391476 );
buf ( n391478 , n391477 );
buf ( n391479 , n391478 );
xor ( n70472 , n391465 , n391479 );
buf ( n391481 , n366402 );
not ( n391482 , n391481 );
buf ( n391483 , n390857 );
not ( n70476 , n391483 );
or ( n391485 , n391482 , n70476 );
not ( n391486 , n342656 );
not ( n70479 , n362537 );
or ( n70480 , n391486 , n70479 );
nand ( n391489 , n63905 , n362534 );
nand ( n391490 , n70480 , n391489 );
buf ( n391491 , n391490 );
buf ( n391492 , n366428 );
nand ( n70485 , n391491 , n391492 );
buf ( n391494 , n70485 );
buf ( n391495 , n391494 );
nand ( n70488 , n391485 , n391495 );
buf ( n391497 , n70488 );
buf ( n391498 , n391497 );
xnor ( n391499 , n70472 , n391498 );
buf ( n391500 , n391499 );
buf ( n391501 , n391500 );
xor ( n391502 , n391464 , n391501 );
buf ( n391503 , n391502 );
buf ( n391504 , n391503 );
not ( n391505 , n391504 );
buf ( n391506 , n391505 );
not ( n70499 , n391506 );
or ( n70500 , n391421 , n70499 );
nand ( n391509 , n391503 , n70411 );
nand ( n391510 , n70500 , n391509 );
not ( n391511 , n390923 );
not ( n70504 , n365227 );
and ( n70505 , n391511 , n70504 );
buf ( n391514 , n342881 );
not ( n391515 , n391514 );
buf ( n391516 , n366676 );
not ( n391517 , n391516 );
or ( n391518 , n391515 , n391517 );
buf ( n391519 , n377990 );
buf ( n391520 , n45065 );
nand ( n391521 , n391519 , n391520 );
buf ( n391522 , n391521 );
buf ( n391523 , n391522 );
nand ( n391524 , n391518 , n391523 );
buf ( n391525 , n391524 );
and ( n391526 , n391525 , n45075 );
nor ( n70519 , n70505 , n391526 );
not ( n391528 , n70519 );
buf ( n391529 , n390841 );
not ( n70522 , n391529 );
buf ( n391531 , n69911 );
nand ( n391532 , n70522 , n391531 );
buf ( n391533 , n391532 );
not ( n70526 , n391533 );
not ( n70527 , n69927 );
or ( n391536 , n70526 , n70527 );
buf ( n391537 , n69911 );
not ( n391538 , n391537 );
buf ( n391539 , n390841 );
nand ( n391540 , n391538 , n391539 );
buf ( n391541 , n391540 );
nand ( n391542 , n391536 , n391541 );
not ( n391543 , n391542 );
or ( n70536 , n391528 , n391543 );
not ( n70537 , n70519 );
not ( n391546 , n391542 );
nand ( n391547 , n70537 , n391546 );
nand ( n70540 , n70536 , n391547 );
buf ( n391549 , n390649 );
not ( n70542 , n391549 );
buf ( n391551 , n70542 );
not ( n391552 , n391551 );
not ( n70545 , n390693 );
or ( n391554 , n391552 , n70545 );
buf ( n391555 , n390696 );
not ( n70548 , n391555 );
buf ( n70549 , n390649 );
buf ( n391558 , n70549 );
not ( n391559 , n391558 );
or ( n70552 , n70548 , n391559 );
buf ( n391561 , n69719 );
nand ( n391562 , n70552 , n391561 );
buf ( n391563 , n391562 );
nand ( n70556 , n391554 , n391563 );
not ( n391565 , n70556 );
and ( n391566 , n70540 , n391565 );
not ( n70559 , n70540 );
and ( n70560 , n70559 , n70556 );
nor ( n391569 , n391566 , n70560 );
not ( n391570 , n391569 );
and ( n70563 , n391510 , n391570 );
not ( n70564 , n391510 );
and ( n70565 , n70564 , n391569 );
nor ( n391574 , n70563 , n70565 );
buf ( n391575 , n391574 );
buf ( n391576 , n390886 );
not ( n70569 , n391576 );
buf ( n391578 , n390963 );
not ( n391579 , n391578 );
or ( n391580 , n70569 , n391579 );
buf ( n391581 , n390963 );
buf ( n391582 , n390886 );
or ( n70575 , n391581 , n391582 );
buf ( n391584 , n390970 );
nand ( n70577 , n70575 , n391584 );
buf ( n391586 , n70577 );
buf ( n391587 , n391586 );
nand ( n391588 , n391580 , n391587 );
buf ( n391589 , n391588 );
buf ( n391590 , n391589 );
xor ( n70583 , n391575 , n391590 );
not ( n391592 , n391180 );
not ( n391593 , n70154 );
or ( n70586 , n391592 , n391593 );
not ( n70587 , n391161 );
and ( n391596 , n70164 , n391168 );
nor ( n391597 , n391596 , n391178 );
not ( n391598 , n391597 );
or ( n70591 , n70587 , n391598 );
not ( n391600 , n70144 );
nand ( n391601 , n70591 , n391600 );
nand ( n70594 , n70586 , n391601 );
buf ( n391603 , n70594 );
xor ( n391604 , n70583 , n391603 );
buf ( n391605 , n391604 );
buf ( n391606 , n391605 );
buf ( n391607 , n391606 );
xnor ( n70600 , n70402 , n391607 );
buf ( n391609 , n70600 );
buf ( n391610 , n391609 );
buf ( n391611 , n70012 );
buf ( n70604 , n391611 );
buf ( n70605 , n70604 );
nor ( n391614 , n70605 , n391010 );
or ( n391615 , n391614 , n391183 );
buf ( n391616 , n391010 );
buf ( n391617 , n70605 );
nand ( n391618 , n391616 , n391617 );
buf ( n391619 , n391618 );
nand ( n70612 , n391615 , n391619 );
not ( n391621 , n70612 );
buf ( n70614 , n391621 );
buf ( n70615 , n70137 );
buf ( n70616 , n391033 );
or ( n70617 , n70615 , n70616 );
buf ( n70618 , n391039 );
nand ( n391627 , n70617 , n70618 );
buf ( n391628 , n391627 );
buf ( n391629 , n391628 );
xor ( n391630 , n390905 , n390932 );
and ( n391631 , n391630 , n390961 );
and ( n70624 , n390905 , n390932 );
or ( n70625 , n391631 , n70624 );
buf ( n391634 , n70625 );
buf ( n391635 , n391634 );
xor ( n391636 , n391629 , n391635 );
buf ( n391637 , n391079 );
buf ( n391638 , n391055 );
or ( n70631 , n391637 , n391638 );
buf ( n391640 , n391144 );
nand ( n391641 , n70631 , n391640 );
buf ( n391642 , n391641 );
buf ( n391643 , n391642 );
buf ( n391644 , n391079 );
buf ( n391645 , n391055 );
nand ( n391646 , n391644 , n391645 );
buf ( n391647 , n391646 );
buf ( n391648 , n391647 );
nand ( n391649 , n391643 , n391648 );
buf ( n391650 , n391649 );
buf ( n391651 , n391650 );
buf ( n391652 , n390954 );
not ( n391653 , n391652 );
buf ( n391654 , n390948 );
not ( n391655 , n391654 );
or ( n391656 , n391653 , n391655 );
and ( n70649 , n366722 , n387355 );
not ( n70650 , n366722 );
and ( n391659 , n70650 , n46397 );
or ( n391660 , n70649 , n391659 );
buf ( n391661 , n391660 );
buf ( n391662 , n365152 );
nand ( n391663 , n391661 , n391662 );
buf ( n391664 , n391663 );
buf ( n391665 , n391664 );
nand ( n70658 , n391656 , n391665 );
buf ( n391667 , n70658 );
buf ( n391668 , n391667 );
xor ( n391669 , n391651 , n391668 );
buf ( n391670 , n49609 );
not ( n70663 , n391670 );
buf ( n391672 , n369769 );
not ( n391673 , n391672 );
buf ( n391674 , n41406 );
not ( n70667 , n391674 );
buf ( n391676 , n70667 );
buf ( n391677 , n391676 );
not ( n391678 , n391677 );
or ( n70671 , n391673 , n391678 );
buf ( n391680 , n365170 );
buf ( n391681 , n369766 );
nand ( n70674 , n391680 , n391681 );
buf ( n391683 , n70674 );
buf ( n391684 , n391683 );
nand ( n70677 , n70671 , n391684 );
buf ( n391686 , n70677 );
buf ( n391687 , n391686 );
not ( n70680 , n391687 );
or ( n391689 , n70663 , n70680 );
or ( n391690 , n363171 , n369769 );
or ( n391691 , n41907 , n369766 );
nand ( n70684 , n391690 , n391691 , n369804 );
buf ( n70685 , n70684 );
nand ( n391694 , n391689 , n70685 );
buf ( n391695 , n391694 );
buf ( n391696 , n391695 );
xor ( n391697 , n391669 , n391696 );
buf ( n391698 , n391697 );
buf ( n391699 , n391698 );
xor ( n70692 , n391636 , n391699 );
buf ( n391701 , n70692 );
buf ( n391702 , n391701 );
not ( n70695 , n69517 );
not ( n70696 , n390469 );
or ( n391705 , n70695 , n70696 );
not ( n391706 , n390451 );
not ( n70699 , n69523 );
or ( n70700 , n391706 , n70699 );
nand ( n70701 , n70700 , n390438 );
nand ( n391710 , n391705 , n70701 );
buf ( n391711 , n69925 );
not ( n70704 , n391711 );
buf ( n391713 , n39208 );
not ( n70706 , n391713 );
or ( n391715 , n70704 , n70706 );
buf ( n70708 , n359312 );
buf ( n391717 , n365980 );
not ( n70710 , n391717 );
buf ( n391719 , n355579 );
not ( n391720 , n391719 );
or ( n70713 , n70710 , n391720 );
buf ( n391722 , n365367 );
buf ( n391723 , n365989 );
nand ( n391724 , n391722 , n391723 );
buf ( n391725 , n391724 );
buf ( n391726 , n391725 );
nand ( n70719 , n70713 , n391726 );
buf ( n391728 , n70719 );
buf ( n391729 , n391728 );
nand ( n70722 , n70708 , n391729 );
buf ( n391731 , n70722 );
buf ( n391732 , n391731 );
nand ( n70725 , n391715 , n391732 );
buf ( n391734 , n70725 );
not ( n70727 , n391734 );
buf ( n391736 , n390722 );
not ( n70729 , n391736 );
buf ( n391738 , n361606 );
not ( n70731 , n391738 );
or ( n70732 , n70729 , n70731 );
nand ( n70733 , n367590 , n369916 );
buf ( n391742 , n70733 );
nand ( n70735 , n70732 , n391742 );
buf ( n391744 , n70735 );
buf ( n391745 , n391744 );
buf ( n391746 , n45983 );
not ( n70739 , n391746 );
buf ( n391748 , n390643 );
not ( n70741 , n391748 );
and ( n70742 , n70739 , n70741 );
buf ( n391751 , n365471 );
not ( n391752 , n391751 );
buf ( n391753 , n364915 );
not ( n391754 , n391753 );
and ( n70747 , n391752 , n391754 );
buf ( n391756 , n362452 );
buf ( n391757 , n364915 );
and ( n70750 , n391756 , n391757 );
nor ( n70751 , n70747 , n70750 );
buf ( n391760 , n70751 );
buf ( n70753 , n391760 );
buf ( n70754 , n366754 );
nor ( n70755 , n70753 , n70754 );
buf ( n70756 , n70755 );
buf ( n70757 , n70756 );
nor ( n70758 , n70742 , n70757 );
buf ( n70759 , n70758 );
buf ( n70760 , n70759 );
nand ( n70761 , n391745 , n70760 );
buf ( n391770 , n70761 );
buf ( n391771 , n391744 );
not ( n70764 , n391771 );
buf ( n391773 , n70764 );
buf ( n391774 , n70759 );
not ( n70767 , n391774 );
buf ( n70768 , n70767 );
nand ( n70769 , n391773 , n70768 );
nand ( n70770 , n391770 , n70769 );
not ( n70771 , n70770 );
or ( n70772 , n70727 , n70771 );
not ( n391781 , n391734 );
nand ( n70774 , n391770 , n70769 , n391781 );
nand ( n391783 , n70772 , n70774 );
buf ( n391784 , n391783 );
not ( n391785 , n391784 );
buf ( n391786 , n391785 );
buf ( n391787 , n391786 );
not ( n70780 , n391787 );
buf ( n391789 , n365115 );
not ( n70782 , n391789 );
buf ( n391791 , n44819 );
not ( n391792 , n391791 );
buf ( n391793 , n370566 );
not ( n70786 , n391793 );
or ( n391795 , n391792 , n70786 );
buf ( n391796 , n42149 );
buf ( n391797 , n364994 );
nand ( n70790 , n391796 , n391797 );
buf ( n391799 , n70790 );
buf ( n391800 , n391799 );
nand ( n70793 , n391795 , n391800 );
buf ( n391802 , n70793 );
buf ( n391803 , n391802 );
not ( n70796 , n391803 );
or ( n391805 , n70782 , n70796 );
buf ( n391806 , n69820 );
buf ( n391807 , n365033 );
nand ( n391808 , n391806 , n391807 );
buf ( n391809 , n391808 );
buf ( n391810 , n391809 );
nand ( n70803 , n391805 , n391810 );
buf ( n391812 , n70803 );
buf ( n391813 , n391812 );
not ( n391814 , n391813 );
buf ( n391815 , n391814 );
buf ( n391816 , n391815 );
not ( n391817 , n391816 );
or ( n70810 , n70780 , n391817 );
buf ( n391819 , n391812 );
buf ( n391820 , n391783 );
nand ( n70813 , n391819 , n391820 );
buf ( n391822 , n70813 );
buf ( n391823 , n391822 );
nand ( n70816 , n70810 , n391823 );
buf ( n391825 , n70816 );
buf ( n391826 , n391825 );
not ( n70819 , n390660 );
not ( n391828 , n70819 );
not ( n391829 , n371300 );
and ( n70822 , n391828 , n391829 );
buf ( n391831 , n46477 );
not ( n391832 , n391831 );
buf ( n391833 , n369282 );
not ( n70826 , n391833 );
or ( n391835 , n391832 , n70826 );
buf ( n391836 , n365757 );
buf ( n391837 , n366683 );
nand ( n391838 , n391836 , n391837 );
buf ( n391839 , n391838 );
buf ( n391840 , n391839 );
nand ( n70833 , n391835 , n391840 );
buf ( n391842 , n70833 );
and ( n70835 , n391842 , n366654 );
nor ( n70836 , n70822 , n70835 );
not ( n70837 , n45345 );
not ( n70838 , n390686 );
or ( n70839 , n70837 , n70838 );
not ( n391848 , n365393 );
nand ( n70841 , n391848 , n365507 );
not ( n391850 , n70841 );
buf ( n391851 , n363119 );
not ( n70844 , n391851 );
buf ( n391853 , n365393 );
nand ( n391854 , n70844 , n391853 );
buf ( n391855 , n391854 );
not ( n391856 , n391855 );
or ( n70849 , n391850 , n391856 );
nand ( n70850 , n70849 , n365954 );
nand ( n391859 , n70839 , n70850 );
not ( n70852 , n391859 );
xor ( n391861 , n70836 , n70852 );
not ( n70854 , n391073 );
not ( n391863 , n359809 );
or ( n391864 , n70854 , n391863 );
buf ( n391865 , n362521 );
buf ( n391866 , n56970 );
not ( n391867 , n391866 );
buf ( n391868 , n361631 );
not ( n70861 , n391868 );
or ( n391870 , n391867 , n70861 );
buf ( n391871 , n45234 );
buf ( n391872 , n377389 );
nand ( n391873 , n391871 , n391872 );
buf ( n391874 , n391873 );
buf ( n391875 , n391874 );
nand ( n70868 , n391870 , n391875 );
buf ( n70869 , n70868 );
buf ( n391878 , n70869 );
nand ( n70871 , n391865 , n391878 );
buf ( n70872 , n70871 );
nand ( n391881 , n391864 , n70872 );
xnor ( n70874 , n391861 , n391881 );
buf ( n391883 , n70874 );
and ( n70876 , n391826 , n391883 );
not ( n391885 , n391826 );
buf ( n391886 , n70874 );
not ( n70879 , n391886 );
buf ( n391888 , n70879 );
buf ( n391889 , n391888 );
and ( n70882 , n391885 , n391889 );
nor ( n391891 , n70876 , n70882 );
buf ( n391892 , n391891 );
xor ( n70885 , n391710 , n391892 );
xor ( n391894 , n390493 , n390507 );
and ( n391895 , n391894 , n390566 );
and ( n70888 , n390493 , n390507 );
or ( n391897 , n391895 , n70888 );
buf ( n391898 , n391897 );
xor ( n70891 , n70885 , n391898 );
buf ( n70892 , n70891 );
not ( n391901 , n70892 );
buf ( n391902 , n391901 );
buf ( n391903 , n391902 );
xor ( n391904 , n391702 , n391903 );
buf ( n391905 , n69526 );
buf ( n391906 , n390568 );
or ( n391907 , n391905 , n391906 );
buf ( n391908 , n391907 );
buf ( n391909 , n391908 );
buf ( n391910 , n69632 );
and ( n391911 , n391909 , n391910 );
and ( n391912 , n390474 , n390569 );
buf ( n391913 , n391912 );
buf ( n391914 , n391913 );
nor ( n70907 , n391911 , n391914 );
buf ( n391916 , n70907 );
buf ( n391917 , n391916 );
not ( n70910 , n391917 );
buf ( n391919 , n70910 );
buf ( n391920 , n391919 );
xnor ( n391921 , n391904 , n391920 );
buf ( n391922 , n391921 );
buf ( n391923 , n391922 );
xor ( n70916 , n70614 , n391923 );
buf ( n391925 , n390603 );
buf ( n391926 , n69636 );
or ( n391927 , n391925 , n391926 );
buf ( n391928 , n391927 );
buf ( n391929 , n391928 );
buf ( n391930 , n390976 );
and ( n391931 , n391929 , n391930 );
and ( n70924 , n390585 , n390604 );
buf ( n391933 , n70924 );
buf ( n70926 , n391933 );
nor ( n70927 , n391931 , n70926 );
buf ( n70928 , n70927 );
buf ( n391937 , n70928 );
xor ( n70930 , n70916 , n391937 );
buf ( n391939 , n70930 );
buf ( n391940 , n391939 );
xor ( n391941 , n391610 , n391940 );
buf ( n391942 , n391186 );
not ( n391943 , n391942 );
buf ( n391944 , n391943 );
buf ( n391945 , n391944 );
buf ( n391946 , n70003 );
not ( n391947 , n391946 );
buf ( n391948 , n391947 );
buf ( n391949 , n391948 );
nand ( n391950 , n391945 , n391949 );
buf ( n391951 , n391950 );
buf ( n391952 , n391951 );
buf ( n391953 , n70188 );
and ( n70946 , n391952 , n391953 );
buf ( n391955 , n391944 );
buf ( n391956 , n391948 );
nor ( n70949 , n391955 , n391956 );
buf ( n391958 , n70949 );
buf ( n391959 , n391958 );
nor ( n391960 , n70946 , n391959 );
buf ( n391961 , n391960 );
buf ( n391962 , n391961 );
xor ( n70955 , n391941 , n391962 );
buf ( n391964 , n70955 );
buf ( n70957 , n391964 );
not ( n391966 , n70957 );
buf ( n391967 , n391966 );
not ( n391968 , n391967 );
or ( n70961 , n70223 , n391968 );
xor ( n391970 , n390981 , n70201 );
xnor ( n70963 , n391970 , n391227 );
not ( n70964 , n70963 );
xor ( n70965 , n389603 , n389620 );
and ( n391974 , n70965 , n390412 );
and ( n391975 , n389603 , n389620 );
or ( n70968 , n391974 , n391975 );
buf ( n391977 , n70968 );
buf ( n391978 , n391977 );
not ( n70971 , n391978 );
buf ( n70972 , n70971 );
nand ( n391981 , n70964 , n70972 );
nand ( n70974 , n70961 , n391981 );
not ( n391983 , n70974 );
nand ( n70975 , n67823 , n69486 , n391983 );
xor ( n391985 , n369168 , n370117 );
xor ( n391986 , n391985 , n370128 );
buf ( n391987 , n391986 );
not ( n70979 , n391987 );
xor ( n70980 , n369139 , n48924 );
xnor ( n391990 , n70980 , n369148 );
not ( n391991 , n391990 );
xor ( n70983 , n369443 , n369669 );
xor ( n70984 , n70983 , n369673 );
buf ( n391994 , n70984 );
buf ( n391995 , n391994 );
not ( n391996 , n391995 );
buf ( n391997 , n391996 );
not ( n70989 , n391997 );
buf ( n391999 , n368478 );
not ( n392000 , n391999 );
buf ( n392001 , n392000 );
buf ( n392002 , n392001 );
not ( n70994 , n392002 );
buf ( n392004 , n371272 );
not ( n392005 , n392004 );
and ( n392006 , n70994 , n392005 );
buf ( n392007 , n365676 );
not ( n392008 , n392007 );
buf ( n392009 , n362288 );
not ( n71001 , n392009 );
or ( n392011 , n392008 , n71001 );
buf ( n392012 , n42149 );
buf ( n392013 , n365673 );
nand ( n392014 , n392012 , n392013 );
buf ( n392015 , n392014 );
buf ( n392016 , n392015 );
nand ( n392017 , n392011 , n392016 );
buf ( n392018 , n392017 );
buf ( n392019 , n392018 );
buf ( n392020 , n45553 );
and ( n392021 , n392019 , n392020 );
nor ( n71013 , n392006 , n392021 );
buf ( n71014 , n71013 );
buf ( n392024 , n71014 );
not ( n392025 , n392024 );
not ( n71017 , n45075 );
not ( n392027 , n369217 );
or ( n71019 , n71017 , n392027 );
not ( n392029 , n342881 );
not ( n71021 , n47193 );
or ( n71022 , n392029 , n71021 );
buf ( n71023 , n367378 );
buf ( n71024 , n365202 );
nand ( n71025 , n71023 , n71024 );
buf ( n71026 , n71025 );
nand ( n392036 , n71022 , n71026 );
nand ( n71028 , n392036 , n365226 );
nand ( n392038 , n71019 , n71028 );
not ( n392039 , n392038 );
buf ( n392040 , n392039 );
not ( n71032 , n392040 );
or ( n392042 , n392025 , n71032 );
xor ( n71034 , n369243 , n369271 );
xor ( n392044 , n71034 , n369300 );
buf ( n392045 , n392044 );
buf ( n392046 , n392045 );
nand ( n392047 , n392042 , n392046 );
buf ( n392048 , n392047 );
buf ( n392049 , n392048 );
buf ( n392050 , n71014 );
not ( n392051 , n392050 );
buf ( n392052 , n392051 );
nand ( n392053 , n392038 , n392052 );
buf ( n392054 , n392053 );
nand ( n392055 , n392049 , n392054 );
buf ( n392056 , n392055 );
not ( n392057 , n342909 );
and ( n392058 , n359778 , n392057 );
not ( n71050 , n359778 );
and ( n392060 , n71050 , n387355 );
nor ( n392061 , n392058 , n392060 );
not ( n71053 , n392061 );
not ( n392063 , n71053 );
not ( n392064 , n45021 );
and ( n392065 , n392063 , n392064 );
and ( n392066 , n49269 , n365152 );
nor ( n71058 , n392065 , n392066 );
buf ( n392068 , n365167 );
not ( n71060 , n392068 );
buf ( n392070 , n368554 );
not ( n392071 , n392070 );
and ( n71063 , n71060 , n392071 );
buf ( n392073 , n40005 );
buf ( n392074 , n368554 );
and ( n392075 , n392073 , n392074 );
nor ( n71067 , n71063 , n392075 );
buf ( n392077 , n71067 );
not ( n71069 , n392077 );
not ( n392079 , n368614 );
and ( n392080 , n71069 , n392079 );
and ( n71072 , n369451 , n387542 );
nor ( n392082 , n392080 , n71072 );
nand ( n392083 , n71058 , n392082 );
not ( n71075 , n392083 );
not ( n392085 , n365115 );
not ( n71077 , n369732 );
or ( n392087 , n392085 , n71077 );
buf ( n71079 , n44819 );
not ( n71080 , n71079 );
buf ( n71081 , n368474 );
not ( n71082 , n71081 );
or ( n71083 , n71080 , n71082 );
buf ( n71084 , n364978 );
buf ( n71085 , n360885 );
nand ( n71086 , n71084 , n71085 );
buf ( n71087 , n71086 );
buf ( n71088 , n71087 );
nand ( n71089 , n71083 , n71088 );
buf ( n71090 , n71089 );
buf ( n392100 , n71090 );
buf ( n392101 , n365033 );
nand ( n392102 , n392100 , n392101 );
buf ( n392103 , n392102 );
nand ( n71095 , n392087 , n392103 );
not ( n392105 , n71095 );
not ( n71097 , n366402 );
not ( n392107 , n391490 );
or ( n71099 , n71097 , n392107 );
nand ( n71100 , n49634 , n366428 );
nand ( n392110 , n71099 , n71100 );
not ( n392111 , n392110 );
buf ( n392112 , n368290 );
not ( n392113 , n392112 );
buf ( n392114 , n365408 );
not ( n71106 , n392114 );
buf ( n392116 , n365507 );
not ( n392117 , n392116 );
or ( n392118 , n71106 , n392117 );
buf ( n392119 , n391855 );
nand ( n392120 , n392118 , n392119 );
buf ( n392121 , n392120 );
buf ( n392122 , n392121 );
not ( n392123 , n392122 );
or ( n392124 , n392113 , n392123 );
buf ( n392125 , n369399 );
buf ( n392126 , n39946 );
nand ( n392127 , n392125 , n392126 );
buf ( n392128 , n392127 );
buf ( n392129 , n392128 );
nand ( n392130 , n392124 , n392129 );
buf ( n392131 , n392130 );
buf ( n392132 , n392131 );
not ( n392133 , n392132 );
buf ( n392134 , n392133 );
nand ( n71126 , n392111 , n392134 );
buf ( n392136 , n71126 );
buf ( n392137 , n70869 );
not ( n71129 , n392137 );
buf ( n392139 , n45795 );
not ( n392140 , n392139 );
or ( n392141 , n71129 , n392140 );
nand ( n71133 , n362521 , n49182 );
buf ( n392143 , n71133 );
nand ( n71135 , n392141 , n392143 );
buf ( n392145 , n71135 );
buf ( n392146 , n392145 );
and ( n71138 , n392136 , n392146 );
and ( n71139 , n392131 , n392110 );
buf ( n392149 , n71139 );
nor ( n71141 , n71138 , n392149 );
buf ( n392151 , n71141 );
buf ( n392152 , n392151 );
not ( n71144 , n392152 );
buf ( n392154 , n71144 );
not ( n71146 , n392154 );
or ( n392156 , n392105 , n71146 );
not ( n392157 , n392151 );
not ( n71149 , n71095 );
not ( n392159 , n71149 );
or ( n392160 , n392157 , n392159 );
buf ( n392161 , n391315 );
not ( n71153 , n392161 );
buf ( n392163 , n45438 );
not ( n392164 , n392163 );
or ( n392165 , n71153 , n392164 );
buf ( n392166 , n41918 );
buf ( n392167 , n369624 );
nand ( n392168 , n392166 , n392167 );
buf ( n392169 , n392168 );
buf ( n71161 , n392169 );
nand ( n392171 , n392165 , n71161 );
buf ( n392172 , n392171 );
buf ( n392173 , n392172 );
not ( n392174 , n369857 );
not ( n392175 , n366751 );
or ( n392176 , n392174 , n392175 );
not ( n71168 , n391760 );
nand ( n71169 , n71168 , n377370 );
nand ( n392179 , n392176 , n71169 );
buf ( n392180 , n392179 );
xor ( n392181 , n392173 , n392180 );
buf ( n392182 , n391728 );
not ( n71174 , n392182 );
buf ( n392184 , n45204 );
not ( n392185 , n392184 );
or ( n71177 , n71174 , n392185 );
nand ( n71178 , n49217 , n46582 );
buf ( n392188 , n71178 );
nand ( n392189 , n71177 , n392188 );
buf ( n392190 , n392189 );
buf ( n392191 , n392190 );
and ( n392192 , n392181 , n392191 );
and ( n392193 , n392173 , n392180 );
or ( n71185 , n392192 , n392193 );
buf ( n392195 , n71185 );
nand ( n392196 , n392160 , n392195 );
nand ( n71188 , n392156 , n392196 );
not ( n71189 , n71188 );
or ( n392199 , n71075 , n71189 );
or ( n392200 , n71058 , n392082 );
nand ( n392201 , n392199 , n392200 );
xor ( n71193 , n392056 , n392201 );
xor ( n71194 , n48869 , n369074 );
xor ( n392204 , n71194 , n369103 );
buf ( n392205 , n392204 );
and ( n392206 , n71193 , n392205 );
and ( n392207 , n392056 , n392201 );
or ( n71199 , n392206 , n392207 );
xor ( n392209 , n49108 , n369312 );
xor ( n392210 , n392209 , n369439 );
xor ( n71202 , n71199 , n392210 );
buf ( n392212 , n49114 );
buf ( n392213 , n369437 );
xor ( n392214 , n392212 , n392213 );
buf ( n392215 , n369432 );
xor ( n71207 , n392214 , n392215 );
buf ( n392217 , n71207 );
not ( n392218 , n392217 );
buf ( n392219 , n369642 );
buf ( n392220 , n49250 );
xor ( n392221 , n392219 , n392220 );
buf ( n392222 , n369477 );
xor ( n71214 , n392221 , n392222 );
buf ( n392224 , n71214 );
buf ( n392225 , n392224 );
buf ( n392226 , n49021 );
buf ( n392227 , n49000 );
xor ( n71219 , n392226 , n392227 );
buf ( n392229 , n71219 );
buf ( n392230 , n392229 );
buf ( n392231 , n369304 );
and ( n71223 , n392230 , n392231 );
not ( n71224 , n392230 );
buf ( n392234 , n369307 );
and ( n392235 , n71224 , n392234 );
nor ( n71227 , n71223 , n392235 );
buf ( n71228 , n71227 );
buf ( n392238 , n71228 );
not ( n71230 , n392238 );
buf ( n392240 , n71230 );
buf ( n392241 , n392240 );
nand ( n392242 , n392225 , n392241 );
buf ( n392243 , n392242 );
not ( n392244 , n392243 );
or ( n392245 , n392218 , n392244 );
buf ( n392246 , n392224 );
not ( n71238 , n392246 );
buf ( n392248 , n71238 );
buf ( n392249 , n392248 );
buf ( n71241 , n71228 );
nand ( n71242 , n392249 , n71241 );
buf ( n392252 , n71242 );
nand ( n71244 , n392245 , n392252 );
and ( n392254 , n71202 , n71244 );
and ( n392255 , n71199 , n392210 );
or ( n71247 , n392254 , n392255 );
buf ( n392257 , n71247 );
not ( n392258 , n392257 );
buf ( n392259 , n392258 );
not ( n71251 , n392259 );
or ( n392261 , n70989 , n71251 );
not ( n392262 , n369648 );
not ( n71254 , n392262 );
not ( n392264 , n369666 );
or ( n392265 , n71254 , n392264 );
nand ( n71257 , n369651 , n369648 );
nand ( n71258 , n392265 , n71257 );
xor ( n392268 , n49455 , n369045 );
and ( n392269 , n71258 , n392268 );
not ( n71261 , n71258 );
not ( n392271 , n392268 );
and ( n392272 , n71261 , n392271 );
nor ( n71264 , n392269 , n392272 );
buf ( n71265 , n71264 );
not ( n392275 , n71265 );
xor ( n392276 , n369708 , n370083 );
xor ( n392277 , n392276 , n370100 );
not ( n71269 , n392277 );
or ( n71270 , n392275 , n71269 );
or ( n392280 , n392277 , n71265 );
not ( n392281 , n49437 );
nand ( n71273 , n369540 , n49362 , n392281 );
nand ( n71274 , n49437 , n49362 , n49364 );
nand ( n71275 , n49364 , n392281 , n369561 );
nand ( n392285 , n369540 , n369561 , n49437 );
nand ( n392286 , n71273 , n71274 , n71275 , n392285 );
not ( n71278 , n392286 );
not ( n392288 , n71278 );
not ( n392289 , n392288 );
not ( n71281 , n369199 );
not ( n392291 , n44915 );
or ( n392292 , n71281 , n392291 );
buf ( n392293 , n39830 );
not ( n71285 , n392293 );
buf ( n392295 , n365052 );
not ( n392296 , n392295 );
and ( n392297 , n71285 , n392296 );
buf ( n392298 , n371416 );
buf ( n392299 , n365052 );
and ( n392300 , n392298 , n392299 );
nor ( n71292 , n392297 , n392300 );
buf ( n392302 , n71292 );
not ( n392303 , n392302 );
nand ( n71295 , n392303 , n47466 );
nand ( n71296 , n392292 , n71295 );
not ( n392306 , n71296 );
or ( n392307 , n392289 , n392306 );
not ( n392308 , n71278 );
not ( n71300 , n71296 );
not ( n71301 , n71300 );
or ( n392311 , n392308 , n71301 );
xor ( n392312 , n49132 , n369366 );
xor ( n392313 , n392312 , n369429 );
nand ( n71305 , n392311 , n392313 );
nand ( n71306 , n392307 , n71305 );
buf ( n392316 , n71306 );
buf ( n392317 , n392316 );
buf ( n392318 , n392317 );
not ( n392319 , n392318 );
xor ( n392320 , n369756 , n369759 );
xor ( n71312 , n392320 , n370079 );
buf ( n392322 , n71312 );
not ( n392323 , n392322 );
or ( n71315 , n392319 , n392323 );
buf ( n392325 , n392322 );
buf ( n392326 , n392318 );
or ( n392327 , n392325 , n392326 );
xor ( n392328 , n369385 , n369409 );
xor ( n71320 , n392328 , n49223 );
buf ( n392330 , n71320 );
not ( n71322 , n392330 );
buf ( n392332 , n369599 );
not ( n392333 , n392332 );
buf ( n392334 , n392333 );
xor ( n71326 , n369607 , n392334 );
xor ( n392336 , n71326 , n369636 );
buf ( n392337 , n392336 );
nand ( n71329 , n369496 , n49306 );
xor ( n71330 , n49335 , n71329 );
xnor ( n392340 , n71330 , n369532 );
buf ( n392341 , n392340 );
nand ( n71333 , n392337 , n392341 );
buf ( n71334 , n71333 );
buf ( n392344 , n71334 );
not ( n392345 , n392344 );
or ( n71337 , n71322 , n392345 );
buf ( n392347 , n392336 );
not ( n392348 , n392347 );
buf ( n392349 , n392348 );
not ( n71341 , n392340 );
nand ( n392351 , n392349 , n71341 );
buf ( n392352 , n392351 );
nand ( n71344 , n71337 , n392352 );
buf ( n392354 , n71344 );
buf ( n392355 , n392354 );
buf ( n392356 , n45492 );
not ( n392357 , n392356 );
buf ( n392358 , n392018 );
not ( n71350 , n392358 );
or ( n71351 , n392357 , n71350 );
buf ( n392361 , n365676 );
not ( n392362 , n392361 );
buf ( n392363 , n362145 );
not ( n71355 , n392363 );
or ( n71356 , n392362 , n71355 );
buf ( n392366 , n370782 );
buf ( n71358 , n365673 );
nand ( n71359 , n392366 , n71358 );
buf ( n392369 , n71359 );
buf ( n392370 , n392369 );
nand ( n71362 , n71356 , n392370 );
buf ( n392372 , n71362 );
buf ( n392373 , n392372 );
buf ( n392374 , n45553 );
nand ( n71366 , n392373 , n392374 );
buf ( n71367 , n71366 );
buf ( n392377 , n71367 );
nand ( n392378 , n71351 , n392377 );
buf ( n392379 , n392378 );
buf ( n392380 , n392379 );
not ( n392381 , n45075 );
not ( n71373 , n392036 );
or ( n392383 , n392381 , n71373 );
and ( n392384 , n40251 , n45065 );
not ( n71376 , n40251 );
and ( n71377 , n71376 , n45060 );
or ( n392387 , n392384 , n71377 );
buf ( n392388 , n392387 );
buf ( n392389 , n45058 );
nand ( n71381 , n392388 , n392389 );
buf ( n392391 , n71381 );
nand ( n392392 , n392383 , n392391 );
buf ( n392393 , n392392 );
xor ( n392394 , n392380 , n392393 );
xor ( n392395 , n369845 , n369870 );
xor ( n71387 , n392395 , n369936 );
buf ( n392397 , n71387 );
buf ( n392398 , n392397 );
and ( n71390 , n392394 , n392398 );
and ( n71391 , n392380 , n392393 );
or ( n392401 , n71390 , n71391 );
buf ( n392402 , n392401 );
buf ( n392403 , n392402 );
xor ( n71395 , n392355 , n392403 );
buf ( n392405 , n368549 );
not ( n392406 , n392405 );
buf ( n392407 , n372458 );
not ( n392408 , n392407 );
or ( n392409 , n392406 , n392408 );
buf ( n392410 , n39867 );
buf ( n392411 , n368554 );
nand ( n392412 , n392410 , n392411 );
buf ( n392413 , n392412 );
buf ( n392414 , n392413 );
nand ( n71406 , n392409 , n392414 );
buf ( n392416 , n71406 );
not ( n392417 , n392416 );
not ( n392418 , n368611 );
or ( n71410 , n392417 , n392418 );
not ( n392420 , n392077 );
nand ( n392421 , n392420 , n387542 );
nand ( n71413 , n71410 , n392421 );
not ( n392423 , n365152 );
not ( n392424 , n392061 );
or ( n71416 , n392423 , n392424 );
buf ( n392426 , n40199 );
buf ( n392427 , n46397 );
and ( n392428 , n392426 , n392427 );
not ( n392429 , n392426 );
buf ( n392430 , n342909 );
and ( n71422 , n392429 , n392430 );
or ( n392432 , n392428 , n71422 );
buf ( n392433 , n392432 );
buf ( n392434 , n392433 );
not ( n71426 , n392434 );
buf ( n392436 , n390954 );
nand ( n392437 , n71426 , n392436 );
buf ( n392438 , n392437 );
nand ( n392439 , n71416 , n392438 );
or ( n392440 , n71413 , n392439 );
or ( n392441 , n363291 , n391280 );
or ( n392442 , n369954 , n365801 );
nand ( n71434 , n392441 , n392442 );
not ( n392444 , n71434 );
not ( n392445 , n70286 );
nand ( n71437 , n41835 , n70287 );
nand ( n71438 , n391318 , n71437 , n391319 , n70292 );
not ( n392448 , n71438 );
or ( n392449 , n392445 , n392448 );
not ( n71441 , n70312 );
nand ( n392451 , n71441 , n391301 );
nand ( n392452 , n392449 , n392451 );
not ( n71444 , n392452 );
or ( n392454 , n392444 , n71444 );
or ( n392455 , n392452 , n71434 );
xor ( n71447 , n369890 , n369902 );
xor ( n392457 , n71447 , n369931 );
buf ( n392458 , n392457 );
nand ( n71450 , n392455 , n392458 );
nand ( n71451 , n392454 , n71450 );
nand ( n392461 , n392440 , n71451 );
buf ( n392462 , n392461 );
buf ( n392463 , n392439 );
buf ( n392464 , n71413 );
nand ( n71456 , n392463 , n392464 );
buf ( n71457 , n71456 );
buf ( n392467 , n71457 );
nand ( n71459 , n392462 , n392467 );
buf ( n392469 , n71459 );
buf ( n71461 , n392469 );
and ( n71462 , n71395 , n71461 );
and ( n71463 , n392355 , n392403 );
or ( n71464 , n71462 , n71463 );
buf ( n71465 , n71464 );
buf ( n392475 , n71465 );
nand ( n71467 , n392327 , n392475 );
buf ( n392477 , n71467 );
nand ( n71469 , n71315 , n392477 );
nand ( n392479 , n392280 , n71469 );
nand ( n392480 , n71270 , n392479 );
nand ( n392481 , n392261 , n392480 );
buf ( n392482 , n391997 );
not ( n392483 , n392482 );
buf ( n392484 , n71247 );
nand ( n71476 , n392483 , n392484 );
buf ( n392486 , n71476 );
and ( n392487 , n392481 , n392486 );
not ( n392488 , n392487 );
and ( n392489 , n391991 , n392488 );
and ( n71481 , n48977 , n369680 );
not ( n392491 , n48977 );
and ( n392492 , n392491 , n370114 );
nor ( n71484 , n71481 , n392492 );
buf ( n392494 , n370110 );
not ( n392495 , n392494 );
buf ( n392496 , n392495 );
and ( n71488 , n71484 , n392496 );
not ( n392498 , n71484 );
buf ( n392499 , n370110 );
and ( n392500 , n392498 , n392499 );
nor ( n71492 , n71488 , n392500 );
not ( n71493 , n71492 );
or ( n392503 , n392489 , n71493 );
nand ( n71495 , n391990 , n392487 );
nand ( n71496 , n392503 , n71495 );
nand ( n71497 , n70979 , n71496 );
buf ( n392507 , n71306 );
buf ( n392508 , n71465 );
xor ( n71500 , n392507 , n392508 );
buf ( n392510 , n392322 );
xnor ( n71502 , n71500 , n392510 );
buf ( n392512 , n71502 );
buf ( n392513 , n392512 );
not ( n392514 , n392513 );
buf ( n392515 , n392514 );
not ( n392516 , n392082 );
not ( n71508 , n71058 );
or ( n392518 , n392516 , n71508 );
nand ( n392519 , n392518 , n392200 );
buf ( n392520 , n392519 );
buf ( n392521 , n71188 );
buf ( n392522 , n392521 );
buf ( n392523 , n392522 );
buf ( n392524 , n392523 );
xnor ( n392525 , n392520 , n392524 );
buf ( n392526 , n392525 );
buf ( n392527 , n392526 );
not ( n71519 , n392527 );
or ( n71520 , n57530 , n377580 );
and ( n392530 , n391342 , n71520 );
buf ( n392531 , n392530 );
not ( n71523 , n392531 );
buf ( n392533 , n392433 );
not ( n392534 , n392533 );
buf ( n392535 , n365155 );
not ( n392536 , n392535 );
and ( n392537 , n392534 , n392536 );
buf ( n392538 , n391660 );
not ( n392539 , n365190 );
buf ( n71531 , n392539 );
and ( n71532 , n392538 , n71531 );
nor ( n71533 , n392537 , n71532 );
buf ( n71534 , n71533 );
buf ( n392544 , n71534 );
not ( n392545 , n392544 );
or ( n71537 , n71523 , n392545 );
buf ( n392547 , n365033 );
not ( n392548 , n392547 );
buf ( n392549 , n391802 );
not ( n71541 , n392549 );
or ( n71542 , n392548 , n71541 );
buf ( n392552 , n71090 );
buf ( n392553 , n365115 );
nand ( n71545 , n392552 , n392553 );
buf ( n392555 , n71545 );
buf ( n392556 , n392555 );
nand ( n392557 , n71542 , n392556 );
buf ( n392558 , n392557 );
buf ( n392559 , n392558 );
nand ( n392560 , n71537 , n392559 );
buf ( n392561 , n392560 );
buf ( n392562 , n71534 );
not ( n392563 , n392562 );
buf ( n392564 , n392530 );
not ( n71556 , n392564 );
buf ( n71557 , n71556 );
buf ( n392567 , n71557 );
nand ( n392568 , n392563 , n392567 );
buf ( n392569 , n392568 );
nand ( n71561 , n392561 , n392569 );
not ( n392571 , n71561 );
not ( n392572 , n392571 );
xor ( n71564 , n71095 , n392154 );
xor ( n392574 , n71564 , n392195 );
not ( n392575 , n392574 );
not ( n71567 , n392575 );
and ( n71568 , n392572 , n71567 );
xor ( n71569 , n392110 , n392134 );
xnor ( n392579 , n71569 , n392145 );
buf ( n392580 , n392579 );
not ( n71572 , n392580 );
buf ( n392582 , n71572 );
buf ( n392583 , n392582 );
not ( n392584 , n392583 );
buf ( n392585 , n391525 );
not ( n392586 , n392585 );
buf ( n392587 , n392586 );
buf ( n392588 , n392587 );
not ( n392589 , n392588 );
buf ( n392590 , n365227 );
not ( n71582 , n392590 );
and ( n71583 , n392589 , n71582 );
buf ( n392593 , n392387 );
buf ( n392594 , n45075 );
and ( n392595 , n392593 , n392594 );
nor ( n71587 , n71583 , n392595 );
buf ( n392597 , n71587 );
buf ( n392598 , n392597 );
not ( n71590 , n392598 );
or ( n392600 , n392584 , n71590 );
xor ( n392601 , n392173 , n392180 );
xor ( n71593 , n392601 , n392191 );
buf ( n392603 , n71593 );
buf ( n392604 , n392603 );
nand ( n71596 , n392600 , n392604 );
buf ( n392606 , n71596 );
not ( n392607 , n392597 );
nand ( n392608 , n392607 , n392579 );
nand ( n392609 , n392606 , n392608 );
nand ( n71601 , n392575 , n392571 );
and ( n392611 , n392609 , n71601 );
nor ( n392612 , n71568 , n392611 );
buf ( n392613 , n392612 );
buf ( n71605 , n392613 );
buf ( n71606 , n71605 );
buf ( n392616 , n71606 );
nand ( n71608 , n71519 , n392616 );
buf ( n392618 , n71608 );
buf ( n392619 , n392618 );
not ( n392620 , n392619 );
xor ( n392621 , n392380 , n392393 );
xor ( n71613 , n392621 , n392398 );
buf ( n392623 , n71613 );
not ( n392624 , n392623 );
not ( n71616 , n49609 );
and ( n71617 , n40090 , n369766 );
not ( n392627 , n40090 );
and ( n392628 , n392627 , n369769 );
or ( n392629 , n71617 , n392628 );
not ( n392630 , n392629 );
or ( n71622 , n71616 , n392630 );
buf ( n392632 , n391686 );
buf ( n392633 , n369804 );
nand ( n71625 , n392632 , n392633 );
buf ( n392635 , n71625 );
nand ( n392636 , n71622 , n392635 );
buf ( n392637 , n392636 );
not ( n71629 , n392637 );
not ( n392639 , n368611 );
not ( n392640 , n391353 );
or ( n71632 , n392639 , n392640 );
not ( n392642 , n368624 );
nand ( n392643 , n392642 , n392416 );
nand ( n71635 , n71632 , n392643 );
not ( n71636 , n71635 );
buf ( n392646 , n71636 );
nand ( n392647 , n71629 , n392646 );
buf ( n392648 , n392647 );
buf ( n392649 , n392648 );
not ( n392650 , n391542 );
not ( n71642 , n70537 );
or ( n71643 , n392650 , n71642 );
not ( n71644 , n70519 );
not ( n392654 , n391546 );
or ( n392655 , n71644 , n392654 );
nand ( n71647 , n392655 , n70556 );
nand ( n71648 , n71643 , n71647 );
buf ( n392658 , n71648 );
and ( n71650 , n392649 , n392658 );
not ( n392660 , n71635 );
not ( n392661 , n392636 );
nor ( n71653 , n392660 , n392661 );
buf ( n392663 , n71653 );
nor ( n392664 , n71650 , n392663 );
buf ( n392665 , n392664 );
nand ( n392666 , n392624 , n392665 );
not ( n392667 , n392666 );
nand ( n71659 , n70276 , n70279 );
not ( n71660 , n71659 );
not ( n392670 , n70313 );
or ( n392671 , n71660 , n392670 );
nand ( n71663 , n70275 , n391272 );
nand ( n392673 , n392671 , n71663 );
not ( n392674 , n44915 );
and ( n71666 , n365052 , n40999 );
not ( n392676 , n365052 );
and ( n71668 , n392676 , n359756 );
or ( n71669 , n71666 , n71668 );
buf ( n392679 , n71669 );
not ( n71671 , n392679 );
buf ( n392681 , n71671 );
not ( n71673 , n392681 );
or ( n71674 , n392674 , n71673 );
nand ( n71675 , n391242 , n47466 );
nand ( n71676 , n71674 , n71675 );
xor ( n71677 , n392673 , n71676 );
not ( n392687 , n71434 );
not ( n392688 , n392687 );
not ( n71680 , n392452 );
or ( n71681 , n392688 , n71680 );
not ( n71682 , n392452 );
nand ( n71683 , n71682 , n71434 );
nand ( n392693 , n71681 , n71683 );
and ( n392694 , n392693 , n392458 );
not ( n392695 , n392693 );
not ( n392696 , n392458 );
and ( n71688 , n392695 , n392696 );
nor ( n392698 , n392694 , n71688 );
and ( n392699 , n71677 , n392698 );
and ( n71691 , n392673 , n71676 );
or ( n71692 , n392699 , n71691 );
not ( n392702 , n71692 );
or ( n392703 , n392667 , n392702 );
buf ( n392704 , n392665 );
not ( n71696 , n392704 );
buf ( n392706 , n71696 );
nand ( n392707 , n392706 , n392623 );
nand ( n392708 , n392703 , n392707 );
buf ( n392709 , n392708 );
not ( n392710 , n392709 );
or ( n392711 , n392620 , n392710 );
buf ( n392712 , n71606 );
not ( n71704 , n392712 );
buf ( n392714 , n392526 );
nand ( n71706 , n71704 , n392714 );
buf ( n392716 , n71706 );
buf ( n392717 , n392716 );
nand ( n71709 , n392711 , n392717 );
buf ( n392719 , n71709 );
buf ( n392720 , n392719 );
buf ( n392721 , n71228 );
buf ( n392722 , n392248 );
xor ( n392723 , n392721 , n392722 );
buf ( n392724 , n392217 );
xnor ( n71716 , n392723 , n392724 );
buf ( n392726 , n71716 );
buf ( n392727 , n392726 );
and ( n392728 , n392720 , n392727 );
not ( n71720 , n392720 );
buf ( n392730 , n392726 );
not ( n392731 , n392730 );
buf ( n392732 , n392731 );
buf ( n392733 , n392732 );
and ( n71725 , n71720 , n392733 );
nor ( n71726 , n392728 , n71725 );
buf ( n392736 , n71726 );
xnor ( n71728 , n392515 , n392736 );
xor ( n71729 , n369820 , n369941 );
xor ( n71730 , n71729 , n370074 );
buf ( n392740 , n71730 );
buf ( n392741 , n392740 );
xor ( n71733 , n370066 , n369990 );
xnor ( n71734 , n71733 , n369964 );
buf ( n71735 , n71734 );
and ( n71736 , n370041 , n49828 );
not ( n71737 , n370041 );
and ( n392747 , n71737 , n370034 );
nor ( n71739 , n71736 , n392747 );
not ( n71740 , n71739 );
not ( n71741 , n71740 );
not ( n392751 , n370050 );
not ( n392752 , n370053 );
and ( n71744 , n392751 , n392752 );
nor ( n392754 , n370059 , n370060 );
nor ( n392755 , n71744 , n392754 );
not ( n71747 , n392755 );
not ( n71748 , n71747 );
or ( n392758 , n71741 , n71748 );
nand ( n392759 , n71739 , n392755 );
nand ( n392760 , n392758 , n392759 );
not ( n71752 , n392760 );
buf ( n392762 , n366654 );
not ( n392763 , n392762 );
buf ( n392764 , n49776 );
not ( n71756 , n392764 );
or ( n392766 , n392763 , n71756 );
buf ( n71758 , n391842 );
buf ( n392768 , n46521 );
nand ( n392769 , n71758 , n392768 );
buf ( n392770 , n392769 );
buf ( n71762 , n392770 );
nand ( n392772 , n392766 , n71762 );
buf ( n392773 , n392772 );
not ( n71765 , n392773 );
not ( n392775 , n71765 );
and ( n392776 , n71752 , n392775 );
nand ( n392777 , n392760 , n71765 );
buf ( n392778 , n391497 );
not ( n392779 , n392778 );
buf ( n392780 , n370034 );
nand ( n71772 , n392779 , n392780 );
buf ( n392782 , n71772 );
buf ( n392783 , n392782 );
buf ( n392784 , n391478 );
and ( n392785 , n392783 , n392784 );
buf ( n392786 , n391497 );
buf ( n392787 , n49828 );
and ( n71779 , n392786 , n392787 );
buf ( n392789 , n71779 );
buf ( n392790 , n392789 );
nor ( n71782 , n392785 , n392790 );
buf ( n392792 , n71782 );
buf ( n392793 , n392792 );
not ( n392794 , n392793 );
buf ( n392795 , n392794 );
and ( n392796 , n392777 , n392795 );
nor ( n392797 , n392776 , n392796 );
buf ( n392798 , n392797 );
nand ( n71790 , n71735 , n392798 );
buf ( n71791 , n71790 );
not ( n392801 , n71791 );
not ( n71793 , n71320 );
not ( n71794 , n71793 );
buf ( n392804 , n392340 );
not ( n71796 , n392804 );
buf ( n392806 , n392349 );
not ( n71798 , n392806 );
or ( n71799 , n71796 , n71798 );
nand ( n71800 , n71341 , n392336 );
buf ( n392810 , n71800 );
nand ( n392811 , n71799 , n392810 );
buf ( n392812 , n392811 );
not ( n392813 , n392812 );
or ( n392814 , n71794 , n392813 );
or ( n71806 , n392812 , n71793 );
nand ( n392816 , n392814 , n71806 );
not ( n392817 , n392816 );
or ( n71809 , n392801 , n392817 );
buf ( n392819 , n71734 );
not ( n392820 , n392819 );
buf ( n392821 , n392797 );
not ( n392822 , n392821 );
buf ( n392823 , n392822 );
buf ( n392824 , n392823 );
nand ( n71816 , n392820 , n392824 );
buf ( n392826 , n71816 );
nand ( n71818 , n71809 , n392826 );
buf ( n392828 , n71818 );
xor ( n71820 , n392741 , n392828 );
xor ( n392830 , n392286 , n71296 );
xor ( n392831 , n392830 , n392313 );
buf ( n392832 , n392831 );
xor ( n392833 , n71820 , n392832 );
buf ( n392834 , n392833 );
not ( n71826 , n392834 );
not ( n71827 , n392612 );
not ( n392837 , n392526 );
not ( n392838 , n392837 );
or ( n392839 , n71827 , n392838 );
not ( n392840 , n392612 );
nand ( n392841 , n392840 , n392526 );
nand ( n71833 , n392839 , n392841 );
and ( n392843 , n71833 , n392708 );
not ( n392844 , n71833 );
not ( n71836 , n392708 );
and ( n71837 , n392844 , n71836 );
nor ( n392847 , n392843 , n71837 );
not ( n392848 , n392847 );
not ( n71840 , n392848 );
or ( n392850 , n71826 , n71840 );
buf ( n392851 , n392834 );
not ( n71843 , n392851 );
buf ( n392853 , n71843 );
buf ( n392854 , n392853 );
not ( n392855 , n392854 );
buf ( n392856 , n392847 );
not ( n392857 , n392856 );
or ( n71849 , n392855 , n392857 );
not ( n71850 , n392609 );
not ( n71851 , n392571 );
and ( n392861 , n71850 , n71851 );
and ( n71853 , n392609 , n392571 );
nor ( n71854 , n392861 , n71853 );
buf ( n392864 , n392574 );
buf ( n392865 , n392864 );
buf ( n392866 , n392865 );
and ( n71858 , n71854 , n392866 );
not ( n71859 , n71854 );
buf ( n392869 , n392866 );
not ( n392870 , n392869 );
buf ( n392871 , n392870 );
and ( n71863 , n71859 , n392871 );
nor ( n392873 , n71858 , n71863 );
buf ( n392874 , n392873 );
buf ( n392875 , n392629 );
buf ( n392876 , n369804 );
and ( n392877 , n392875 , n392876 );
buf ( n392878 , n369777 );
not ( n392879 , n392878 );
buf ( n392880 , n369813 );
nor ( n392881 , n392879 , n392880 );
buf ( n392882 , n392881 );
buf ( n392883 , n392882 );
nor ( n71875 , n392877 , n392883 );
buf ( n71876 , n71875 );
buf ( n392886 , n71876 );
not ( n392887 , n392886 );
buf ( n392888 , n392887 );
buf ( n392889 , n45492 );
not ( n392890 , n392889 );
buf ( n392891 , n392372 );
not ( n71883 , n392891 );
or ( n71884 , n392890 , n71883 );
buf ( n392894 , n391436 );
buf ( n392895 , n45553 );
nand ( n392896 , n392894 , n392895 );
buf ( n392897 , n392896 );
buf ( n71889 , n392897 );
nand ( n392899 , n71884 , n71889 );
buf ( n392900 , n392899 );
buf ( n392901 , n392900 );
not ( n392902 , n392901 );
buf ( n71894 , n70836 );
not ( n71895 , n71894 );
not ( n71896 , n71895 );
not ( n392906 , n391859 );
or ( n71898 , n71896 , n392906 );
not ( n71899 , n70852 );
not ( n71900 , n71894 );
or ( n392910 , n71899 , n71900 );
nand ( n392911 , n392910 , n391881 );
nand ( n71903 , n71898 , n392911 );
buf ( n392913 , n71903 );
not ( n71905 , n392913 );
or ( n392915 , n392902 , n71905 );
or ( n71907 , n71903 , n392900 );
not ( n71908 , n70768 );
not ( n71909 , n391744 );
or ( n71910 , n71908 , n71909 );
not ( n71911 , n70759 );
not ( n392921 , n391773 );
or ( n71913 , n71911 , n392921 );
nand ( n392923 , n71913 , n391734 );
nand ( n392924 , n71910 , n392923 );
nand ( n71916 , n71907 , n392924 );
buf ( n71917 , n71916 );
nand ( n392927 , n392915 , n71917 );
buf ( n392928 , n392927 );
xor ( n71920 , n392888 , n392928 );
not ( n392930 , n71669 );
not ( n392931 , n44913 );
and ( n392932 , n392930 , n392931 );
buf ( n392933 , n392302 );
buf ( n392934 , n365083 );
nor ( n392935 , n392933 , n392934 );
buf ( n392936 , n392935 );
nor ( n71928 , n392932 , n392936 );
and ( n392938 , n71920 , n71928 );
not ( n392939 , n71920 );
buf ( n392940 , n71928 );
not ( n71932 , n392940 );
buf ( n392942 , n71932 );
and ( n392943 , n392939 , n392942 );
nor ( n71935 , n392938 , n392943 );
buf ( n392945 , n71935 );
nand ( n392946 , n392874 , n392945 );
buf ( n392947 , n392946 );
buf ( n392948 , n392947 );
not ( n392949 , n71903 );
not ( n71941 , n392949 );
and ( n71942 , n392924 , n392900 );
not ( n392952 , n392924 );
not ( n392953 , n392900 );
and ( n392954 , n392952 , n392953 );
nor ( n71946 , n71942 , n392954 );
not ( n392956 , n71946 );
or ( n392957 , n71941 , n392956 );
or ( n71949 , n71946 , n392949 );
nand ( n71950 , n392957 , n71949 );
buf ( n392960 , n71950 );
xor ( n392961 , n391651 , n391668 );
and ( n392962 , n392961 , n391696 );
and ( n392963 , n391651 , n391668 );
or ( n71955 , n392962 , n392963 );
buf ( n392965 , n71955 );
buf ( n392966 , n392965 );
xor ( n71958 , n392960 , n392966 );
xor ( n71959 , n392597 , n392603 );
xnor ( n392969 , n71959 , n392579 );
buf ( n392970 , n392969 );
and ( n71962 , n71958 , n392970 );
and ( n392972 , n392960 , n392966 );
or ( n392973 , n71962 , n392972 );
buf ( n392974 , n392973 );
buf ( n392975 , n392974 );
and ( n392976 , n392948 , n392975 );
buf ( n392977 , n392873 );
buf ( n392978 , n71935 );
nor ( n71970 , n392977 , n392978 );
buf ( n71971 , n71970 );
buf ( n392981 , n71971 );
nor ( n71973 , n392976 , n392981 );
buf ( n392983 , n71973 );
buf ( n392984 , n392983 );
not ( n71976 , n392984 );
buf ( n392986 , n71976 );
buf ( n392987 , n392986 );
nand ( n71979 , n71849 , n392987 );
buf ( n392989 , n71979 );
nand ( n392990 , n392850 , n392989 );
xor ( n392991 , n392355 , n392403 );
xor ( n392992 , n392991 , n71461 );
buf ( n392993 , n392992 );
not ( n392994 , n392993 );
not ( n392995 , n392994 );
not ( n71987 , n392995 );
not ( n71988 , n392052 );
not ( n392998 , n392039 );
or ( n71990 , n71988 , n392998 );
nand ( n71991 , n71014 , n392038 );
nand ( n71992 , n71990 , n71991 );
xor ( n393002 , n392045 , n71992 );
not ( n71994 , n393002 );
not ( n393004 , n71994 );
xor ( n71996 , n369753 , n369744 );
xnor ( n71997 , n71996 , n49510 );
buf ( n393007 , n71997 );
not ( n393008 , n393007 );
buf ( n393009 , n393008 );
not ( n393010 , n393009 );
or ( n393011 , n393004 , n393010 );
buf ( n393012 , n393002 );
buf ( n393013 , n71997 );
nand ( n393014 , n393012 , n393013 );
buf ( n393015 , n393014 );
nand ( n393016 , n393011 , n393015 );
buf ( n393017 , n71876 );
not ( n72009 , n393017 );
buf ( n393019 , n71928 );
not ( n72011 , n393019 );
or ( n72012 , n72009 , n72011 );
buf ( n393022 , n392928 );
nand ( n72014 , n72012 , n393022 );
buf ( n393024 , n72014 );
buf ( n393025 , n393024 );
buf ( n393026 , n392888 );
buf ( n393027 , n392942 );
nand ( n72019 , n393026 , n393027 );
buf ( n393029 , n72019 );
buf ( n393030 , n393029 );
nand ( n72022 , n393025 , n393030 );
buf ( n393032 , n72022 );
buf ( n393033 , n393032 );
not ( n393034 , n393033 );
buf ( n393035 , n393034 );
and ( n393036 , n393016 , n393035 );
not ( n393037 , n393016 );
and ( n72029 , n393037 , n393032 );
nor ( n393039 , n393036 , n72029 );
not ( n393040 , n393039 );
not ( n72032 , n393040 );
or ( n72033 , n71987 , n72032 );
not ( n393043 , n392994 );
not ( n393044 , n393039 );
or ( n393045 , n393043 , n393044 );
buf ( n393046 , n391441 );
not ( n393047 , n393046 );
buf ( n393048 , n393047 );
buf ( n393049 , n393048 );
not ( n72041 , n393049 );
buf ( n393051 , n391500 );
not ( n393052 , n393051 );
or ( n72044 , n72041 , n393052 );
buf ( n393054 , n391462 );
nand ( n72046 , n72044 , n393054 );
buf ( n393056 , n72046 );
buf ( n393057 , n393056 );
buf ( n393058 , n391500 );
not ( n72050 , n393058 );
buf ( n393060 , n391441 );
nand ( n393061 , n72050 , n393060 );
buf ( n393062 , n393061 );
buf ( n393063 , n393062 );
nand ( n393064 , n393057 , n393063 );
buf ( n393065 , n393064 );
buf ( n393066 , n393065 );
buf ( n72058 , n392760 );
not ( n72059 , n72058 );
xnor ( n72060 , n392792 , n392773 );
not ( n72061 , n72060 );
or ( n72062 , n72059 , n72061 );
or ( n72063 , n72060 , n72058 );
nand ( n393073 , n72062 , n72063 );
buf ( n393074 , n393073 );
xor ( n72066 , n393066 , n393074 );
buf ( n393076 , n391812 );
not ( n393077 , n393076 );
buf ( n393078 , n391888 );
not ( n72070 , n393078 );
or ( n72071 , n393077 , n72070 );
buf ( n393081 , n391815 );
not ( n72073 , n393081 );
buf ( n393083 , n70874 );
not ( n393084 , n393083 );
or ( n72076 , n72073 , n393084 );
buf ( n393086 , n391786 );
nand ( n72078 , n72076 , n393086 );
buf ( n393088 , n72078 );
buf ( n393089 , n393088 );
nand ( n72081 , n72071 , n393089 );
buf ( n393091 , n72081 );
buf ( n393092 , n393091 );
and ( n72084 , n72066 , n393092 );
and ( n393094 , n393066 , n393074 );
or ( n72086 , n72084 , n393094 );
buf ( n393096 , n72086 );
xor ( n72088 , n392439 , n71413 );
xnor ( n72089 , n72088 , n71451 );
not ( n72090 , n72089 );
nor ( n72091 , n393096 , n72090 );
not ( n393101 , n392816 );
not ( n72093 , n393101 );
not ( n72094 , n72093 );
not ( n72095 , n392797 );
not ( n72096 , n71734 );
not ( n72097 , n72096 );
or ( n72098 , n72095 , n72097 );
nand ( n72099 , n71734 , n392823 );
nand ( n72100 , n72098 , n72099 );
not ( n72101 , n72100 );
or ( n72102 , n72094 , n72101 );
or ( n72103 , n72093 , n72100 );
nand ( n72104 , n72102 , n72103 );
or ( n72105 , n72091 , n72104 );
nand ( n72106 , n393096 , n72090 );
nand ( n72107 , n72105 , n72106 );
nand ( n72108 , n393045 , n72107 );
nand ( n72109 , n72033 , n72108 );
not ( n72110 , n72109 );
xor ( n72111 , n392056 , n392201 );
xor ( n72112 , n72111 , n392205 );
buf ( n393122 , n72112 );
buf ( n393123 , n393009 );
not ( n72115 , n393123 );
not ( n393125 , n393002 );
not ( n393126 , n393125 );
buf ( n393127 , n393126 );
not ( n393128 , n393127 );
or ( n72120 , n72115 , n393128 );
buf ( n393130 , n393125 );
not ( n72122 , n393130 );
buf ( n393132 , n71997 );
not ( n393133 , n393132 );
or ( n393134 , n72122 , n393133 );
buf ( n393135 , n393032 );
nand ( n393136 , n393134 , n393135 );
buf ( n393137 , n393136 );
buf ( n393138 , n393137 );
nand ( n393139 , n72120 , n393138 );
buf ( n393140 , n393139 );
buf ( n393141 , n393140 );
xor ( n72133 , n393122 , n393141 );
buf ( n393143 , n72133 );
buf ( n393144 , n393143 );
xor ( n393145 , n392741 , n392828 );
and ( n72137 , n393145 , n392832 );
and ( n72138 , n392741 , n392828 );
or ( n393148 , n72137 , n72138 );
buf ( n393149 , n393148 );
buf ( n393150 , n393149 );
and ( n393151 , n393144 , n393150 );
not ( n393152 , n393144 );
buf ( n393153 , n393149 );
not ( n393154 , n393153 );
buf ( n393155 , n393154 );
buf ( n393156 , n393155 );
and ( n72148 , n393152 , n393156 );
nor ( n393158 , n393151 , n72148 );
buf ( n393159 , n393158 );
not ( n72151 , n393159 );
not ( n393161 , n72151 );
or ( n393162 , n72110 , n393161 );
not ( n72154 , n392995 );
not ( n72155 , n393040 );
or ( n72156 , n72154 , n72155 );
nand ( n72157 , n72156 , n72108 );
not ( n72158 , n72157 );
nand ( n72159 , n72158 , n393159 );
nand ( n72160 , n393162 , n72159 );
xnor ( n72161 , n392990 , n72160 );
buf ( n393171 , n72161 );
not ( n72163 , n393171 );
buf ( n393173 , n72163 );
xor ( n72165 , n71728 , n393173 );
xor ( n72166 , n392994 , n393040 );
xnor ( n393176 , n72166 , n72107 );
not ( n72168 , n393176 );
not ( n72169 , n72168 );
buf ( n393179 , n392853 );
not ( n393180 , n393179 );
buf ( n393181 , n392986 );
not ( n72173 , n393181 );
or ( n393183 , n393180 , n72173 );
buf ( n393184 , n392983 );
buf ( n393185 , n392834 );
nand ( n72177 , n393184 , n393185 );
buf ( n393187 , n72177 );
buf ( n393188 , n393187 );
nand ( n72180 , n393183 , n393188 );
buf ( n393190 , n72180 );
buf ( n393191 , n393190 );
buf ( n72183 , n392847 );
buf ( n393193 , n72183 );
and ( n393194 , n393191 , n393193 );
not ( n72186 , n393191 );
not ( n393196 , n72183 );
buf ( n393197 , n393196 );
and ( n72189 , n72186 , n393197 );
nor ( n393199 , n393194 , n72189 );
buf ( n393200 , n393199 );
not ( n393201 , n393200 );
or ( n72193 , n72169 , n393201 );
buf ( n393203 , n390543 );
buf ( n393204 , n391250 );
nand ( n72196 , n393203 , n393204 );
buf ( n72197 , n72196 );
buf ( n393207 , n72197 );
buf ( n393208 , n69614 );
and ( n72200 , n393207 , n393208 );
buf ( n393210 , n391263 );
not ( n393211 , n393210 );
buf ( n393212 , n393211 );
buf ( n393213 , n393212 );
nor ( n393214 , n72200 , n393213 );
buf ( n393215 , n393214 );
buf ( n393216 , n393215 );
not ( n72208 , n393216 );
buf ( n393218 , n70236 );
not ( n72210 , n393218 );
or ( n393220 , n72208 , n72210 );
buf ( n393221 , n391326 );
nand ( n72213 , n393220 , n393221 );
buf ( n393223 , n72213 );
buf ( n393224 , n393223 );
buf ( n393225 , n393215 );
not ( n393226 , n393225 );
buf ( n72218 , n391247 );
nand ( n72219 , n393226 , n72218 );
buf ( n72220 , n72219 );
buf ( n393230 , n72220 );
nand ( n72222 , n393224 , n393230 );
buf ( n72223 , n72222 );
buf ( n393233 , n72223 );
buf ( n393234 , n71534 );
not ( n72226 , n393234 );
buf ( n393236 , n392558 );
not ( n393237 , n393236 );
or ( n72229 , n72226 , n393237 );
buf ( n393239 , n71534 );
buf ( n393240 , n392558 );
or ( n72232 , n393239 , n393240 );
nand ( n393242 , n72229 , n72232 );
buf ( n393243 , n393242 );
buf ( n393244 , n393243 );
buf ( n393245 , n71557 );
and ( n72237 , n393244 , n393245 );
not ( n393247 , n393244 );
buf ( n393248 , n392530 );
and ( n393249 , n393247 , n393248 );
nor ( n393250 , n72237 , n393249 );
buf ( n393251 , n393250 );
buf ( n393252 , n393251 );
xor ( n393253 , n393233 , n393252 );
xor ( n72245 , n391347 , n391361 );
and ( n393255 , n72245 , n391382 );
and ( n393256 , n391347 , n391361 );
or ( n72248 , n393255 , n393256 );
buf ( n393258 , n72248 );
buf ( n393259 , n393258 );
and ( n72251 , n393253 , n393259 );
and ( n393261 , n393233 , n393252 );
or ( n72253 , n72251 , n393261 );
buf ( n393263 , n72253 );
buf ( n393264 , n393263 );
buf ( n393265 , n392623 );
buf ( n393266 , n392706 );
xor ( n393267 , n393265 , n393266 );
buf ( n393268 , n71692 );
xor ( n72260 , n393267 , n393268 );
buf ( n393270 , n72260 );
buf ( n393271 , n393270 );
xor ( n72263 , n393264 , n393271 );
xor ( n393273 , n393066 , n393074 );
xor ( n72265 , n393273 , n393092 );
buf ( n393275 , n72265 );
buf ( n72267 , n71648 );
not ( n393277 , n72267 );
buf ( n393278 , n393277 );
not ( n393279 , n393278 );
not ( n393280 , n71635 );
not ( n72272 , n392661 );
or ( n393282 , n393280 , n72272 );
nand ( n72274 , n392636 , n71636 );
nand ( n72275 , n393282 , n72274 );
not ( n72276 , n72275 );
not ( n72277 , n72276 );
or ( n393287 , n393279 , n72277 );
not ( n72279 , n393278 );
nand ( n393289 , n72279 , n72275 );
nand ( n72281 , n393287 , n393289 );
not ( n72282 , n72281 );
or ( n393292 , n393275 , n72282 );
not ( n393293 , n391506 );
nand ( n72285 , n393293 , n391569 );
buf ( n393295 , n72285 );
buf ( n393296 , n70411 );
and ( n72288 , n393295 , n393296 );
buf ( n393298 , n391503 );
nor ( n72290 , n393298 , n391569 );
buf ( n393300 , n72290 );
nor ( n393301 , n72288 , n393300 );
buf ( n393302 , n393301 );
buf ( n393303 , n393302 );
not ( n393304 , n393303 );
buf ( n393305 , n393304 );
nand ( n72297 , n393292 , n393305 );
buf ( n393307 , n72297 );
nand ( n72299 , n393275 , n72282 );
buf ( n393309 , n72299 );
nand ( n72301 , n393307 , n393309 );
buf ( n393311 , n72301 );
buf ( n393312 , n393311 );
and ( n393313 , n72263 , n393312 );
and ( n72305 , n393264 , n393271 );
or ( n72306 , n393313 , n72305 );
buf ( n393316 , n72306 );
nand ( n393317 , n72193 , n393316 );
buf ( n393318 , n393317 );
not ( n393319 , n72168 );
buf ( n393320 , n393200 );
not ( n72312 , n393320 );
buf ( n72313 , n72312 );
nand ( n393323 , n393319 , n72313 );
buf ( n393324 , n393323 );
nand ( n393325 , n393318 , n393324 );
buf ( n393326 , n393325 );
xnor ( n72318 , n72165 , n393326 );
not ( n393328 , n72090 );
not ( n72320 , n393096 );
not ( n72321 , n72320 );
or ( n393331 , n393328 , n72321 );
nand ( n393332 , n393096 , n72089 );
nand ( n72324 , n393331 , n393332 );
and ( n393334 , n72324 , n72104 );
not ( n393335 , n72324 );
not ( n72327 , n72104 );
and ( n393337 , n393335 , n72327 );
nor ( n393338 , n393334 , n393337 );
buf ( n393339 , n393338 );
xor ( n72331 , n71935 , n392974 );
xnor ( n393341 , n72331 , n392873 );
buf ( n393342 , n393341 );
xor ( n393343 , n393339 , n393342 );
xor ( n72335 , n392673 , n71676 );
xor ( n393345 , n72335 , n392698 );
buf ( n393346 , n393345 );
not ( n72338 , n391710 );
or ( n72339 , n391892 , n72338 );
buf ( n393349 , n72339 );
not ( n393350 , n72338 );
not ( n393351 , n391892 );
or ( n72343 , n393350 , n393351 );
nand ( n393353 , n72343 , n391898 );
buf ( n393354 , n393353 );
nand ( n72346 , n393349 , n393354 );
buf ( n393356 , n72346 );
buf ( n393357 , n393356 );
or ( n72349 , n393346 , n393357 );
xor ( n72350 , n391629 , n391635 );
and ( n72351 , n72350 , n391699 );
and ( n393361 , n391629 , n391635 );
or ( n393362 , n72351 , n393361 );
buf ( n393363 , n393362 );
buf ( n72355 , n393363 );
nand ( n393365 , n72349 , n72355 );
buf ( n393366 , n393365 );
buf ( n393367 , n393366 );
buf ( n393368 , n393356 );
buf ( n393369 , n393345 );
nand ( n393370 , n393368 , n393369 );
buf ( n393371 , n393370 );
buf ( n393372 , n393371 );
and ( n393373 , n393367 , n393372 );
buf ( n393374 , n393373 );
buf ( n393375 , n393374 );
and ( n393376 , n393343 , n393375 );
and ( n72368 , n393339 , n393342 );
or ( n72369 , n393376 , n72368 );
buf ( n393379 , n72369 );
xor ( n72371 , n392960 , n392966 );
xor ( n72372 , n72371 , n392970 );
buf ( n393382 , n72372 );
buf ( n393383 , n393382 );
not ( n72375 , n393383 );
buf ( n393385 , n72375 );
buf ( n393386 , n393385 );
not ( n72378 , n393386 );
xor ( n72379 , n393233 , n393252 );
xor ( n72380 , n72379 , n393259 );
buf ( n393390 , n72380 );
buf ( n393391 , n393390 );
not ( n393392 , n393391 );
buf ( n393393 , n393392 );
buf ( n393394 , n393393 );
not ( n393395 , n393394 );
or ( n393396 , n72378 , n393395 );
xor ( n72388 , n391328 , n391385 );
and ( n72389 , n72388 , n391400 );
and ( n393399 , n391328 , n391385 );
or ( n393400 , n72389 , n393399 );
buf ( n393401 , n393400 );
buf ( n393402 , n393401 );
nand ( n393403 , n393396 , n393402 );
buf ( n393404 , n393403 );
buf ( n393405 , n393404 );
buf ( n393406 , n393390 );
buf ( n393407 , n393382 );
nand ( n393408 , n393406 , n393407 );
buf ( n393409 , n393408 );
buf ( n393410 , n393409 );
nand ( n72402 , n393405 , n393410 );
buf ( n393412 , n72402 );
xor ( n393413 , n393264 , n393271 );
xor ( n72405 , n393413 , n393312 );
buf ( n393415 , n72405 );
or ( n393416 , n393412 , n393415 );
buf ( n393417 , n393305 );
not ( n72409 , n393417 );
buf ( n393419 , n72281 );
not ( n393420 , n393419 );
or ( n393421 , n72409 , n393420 );
not ( n72413 , n72281 );
nand ( n393423 , n393302 , n72413 );
buf ( n393424 , n393423 );
nand ( n72416 , n393421 , n393424 );
buf ( n393426 , n72416 );
buf ( n393427 , n393426 );
buf ( n72419 , n393275 );
not ( n72420 , n72419 );
buf ( n393430 , n72420 );
buf ( n72422 , n393430 );
and ( n72423 , n393427 , n72422 );
not ( n393433 , n393427 );
buf ( n72425 , n393275 );
and ( n72426 , n393433 , n72425 );
nor ( n393436 , n72423 , n72426 );
buf ( n393437 , n393436 );
buf ( n393438 , n393437 );
not ( n72430 , n393438 );
buf ( n393440 , n72430 );
buf ( n393441 , n393440 );
not ( n72433 , n393441 );
buf ( n393443 , n393345 );
buf ( n393444 , n393363 );
xor ( n393445 , n393443 , n393444 );
buf ( n393446 , n393356 );
xnor ( n393447 , n393445 , n393446 );
buf ( n393448 , n393447 );
not ( n72440 , n393448 );
buf ( n393450 , n72440 );
not ( n393451 , n393450 );
or ( n393452 , n72433 , n393451 );
buf ( n393453 , n393437 );
not ( n72445 , n393453 );
buf ( n393455 , n393448 );
not ( n72447 , n393455 );
or ( n393457 , n72445 , n72447 );
xor ( n393458 , n391575 , n391590 );
and ( n72450 , n393458 , n391603 );
and ( n393460 , n391575 , n391590 );
or ( n393461 , n72450 , n393460 );
buf ( n393462 , n393461 );
buf ( n393463 , n393462 );
nand ( n393464 , n393457 , n393463 );
buf ( n393465 , n393464 );
buf ( n393466 , n393465 );
nand ( n393467 , n393452 , n393466 );
buf ( n393468 , n393467 );
nand ( n393469 , n393416 , n393468 );
nand ( n72461 , n393415 , n393412 );
and ( n72462 , n393469 , n72461 );
xor ( n393472 , n393379 , n72462 );
not ( n393473 , n393316 );
not ( n393474 , n393473 );
not ( n72466 , n393176 );
or ( n393476 , n393474 , n72466 );
nand ( n393477 , n72168 , n393316 );
nand ( n72469 , n393476 , n393477 );
and ( n72470 , n72469 , n393200 );
not ( n393480 , n72469 );
and ( n393481 , n393480 , n72313 );
nor ( n72473 , n72470 , n393481 );
and ( n72474 , n393472 , n72473 );
and ( n393484 , n393379 , n72462 );
or ( n393485 , n72474 , n393484 );
nand ( n72477 , n72318 , n393485 );
nand ( n72478 , n71497 , n72477 );
xor ( n72479 , n71264 , n71469 );
xnor ( n393489 , n72479 , n392277 );
not ( n393490 , n393159 );
nand ( n72482 , n393490 , n72158 );
not ( n72483 , n72482 );
not ( n72484 , n392990 );
or ( n393494 , n72483 , n72484 );
not ( n393495 , n393490 );
nand ( n72487 , n393495 , n72109 );
nand ( n393497 , n393494 , n72487 );
buf ( n393498 , n393497 );
not ( n393499 , n393498 );
buf ( n393500 , n393499 );
xor ( n72492 , n393489 , n393500 );
buf ( n393502 , n393140 );
buf ( n393503 , n72112 );
or ( n72495 , n393502 , n393503 );
buf ( n393505 , n72495 );
not ( n393506 , n393505 );
not ( n393507 , n393149 );
or ( n72499 , n393506 , n393507 );
and ( n393509 , n393122 , n393141 );
buf ( n393510 , n393509 );
not ( n72502 , n393510 );
nand ( n72503 , n72499 , n72502 );
not ( n393513 , n72503 );
xor ( n393514 , n71199 , n392210 );
xor ( n72506 , n393514 , n71244 );
and ( n393516 , n393513 , n72506 );
not ( n393517 , n393513 );
not ( n72509 , n72506 );
and ( n72510 , n393517 , n72509 );
nor ( n393520 , n393516 , n72510 );
not ( n393521 , n392515 );
not ( n393522 , n392732 );
or ( n72514 , n393521 , n393522 );
buf ( n393524 , n392726 );
not ( n393525 , n393524 );
buf ( n393526 , n392512 );
not ( n72518 , n393526 );
or ( n72519 , n393525 , n72518 );
buf ( n393529 , n392719 );
nand ( n393530 , n72519 , n393529 );
buf ( n393531 , n393530 );
nand ( n393532 , n72514 , n393531 );
and ( n393533 , n393520 , n393532 );
not ( n72525 , n393520 );
not ( n393535 , n393532 );
and ( n393536 , n72525 , n393535 );
nor ( n72528 , n393533 , n393536 );
and ( n72529 , n72492 , n72528 );
and ( n393539 , n393489 , n393500 );
or ( n393540 , n72529 , n393539 );
not ( n393541 , n393540 );
buf ( n393542 , n369689 );
buf ( n393543 , n49900 );
xor ( n393544 , n393542 , n393543 );
buf ( n393545 , n370107 );
xnor ( n72537 , n393544 , n393545 );
buf ( n72538 , n72537 );
buf ( n393548 , n72538 );
nand ( n72540 , n72509 , n393513 );
and ( n72541 , n72540 , n393532 );
not ( n72542 , n72506 );
nor ( n393552 , n72542 , n393513 );
nor ( n393553 , n72541 , n393552 );
buf ( n393554 , n393553 );
xor ( n72546 , n393548 , n393554 );
buf ( n393556 , n71247 );
not ( n393557 , n393556 );
buf ( n393558 , n391997 );
not ( n393559 , n393558 );
or ( n393560 , n393557 , n393559 );
buf ( n393561 , n391994 );
buf ( n393562 , n392259 );
nand ( n393563 , n393561 , n393562 );
buf ( n393564 , n393563 );
buf ( n393565 , n393564 );
nand ( n393566 , n393560 , n393565 );
buf ( n393567 , n393566 );
buf ( n393568 , n393567 );
buf ( n393569 , n392480 );
not ( n393570 , n393569 );
buf ( n393571 , n393570 );
buf ( n393572 , n393571 );
and ( n393573 , n393568 , n393572 );
not ( n72565 , n393568 );
buf ( n393575 , n392480 );
and ( n393576 , n72565 , n393575 );
nor ( n72568 , n393573 , n393576 );
buf ( n393578 , n72568 );
buf ( n393579 , n393578 );
xor ( n72571 , n72546 , n393579 );
buf ( n393581 , n72571 );
not ( n393582 , n393581 );
or ( n393583 , n393541 , n393582 );
xor ( n72575 , n393489 , n393500 );
xor ( n393585 , n72575 , n72528 );
not ( n393586 , n72161 );
buf ( n393587 , n71728 );
not ( n72579 , n393587 );
buf ( n393589 , n72579 );
not ( n393590 , n393589 );
and ( n72582 , n393586 , n393590 );
buf ( n393592 , n71728 );
not ( n393593 , n393592 );
buf ( n393594 , n72161 );
nand ( n72586 , n393593 , n393594 );
buf ( n393596 , n72586 );
and ( n72588 , n393596 , n393326 );
nor ( n393598 , n72582 , n72588 );
nand ( n393599 , n393585 , n393598 );
nand ( n72591 , n393583 , n393599 );
not ( n72592 , n72591 );
xor ( n72593 , n391991 , n392488 );
xor ( n393603 , n71492 , n72593 );
xor ( n393604 , n393548 , n393554 );
and ( n72596 , n393604 , n393579 );
and ( n72597 , n393548 , n393554 );
or ( n72598 , n72596 , n72597 );
buf ( n72599 , n72598 );
nand ( n72600 , n393603 , n72599 );
nand ( n72601 , n72592 , n72600 );
nor ( n72602 , n72478 , n72601 );
nand ( n72603 , n391967 , n391230 );
buf ( n393613 , n69484 );
not ( n72605 , n393613 );
buf ( n393615 , n72605 );
nand ( n393616 , n72603 , n393615 , n391981 );
nand ( n393617 , n72602 , n393616 );
not ( n72609 , n393617 );
and ( n393619 , n390428 , n389596 );
buf ( n393620 , n68665 );
buf ( n393621 , n389590 );
nand ( n72613 , n393620 , n393621 );
buf ( n72614 , n72613 );
buf ( n393624 , n72614 );
buf ( n393625 , n393624 );
buf ( n393626 , n393625 );
buf ( n393627 , n393626 );
nand ( n393628 , n388709 , n67818 );
buf ( n393629 , n393628 );
buf ( n72621 , n393629 );
buf ( n72622 , n72621 );
buf ( n393632 , n72622 );
nand ( n393633 , n393627 , n393632 );
buf ( n393634 , n393633 );
nand ( n72626 , n393619 , n391983 , n393634 );
nand ( n393636 , n391977 , n70963 );
not ( n393637 , n393636 );
nand ( n72629 , n72603 , n393637 );
xor ( n72630 , n393379 , n72462 );
xor ( n393640 , n72630 , n72473 );
xor ( n393641 , n393339 , n393342 );
xor ( n393642 , n393641 , n393375 );
buf ( n393643 , n393642 );
buf ( n393644 , n391605 );
buf ( n393645 , n391402 );
or ( n72637 , n393644 , n393645 );
buf ( n393647 , n391408 );
nand ( n393648 , n72637 , n393647 );
buf ( n393649 , n393648 );
buf ( n393650 , n393649 );
buf ( n393651 , n391605 );
buf ( n393652 , n391402 );
nand ( n393653 , n393651 , n393652 );
buf ( n393654 , n393653 );
buf ( n393655 , n393654 );
nand ( n72647 , n393650 , n393655 );
buf ( n393657 , n72647 );
not ( n393658 , n393657 );
buf ( n393659 , n391919 );
not ( n72651 , n393659 );
buf ( n393661 , n391902 );
not ( n72653 , n393661 );
or ( n72654 , n72651 , n72653 );
buf ( n72655 , n391916 );
not ( n72656 , n72655 );
buf ( n393666 , n70891 );
not ( n393667 , n393666 );
or ( n72659 , n72656 , n393667 );
buf ( n72660 , n391701 );
nand ( n393670 , n72659 , n72660 );
buf ( n393671 , n393670 );
buf ( n393672 , n393671 );
nand ( n393673 , n72654 , n393672 );
buf ( n393674 , n393673 );
not ( n72666 , n393674 );
buf ( n393676 , n393385 );
not ( n393677 , n393676 );
buf ( n393678 , n393390 );
not ( n72670 , n393678 );
or ( n393680 , n393677 , n72670 );
buf ( n393681 , n393393 );
buf ( n393682 , n393382 );
nand ( n72674 , n393681 , n393682 );
buf ( n72675 , n72674 );
buf ( n393685 , n72675 );
nand ( n72677 , n393680 , n393685 );
buf ( n393687 , n72677 );
not ( n393688 , n393401 );
not ( n393689 , n393688 );
or ( n393690 , n393687 , n393689 );
nand ( n72682 , n393689 , n393687 );
nand ( n393692 , n393690 , n72682 );
nand ( n393693 , n72666 , n393692 );
not ( n72685 , n393693 );
or ( n72686 , n393658 , n72685 );
not ( n393696 , n393692 );
nand ( n393697 , n393696 , n393674 );
nand ( n393698 , n72686 , n393697 );
not ( n72690 , n393698 );
xor ( n393700 , n393643 , n72690 );
buf ( n393701 , n393412 );
buf ( n393702 , n393415 );
xor ( n72694 , n393701 , n393702 );
buf ( n393704 , n393468 );
xnor ( n393705 , n72694 , n393704 );
buf ( n393706 , n393705 );
and ( n72698 , n393700 , n393706 );
and ( n72699 , n393643 , n72690 );
or ( n393709 , n72698 , n72699 );
nand ( n393710 , n393640 , n393709 );
buf ( n393711 , n70221 );
not ( n72703 , n393711 );
buf ( n393713 , n72703 );
nand ( n393714 , n393713 , n391964 );
and ( n72706 , n393710 , n393714 );
buf ( n393716 , n393437 );
not ( n72708 , n393716 );
buf ( n393718 , n72440 );
not ( n72710 , n393718 );
or ( n72711 , n72708 , n72710 );
buf ( n393721 , n393448 );
buf ( n393722 , n393440 );
nand ( n72714 , n393721 , n393722 );
buf ( n393724 , n72714 );
buf ( n393725 , n393724 );
nand ( n72717 , n72711 , n393725 );
buf ( n393727 , n72717 );
buf ( n393728 , n393727 );
buf ( n393729 , n393462 );
not ( n72721 , n393729 );
buf ( n393731 , n72721 );
buf ( n393732 , n393731 );
and ( n72724 , n393728 , n393732 );
not ( n72725 , n393728 );
buf ( n393735 , n393462 );
and ( n393736 , n72725 , n393735 );
nor ( n72728 , n72724 , n393736 );
buf ( n393738 , n72728 );
xor ( n72730 , n70614 , n391923 );
and ( n72731 , n72730 , n391937 );
and ( n72732 , n70614 , n391923 );
or ( n393742 , n72731 , n72732 );
buf ( n393743 , n393742 );
xor ( n393744 , n393738 , n393743 );
not ( n72736 , n393688 );
not ( n72737 , n393687 );
not ( n393747 , n72737 );
or ( n393748 , n72736 , n393747 );
nand ( n72740 , n393748 , n72682 );
xor ( n393750 , n393674 , n72740 );
xor ( n393751 , n393750 , n393657 );
xor ( n72743 , n393744 , n393751 );
xor ( n393753 , n391610 , n391940 );
and ( n393754 , n393753 , n391962 );
and ( n72746 , n391610 , n391940 );
or ( n393756 , n393754 , n72746 );
buf ( n393757 , n393756 );
nand ( n72749 , n72743 , n393757 );
xor ( n393759 , n393643 , n72690 );
xor ( n72751 , n393759 , n393706 );
buf ( n393761 , n72751 );
xor ( n72753 , n393738 , n393743 );
and ( n393763 , n72753 , n393751 );
and ( n72755 , n393738 , n393743 );
or ( n393765 , n393763 , n72755 );
buf ( n393766 , n393765 );
nand ( n72758 , n393761 , n393766 );
buf ( n393768 , n72758 );
nand ( n393769 , n72749 , n393768 );
not ( n72761 , n393769 );
nand ( n393771 , n72629 , n72706 , n72761 );
not ( n72763 , n393771 );
nand ( n393773 , n70975 , n72609 , n72626 , n72763 );
nor ( n393774 , n72743 , n393757 );
not ( n72766 , n393774 );
not ( n393776 , n393768 );
or ( n393777 , n72766 , n393776 );
not ( n72769 , n72751 );
not ( n72770 , n393765 );
nand ( n393780 , n72769 , n72770 );
nand ( n72772 , n393777 , n393780 );
buf ( n393782 , n393640 );
not ( n72774 , n393782 );
buf ( n393784 , n72774 );
buf ( n393785 , n393784 );
buf ( n72777 , n393709 );
not ( n393787 , n72777 );
buf ( n393788 , n393787 );
buf ( n393789 , n393788 );
and ( n393790 , n393785 , n393789 );
buf ( n393791 , n393790 );
nor ( n393792 , n72772 , n393791 );
not ( n393793 , n393485 );
not ( n393794 , n72318 );
or ( n72786 , n393793 , n393794 );
nand ( n393796 , n72786 , n393710 );
not ( n393797 , n393796 );
not ( n72789 , n393797 );
nor ( n393799 , n393792 , n72789 );
buf ( n393800 , n393799 );
buf ( n393801 , n393603 );
not ( n72793 , n393801 );
buf ( n393803 , n72793 );
not ( n393804 , n393803 );
buf ( n393805 , n72599 );
not ( n72797 , n393805 );
buf ( n393807 , n72797 );
not ( n393808 , n393807 );
or ( n72800 , n393804 , n393808 );
buf ( n393810 , n71496 );
not ( n393811 , n393810 );
buf ( n393812 , n391987 );
nand ( n393813 , n393811 , n393812 );
buf ( n393814 , n393813 );
nand ( n393815 , n72800 , n393814 );
not ( n72807 , n393815 );
nand ( n72808 , n393581 , n393540 );
not ( n393818 , n72808 );
buf ( n393819 , n393585 );
not ( n393820 , n393819 );
buf ( n393821 , n393820 );
buf ( n393822 , n393598 );
not ( n393823 , n393822 );
buf ( n393824 , n393823 );
nand ( n72816 , n393821 , n393824 );
not ( n393826 , n72816 );
not ( n393827 , n393826 );
or ( n72819 , n393818 , n393827 );
not ( n393829 , n393581 );
not ( n393830 , n393540 );
nand ( n393831 , n393829 , n393830 );
nand ( n72823 , n72819 , n393831 );
buf ( n393833 , n72823 );
not ( n393834 , n393833 );
buf ( n393835 , n393834 );
buf ( n393836 , n72318 );
buf ( n393837 , n393485 );
or ( n72829 , n393836 , n393837 );
buf ( n393839 , n72829 );
nand ( n393840 , n72807 , n393835 , n393839 );
buf ( n72832 , n393840 );
or ( n72833 , n393800 , n72832 );
nor ( n72834 , n72823 , n393815 );
not ( n72835 , n72592 );
and ( n393845 , n72834 , n72835 );
not ( n393846 , n391987 );
nand ( n72838 , n393846 , n71496 );
nand ( n393848 , n72838 , n72600 );
and ( n393849 , n393848 , n393814 );
nor ( n72841 , n393845 , n393849 );
buf ( n393851 , n72841 );
nand ( n393852 , n72833 , n393851 );
buf ( n393853 , n393852 );
nand ( n393854 , n393773 , n393853 );
not ( n72846 , n393854 );
or ( n72847 , n375852 , n72846 );
buf ( n393857 , n377580 );
not ( n72849 , n393857 );
buf ( n393859 , n377585 );
buf ( n393860 , n361716 );
and ( n393861 , n393859 , n393860 );
not ( n72853 , n393859 );
buf ( n393863 , n51996 );
and ( n393864 , n72853 , n393863 );
nor ( n72856 , n393861 , n393864 );
buf ( n393866 , n72856 );
buf ( n393867 , n393866 );
not ( n72859 , n393867 );
or ( n393869 , n72849 , n72859 );
xnor ( n72861 , n377585 , n386701 );
buf ( n393871 , n72861 );
buf ( n393872 , n57530 );
nand ( n72864 , n393871 , n393872 );
buf ( n393874 , n72864 );
buf ( n393875 , n393874 );
nand ( n72867 , n393869 , n393875 );
buf ( n72868 , n72867 );
buf ( n393878 , n72868 );
buf ( n393879 , n369804 );
not ( n393880 , n393879 );
buf ( n72872 , n369763 );
not ( n393882 , n72872 );
buf ( n393883 , n393882 );
buf ( n393884 , n393883 );
not ( n393885 , n393884 );
buf ( n393886 , n363041 );
not ( n393887 , n393886 );
or ( n393888 , n393885 , n393887 );
not ( n72880 , n45152 );
buf ( n393890 , n72880 );
buf ( n393891 , n369763 );
nand ( n393892 , n393890 , n393891 );
buf ( n393893 , n393892 );
buf ( n393894 , n393893 );
nand ( n72886 , n393888 , n393894 );
buf ( n393896 , n72886 );
buf ( n393897 , n393896 );
not ( n393898 , n393897 );
or ( n72890 , n393880 , n393898 );
buf ( n393900 , n393883 );
not ( n393901 , n393900 );
buf ( n393902 , n366187 );
not ( n393903 , n393902 );
or ( n393904 , n393901 , n393903 );
buf ( n393905 , n386390 );
buf ( n393906 , n369763 );
nand ( n393907 , n393905 , n393906 );
buf ( n393908 , n393907 );
buf ( n393909 , n393908 );
nand ( n393910 , n393904 , n393909 );
buf ( n393911 , n393910 );
buf ( n393912 , n393911 );
buf ( n393913 , n49609 );
nand ( n72905 , n393912 , n393913 );
buf ( n393915 , n72905 );
buf ( n393916 , n393915 );
nand ( n72908 , n72890 , n393916 );
buf ( n72909 , n72908 );
buf ( n393919 , n72909 );
not ( n72911 , n393919 );
buf ( n393921 , n368608 );
not ( n393922 , n393921 );
buf ( n393923 , n368549 );
not ( n72915 , n393923 );
buf ( n393925 , n44661 );
not ( n393926 , n393925 );
or ( n72918 , n72915 , n393926 );
buf ( n393928 , n364827 );
buf ( n393929 , n380424 );
nand ( n72921 , n393928 , n393929 );
buf ( n393931 , n72921 );
buf ( n393932 , n393931 );
nand ( n393933 , n72918 , n393932 );
buf ( n393934 , n393933 );
buf ( n393935 , n393934 );
not ( n393936 , n393935 );
or ( n72928 , n393922 , n393936 );
buf ( n72929 , n368549 );
not ( n72930 , n72929 );
buf ( n393940 , n364855 );
not ( n393941 , n393940 );
or ( n72933 , n72930 , n393941 );
buf ( n393943 , n351367 );
buf ( n393944 , n380424 );
nand ( n393945 , n393943 , n393944 );
buf ( n393946 , n393945 );
buf ( n393947 , n393946 );
nand ( n393948 , n72933 , n393947 );
buf ( n393949 , n393948 );
buf ( n393950 , n393949 );
buf ( n393951 , n387542 );
nand ( n393952 , n393950 , n393951 );
buf ( n393953 , n393952 );
buf ( n393954 , n393953 );
nand ( n72946 , n72928 , n393954 );
buf ( n393956 , n72946 );
buf ( n393957 , n393956 );
not ( n72949 , n393957 );
or ( n393959 , n72911 , n72949 );
buf ( n393960 , n72909 );
buf ( n393961 , n393956 );
or ( n393962 , n393960 , n393961 );
buf ( n393963 , n365226 );
not ( n72955 , n393963 );
buf ( n393965 , n342879 );
not ( n393966 , n393965 );
buf ( n393967 , n382496 );
not ( n393968 , n393967 );
or ( n393969 , n393966 , n393968 );
buf ( n393970 , n31231 );
not ( n72962 , n65351 );
buf ( n393972 , n72962 );
nand ( n393973 , n393970 , n393972 );
buf ( n393974 , n393973 );
buf ( n393975 , n393974 );
nand ( n393976 , n393969 , n393975 );
buf ( n393977 , n393976 );
buf ( n393978 , n393977 );
not ( n393979 , n393978 );
or ( n393980 , n72955 , n393979 );
buf ( n393981 , n386047 );
buf ( n393982 , n45075 );
nand ( n393983 , n393981 , n393982 );
buf ( n393984 , n393983 );
buf ( n393985 , n393984 );
nand ( n393986 , n393980 , n393985 );
buf ( n393987 , n393986 );
buf ( n393988 , n393987 );
xor ( n72980 , n386067 , n386084 );
xor ( n72981 , n72980 , n386115 );
buf ( n393991 , n72981 );
buf ( n72983 , n393991 );
xor ( n72984 , n393988 , n72983 );
buf ( n393994 , n365108 );
not ( n393995 , n393994 );
buf ( n393996 , n386108 );
not ( n72988 , n393996 );
or ( n393998 , n393995 , n72988 );
buf ( n72990 , n386091 );
buf ( n394000 , n364975 );
not ( n72992 , n394000 );
buf ( n394002 , n31124 );
not ( n394003 , n394002 );
buf ( n394004 , n394003 );
buf ( n394005 , n394004 );
not ( n394006 , n394005 );
or ( n72998 , n72992 , n394006 );
buf ( n394008 , n351160 );
buf ( n394009 , n386102 );
nand ( n73001 , n394008 , n394009 );
buf ( n394011 , n73001 );
buf ( n394012 , n394011 );
nand ( n73004 , n72998 , n394012 );
buf ( n394014 , n73004 );
buf ( n394015 , n394014 );
nand ( n73007 , n72990 , n394015 );
buf ( n394017 , n73007 );
buf ( n394018 , n394017 );
nand ( n394019 , n393998 , n394018 );
buf ( n394020 , n394019 );
buf ( n394021 , n394020 );
not ( n73013 , n380901 );
buf ( n394023 , n365393 );
not ( n73015 , n394023 );
buf ( n394025 , n366659 );
not ( n394026 , n394025 );
or ( n394027 , n73015 , n394026 );
buf ( n394028 , n365393 );
not ( n394029 , n394028 );
buf ( n394030 , n342617 );
nand ( n73022 , n394029 , n394030 );
buf ( n73023 , n73022 );
buf ( n394033 , n73023 );
nand ( n73025 , n394027 , n394033 );
buf ( n394035 , n73025 );
not ( n73027 , n394035 );
or ( n73028 , n73013 , n73027 );
buf ( n394038 , n351345 );
not ( n73030 , n394038 );
buf ( n394040 , n366659 );
not ( n73032 , n394040 );
or ( n394042 , n73030 , n73032 );
buf ( n394043 , n342617 );
not ( n394044 , n351345 );
buf ( n394045 , n394044 );
nand ( n394046 , n394043 , n394045 );
buf ( n394047 , n394046 );
buf ( n394048 , n394047 );
nand ( n73040 , n394042 , n394048 );
buf ( n394050 , n73040 );
buf ( n394051 , n394050 );
buf ( n394052 , n375920 );
nand ( n394053 , n394051 , n394052 );
buf ( n394054 , n394053 );
nand ( n73046 , n73028 , n394054 );
buf ( n394056 , n73046 );
xor ( n394057 , n394021 , n394056 );
buf ( n394058 , n45075 );
not ( n73050 , n394058 );
buf ( n394060 , n393977 );
not ( n394061 , n394060 );
or ( n394062 , n73050 , n394061 );
and ( n73054 , n31193 , n72962 );
not ( n394064 , n31193 );
not ( n394065 , n65349 );
not ( n394066 , n394065 );
and ( n73058 , n394064 , n394066 );
or ( n394068 , n73054 , n73058 );
buf ( n394069 , n394068 );
buf ( n394070 , n365226 );
nand ( n394071 , n394069 , n394070 );
buf ( n394072 , n394071 );
buf ( n394073 , n394072 );
nand ( n394074 , n394062 , n394073 );
buf ( n394075 , n394074 );
buf ( n394076 , n394075 );
and ( n394077 , n394057 , n394076 );
and ( n394078 , n394021 , n394056 );
or ( n73070 , n394077 , n394078 );
buf ( n394080 , n73070 );
buf ( n394081 , n394080 );
xor ( n73073 , n72984 , n394081 );
buf ( n394083 , n73073 );
buf ( n394084 , n394083 );
nand ( n394085 , n393962 , n394084 );
buf ( n394086 , n394085 );
buf ( n394087 , n394086 );
nand ( n394088 , n393959 , n394087 );
buf ( n394089 , n394088 );
buf ( n394090 , n394089 );
xor ( n394091 , n393878 , n394090 );
buf ( n394092 , n379515 );
buf ( n394093 , n366277 );
and ( n394094 , n394092 , n394093 );
not ( n394095 , n394092 );
buf ( n394096 , n360610 );
and ( n73088 , n394095 , n394096 );
nor ( n394098 , n394094 , n73088 );
buf ( n394099 , n394098 );
buf ( n394100 , n394099 );
not ( n394101 , n394100 );
buf ( n394102 , n46113 );
not ( n73094 , n394102 );
or ( n73095 , n394101 , n73094 );
buf ( n394105 , n377094 );
buf ( n394106 , n360610 );
and ( n73098 , n394105 , n394106 );
not ( n394108 , n394105 );
buf ( n73100 , n45270 );
and ( n394110 , n394108 , n73100 );
nor ( n73102 , n73098 , n394110 );
buf ( n394112 , n73102 );
buf ( n394113 , n394112 );
buf ( n73105 , n366757 );
buf ( n394115 , n73105 );
nand ( n394116 , n394113 , n394115 );
buf ( n394117 , n394116 );
buf ( n394118 , n394117 );
nand ( n394119 , n73095 , n394118 );
buf ( n394120 , n394119 );
buf ( n394121 , n394120 );
and ( n394122 , n394091 , n394121 );
and ( n73114 , n393878 , n394090 );
or ( n394124 , n394122 , n73114 );
buf ( n394125 , n394124 );
not ( n73117 , n394125 );
not ( n73118 , n73117 );
buf ( n394128 , n377757 );
not ( n73120 , n394128 );
buf ( n394130 , n366086 );
not ( n394131 , n394130 );
or ( n394132 , n73120 , n394131 );
buf ( n394133 , n369577 );
buf ( n394134 , n378886 );
nand ( n394135 , n394133 , n394134 );
buf ( n394136 , n394135 );
buf ( n394137 , n394136 );
nand ( n394138 , n394132 , n394137 );
buf ( n394139 , n394138 );
buf ( n73131 , n394139 );
not ( n73132 , n73131 );
buf ( n73133 , n361606 );
not ( n73134 , n73133 );
or ( n73135 , n73132 , n73134 );
buf ( n73136 , n385843 );
buf ( n73137 , n367590 );
nand ( n73138 , n73136 , n73137 );
buf ( n73139 , n73138 );
buf ( n73140 , n73139 );
nand ( n73141 , n73135 , n73140 );
buf ( n73142 , n73141 );
buf ( n394152 , n73142 );
not ( n73144 , n394152 );
buf ( n394154 , n22956 );
buf ( n394155 , n352209 );
and ( n394156 , n394154 , n394155 );
not ( n394157 , n394154 );
buf ( n394158 , n386359 );
and ( n73150 , n394157 , n394158 );
nor ( n394160 , n394156 , n73150 );
buf ( n394161 , n394160 );
not ( n73153 , n394161 );
not ( n394163 , n45014 );
not ( n394164 , n394163 );
and ( n73156 , n73153 , n394164 );
buf ( n394166 , n57280 );
not ( n394167 , n394166 );
not ( n73159 , n352192 );
buf ( n394169 , n73159 );
not ( n394170 , n394169 );
or ( n73162 , n394167 , n394170 );
buf ( n394172 , n352192 );
buf ( n394173 , n377728 );
nand ( n73165 , n394172 , n394173 );
buf ( n394175 , n73165 );
buf ( n394176 , n394175 );
nand ( n73168 , n73162 , n394176 );
buf ( n394178 , n73168 );
and ( n73170 , n394178 , n365152 );
nor ( n73171 , n73156 , n73170 );
buf ( n73172 , n73171 );
buf ( n394182 , n48502 );
not ( n73174 , n394182 );
not ( n394184 , n377712 );
not ( n394185 , n377389 );
and ( n73177 , n394184 , n394185 );
buf ( n394187 , n362417 );
buf ( n394188 , n377389 );
and ( n394189 , n394187 , n394188 );
buf ( n394190 , n394189 );
nor ( n394191 , n73177 , n394190 );
buf ( n394192 , n394191 );
not ( n73184 , n394192 );
and ( n394194 , n73174 , n73184 );
buf ( n394195 , n386131 );
buf ( n394196 , n67754 );
nor ( n73188 , n394195 , n394196 );
buf ( n394198 , n73188 );
buf ( n394199 , n394198 );
nor ( n73191 , n394194 , n394199 );
buf ( n394201 , n73191 );
buf ( n394202 , n394201 );
xor ( n394203 , n73172 , n394202 );
buf ( n394204 , n386119 );
buf ( n394205 , n386054 );
xor ( n73197 , n394204 , n394205 );
buf ( n394207 , n386032 );
not ( n394208 , n394207 );
xor ( n394209 , n73197 , n394208 );
buf ( n394210 , n394209 );
buf ( n394211 , n394210 );
and ( n394212 , n394203 , n394211 );
and ( n73204 , n73172 , n394202 );
or ( n394214 , n394212 , n73204 );
buf ( n394215 , n394214 );
buf ( n394216 , n394215 );
not ( n394217 , n394216 );
and ( n73209 , n73144 , n394217 );
buf ( n394219 , n73142 );
buf ( n394220 , n394215 );
and ( n394221 , n394219 , n394220 );
nor ( n73213 , n73209 , n394221 );
buf ( n73214 , n73213 );
not ( n394224 , n65193 );
not ( n73216 , n361060 );
or ( n394226 , n394224 , n73216 );
buf ( n394227 , n378856 );
not ( n73219 , n394227 );
buf ( n394229 , n45116 );
not ( n73221 , n394229 );
or ( n394231 , n73219 , n73221 );
buf ( n394232 , n365266 );
buf ( n394233 , n378847 );
nand ( n394234 , n394232 , n394233 );
buf ( n394235 , n394234 );
buf ( n394236 , n394235 );
nand ( n73228 , n394231 , n394236 );
buf ( n394238 , n73228 );
nand ( n394239 , n365279 , n394238 );
nand ( n394240 , n394226 , n394239 );
and ( n394241 , n73214 , n394240 );
not ( n73233 , n73214 );
not ( n394243 , n394240 );
and ( n73235 , n73233 , n394243 );
nor ( n73236 , n394241 , n73235 );
buf ( n394246 , n73236 );
not ( n73238 , n394246 );
buf ( n394248 , n73238 );
buf ( n394249 , n394248 );
not ( n73241 , n394249 );
buf ( n394251 , n58923 );
not ( n394252 , n394251 );
buf ( n394253 , n379371 );
not ( n394254 , n394253 );
buf ( n394255 , n360851 );
not ( n73247 , n394255 );
or ( n394257 , n394254 , n73247 );
buf ( n73249 , n379380 );
buf ( n73250 , n362458 );
nand ( n73251 , n73249 , n73250 );
buf ( n73252 , n73251 );
buf ( n73253 , n73252 );
nand ( n73254 , n394257 , n73253 );
buf ( n73255 , n73254 );
buf ( n394265 , n73255 );
not ( n394266 , n394265 );
or ( n73258 , n394252 , n394266 );
buf ( n394268 , n58867 );
buf ( n394269 , n379371 );
not ( n394270 , n394269 );
buf ( n394271 , n360886 );
not ( n394272 , n394271 );
or ( n394273 , n394270 , n394272 );
buf ( n394274 , n390918 );
buf ( n394275 , n379380 );
nand ( n394276 , n394274 , n394275 );
buf ( n394277 , n394276 );
buf ( n394278 , n394277 );
nand ( n394279 , n394273 , n394278 );
buf ( n394280 , n394279 );
buf ( n394281 , n394280 );
nand ( n394282 , n394268 , n394281 );
buf ( n394283 , n394282 );
buf ( n394284 , n394283 );
nand ( n73276 , n73258 , n394284 );
buf ( n394286 , n73276 );
buf ( n394287 , n394286 );
not ( n73279 , n394287 );
buf ( n394289 , n73279 );
buf ( n394290 , n394289 );
not ( n73282 , n394290 );
or ( n73283 , n73241 , n73282 );
buf ( n394293 , n73236 );
buf ( n394294 , n394286 );
nand ( n73286 , n394293 , n394294 );
buf ( n394296 , n73286 );
buf ( n394297 , n394296 );
nand ( n394298 , n73283 , n394297 );
buf ( n394299 , n394298 );
not ( n73291 , n394299 );
not ( n394301 , n73291 );
or ( n73293 , n73118 , n394301 );
not ( n73294 , n73117 );
nand ( n73295 , n73294 , n394299 );
nand ( n73296 , n73293 , n73295 );
not ( n73297 , n73296 );
buf ( n394307 , n73297 );
not ( n73299 , n394307 );
xor ( n73300 , n386019 , n386122 );
xor ( n73301 , n73300 , n386144 );
buf ( n394311 , n73301 );
buf ( n394312 , n394311 );
xor ( n73304 , n393988 , n72983 );
and ( n394314 , n73304 , n394081 );
and ( n73306 , n393988 , n72983 );
or ( n394316 , n394314 , n73306 );
buf ( n394317 , n394316 );
buf ( n394318 , n394317 );
buf ( n394319 , n44915 );
not ( n394320 , n394319 );
buf ( n394321 , n365041 );
not ( n394322 , n394321 );
buf ( n394323 , n44661 );
not ( n394324 , n394323 );
or ( n394325 , n394322 , n394324 );
buf ( n394326 , n31072 );
buf ( n394327 , n380497 );
nand ( n394328 , n394326 , n394327 );
buf ( n394329 , n394328 );
buf ( n394330 , n394329 );
nand ( n394331 , n394325 , n394330 );
buf ( n394332 , n394331 );
buf ( n394333 , n394332 );
not ( n394334 , n394333 );
or ( n394335 , n394320 , n394334 );
buf ( n394336 , n365041 );
not ( n394337 , n394336 );
buf ( n394338 , n44638 );
not ( n394339 , n394338 );
or ( n394340 , n394337 , n394339 );
buf ( n394341 , n364804 );
buf ( n394342 , n380497 );
nand ( n394343 , n394341 , n394342 );
buf ( n394344 , n394343 );
buf ( n394345 , n394344 );
nand ( n394346 , n394340 , n394345 );
buf ( n394347 , n394346 );
buf ( n394348 , n394347 );
buf ( n394349 , n47466 );
nand ( n73317 , n394348 , n394349 );
buf ( n394351 , n73317 );
buf ( n394352 , n394351 );
nand ( n394353 , n394335 , n394352 );
buf ( n394354 , n394353 );
buf ( n394355 , n394354 );
xor ( n394356 , n394318 , n394355 );
buf ( n394357 , n360562 );
not ( n394358 , n394357 );
buf ( n394359 , n367600 );
not ( n73327 , n394359 );
or ( n73328 , n394358 , n73327 );
buf ( n394362 , n378098 );
nand ( n73330 , n73328 , n394362 );
buf ( n394364 , n73330 );
buf ( n394365 , n394364 );
buf ( n394366 , n366151 );
buf ( n394367 , n365569 );
buf ( n394368 , n40461 );
nand ( n394369 , n394367 , n394368 );
buf ( n394370 , n394369 );
buf ( n394371 , n394370 );
and ( n394372 , n394365 , n394366 , n394371 );
buf ( n394373 , n394372 );
buf ( n394374 , n394373 );
and ( n73342 , n394356 , n394374 );
and ( n73343 , n394318 , n394355 );
or ( n73344 , n73342 , n73343 );
buf ( n394378 , n73344 );
buf ( n394379 , n394378 );
xor ( n73347 , n394312 , n394379 );
buf ( n394381 , n394112 );
not ( n73349 , n394381 );
buf ( n394383 , n46557 );
not ( n73351 , n394383 );
or ( n73352 , n73349 , n73351 );
buf ( n394386 , n377068 );
not ( n73354 , n394386 );
buf ( n394388 , n365468 );
not ( n394389 , n394388 );
or ( n73357 , n73354 , n394389 );
buf ( n394391 , n362452 );
buf ( n394392 , n377071 );
nand ( n73360 , n394391 , n394392 );
buf ( n73361 , n73360 );
buf ( n73362 , n73361 );
nand ( n73363 , n73357 , n73362 );
buf ( n73364 , n73363 );
buf ( n73365 , n73364 );
buf ( n394399 , n360577 );
nand ( n73367 , n73365 , n394399 );
buf ( n394401 , n73367 );
buf ( n394402 , n394401 );
nand ( n394403 , n73352 , n394402 );
buf ( n394404 , n394403 );
buf ( n394405 , n394404 );
xor ( n394406 , n73347 , n394405 );
buf ( n394407 , n394406 );
buf ( n394408 , n380356 );
not ( n394409 , n394408 );
buf ( n394410 , n380368 );
not ( n73378 , n394410 );
buf ( n394412 , n366725 );
not ( n73380 , n394412 );
or ( n73381 , n73378 , n73380 );
nand ( n73382 , n59867 , n366722 );
buf ( n394416 , n73382 );
nand ( n73384 , n73381 , n394416 );
buf ( n394418 , n73384 );
buf ( n394419 , n394418 );
not ( n73387 , n394419 );
or ( n73388 , n394409 , n73387 );
buf ( n73389 , n380368 );
not ( n73390 , n73389 );
buf ( n73391 , n69990 );
not ( n73392 , n73391 );
or ( n73393 , n73390 , n73392 );
buf ( n394427 , n40251 );
buf ( n394428 , n384667 );
nand ( n394429 , n394427 , n394428 );
buf ( n394430 , n394429 );
buf ( n394431 , n394430 );
nand ( n394432 , n73393 , n394431 );
buf ( n394433 , n394432 );
buf ( n394434 , n394433 );
buf ( n394435 , n380407 );
nand ( n394436 , n394434 , n394435 );
buf ( n394437 , n394436 );
buf ( n394438 , n394437 );
nand ( n394439 , n73388 , n394438 );
buf ( n394440 , n394439 );
and ( n73408 , n394407 , n394440 );
not ( n394442 , n394407 );
not ( n394443 , n394440 );
and ( n73411 , n394442 , n394443 );
or ( n394445 , n73408 , n73411 );
buf ( n394446 , n379841 );
not ( n73414 , n394446 );
buf ( n394448 , n366407 );
not ( n73416 , n394448 );
or ( n73417 , n73414 , n73416 );
buf ( n73418 , n362285 );
buf ( n394452 , n379847 );
nand ( n73420 , n73418 , n394452 );
buf ( n394454 , n73420 );
buf ( n394455 , n394454 );
nand ( n394456 , n73417 , n394455 );
buf ( n394457 , n394456 );
buf ( n394458 , n394457 );
buf ( n394459 , n379890 );
and ( n73427 , n394458 , n394459 );
buf ( n394461 , n379841 );
not ( n73429 , n394461 );
buf ( n394463 , n45718 );
not ( n394464 , n394463 );
or ( n394465 , n73429 , n394464 );
buf ( n394466 , n362136 );
buf ( n394467 , n379847 );
nand ( n394468 , n394466 , n394467 );
buf ( n394469 , n394468 );
buf ( n394470 , n394469 );
nand ( n394471 , n394465 , n394470 );
buf ( n394472 , n394471 );
buf ( n394473 , n394472 );
not ( n73441 , n394473 );
buf ( n394475 , n59424 );
nor ( n73443 , n73441 , n394475 );
buf ( n394477 , n73443 );
buf ( n394478 , n394477 );
nor ( n73446 , n73427 , n394478 );
buf ( n394480 , n73446 );
buf ( n394481 , n394480 );
not ( n73449 , n394481 );
buf ( n394483 , n73449 );
buf ( n394484 , n394483 );
and ( n73452 , n394445 , n394484 );
not ( n394486 , n394445 );
and ( n394487 , n394486 , n394480 );
nor ( n73455 , n73452 , n394487 );
not ( n394489 , n73455 );
buf ( n394490 , n394489 );
not ( n394491 , n394490 );
or ( n73459 , n73299 , n394491 );
buf ( n394493 , n73296 );
not ( n394494 , n394493 );
buf ( n394495 , n73455 );
not ( n394496 , n394495 );
or ( n394497 , n394494 , n394496 );
not ( n73465 , n49669 );
buf ( n394499 , n377712 );
not ( n394500 , n394499 );
buf ( n394501 , n377352 );
not ( n394502 , n394501 );
and ( n73470 , n394500 , n394502 );
buf ( n394504 , n45595 );
buf ( n394505 , n377352 );
and ( n73473 , n394504 , n394505 );
nor ( n73474 , n73470 , n73473 );
buf ( n394508 , n73474 );
not ( n73476 , n394508 );
not ( n73477 , n73476 );
or ( n73478 , n73465 , n73477 );
not ( n73479 , n362386 );
or ( n73480 , n73479 , n394191 );
nand ( n73481 , n73478 , n73480 );
buf ( n394515 , n47466 );
not ( n394516 , n394515 );
buf ( n394517 , n365041 );
not ( n394518 , n394517 );
buf ( n394519 , n73159 );
not ( n73487 , n394519 );
or ( n394521 , n394518 , n73487 );
buf ( n394522 , n391133 );
buf ( n394523 , n365052 );
nand ( n73491 , n394522 , n394523 );
buf ( n394525 , n73491 );
buf ( n394526 , n394525 );
nand ( n394527 , n394521 , n394526 );
buf ( n394528 , n394527 );
buf ( n394529 , n394528 );
not ( n394530 , n394529 );
or ( n73498 , n394516 , n394530 );
buf ( n394532 , n394347 );
buf ( n394533 , n44915 );
nand ( n394534 , n394532 , n394533 );
buf ( n394535 , n394534 );
buf ( n394536 , n394535 );
nand ( n394537 , n73498 , n394536 );
buf ( n394538 , n394537 );
or ( n394539 , n73481 , n394538 );
not ( n394540 , n375896 );
not ( n73508 , n394050 );
or ( n394542 , n394540 , n73508 );
buf ( n394543 , n385966 );
not ( n73511 , n394543 );
buf ( n394545 , n375920 );
nand ( n73513 , n73511 , n394545 );
buf ( n394547 , n73513 );
nand ( n73515 , n394542 , n394547 );
xor ( n73516 , n384128 , n384131 );
xor ( n394550 , n73516 , n384136 );
xor ( n394551 , n384282 , n63839 );
xor ( n73519 , n394550 , n394551 );
buf ( n394553 , n73519 );
buf ( n394554 , n60054 );
buf ( n394555 , n380844 );
and ( n394556 , n394554 , n394555 );
not ( n394557 , n394554 );
buf ( n394558 , n380838 );
and ( n73526 , n394557 , n394558 );
nor ( n394560 , n394556 , n73526 );
buf ( n394561 , n394560 );
buf ( n394562 , n394561 );
buf ( n394563 , n380581 );
or ( n394564 , n394562 , n394563 );
buf ( n394565 , n384327 );
buf ( n394566 , n378453 );
or ( n73534 , n394565 , n394566 );
nand ( n73535 , n394564 , n73534 );
buf ( n394569 , n73535 );
buf ( n394570 , n376971 );
buf ( n394571 , n384343 );
and ( n394572 , n394570 , n394571 );
buf ( n394573 , n376993 );
buf ( n394574 , n384089 );
and ( n73542 , n394573 , n394574 );
nor ( n73543 , n394572 , n73542 );
buf ( n394577 , n73543 );
buf ( n394578 , n394577 );
buf ( n394579 , n384354 );
or ( n394580 , n394578 , n394579 );
buf ( n73548 , n384350 );
buf ( n394582 , n384082 );
or ( n394583 , n73548 , n394582 );
nand ( n394584 , n394580 , n394583 );
buf ( n394585 , n394584 );
xor ( n73553 , n394569 , n394585 );
buf ( n394587 , n62243 );
buf ( n394588 , n378372 );
and ( n394589 , n394587 , n394588 );
not ( n73557 , n394587 );
buf ( n394591 , n378368 );
and ( n394592 , n73557 , n394591 );
nor ( n73560 , n394589 , n394592 );
buf ( n394594 , n73560 );
buf ( n394595 , n394594 );
buf ( n394596 , n382849 );
or ( n394597 , n394595 , n394596 );
buf ( n394598 , n63651 );
buf ( n394599 , n384157 );
or ( n394600 , n394598 , n394599 );
nand ( n73568 , n394597 , n394600 );
buf ( n394602 , n73568 );
and ( n73570 , n73553 , n394602 );
and ( n73571 , n394569 , n394585 );
or ( n394605 , n73570 , n73571 );
buf ( n394606 , n394605 );
buf ( n394607 , n384205 );
not ( n394608 , n394607 );
buf ( n394609 , n384178 );
not ( n73577 , n394609 );
or ( n394611 , n394608 , n73577 );
buf ( n394612 , n384208 );
nand ( n73580 , n394611 , n394612 );
buf ( n394614 , n73580 );
buf ( n394615 , n394614 );
xor ( n73583 , n394606 , n394615 );
buf ( n394617 , n62202 );
buf ( n394618 , n57800 );
and ( n73586 , n394617 , n394618 );
buf ( n394620 , n382803 );
buf ( n394621 , n376903 );
and ( n394622 , n394620 , n394621 );
nor ( n73590 , n73586 , n394622 );
buf ( n73591 , n73590 );
buf ( n394625 , n73591 );
buf ( n394626 , n378341 );
or ( n394627 , n394625 , n394626 );
buf ( n394628 , n63726 );
buf ( n394629 , n378424 );
or ( n73597 , n394628 , n394629 );
nand ( n394631 , n394627 , n73597 );
buf ( n394632 , n394631 );
buf ( n394633 , n394632 );
buf ( n394634 , n384380 );
buf ( n394635 , n376866 );
and ( n73603 , n394634 , n394635 );
buf ( n394637 , n384386 );
buf ( n394638 , n382743 );
and ( n394639 , n394637 , n394638 );
nor ( n394640 , n73603 , n394639 );
buf ( n394641 , n394640 );
buf ( n394642 , n394641 );
buf ( n394643 , n376924 );
or ( n73611 , n394642 , n394643 );
buf ( n394645 , n63800 );
buf ( n394646 , n56517 );
or ( n394647 , n394645 , n394646 );
nand ( n73615 , n73611 , n394647 );
buf ( n73616 , n73615 );
buf ( n394650 , n73616 );
nand ( n73618 , n376696 , n376698 );
not ( n394652 , n56028 );
not ( n394653 , n394652 );
not ( n73621 , n376690 );
or ( n394655 , n394653 , n73621 );
not ( n73623 , n376695 );
nand ( n394657 , n394655 , n73623 );
xnor ( n73625 , n73618 , n394657 );
buf ( n394659 , n73625 );
buf ( n394660 , n376990 );
and ( n73628 , n394659 , n394660 );
buf ( n394662 , n73625 );
not ( n73630 , n394662 );
buf ( n73631 , n73630 );
buf ( n394665 , n73631 );
buf ( n394666 , n376997 );
and ( n73634 , n394665 , n394666 );
buf ( n394668 , n377003 );
nor ( n73636 , n73628 , n73634 , n394668 );
buf ( n394670 , n73636 );
buf ( n394671 , n394670 );
or ( n394672 , n394650 , n394671 );
buf ( n394673 , n394672 );
buf ( n394674 , n394673 );
xor ( n394675 , n394633 , n394674 );
buf ( n394676 , n380651 );
buf ( n394677 , n380817 );
and ( n73645 , n394676 , n394677 );
buf ( n394679 , n380657 );
buf ( n394680 , n63664 );
and ( n394681 , n394679 , n394680 );
nor ( n73649 , n73645 , n394681 );
buf ( n394683 , n73649 );
buf ( n394684 , n394683 );
buf ( n394685 , n60313 );
or ( n394686 , n394684 , n394685 );
buf ( n394687 , n63668 );
buf ( n394688 , n380733 );
or ( n73656 , n394687 , n394688 );
nand ( n73657 , n394686 , n73656 );
buf ( n394691 , n73657 );
buf ( n394692 , n394691 );
and ( n394693 , n394675 , n394692 );
and ( n394694 , n394633 , n394674 );
or ( n73662 , n394693 , n394694 );
buf ( n394696 , n73662 );
buf ( n394697 , n394696 );
and ( n394698 , n73583 , n394697 );
and ( n73666 , n394606 , n394615 );
or ( n73667 , n394698 , n73666 );
buf ( n394701 , n73667 );
xor ( n394702 , n384251 , n384268 );
xor ( n73670 , n394702 , n384273 );
buf ( n394704 , n73670 );
xor ( n394705 , n394701 , n394704 );
xor ( n73673 , n384339 , n384461 );
xor ( n394707 , n73673 , n384466 );
buf ( n394708 , n394707 );
and ( n73676 , n394705 , n394708 );
and ( n394710 , n394701 , n394704 );
or ( n73678 , n73676 , n394710 );
xor ( n394712 , n384470 , n384473 );
xor ( n73680 , n394712 , n63836 );
and ( n73681 , n73678 , n73680 );
xor ( n394715 , n384360 , n384377 );
xor ( n73683 , n394715 , n384456 );
buf ( n394717 , n73683 );
xor ( n394718 , n384301 , n384318 );
xor ( n394719 , n394718 , n384335 );
and ( n394720 , n394717 , n394719 );
buf ( n394721 , n376743 );
buf ( n394722 , n384421 );
not ( n394723 , n394722 );
buf ( n394724 , n394723 );
buf ( n394725 , n394724 );
and ( n394726 , n394721 , n394725 );
buf ( n394727 , n376871 );
buf ( n394728 , n394724 );
not ( n394729 , n394728 );
buf ( n394730 , n394729 );
buf ( n394731 , n394730 );
and ( n73699 , n394727 , n394731 );
nor ( n394733 , n394726 , n73699 );
buf ( n394734 , n394733 );
buf ( n394735 , n394734 );
buf ( n394736 , n384414 );
or ( n394737 , n394735 , n394736 );
buf ( n394738 , n384429 );
nand ( n394739 , n394737 , n394738 );
buf ( n394740 , n394739 );
buf ( n394741 , n394740 );
buf ( n394742 , n63406 );
buf ( n394743 , n57800 );
and ( n73711 , n394742 , n394743 );
buf ( n394745 , n384054 );
buf ( n394746 , n376903 );
and ( n394747 , n394745 , n394746 );
nor ( n73715 , n73711 , n394747 );
buf ( n73716 , n73715 );
buf ( n394750 , n73716 );
buf ( n394751 , n378341 );
or ( n73719 , n394750 , n394751 );
buf ( n394753 , n73591 );
buf ( n394754 , n378424 );
or ( n73722 , n394753 , n394754 );
nand ( n73723 , n73719 , n73722 );
buf ( n394757 , n73723 );
buf ( n394758 , n394757 );
xor ( n73726 , n394741 , n394758 );
buf ( n394760 , n378468 );
not ( n73728 , n394760 );
buf ( n394762 , n382596 );
buf ( n394763 , n60054 );
or ( n73731 , n394762 , n394763 );
buf ( n394765 , n61992 );
buf ( n394766 , n380570 );
or ( n73734 , n394765 , n394766 );
nand ( n394768 , n73731 , n73734 );
buf ( n394769 , n394768 );
buf ( n394770 , n394769 );
not ( n394771 , n394770 );
or ( n73739 , n73728 , n394771 );
buf ( n394773 , n394561 );
not ( n394774 , n58009 );
buf ( n394775 , n394774 );
or ( n73743 , n394773 , n394775 );
nand ( n73744 , n73739 , n73743 );
buf ( n394778 , n73744 );
buf ( n394779 , n394778 );
and ( n73747 , n73726 , n394779 );
and ( n394781 , n394741 , n394758 );
or ( n394782 , n73747 , n394781 );
buf ( n394783 , n394782 );
xor ( n73751 , n384393 , n384433 );
xor ( n394785 , n73751 , n384451 );
buf ( n394786 , n394785 );
xor ( n73754 , n394783 , n394786 );
buf ( n394788 , n384343 );
buf ( n73756 , n57747 );
and ( n73757 , n394788 , n73756 );
not ( n394791 , n394788 );
buf ( n394792 , n57754 );
and ( n394793 , n394791 , n394792 );
nor ( n73761 , n73757 , n394793 );
buf ( n394795 , n73761 );
buf ( n394796 , n394795 );
buf ( n394797 , n384354 );
or ( n394798 , n394796 , n394797 );
buf ( n394799 , n394577 );
buf ( n394800 , n384082 );
or ( n394801 , n394799 , n394800 );
nand ( n394802 , n394798 , n394801 );
buf ( n394803 , n394802 );
buf ( n394804 , n394803 );
not ( n394805 , n376399 );
nand ( n73773 , n394805 , n56294 );
not ( n394807 , n376427 );
not ( n394808 , n376690 );
or ( n394809 , n394807 , n394808 );
nand ( n73777 , n394809 , n376692 );
or ( n394811 , n73773 , n73777 );
nand ( n394812 , n73777 , n73773 );
nand ( n73780 , n394811 , n394812 );
buf ( n394814 , n73780 );
not ( n394815 , n394814 );
buf ( n394816 , n394815 );
buf ( n394817 , n394816 );
buf ( n394818 , n376997 );
or ( n73786 , n394817 , n394818 );
buf ( n394820 , n73780 );
buf ( n394821 , n376990 );
or ( n73789 , n394820 , n394821 );
buf ( n394823 , n377003 );
not ( n73791 , n394823 );
buf ( n394825 , n73791 );
buf ( n394826 , n394825 );
nand ( n73794 , n73786 , n73789 , n394826 );
buf ( n394828 , n73794 );
buf ( n394829 , n394828 );
buf ( n394830 , n384408 );
or ( n73798 , n320439 , n591 );
nand ( n394832 , n73798 , n376779 );
buf ( n394833 , n394832 );
not ( n394834 , n394833 );
buf ( n394835 , n394834 );
buf ( n394836 , n394835 );
nand ( n394837 , n394830 , n394836 );
buf ( n394838 , n394837 );
buf ( n394839 , n394838 );
buf ( n394840 , n63765 );
buf ( n394841 , n394840 );
not ( n73809 , n394841 );
buf ( n394843 , n394832 );
nand ( n394844 , n73809 , n394843 );
buf ( n394845 , n394844 );
buf ( n394846 , n394845 );
nand ( n394847 , n394839 , n394846 );
buf ( n394848 , n394847 );
buf ( n394849 , n394848 );
nand ( n394850 , n394829 , n394849 );
buf ( n394851 , n394850 );
buf ( n394852 , n394851 );
xor ( n394853 , n394804 , n394852 );
buf ( n394854 , n380735 );
not ( n73822 , n394854 );
buf ( n394856 , n60171 );
buf ( n394857 , n63664 );
or ( n394858 , n394856 , n394857 );
buf ( n394859 , n380680 );
buf ( n394860 , n380817 );
or ( n394861 , n394859 , n394860 );
nand ( n394862 , n394858 , n394861 );
buf ( n394863 , n394862 );
buf ( n394864 , n394863 );
not ( n73832 , n394864 );
or ( n394866 , n73822 , n73832 );
buf ( n394867 , n394683 );
buf ( n394868 , n380733 );
or ( n394869 , n394867 , n394868 );
nand ( n394870 , n394866 , n394869 );
buf ( n394871 , n394870 );
buf ( n394872 , n394871 );
and ( n394873 , n394853 , n394872 );
and ( n394874 , n394804 , n394852 );
or ( n73842 , n394873 , n394874 );
buf ( n394876 , n73842 );
and ( n394877 , n73754 , n394876 );
and ( n73845 , n394783 , n394786 );
or ( n394879 , n394877 , n73845 );
xor ( n73847 , n384301 , n384318 );
xor ( n394881 , n73847 , n384335 );
and ( n394882 , n394879 , n394881 );
and ( n73850 , n394717 , n394879 );
or ( n73851 , n394720 , n394882 , n73850 );
xor ( n394885 , n394701 , n394704 );
xor ( n73853 , n394885 , n394708 );
and ( n73854 , n73851 , n73853 );
xor ( n394888 , n394633 , n394674 );
xor ( n394889 , n394888 , n394692 );
buf ( n394890 , n394889 );
xor ( n73858 , n394569 , n394585 );
xor ( n394892 , n73858 , n394602 );
and ( n394893 , n394890 , n394892 );
buf ( n394894 , n394670 );
not ( n394895 , n394894 );
buf ( n394896 , n73616 );
not ( n73864 , n394896 );
or ( n394898 , n394895 , n73864 );
buf ( n394899 , n394673 );
nand ( n73867 , n394898 , n394899 );
buf ( n394901 , n73867 );
buf ( n394902 , n60089 );
buf ( n394903 , n382835 );
and ( n73871 , n394902 , n394903 );
buf ( n394905 , n60094 );
buf ( n394906 , n62243 );
and ( n73874 , n394905 , n394906 );
nor ( n73875 , n73871 , n73874 );
buf ( n394909 , n73875 );
buf ( n394910 , n394909 );
buf ( n394911 , n382849 );
or ( n394912 , n394910 , n394911 );
buf ( n394913 , n394594 );
buf ( n394914 , n384157 );
or ( n73882 , n394913 , n394914 );
nand ( n73883 , n394912 , n73882 );
buf ( n394917 , n73883 );
xor ( n394918 , n394901 , n394917 );
buf ( n394919 , n63549 );
buf ( n394920 , n57800 );
and ( n394921 , n394919 , n394920 );
buf ( n394922 , n384199 );
buf ( n394923 , n378284 );
and ( n394924 , n394922 , n394923 );
nor ( n394925 , n394921 , n394924 );
buf ( n394926 , n394925 );
buf ( n394927 , n394926 );
buf ( n394928 , n378341 );
or ( n394929 , n394927 , n394928 );
buf ( n394930 , n73716 );
buf ( n394931 , n378424 );
or ( n394932 , n394930 , n394931 );
nand ( n73900 , n394929 , n394932 );
buf ( n73901 , n73900 );
buf ( n394935 , n73625 );
buf ( n394936 , n376866 );
and ( n73904 , n394935 , n394936 );
buf ( n394938 , n73631 );
buf ( n394939 , n382743 );
and ( n73907 , n394938 , n394939 );
nor ( n73908 , n73904 , n73907 );
buf ( n394942 , n73908 );
buf ( n394943 , n394942 );
buf ( n394944 , n376924 );
or ( n73912 , n394943 , n394944 );
buf ( n394946 , n394641 );
buf ( n394947 , n56517 );
or ( n73915 , n394946 , n394947 );
nand ( n73916 , n73912 , n73915 );
buf ( n394950 , n73916 );
xor ( n73918 , n73901 , n394950 );
buf ( n394952 , n58009 );
not ( n394953 , n394952 );
buf ( n394954 , n394769 );
not ( n73922 , n394954 );
or ( n73923 , n394953 , n73922 );
buf ( n394957 , n62202 );
buf ( n394958 , n380570 );
and ( n73926 , n394957 , n394958 );
buf ( n394960 , n382803 );
buf ( n394961 , n60054 );
and ( n73929 , n394960 , n394961 );
nor ( n73930 , n73926 , n73929 );
buf ( n394964 , n73930 );
buf ( n394965 , n394964 );
buf ( n394966 , n380581 );
or ( n73934 , n394965 , n394966 );
nand ( n73935 , n73923 , n73934 );
buf ( n394969 , n73935 );
and ( n394970 , n73918 , n394969 );
and ( n73938 , n73901 , n394950 );
or ( n394972 , n394970 , n73938 );
and ( n394973 , n394918 , n394972 );
and ( n73941 , n394901 , n394917 );
or ( n394975 , n394973 , n73941 );
xor ( n73943 , n394569 , n394585 );
xor ( n73944 , n73943 , n394602 );
and ( n73945 , n394975 , n73944 );
and ( n394979 , n394890 , n394975 );
or ( n394980 , n394893 , n73945 , n394979 );
xor ( n73948 , n394606 , n394615 );
xor ( n394982 , n73948 , n394697 );
buf ( n394983 , n394982 );
xor ( n73951 , n394980 , n394983 );
xor ( n73952 , n384301 , n384318 );
xor ( n73953 , n73952 , n384335 );
xor ( n73954 , n394717 , n394879 );
xor ( n73955 , n73953 , n73954 );
and ( n394989 , n73951 , n73955 );
and ( n73957 , n394980 , n394983 );
or ( n73958 , n394989 , n73957 );
xor ( n394992 , n394701 , n394704 );
xor ( n394993 , n394992 , n394708 );
and ( n394994 , n73958 , n394993 );
and ( n394995 , n73851 , n73958 );
or ( n73963 , n73854 , n394994 , n394995 );
xor ( n394997 , n384470 , n384473 );
xor ( n394998 , n394997 , n63836 );
and ( n73966 , n73963 , n394998 );
and ( n73967 , n73678 , n73963 );
or ( n395001 , n73681 , n73966 , n73967 );
buf ( n395002 , n395001 );
xor ( n395003 , n394553 , n395002 );
buf ( n395004 , n45802 );
not ( n395005 , n395004 );
buf ( n395006 , n61903 );
not ( n73974 , n395006 );
or ( n73975 , n395005 , n73974 );
buf ( n395009 , n22619 );
buf ( n395010 , n60751 );
nand ( n73978 , n395009 , n395010 );
buf ( n395012 , n73978 );
buf ( n395013 , n395012 );
nand ( n395014 , n73975 , n395013 );
buf ( n395015 , n395014 );
buf ( n73983 , n395015 );
not ( n73984 , n73983 );
buf ( n395018 , n384501 );
not ( n73986 , n395018 );
or ( n395020 , n73984 , n73986 );
buf ( n395021 , n386071 );
buf ( n395022 , n56794 );
nand ( n73990 , n395021 , n395022 );
buf ( n395024 , n73990 );
buf ( n395025 , n395024 );
nand ( n73993 , n395020 , n395025 );
buf ( n395027 , n73993 );
buf ( n395028 , n395027 );
and ( n73996 , n395003 , n395028 );
and ( n73997 , n394553 , n395002 );
or ( n395031 , n73996 , n73997 );
buf ( n395032 , n395031 );
xor ( n395033 , n73515 , n395032 );
buf ( n395034 , n50782 );
not ( n74002 , n395034 );
buf ( n395036 , n48458 );
not ( n395037 , n395036 );
buf ( n395038 , n395037 );
buf ( n395039 , n395038 );
buf ( n395040 , n375944 );
and ( n395041 , n395039 , n395040 );
not ( n395042 , n395039 );
buf ( n395043 , n342654 );
and ( n395044 , n395042 , n395043 );
nor ( n395045 , n395041 , n395044 );
buf ( n395046 , n395045 );
buf ( n395047 , n395046 );
not ( n395048 , n395047 );
and ( n74016 , n74002 , n395048 );
buf ( n395050 , n65331 );
buf ( n395051 , n377168 );
nor ( n395052 , n395050 , n395051 );
buf ( n395053 , n395052 );
buf ( n395054 , n395053 );
nor ( n395055 , n74016 , n395054 );
buf ( n395056 , n395055 );
xnor ( n74024 , n395033 , n395056 );
and ( n74025 , n394539 , n74024 );
and ( n395059 , n73481 , n394538 );
nor ( n395060 , n74025 , n395059 );
buf ( n395061 , n395060 );
not ( n395062 , n395061 );
buf ( n395063 , n395062 );
buf ( n395064 , n395063 );
not ( n395065 , n395064 );
buf ( n395066 , n369577 );
not ( n74034 , n395066 );
buf ( n395068 , n377146 );
not ( n395069 , n395068 );
and ( n395070 , n74034 , n395069 );
buf ( n395071 , n45908 );
buf ( n395072 , n377146 );
and ( n395073 , n395071 , n395072 );
nor ( n74041 , n395070 , n395073 );
buf ( n395075 , n74041 );
buf ( n395076 , n395075 );
not ( n395077 , n395076 );
buf ( n395078 , n395077 );
buf ( n395079 , n395078 );
not ( n395080 , n395079 );
buf ( n395081 , n364849 );
not ( n395082 , n395081 );
or ( n395083 , n395080 , n395082 );
buf ( n395084 , n394139 );
buf ( n395085 , n50987 );
nand ( n395086 , n395084 , n395085 );
buf ( n395087 , n395086 );
buf ( n395088 , n395087 );
nand ( n395089 , n395083 , n395088 );
buf ( n395090 , n395089 );
buf ( n395091 , n395090 );
not ( n74059 , n395091 );
buf ( n74060 , n74059 );
buf ( n395094 , n74060 );
not ( n395095 , n395094 );
or ( n395096 , n395065 , n395095 );
buf ( n395097 , n395090 );
buf ( n395098 , n395060 );
nand ( n395099 , n395097 , n395098 );
buf ( n395100 , n395099 );
buf ( n395101 , n395100 );
nand ( n395102 , n395096 , n395101 );
buf ( n395103 , n395102 );
buf ( n395104 , n395103 );
buf ( n395105 , n377068 );
not ( n395106 , n395105 );
buf ( n395107 , n45116 );
not ( n395108 , n395107 );
or ( n74076 , n395106 , n395108 );
not ( n74077 , n64636 );
buf ( n395111 , n74077 );
buf ( n395112 , n377071 );
nand ( n74080 , n395111 , n395112 );
buf ( n395114 , n74080 );
buf ( n395115 , n395114 );
nand ( n395116 , n74076 , n395115 );
buf ( n395117 , n395116 );
buf ( n395118 , n395117 );
not ( n395119 , n395118 );
buf ( n395120 , n365279 );
not ( n74088 , n395120 );
or ( n74089 , n395119 , n74088 );
buf ( n395123 , n361060 );
buf ( n395124 , n394238 );
nand ( n74092 , n395123 , n395124 );
buf ( n395126 , n74092 );
buf ( n395127 , n395126 );
nand ( n395128 , n74089 , n395127 );
buf ( n395129 , n395128 );
buf ( n395130 , n395129 );
buf ( n395131 , n395130 );
buf ( n395132 , n395131 );
buf ( n395133 , n395132 );
xor ( n395134 , n395104 , n395133 );
buf ( n395135 , n395134 );
not ( n74103 , n395135 );
buf ( n395137 , n394433 );
buf ( n395138 , n380356 );
and ( n395139 , n395137 , n395138 );
buf ( n395140 , n380368 );
not ( n74108 , n395140 );
buf ( n395142 , n366676 );
not ( n395143 , n395142 );
or ( n74111 , n74108 , n395143 );
buf ( n395145 , n377990 );
buf ( n395146 , n384667 );
nand ( n395147 , n395145 , n395146 );
buf ( n395148 , n395147 );
buf ( n395149 , n395148 );
nand ( n74117 , n74111 , n395149 );
buf ( n74118 , n74117 );
buf ( n395152 , n74118 );
not ( n74120 , n395152 );
buf ( n395154 , n385064 );
nor ( n395155 , n74120 , n395154 );
buf ( n395156 , n395155 );
buf ( n395157 , n395156 );
nor ( n395158 , n395139 , n395157 );
buf ( n395159 , n395158 );
nand ( n74127 , n74103 , n395159 );
not ( n395161 , n74127 );
buf ( n395162 , n385974 );
not ( n74130 , n395162 );
buf ( n395164 , n386003 );
not ( n395165 , n395164 );
or ( n395166 , n74130 , n395165 );
buf ( n395167 , n386003 );
buf ( n395168 , n385974 );
or ( n395169 , n395167 , n395168 );
nand ( n74137 , n395166 , n395169 );
buf ( n395171 , n74137 );
buf ( n395172 , n395171 );
buf ( n395173 , n386012 );
not ( n395174 , n395173 );
buf ( n395175 , n395174 );
buf ( n395176 , n395175 );
and ( n395177 , n395172 , n395176 );
not ( n74145 , n395172 );
buf ( n395179 , n386012 );
and ( n395180 , n74145 , n395179 );
nor ( n74148 , n395177 , n395180 );
buf ( n395182 , n74148 );
buf ( n395183 , n368994 );
not ( n395184 , n395183 );
buf ( n395185 , n381286 );
not ( n74153 , n395185 );
or ( n395187 , n395184 , n74153 );
buf ( n395188 , n46693 );
buf ( n395189 , n385238 );
nand ( n74157 , n395188 , n395189 );
buf ( n74158 , n74157 );
buf ( n395192 , n74158 );
nand ( n74160 , n395187 , n395192 );
buf ( n395194 , n74160 );
buf ( n395195 , n395194 );
not ( n395196 , n395195 );
buf ( n395197 , n363429 );
not ( n74165 , n395197 );
or ( n395199 , n395196 , n74165 );
buf ( n395200 , n65034 );
buf ( n395201 , n57228 );
nand ( n74169 , n395200 , n395201 );
buf ( n395203 , n74169 );
buf ( n395204 , n395203 );
nand ( n74172 , n395199 , n395204 );
buf ( n395206 , n74172 );
xor ( n395207 , n395182 , n395206 );
not ( n74175 , n395056 );
not ( n74176 , n73515 );
not ( n74177 , n74176 );
and ( n74178 , n74175 , n74177 );
nand ( n74179 , n395056 , n74176 );
and ( n395213 , n74179 , n395032 );
nor ( n395214 , n74178 , n395213 );
xor ( n395215 , n395207 , n395214 );
buf ( n395216 , n395215 );
buf ( n395217 , n49609 );
not ( n395218 , n395217 );
and ( n395219 , n366077 , n369769 );
not ( n74187 , n366077 );
and ( n74188 , n74187 , n369766 );
or ( n395222 , n395219 , n74188 );
buf ( n395223 , n395222 );
not ( n395224 , n395223 );
or ( n74192 , n395218 , n395224 );
buf ( n395226 , n393911 );
buf ( n395227 , n369804 );
nand ( n74195 , n395226 , n395227 );
buf ( n395229 , n74195 );
buf ( n395230 , n395229 );
nand ( n395231 , n74192 , n395230 );
buf ( n395232 , n395231 );
buf ( n395233 , n395232 );
xor ( n74201 , n395216 , n395233 );
buf ( n395235 , n58984 );
not ( n74203 , n395235 );
buf ( n395237 , n44634 );
not ( n395238 , n395237 );
or ( n74206 , n74203 , n395238 );
buf ( n395240 , n45455 );
buf ( n395241 , n379482 );
nand ( n395242 , n395240 , n395241 );
buf ( n395243 , n395242 );
buf ( n74211 , n395243 );
nand ( n395245 , n74206 , n74211 );
buf ( n395246 , n395245 );
buf ( n395247 , n395246 );
not ( n395248 , n395247 );
buf ( n395249 , n362030 );
not ( n395250 , n395249 );
or ( n74218 , n395248 , n395250 );
buf ( n395252 , n41918 );
buf ( n395253 , n377122 );
not ( n395254 , n395253 );
buf ( n395255 , n44634 );
not ( n74223 , n395255 );
or ( n74224 , n395254 , n74223 );
buf ( n395258 , n45455 );
buf ( n395259 , n57463 );
nand ( n74227 , n395258 , n395259 );
buf ( n395261 , n74227 );
buf ( n395262 , n395261 );
nand ( n74230 , n74224 , n395262 );
buf ( n395264 , n74230 );
buf ( n395265 , n395264 );
nand ( n74233 , n395252 , n395265 );
buf ( n395267 , n74233 );
buf ( n395268 , n395267 );
nand ( n74236 , n74218 , n395268 );
buf ( n395270 , n74236 );
buf ( n395271 , n395270 );
xor ( n74239 , n74201 , n395271 );
buf ( n395273 , n74239 );
not ( n395274 , n395273 );
or ( n395275 , n395161 , n395274 );
buf ( n395276 , n395159 );
not ( n74244 , n395276 );
buf ( n395278 , n395135 );
nand ( n395279 , n74244 , n395278 );
buf ( n395280 , n395279 );
nand ( n74248 , n395275 , n395280 );
buf ( n395282 , n74248 );
nand ( n395283 , n394497 , n395282 );
buf ( n395284 , n395283 );
buf ( n395285 , n395284 );
nand ( n395286 , n73459 , n395285 );
buf ( n395287 , n395286 );
buf ( n395288 , n395287 );
buf ( n395289 , n383713 );
buf ( n395290 , n383722 );
xor ( n395291 , n395289 , n395290 );
buf ( n395292 , n63047 );
xnor ( n395293 , n395291 , n395292 );
buf ( n395294 , n395293 );
buf ( n395295 , n395294 );
buf ( n395296 , n377580 );
not ( n74264 , n395296 );
buf ( n395298 , n385674 );
not ( n395299 , n395298 );
or ( n395300 , n74264 , n395299 );
and ( n395301 , n377585 , n365760 );
not ( n74269 , n377585 );
and ( n395303 , n74269 , n361667 );
or ( n395304 , n395301 , n395303 );
buf ( n395305 , n395304 );
buf ( n395306 , n57530 );
nand ( n395307 , n395305 , n395306 );
buf ( n395308 , n395307 );
buf ( n395309 , n395308 );
nand ( n74277 , n395300 , n395309 );
buf ( n395311 , n74277 );
buf ( n74279 , n395311 );
xor ( n74280 , n395295 , n74279 );
buf ( n395314 , n395264 );
not ( n395315 , n395314 );
buf ( n395316 , n366046 );
not ( n395317 , n395316 );
or ( n395318 , n395315 , n395317 );
buf ( n395319 , n371063 );
buf ( n395320 , n385913 );
nand ( n395321 , n395319 , n395320 );
buf ( n395322 , n395321 );
buf ( n395323 , n395322 );
nand ( n74291 , n395318 , n395323 );
buf ( n395325 , n74291 );
not ( n395326 , n395325 );
buf ( n395327 , n359312 );
buf ( n395328 , n378098 );
nand ( n395329 , n395327 , n395328 );
buf ( n395330 , n395329 );
buf ( n395331 , n395330 );
not ( n395332 , n395331 );
buf ( n395333 , n395332 );
not ( n74301 , n395333 );
or ( n395335 , n395326 , n74301 );
buf ( n395336 , n395325 );
buf ( n395337 , n395333 );
nor ( n74305 , n395336 , n395337 );
buf ( n74306 , n74305 );
buf ( n395340 , n395206 );
not ( n74308 , n395340 );
buf ( n395342 , n74308 );
buf ( n395343 , n395342 );
not ( n74311 , n395343 );
buf ( n395345 , n395214 );
not ( n395346 , n395345 );
or ( n395347 , n74311 , n395346 );
buf ( n74315 , n395182 );
not ( n395349 , n74315 );
buf ( n395350 , n395349 );
buf ( n395351 , n395350 );
nand ( n395352 , n395347 , n395351 );
buf ( n395353 , n395352 );
buf ( n395354 , n395353 );
buf ( n395355 , n395214 );
not ( n395356 , n395355 );
buf ( n395357 , n395206 );
nand ( n395358 , n395356 , n395357 );
buf ( n395359 , n395358 );
buf ( n395360 , n395359 );
nand ( n74328 , n395354 , n395360 );
buf ( n74329 , n74328 );
buf ( n395363 , n74329 );
not ( n74331 , n395363 );
buf ( n395365 , n74331 );
or ( n395366 , n74306 , n395365 );
nand ( n74334 , n395335 , n395366 );
buf ( n395368 , n74334 );
xor ( n395369 , n74280 , n395368 );
buf ( n395370 , n395369 );
buf ( n395371 , n395370 );
not ( n74339 , n394248 );
not ( n74340 , n394286 );
or ( n395374 , n74339 , n74340 );
not ( n395375 , n394289 );
not ( n74343 , n73236 );
or ( n395377 , n395375 , n74343 );
nand ( n74345 , n395377 , n394125 );
nand ( n395379 , n395374 , n74345 );
buf ( n395380 , n395379 );
xor ( n74348 , n395371 , n395380 );
not ( n395382 , n394440 );
not ( n395383 , n394483 );
or ( n74351 , n395382 , n395383 );
not ( n395385 , n394480 );
not ( n395386 , n394443 );
or ( n74354 , n395385 , n395386 );
nand ( n74355 , n74354 , n394407 );
nand ( n395389 , n74351 , n74355 );
buf ( n395390 , n395389 );
xor ( n395391 , n74348 , n395390 );
buf ( n395392 , n395391 );
buf ( n395393 , n395392 );
or ( n395394 , n395288 , n395393 );
buf ( n395395 , n58871 );
not ( n74363 , n395395 );
buf ( n395397 , n379371 );
not ( n74365 , n395397 );
buf ( n395399 , n370566 );
not ( n395400 , n395399 );
or ( n74368 , n74365 , n395400 );
buf ( n395402 , n42149 );
buf ( n395403 , n379380 );
nand ( n395404 , n395402 , n395403 );
buf ( n395405 , n395404 );
buf ( n395406 , n395405 );
nand ( n74374 , n74368 , n395406 );
buf ( n395408 , n74374 );
buf ( n395409 , n395408 );
not ( n395410 , n395409 );
or ( n74378 , n74363 , n395410 );
buf ( n395412 , n394280 );
buf ( n395413 , n58923 );
nand ( n395414 , n395412 , n395413 );
buf ( n395415 , n395414 );
buf ( n395416 , n395415 );
nand ( n74384 , n74378 , n395416 );
buf ( n395418 , n74384 );
xor ( n74386 , n393878 , n394090 );
xor ( n74387 , n74386 , n394121 );
buf ( n395421 , n74387 );
xor ( n74389 , n395418 , n395421 );
buf ( n395423 , n41882 );
not ( n74391 , n395423 );
buf ( n395425 , n377068 );
buf ( n395426 , n44634 );
and ( n395427 , n395425 , n395426 );
not ( n74395 , n395425 );
buf ( n395429 , n41892 );
and ( n74397 , n74395 , n395429 );
nor ( n395431 , n395427 , n74397 );
buf ( n395432 , n395431 );
buf ( n395433 , n395432 );
not ( n74401 , n395433 );
and ( n74402 , n74391 , n74401 );
buf ( n395436 , n378856 );
buf ( n395437 , n44634 );
and ( n74405 , n395436 , n395437 );
not ( n74406 , n395436 );
buf ( n395440 , n41892 );
and ( n74408 , n74406 , n395440 );
nor ( n395442 , n74405 , n74408 );
buf ( n395443 , n395442 );
buf ( n395444 , n395443 );
buf ( n395445 , n365619 );
nor ( n74413 , n395444 , n395445 );
buf ( n74414 , n74413 );
buf ( n395448 , n74414 );
nor ( n74416 , n74402 , n395448 );
buf ( n74417 , n74416 );
buf ( n395451 , n74417 );
not ( n74419 , n395451 );
buf ( n395453 , n74419 );
buf ( n395454 , n395453 );
not ( n74422 , n395454 );
buf ( n395456 , n361971 );
not ( n74424 , n395456 );
buf ( n395458 , n377146 );
buf ( n395459 , n364744 );
and ( n395460 , n395458 , n395459 );
not ( n74428 , n395458 );
buf ( n395462 , n364783 );
and ( n395463 , n74428 , n395462 );
nor ( n74431 , n395460 , n395463 );
buf ( n74432 , n74431 );
buf ( n395466 , n74432 );
not ( n74434 , n395466 );
and ( n395468 , n74424 , n74434 );
buf ( n395469 , n377757 );
buf ( n395470 , n367248 );
and ( n395471 , n395469 , n395470 );
not ( n395472 , n395469 );
buf ( n395473 , n361911 );
and ( n74441 , n395472 , n395473 );
nor ( n395475 , n395471 , n74441 );
buf ( n395476 , n395475 );
buf ( n395477 , n395476 );
buf ( n395478 , n369896 );
nor ( n74446 , n395477 , n395478 );
buf ( n395480 , n74446 );
buf ( n395481 , n395480 );
nor ( n74449 , n395468 , n395481 );
buf ( n395483 , n74449 );
buf ( n395484 , n395483 );
not ( n74452 , n395484 );
buf ( n395486 , n74452 );
buf ( n395487 , n395486 );
not ( n74455 , n395487 );
or ( n395489 , n74422 , n74455 );
buf ( n395490 , n74417 );
not ( n395491 , n395490 );
buf ( n395492 , n395483 );
not ( n395493 , n395492 );
or ( n395494 , n395491 , n395493 );
buf ( n395495 , n365152 );
not ( n74463 , n395495 );
buf ( n395497 , n22955 );
buf ( n395498 , n395497 );
not ( n74466 , n395498 );
buf ( n395500 , n377297 );
not ( n395501 , n395500 );
or ( n74469 , n74466 , n395501 );
buf ( n395503 , n351291 );
buf ( n395504 , n342908 );
nand ( n395505 , n395503 , n395504 );
buf ( n395506 , n395505 );
buf ( n395507 , n395506 );
nand ( n395508 , n74469 , n395507 );
buf ( n395509 , n395508 );
buf ( n395510 , n395509 );
not ( n395511 , n395510 );
or ( n74479 , n74463 , n395511 );
buf ( n74480 , n57280 );
not ( n74481 , n74480 );
buf ( n74482 , n375886 );
not ( n74483 , n74482 );
or ( n74484 , n74481 , n74483 );
buf ( n395518 , n365440 );
buf ( n395519 , n342908 );
nand ( n74487 , n395518 , n395519 );
buf ( n395521 , n74487 );
buf ( n395522 , n395521 );
nand ( n395523 , n74484 , n395522 );
buf ( n395524 , n395523 );
buf ( n395525 , n395524 );
buf ( n395526 , n45014 );
nand ( n74494 , n395525 , n395526 );
buf ( n395528 , n74494 );
buf ( n395529 , n395528 );
nand ( n74497 , n74479 , n395529 );
buf ( n395531 , n74497 );
buf ( n395532 , n395531 );
buf ( n395533 , n365722 );
buf ( n395534 , n351345 );
not ( n74502 , n395534 );
buf ( n395536 , n61903 );
not ( n395537 , n395536 );
or ( n395538 , n74502 , n395537 );
buf ( n395539 , n61903 );
not ( n395540 , n395539 );
buf ( n395541 , n395540 );
buf ( n395542 , n395541 );
buf ( n395543 , n394044 );
nand ( n395544 , n395542 , n395543 );
buf ( n395545 , n395544 );
buf ( n395546 , n395545 );
nand ( n395547 , n395538 , n395546 );
buf ( n395548 , n395547 );
buf ( n395549 , n395548 );
not ( n74517 , n395549 );
buf ( n395551 , n74517 );
buf ( n395552 , n395551 );
or ( n74520 , n395533 , n395552 );
buf ( n395554 , n395015 );
not ( n74522 , n395554 );
buf ( n395556 , n74522 );
buf ( n395557 , n395556 );
buf ( n395558 , n56794 );
not ( n395559 , n395558 );
buf ( n395560 , n395559 );
buf ( n395561 , n395560 );
or ( n74529 , n395557 , n395561 );
nand ( n395563 , n74520 , n74529 );
buf ( n395564 , n395563 );
buf ( n395565 , n395564 );
xor ( n74533 , n394701 , n394704 );
xor ( n395567 , n74533 , n394708 );
xor ( n395568 , n73851 , n73958 );
xor ( n74536 , n395567 , n395568 );
buf ( n395570 , n74536 );
buf ( n395571 , n380651 );
buf ( n395572 , n382835 );
and ( n395573 , n395571 , n395572 );
buf ( n395574 , n380657 );
buf ( n395575 , n62243 );
and ( n74543 , n395574 , n395575 );
nor ( n395577 , n395573 , n74543 );
buf ( n395578 , n395577 );
buf ( n395579 , n395578 );
buf ( n395580 , n382849 );
or ( n74548 , n395579 , n395580 );
buf ( n395582 , n394909 );
buf ( n395583 , n384157 );
or ( n74551 , n395582 , n395583 );
nand ( n74552 , n74548 , n74551 );
buf ( n395586 , n74552 );
buf ( n395587 , n394828 );
buf ( n395588 , n394848 );
or ( n395589 , n395587 , n395588 );
buf ( n395590 , n394851 );
nand ( n74558 , n395589 , n395590 );
buf ( n395592 , n74558 );
xor ( n74560 , n395586 , n395592 );
buf ( n395594 , n380730 );
not ( n395595 , n395594 );
buf ( n395596 , n394863 );
not ( n395597 , n395596 );
or ( n395598 , n395595 , n395597 );
buf ( n395599 , n380838 );
buf ( n395600 , n380817 );
and ( n74568 , n395599 , n395600 );
buf ( n395602 , n380844 );
buf ( n395603 , n57983 );
and ( n74571 , n395602 , n395603 );
nor ( n395605 , n74568 , n74571 );
buf ( n395606 , n395605 );
buf ( n395607 , n395606 );
buf ( n395608 , n60313 );
or ( n74576 , n395607 , n395608 );
nand ( n395610 , n395598 , n74576 );
buf ( n395611 , n395610 );
and ( n74579 , n74560 , n395611 );
and ( n395613 , n395586 , n395592 );
or ( n74581 , n74579 , n395613 );
buf ( n395615 , n74581 );
xor ( n74583 , n394741 , n394758 );
xor ( n395617 , n74583 , n394779 );
buf ( n395618 , n395617 );
buf ( n395619 , n395618 );
xor ( n74587 , n395615 , n395619 );
buf ( n395621 , n376971 );
buf ( n395622 , n394724 );
and ( n395623 , n395621 , n395622 );
buf ( n395624 , n376993 );
buf ( n395625 , n394730 );
and ( n395626 , n395624 , n395625 );
nor ( n74594 , n395623 , n395626 );
buf ( n74595 , n74594 );
buf ( n395629 , n74595 );
buf ( n395630 , n384414 );
or ( n395631 , n395629 , n395630 );
buf ( n395632 , n394734 );
buf ( n395633 , n384411 );
not ( n395634 , n395633 );
buf ( n395635 , n395634 );
buf ( n395636 , n395635 );
or ( n395637 , n395632 , n395636 );
nand ( n395638 , n395631 , n395637 );
buf ( n395639 , n395638 );
buf ( n395640 , n395639 );
not ( n395641 , n384343 );
not ( n74609 , n378372 );
or ( n74610 , n395641 , n74609 );
or ( n74611 , n378372 , n384343 );
nand ( n395645 , n74610 , n74611 );
buf ( n395646 , n395645 );
buf ( n395647 , n384354 );
or ( n74615 , n395646 , n395647 );
buf ( n395649 , n394795 );
buf ( n395650 , n384082 );
or ( n395651 , n395649 , n395650 );
nand ( n395652 , n74615 , n395651 );
buf ( n395653 , n395652 );
buf ( n395654 , n395653 );
xor ( n395655 , n395640 , n395654 );
buf ( n395656 , n382743 );
buf ( n395657 , n73780 );
and ( n395658 , n395656 , n395657 );
not ( n74626 , n395656 );
buf ( n395660 , n394816 );
and ( n395661 , n74626 , n395660 );
nor ( n74629 , n395658 , n395661 );
buf ( n74630 , n74629 );
buf ( n395664 , n74630 );
not ( n74632 , n395664 );
buf ( n74633 , n74632 );
buf ( n395667 , n74633 );
buf ( n395668 , n376924 );
or ( n395669 , n395667 , n395668 );
buf ( n395670 , n394942 );
buf ( n395671 , n56517 );
or ( n395672 , n395670 , n395671 );
nand ( n395673 , n395669 , n395672 );
buf ( n395674 , n395673 );
buf ( n395675 , n395674 );
and ( n395676 , n376427 , n376692 );
xor ( n74644 , n395676 , n376690 );
buf ( n395678 , n74644 );
buf ( n395679 , n376990 );
and ( n74647 , n395678 , n395679 );
buf ( n395681 , n74644 );
not ( n395682 , n395681 );
buf ( n395683 , n395682 );
buf ( n395684 , n395683 );
buf ( n395685 , n376997 );
and ( n395686 , n395684 , n395685 );
buf ( n395687 , n377003 );
nor ( n395688 , n74647 , n395686 , n395687 );
buf ( n395689 , n395688 );
buf ( n395690 , n395689 );
xor ( n395691 , n395675 , n395690 );
buf ( n395692 , n378468 );
not ( n395693 , n395692 );
buf ( n395694 , n63406 );
buf ( n395695 , n380570 );
and ( n395696 , n395694 , n395695 );
buf ( n395697 , n384054 );
buf ( n395698 , n60054 );
and ( n395699 , n395697 , n395698 );
nor ( n395700 , n395696 , n395699 );
buf ( n395701 , n395700 );
buf ( n395702 , n395701 );
not ( n395703 , n395702 );
buf ( n395704 , n395703 );
buf ( n395705 , n395704 );
not ( n395706 , n395705 );
or ( n74674 , n395693 , n395706 );
buf ( n395708 , n394964 );
buf ( n395709 , n394774 );
or ( n74677 , n395708 , n395709 );
nand ( n395711 , n74674 , n74677 );
buf ( n395712 , n395711 );
buf ( n395713 , n395712 );
and ( n74681 , n395691 , n395713 );
and ( n74682 , n395675 , n395690 );
or ( n74683 , n74681 , n74682 );
buf ( n395717 , n74683 );
buf ( n395718 , n395717 );
and ( n74686 , n395655 , n395718 );
and ( n74687 , n395640 , n395654 );
or ( n74688 , n74686 , n74687 );
buf ( n395722 , n74688 );
buf ( n395723 , n395722 );
and ( n74691 , n74587 , n395723 );
and ( n74692 , n395615 , n395619 );
or ( n395726 , n74691 , n74692 );
buf ( n395727 , n395726 );
xor ( n395728 , n394783 , n394786 );
xor ( n74696 , n395728 , n394876 );
and ( n395730 , n395727 , n74696 );
xor ( n74698 , n394569 , n394585 );
xor ( n395732 , n74698 , n394602 );
xor ( n74700 , n394890 , n394975 );
xor ( n74701 , n395732 , n74700 );
xor ( n395735 , n394783 , n394786 );
xor ( n74703 , n395735 , n394876 );
and ( n395737 , n74701 , n74703 );
and ( n74705 , n395727 , n74701 );
or ( n395739 , n395730 , n395737 , n74705 );
xor ( n395740 , n394980 , n394983 );
xor ( n74708 , n395740 , n73955 );
and ( n395742 , n395739 , n74708 );
xor ( n395743 , n395615 , n395619 );
xor ( n74711 , n395743 , n395723 );
buf ( n395745 , n74711 );
xor ( n395746 , n395675 , n395690 );
xor ( n395747 , n395746 , n395713 );
buf ( n395748 , n395747 );
buf ( n395749 , n395748 );
buf ( n395750 , n60089 );
buf ( n395751 , n384343 );
and ( n395752 , n395750 , n395751 );
buf ( n395753 , n60094 );
buf ( n395754 , n384089 );
and ( n395755 , n395753 , n395754 );
nor ( n395756 , n395752 , n395755 );
buf ( n395757 , n395756 );
buf ( n395758 , n395757 );
buf ( n395759 , n384354 );
or ( n395760 , n395758 , n395759 );
buf ( n395761 , n395645 );
buf ( n395762 , n384082 );
or ( n395763 , n395761 , n395762 );
nand ( n74731 , n395760 , n395763 );
buf ( n395765 , n74731 );
buf ( n395766 , n395765 );
xor ( n74734 , n395749 , n395766 );
or ( n395768 , n394774 , n395701 );
not ( n395769 , n380581 );
and ( n74737 , n63549 , n60054 );
not ( n395771 , n63549 );
and ( n395772 , n395771 , n57789 );
nor ( n74740 , n74737 , n395772 );
nand ( n395774 , n395769 , n74740 );
nand ( n395775 , n395768 , n395774 );
buf ( n395776 , n73625 );
buf ( n395777 , n57800 );
and ( n395778 , n395776 , n395777 );
buf ( n74746 , n73631 );
buf ( n395780 , n376903 );
and ( n395781 , n74746 , n395780 );
nor ( n395782 , n395778 , n395781 );
buf ( n395783 , n395782 );
buf ( n395784 , n395783 );
buf ( n395785 , n378341 );
or ( n74753 , n395784 , n395785 );
buf ( n395787 , n384380 );
buf ( n395788 , n57800 );
and ( n74756 , n395787 , n395788 );
buf ( n395790 , n384386 );
buf ( n395791 , n378284 );
and ( n395792 , n395790 , n395791 );
nor ( n74760 , n74756 , n395792 );
buf ( n395794 , n74760 );
buf ( n395795 , n395794 );
buf ( n395796 , n378424 );
or ( n74764 , n395795 , n395796 );
nand ( n395798 , n74753 , n74764 );
buf ( n395799 , n395798 );
xor ( n74767 , n395775 , n395799 );
not ( n395801 , n56087 );
not ( n395802 , n395801 );
not ( n74770 , n56280 );
or ( n395804 , n395802 , n74770 );
nand ( n74772 , n395804 , n56284 );
not ( n74773 , n56062 );
nand ( n395807 , n74773 , n376687 );
or ( n74775 , n74772 , n395807 );
nand ( n395809 , n74772 , n395807 );
nand ( n395810 , n74775 , n395809 );
buf ( n395811 , n395810 );
buf ( n395812 , n376990 );
and ( n74780 , n395811 , n395812 );
buf ( n395814 , n395810 );
not ( n395815 , n395814 );
buf ( n395816 , n395815 );
buf ( n395817 , n395816 );
buf ( n395818 , n376997 );
and ( n74786 , n395817 , n395818 );
buf ( n395820 , n377003 );
nor ( n74788 , n74780 , n74786 , n395820 );
buf ( n395822 , n74788 );
buf ( n395823 , n395822 );
not ( n74791 , n56517 );
buf ( n395825 , n74791 );
not ( n74793 , n395825 );
buf ( n395827 , n74630 );
not ( n395828 , n395827 );
or ( n395829 , n74793 , n395828 );
buf ( n395830 , n74644 );
buf ( n395831 , n376866 );
and ( n395832 , n395830 , n395831 );
buf ( n395833 , n395683 );
buf ( n395834 , n382743 );
and ( n395835 , n395833 , n395834 );
nor ( n395836 , n395832 , n395835 );
buf ( n395837 , n395836 );
buf ( n395838 , n395837 );
buf ( n395839 , n376924 );
or ( n74807 , n395838 , n395839 );
nand ( n395841 , n395829 , n74807 );
buf ( n395842 , n395841 );
buf ( n395843 , n395842 );
xor ( n395844 , n395823 , n395843 );
buf ( n395845 , n395844 );
and ( n74813 , n74767 , n395845 );
and ( n74814 , n395775 , n395799 );
or ( n74815 , n74813 , n74814 );
buf ( n395849 , n74815 );
and ( n74817 , n74734 , n395849 );
and ( n395851 , n395749 , n395766 );
or ( n74819 , n74817 , n395851 );
buf ( n395853 , n74819 );
xor ( n74821 , n395586 , n395592 );
xor ( n74822 , n74821 , n395611 );
and ( n395856 , n395853 , n74822 );
xor ( n74824 , n395640 , n395654 );
xor ( n395858 , n74824 , n395718 );
buf ( n395859 , n395858 );
xor ( n74827 , n395586 , n395592 );
xor ( n395861 , n74827 , n395611 );
and ( n395862 , n395859 , n395861 );
and ( n74830 , n395853 , n395859 );
or ( n395864 , n395856 , n395862 , n74830 );
xor ( n395865 , n395745 , n395864 );
xor ( n74833 , n394901 , n394917 );
xor ( n395867 , n74833 , n394972 );
xor ( n395868 , n394804 , n394852 );
xor ( n395869 , n395868 , n394872 );
buf ( n395870 , n395869 );
and ( n395871 , n395823 , n395843 );
buf ( n395872 , n395871 );
buf ( n395873 , n395872 );
buf ( n395874 , n395794 );
buf ( n395875 , n378341 );
or ( n74843 , n395874 , n395875 );
buf ( n395877 , n394926 );
buf ( n395878 , n378424 );
or ( n395879 , n395877 , n395878 );
nand ( n74847 , n74843 , n395879 );
buf ( n74848 , n74847 );
buf ( n395882 , n74848 );
xor ( n74850 , n395873 , n395882 );
buf ( n395884 , n376743 );
buf ( n395885 , n394840 );
and ( n74853 , n395884 , n395885 );
buf ( n395887 , n376871 );
buf ( n395888 , n394840 );
not ( n74856 , n395888 );
buf ( n395890 , n74856 );
buf ( n395891 , n395890 );
and ( n74859 , n395887 , n395891 );
nor ( n395893 , n74853 , n74859 );
buf ( n395894 , n395893 );
buf ( n395895 , n395894 );
buf ( n395896 , n394838 );
or ( n395897 , n395895 , n395896 );
buf ( n395898 , n394845 );
nand ( n74866 , n395897 , n395898 );
buf ( n395900 , n74866 );
buf ( n395901 , n395900 );
and ( n74869 , n74850 , n395901 );
and ( n74870 , n395873 , n395882 );
or ( n395904 , n74869 , n74870 );
buf ( n395905 , n395904 );
xor ( n395906 , n73901 , n394950 );
xor ( n74874 , n395906 , n394969 );
and ( n74875 , n395905 , n74874 );
buf ( n395909 , n57747 );
buf ( n395910 , n394724 );
and ( n395911 , n395909 , n395910 );
buf ( n395912 , n57754 );
buf ( n395913 , n394730 );
and ( n74881 , n395912 , n395913 );
nor ( n74882 , n395911 , n74881 );
buf ( n395916 , n74882 );
buf ( n395917 , n395916 );
buf ( n395918 , n384414 );
or ( n395919 , n395917 , n395918 );
buf ( n395920 , n74595 );
buf ( n395921 , n395635 );
or ( n74889 , n395920 , n395921 );
nand ( n395923 , n395919 , n74889 );
buf ( n395924 , n395923 );
buf ( n395925 , n395924 );
buf ( n395926 , n61992 );
buf ( n395927 , n380817 );
and ( n74895 , n395926 , n395927 );
buf ( n395929 , n382596 );
buf ( n395930 , n57983 );
and ( n74898 , n395929 , n395930 );
nor ( n395932 , n74895 , n74898 );
buf ( n395933 , n395932 );
buf ( n395934 , n395933 );
buf ( n395935 , n60313 );
or ( n395936 , n395934 , n395935 );
buf ( n395937 , n395606 );
buf ( n395938 , n380733 );
or ( n395939 , n395937 , n395938 );
nand ( n395940 , n395936 , n395939 );
buf ( n395941 , n395940 );
buf ( n395942 , n395941 );
xor ( n395943 , n395925 , n395942 );
not ( n74911 , n382655 );
not ( n395945 , n62243 );
not ( n74913 , n60171 );
or ( n74914 , n395945 , n74913 );
nand ( n74915 , n382835 , n380680 );
nand ( n74916 , n74914 , n74915 );
not ( n395950 , n74916 );
or ( n395951 , n74911 , n395950 );
or ( n395952 , n395578 , n384157 );
nand ( n74920 , n395951 , n395952 );
buf ( n395954 , n74920 );
and ( n395955 , n395943 , n395954 );
and ( n74923 , n395925 , n395942 );
or ( n74924 , n395955 , n74923 );
buf ( n395958 , n74924 );
xor ( n395959 , n73901 , n394950 );
xor ( n74927 , n395959 , n394969 );
and ( n395961 , n395958 , n74927 );
and ( n74929 , n395905 , n395958 );
or ( n74930 , n74875 , n395961 , n74929 );
xor ( n395964 , n395870 , n74930 );
xor ( n74932 , n395867 , n395964 );
and ( n395966 , n395865 , n74932 );
and ( n74934 , n395745 , n395864 );
or ( n74935 , n395966 , n74934 );
buf ( n74936 , n74935 );
xor ( n395970 , n394901 , n394917 );
xor ( n74938 , n395970 , n394972 );
and ( n395972 , n395870 , n74938 );
xor ( n395973 , n394901 , n394917 );
xor ( n74941 , n395973 , n394972 );
and ( n395975 , n74930 , n74941 );
and ( n395976 , n395870 , n74930 );
or ( n395977 , n395972 , n395975 , n395976 );
buf ( n395978 , n395977 );
xor ( n395979 , n74936 , n395978 );
xor ( n395980 , n394783 , n394786 );
xor ( n74948 , n395980 , n394876 );
xor ( n395982 , n395727 , n74701 );
xor ( n395983 , n74948 , n395982 );
buf ( n395984 , n395983 );
and ( n395985 , n395979 , n395984 );
and ( n395986 , n74936 , n395978 );
or ( n74954 , n395985 , n395986 );
buf ( n395988 , n74954 );
xor ( n395989 , n394980 , n394983 );
xor ( n74957 , n395989 , n73955 );
and ( n74958 , n395988 , n74957 );
and ( n395992 , n395739 , n395988 );
or ( n395993 , n395742 , n74958 , n395992 );
buf ( n395994 , n395993 );
xor ( n395995 , n395570 , n395994 );
not ( n395996 , n365108 );
buf ( n395997 , n386093 );
not ( n74965 , n395997 );
buf ( n395999 , n364900 );
not ( n74967 , n395999 );
or ( n74968 , n74965 , n74967 );
buf ( n396002 , n364975 );
not ( n396003 , n396002 );
buf ( n396004 , n396003 );
buf ( n396005 , n396004 );
buf ( n396006 , n352268 );
nand ( n74974 , n396005 , n396006 );
buf ( n396008 , n74974 );
buf ( n396009 , n396008 );
nand ( n396010 , n74968 , n396009 );
buf ( n396011 , n396010 );
not ( n396012 , n396011 );
or ( n396013 , n395996 , n396012 );
buf ( n74975 , n31093 );
not ( n74976 , n74975 );
buf ( n74977 , n74976 );
buf ( n396017 , n74977 );
not ( n396018 , n396017 );
buf ( n396019 , n396018 );
not ( n396020 , n396019 );
not ( n396021 , n396004 );
or ( n396022 , n396020 , n396021 );
buf ( n396023 , n364975 );
buf ( n396024 , n60751 );
nand ( n396025 , n396023 , n396024 );
buf ( n396026 , n396025 );
nand ( n396027 , n396022 , n396026 );
nand ( n396028 , n386091 , n396027 );
nand ( n396029 , n396013 , n396028 );
buf ( n396030 , n396029 );
and ( n396031 , n395995 , n396030 );
and ( n74978 , n395570 , n395994 );
or ( n74979 , n396031 , n74978 );
buf ( n396034 , n74979 );
buf ( n396035 , n396034 );
xor ( n396036 , n395565 , n396035 );
buf ( n396037 , n395038 );
not ( n396038 , n396037 );
buf ( n396039 , n366659 );
not ( n396040 , n396039 );
or ( n396041 , n396038 , n396040 );
buf ( n396042 , n375914 );
buf ( n74989 , n48458 );
nand ( n74990 , n396042 , n74989 );
buf ( n396045 , n74990 );
buf ( n396046 , n396045 );
nand ( n74993 , n396041 , n396046 );
buf ( n396048 , n74993 );
buf ( n396049 , n396048 );
not ( n396050 , n396049 );
buf ( n396051 , n375896 );
not ( n396052 , n396051 );
or ( n396053 , n396050 , n396052 );
buf ( n396054 , n394035 );
buf ( n396055 , n375920 );
nand ( n396056 , n396054 , n396055 );
buf ( n396057 , n396056 );
buf ( n396058 , n396057 );
nand ( n396059 , n396053 , n396058 );
buf ( n396060 , n396059 );
buf ( n396061 , n396060 );
and ( n396062 , n396036 , n396061 );
and ( n75009 , n395565 , n396035 );
or ( n75010 , n396062 , n75009 );
buf ( n396065 , n75010 );
buf ( n396066 , n396065 );
xor ( n75013 , n395532 , n396066 );
xor ( n396068 , n394021 , n394056 );
xor ( n75015 , n396068 , n394076 );
buf ( n396070 , n75015 );
buf ( n396071 , n396070 );
xor ( n396072 , n75013 , n396071 );
buf ( n396073 , n396072 );
buf ( n396074 , n396073 );
nand ( n396075 , n395494 , n396074 );
buf ( n396076 , n396075 );
buf ( n396077 , n396076 );
nand ( n396078 , n395489 , n396077 );
buf ( n396079 , n396078 );
buf ( n75026 , n396079 );
not ( n75027 , n75026 );
buf ( n75028 , n75027 );
buf ( n396083 , n75028 );
not ( n396084 , n396083 );
buf ( n396085 , n69397 );
buf ( n396086 , n379841 );
and ( n396087 , n396085 , n396086 );
buf ( n396088 , n374178 );
buf ( n396089 , n379847 );
and ( n396090 , n396088 , n396089 );
nor ( n75037 , n396087 , n396090 );
buf ( n75038 , n75037 );
buf ( n396093 , n75038 );
not ( n75040 , n396093 );
buf ( n396095 , n379893 );
not ( n75042 , n396095 );
and ( n396097 , n75040 , n75042 );
buf ( n396098 , n379841 );
not ( n396099 , n396098 );
buf ( n396100 , n41615 );
not ( n75045 , n396100 );
or ( n396102 , n396099 , n75045 );
buf ( n396103 , n41616 );
buf ( n396104 , n379847 );
nand ( n396105 , n396103 , n396104 );
buf ( n396106 , n396105 );
buf ( n396107 , n396106 );
nand ( n396108 , n396102 , n396107 );
buf ( n396109 , n396108 );
buf ( n396110 , n396109 );
buf ( n396111 , n379916 );
and ( n396112 , n396110 , n396111 );
nor ( n396113 , n396097 , n396112 );
buf ( n396114 , n396113 );
buf ( n396115 , n396114 );
not ( n396116 , n396115 );
or ( n396117 , n396084 , n396116 );
buf ( n396118 , n377353 );
not ( n75048 , n396118 );
buf ( n396120 , n381286 );
not ( n396121 , n396120 );
or ( n396122 , n75048 , n396121 );
buf ( n396123 , n22768 );
not ( n396124 , n396123 );
buf ( n396125 , n377352 );
nand ( n396126 , n396124 , n396125 );
buf ( n396127 , n396126 );
buf ( n396128 , n396127 );
nand ( n396129 , n396122 , n396128 );
buf ( n396130 , n396129 );
buf ( n396131 , n396130 );
not ( n396132 , n396131 );
buf ( n396133 , n363429 );
not ( n396134 , n396133 );
or ( n396135 , n396132 , n396134 );
buf ( n396136 , n390220 );
not ( n396137 , n396136 );
buf ( n396138 , n56970 );
not ( n396139 , n396138 );
buf ( n396140 , n342718 );
not ( n396141 , n396140 );
or ( n396142 , n396139 , n396141 );
buf ( n396143 , n386354 );
buf ( n396144 , n377389 );
nand ( n396145 , n396143 , n396144 );
buf ( n396146 , n396145 );
buf ( n396147 , n396146 );
nand ( n396148 , n396142 , n396147 );
buf ( n396149 , n396148 );
buf ( n396150 , n396149 );
nand ( n396151 , n396137 , n396150 );
buf ( n396152 , n396151 );
buf ( n396153 , n396152 );
nand ( n396154 , n396135 , n396153 );
buf ( n396155 , n396154 );
buf ( n396156 , n396155 );
buf ( n396157 , n44915 );
not ( n396158 , n396157 );
buf ( n396159 , n365041 );
not ( n75063 , n396159 );
buf ( n396161 , n365259 );
not ( n396162 , n396161 );
or ( n75066 , n75063 , n396162 );
buf ( n396164 , n386359 );
not ( n75068 , n396164 );
buf ( n396166 , n380497 );
nand ( n396167 , n75068 , n396166 );
buf ( n396168 , n396167 );
buf ( n396169 , n396168 );
nand ( n396170 , n75066 , n396169 );
buf ( n396171 , n396170 );
buf ( n396172 , n396171 );
not ( n396173 , n396172 );
or ( n396174 , n396158 , n396173 );
buf ( n396175 , n365041 );
not ( n75076 , n396175 );
buf ( n396177 , n377297 );
not ( n396178 , n396177 );
or ( n75079 , n75076 , n396178 );
buf ( n396180 , n377301 );
buf ( n396181 , n380497 );
nand ( n75082 , n396180 , n396181 );
buf ( n75083 , n75082 );
buf ( n396184 , n75083 );
nand ( n75085 , n75079 , n396184 );
buf ( n396186 , n75085 );
buf ( n396187 , n396186 );
buf ( n396188 , n47466 );
nand ( n75089 , n396187 , n396188 );
buf ( n75090 , n75089 );
buf ( n396191 , n75090 );
nand ( n75092 , n396174 , n396191 );
buf ( n396193 , n75092 );
buf ( n396194 , n396193 );
xor ( n396195 , n396156 , n396194 );
xor ( n75096 , n384470 , n384473 );
xor ( n396197 , n75096 , n63836 );
xor ( n396198 , n73678 , n73963 );
xor ( n75099 , n396197 , n396198 );
buf ( n396200 , n75099 );
buf ( n396201 , n365108 );
not ( n75102 , n396201 );
buf ( n396203 , n394014 );
not ( n396204 , n396203 );
or ( n396205 , n75102 , n396204 );
buf ( n396206 , n365021 );
buf ( n396207 , n396011 );
nand ( n396208 , n396206 , n396207 );
buf ( n396209 , n396208 );
buf ( n396210 , n396209 );
nand ( n396211 , n396205 , n396210 );
buf ( n396212 , n396211 );
buf ( n396213 , n396212 );
xor ( n396214 , n396200 , n396213 );
buf ( n396215 , n365242 );
not ( n396216 , n396215 );
buf ( n396217 , n394068 );
not ( n396218 , n396217 );
or ( n396219 , n396216 , n396218 );
buf ( n396220 , n65351 );
not ( n396221 , n396220 );
buf ( n396222 , n381220 );
not ( n396223 , n396222 );
or ( n396224 , n396221 , n396223 );
buf ( n396225 , n351195 );
buf ( n396226 , n386040 );
nand ( n396227 , n396225 , n396226 );
buf ( n75110 , n396227 );
buf ( n396229 , n75110 );
nand ( n75112 , n396224 , n396229 );
buf ( n396231 , n75112 );
buf ( n396232 , n396231 );
buf ( n396233 , n45055 );
nand ( n396234 , n396232 , n396233 );
buf ( n396235 , n396234 );
buf ( n396236 , n396235 );
nand ( n75118 , n396219 , n396236 );
buf ( n396238 , n75118 );
buf ( n396239 , n396238 );
xor ( n75121 , n396214 , n396239 );
buf ( n396241 , n75121 );
buf ( n396242 , n396241 );
buf ( n396243 , n365152 );
not ( n75125 , n396243 );
buf ( n396245 , n395524 );
not ( n75127 , n396245 );
or ( n396247 , n75125 , n75127 );
buf ( n396248 , n395497 );
not ( n396249 , n396248 );
buf ( n396250 , n375873 );
not ( n75132 , n396250 );
or ( n396252 , n396249 , n75132 );
buf ( n396253 , n382496 );
buf ( n396254 , n395497 );
or ( n396255 , n396253 , n396254 );
buf ( n396256 , n396255 );
buf ( n396257 , n396256 );
nand ( n396258 , n396252 , n396257 );
buf ( n396259 , n396258 );
buf ( n396260 , n396259 );
buf ( n396261 , n45014 );
nand ( n396262 , n396260 , n396261 );
buf ( n396263 , n396262 );
buf ( n396264 , n396263 );
nand ( n75146 , n396247 , n396264 );
buf ( n396266 , n75146 );
buf ( n396267 , n396266 );
xor ( n75149 , n396242 , n396267 );
buf ( n396269 , n49178 );
not ( n75151 , n396269 );
buf ( n396271 , n56849 );
not ( n396272 , n396271 );
or ( n75154 , n75151 , n396272 );
buf ( n396274 , n58073 );
not ( n75156 , n396274 );
buf ( n396276 , n369374 );
nand ( n396277 , n75156 , n396276 );
buf ( n396278 , n396277 );
buf ( n396279 , n396278 );
nand ( n396280 , n75154 , n396279 );
buf ( n396281 , n396280 );
buf ( n396282 , n396281 );
not ( n75164 , n396282 );
buf ( n396284 , n366399 );
not ( n396285 , n396284 );
or ( n396286 , n75164 , n396285 );
buf ( n396287 , n368994 );
not ( n396288 , n396287 );
not ( n396289 , n56849 );
buf ( n396290 , n396289 );
not ( n396291 , n396290 );
or ( n396292 , n396288 , n396291 );
buf ( n396293 , n386807 );
buf ( n396294 , n385238 );
nand ( n396295 , n396293 , n396294 );
buf ( n396296 , n396295 );
buf ( n396297 , n396296 );
nand ( n396298 , n396292 , n396297 );
buf ( n396299 , n396298 );
buf ( n396300 , n396299 );
buf ( n396301 , n377271 );
nand ( n396302 , n396300 , n396301 );
buf ( n396303 , n396302 );
buf ( n396304 , n396303 );
nand ( n396305 , n396286 , n396304 );
buf ( n396306 , n396305 );
buf ( n396307 , n396306 );
xor ( n396308 , n75149 , n396307 );
buf ( n396309 , n396308 );
buf ( n396310 , n396309 );
and ( n396311 , n396195 , n396310 );
and ( n75193 , n396156 , n396194 );
or ( n396313 , n396311 , n75193 );
buf ( n396314 , n396313 );
not ( n75196 , n396314 );
buf ( n75197 , n75196 );
not ( n75198 , n75197 );
not ( n396318 , n370050 );
and ( n75200 , n56687 , n367600 );
not ( n75201 , n56687 );
and ( n396321 , n75201 , n74077 );
or ( n396322 , n75200 , n396321 );
not ( n75204 , n396322 );
and ( n396324 , n396318 , n75204 );
buf ( n396325 , n379515 );
buf ( n396326 , n372230 );
and ( n396327 , n396325 , n396326 );
not ( n396328 , n396325 );
buf ( n396329 , n361026 );
and ( n396330 , n396328 , n396329 );
nor ( n75212 , n396327 , n396330 );
buf ( n396332 , n75212 );
nor ( n396333 , n396332 , n370060 );
nor ( n396334 , n396324 , n396333 );
buf ( n396335 , n396334 );
not ( n396336 , n396335 );
or ( n396337 , n75198 , n396336 );
buf ( n396338 , n377268 );
nor ( n396339 , n370984 , n50779 );
buf ( n396340 , n396339 );
xor ( n75222 , n56970 , n22707 );
buf ( n396342 , n75222 );
not ( n75224 , n396342 );
and ( n396344 , n396340 , n75224 );
buf ( n396345 , n396344 );
buf ( n396346 , n396345 );
and ( n75228 , n396338 , n396346 );
not ( n75229 , n396338 );
buf ( n396349 , n396281 );
and ( n75231 , n75229 , n396349 );
nor ( n75232 , n75228 , n75231 );
buf ( n396352 , n75232 );
buf ( n396353 , n396352 );
not ( n396354 , n396353 );
buf ( n396355 , n396354 );
buf ( n396356 , n396355 );
not ( n75238 , n396356 );
buf ( n396358 , n395038 );
not ( n396359 , n396358 );
buf ( n396360 , n366639 );
not ( n75242 , n396360 );
or ( n396362 , n396359 , n75242 );
buf ( n396363 , n342564 );
buf ( n396364 , n48458 );
nand ( n396365 , n396363 , n396364 );
buf ( n396366 , n396365 );
buf ( n396367 , n396366 );
nand ( n396368 , n396362 , n396367 );
buf ( n396369 , n396368 );
buf ( n396370 , n396369 );
not ( n396371 , n396370 );
buf ( n396372 , n45544 );
not ( n75254 , n396372 );
buf ( n75255 , n75254 );
buf ( n396375 , n75255 );
not ( n75257 , n396375 );
or ( n396377 , n396371 , n75257 );
buf ( n396378 , n365390 );
not ( n75260 , n396378 );
buf ( n396380 , n366639 );
not ( n75262 , n396380 );
or ( n396382 , n75260 , n75262 );
buf ( n75264 , n342564 );
buf ( n396384 , n365387 );
nand ( n396385 , n75264 , n396384 );
buf ( n396386 , n396385 );
buf ( n396387 , n396386 );
nand ( n396388 , n396382 , n396387 );
buf ( n396389 , n396388 );
buf ( n396390 , n396389 );
buf ( n396391 , n45491 );
nand ( n396392 , n396390 , n396391 );
buf ( n396393 , n396392 );
buf ( n396394 , n396393 );
nand ( n75276 , n396377 , n396394 );
buf ( n396396 , n75276 );
buf ( n396397 , n396396 );
not ( n75279 , n396397 );
buf ( n396399 , n365183 );
not ( n75281 , n396399 );
buf ( n396401 , n45050 );
buf ( n75283 , n396401 );
not ( n396403 , n75283 );
xor ( n75285 , n396403 , n351195 );
buf ( n75286 , n75285 );
not ( n75287 , n75286 );
or ( n75288 , n75281 , n75287 );
xor ( n396408 , n31193 , n396403 );
buf ( n396409 , n396408 );
buf ( n396410 , n365152 );
nand ( n396411 , n396409 , n396410 );
buf ( n396412 , n396411 );
buf ( n396413 , n396412 );
nand ( n396414 , n75288 , n396413 );
buf ( n396415 , n396414 );
buf ( n396416 , n396415 );
not ( n75298 , n396416 );
buf ( n396418 , n75298 );
buf ( n75300 , n396418 );
nand ( n75301 , n75279 , n75300 );
buf ( n75302 , n75301 );
xor ( n396422 , n74936 , n395978 );
xor ( n75304 , n396422 , n395984 );
buf ( n396424 , n75304 );
buf ( n396425 , n396424 );
not ( n75307 , n396425 );
not ( n75308 , n365224 );
buf ( n396428 , n65349 );
buf ( n396429 , n31093 );
and ( n396430 , n396428 , n396429 );
not ( n396431 , n396428 );
buf ( n396432 , n74977 );
and ( n75314 , n396431 , n396432 );
or ( n75315 , n396430 , n75314 );
buf ( n396435 , n75315 );
not ( n75317 , n396435 );
and ( n75318 , n75308 , n75317 );
not ( n396438 , n65349 );
not ( n396439 , n32234 );
or ( n75321 , n396438 , n396439 );
not ( n396441 , n386040 );
or ( n75323 , n32234 , n396441 );
nand ( n75324 , n75321 , n75323 );
and ( n396444 , n75324 , n365242 );
nor ( n75326 , n75318 , n396444 );
buf ( n75327 , n75326 );
nand ( n75328 , n75307 , n75327 );
buf ( n75329 , n75328 );
buf ( n396449 , n75329 );
xor ( n75331 , n73901 , n394950 );
xor ( n396451 , n75331 , n394969 );
xor ( n396452 , n395905 , n395958 );
xor ( n396453 , n396451 , n396452 );
buf ( n396454 , n396453 );
buf ( n396455 , n380651 );
buf ( n396456 , n384343 );
and ( n75338 , n396455 , n396456 );
buf ( n396458 , n380657 );
buf ( n396459 , n384089 );
and ( n75341 , n396458 , n396459 );
nor ( n396461 , n75338 , n75341 );
buf ( n396462 , n396461 );
buf ( n396463 , n396462 );
buf ( n396464 , n384354 );
or ( n396465 , n396463 , n396464 );
buf ( n396466 , n395757 );
buf ( n396467 , n384082 );
or ( n75349 , n396466 , n396467 );
nand ( n75350 , n396465 , n75349 );
buf ( n396470 , n75350 );
buf ( n396471 , n396470 );
not ( n75353 , n394832 );
not ( n396473 , n395894 );
not ( n396474 , n396473 );
or ( n75356 , n75353 , n396474 );
and ( n396476 , n376993 , n395890 );
not ( n396477 , n376993 );
and ( n75359 , n396477 , n394840 );
or ( n75360 , n396476 , n75359 );
not ( n396480 , n394838 );
nand ( n396481 , n75360 , n396480 );
nand ( n75363 , n75356 , n396481 );
buf ( n396483 , n75363 );
xor ( n75365 , n396471 , n396483 );
buf ( n396485 , n384380 );
buf ( n396486 , n57789 );
and ( n75368 , n396485 , n396486 );
buf ( n396488 , n384386 );
buf ( n396489 , n60054 );
and ( n396490 , n396488 , n396489 );
nor ( n75372 , n75368 , n396490 );
buf ( n396492 , n75372 );
or ( n396493 , n396492 , n380581 );
not ( n396494 , n394774 );
nand ( n75376 , n396494 , n74740 );
nand ( n396496 , n396493 , n75376 );
buf ( n396497 , n396496 );
or ( n75379 , n73773 , n73777 );
nand ( n396499 , n75379 , n394812 );
buf ( n396500 , n396499 );
buf ( n396501 , n57800 );
and ( n396502 , n396500 , n396501 );
buf ( n396503 , n394816 );
buf ( n396504 , n376903 );
and ( n75386 , n396503 , n396504 );
nor ( n396506 , n396502 , n75386 );
buf ( n396507 , n396506 );
buf ( n396508 , n396507 );
buf ( n396509 , n378341 );
or ( n396510 , n396508 , n396509 );
buf ( n396511 , n395783 );
buf ( n396512 , n378424 );
or ( n75394 , n396511 , n396512 );
nand ( n396514 , n396510 , n75394 );
buf ( n396515 , n396514 );
buf ( n396516 , n396515 );
xor ( n396517 , n396497 , n396516 );
buf ( n396518 , n380735 );
not ( n396519 , n396518 );
buf ( n396520 , n384054 );
buf ( n396521 , n57983 );
or ( n396522 , n396520 , n396521 );
buf ( n396523 , n63406 );
buf ( n396524 , n380817 );
or ( n75406 , n396523 , n396524 );
nand ( n396526 , n396522 , n75406 );
buf ( n396527 , n396526 );
buf ( n396528 , n396527 );
not ( n75410 , n396528 );
or ( n75411 , n396519 , n75410 );
buf ( n396531 , n382795 );
buf ( n396532 , n380817 );
and ( n75414 , n396531 , n396532 );
buf ( n396534 , n382803 );
buf ( n396535 , n63664 );
and ( n75417 , n396534 , n396535 );
nor ( n75418 , n75414 , n75417 );
buf ( n396538 , n75418 );
buf ( n396539 , n396538 );
buf ( n396540 , n380733 );
or ( n396541 , n396539 , n396540 );
nand ( n396542 , n75411 , n396541 );
buf ( n396543 , n396542 );
buf ( n396544 , n396543 );
and ( n396545 , n396517 , n396544 );
and ( n396546 , n396497 , n396516 );
or ( n396547 , n396545 , n396546 );
buf ( n396548 , n396547 );
buf ( n396549 , n396548 );
and ( n396550 , n75365 , n396549 );
and ( n396551 , n396471 , n396483 );
or ( n396552 , n396550 , n396551 );
buf ( n396553 , n396552 );
buf ( n396554 , n396553 );
xor ( n396555 , n395873 , n395882 );
xor ( n396556 , n396555 , n395901 );
buf ( n396557 , n396556 );
buf ( n396558 , n396557 );
xor ( n396559 , n396554 , n396558 );
buf ( n396560 , n396538 );
buf ( n396561 , n60313 );
or ( n396562 , n396560 , n396561 );
buf ( n396563 , n395933 );
buf ( n396564 , n380733 );
or ( n396565 , n396563 , n396564 );
nand ( n396566 , n396562 , n396565 );
buf ( n396567 , n396566 );
buf ( n396568 , n396567 );
buf ( n396569 , n382743 );
buf ( n396570 , n395810 );
and ( n396571 , n396569 , n396570 );
not ( n75433 , n396569 );
buf ( n396573 , n395816 );
and ( n396574 , n75433 , n396573 );
nor ( n75436 , n396571 , n396574 );
buf ( n396576 , n75436 );
buf ( n75438 , n396576 );
not ( n75439 , n75438 );
buf ( n396579 , n75439 );
buf ( n396580 , n396579 );
buf ( n396581 , n376924 );
or ( n75443 , n396580 , n396581 );
buf ( n396583 , n395837 );
buf ( n396584 , n56517 );
or ( n75446 , n396583 , n396584 );
nand ( n396586 , n75443 , n75446 );
buf ( n396587 , n396586 );
buf ( n75449 , n396587 );
and ( n396589 , n395801 , n56284 );
xor ( n75451 , n396589 , n56280 );
buf ( n396591 , n75451 );
buf ( n396592 , n376990 );
and ( n396593 , n396591 , n396592 );
buf ( n396594 , n75451 );
not ( n75456 , n396594 );
buf ( n396596 , n75456 );
buf ( n396597 , n396596 );
buf ( n396598 , n376997 );
and ( n396599 , n396597 , n396598 );
buf ( n396600 , n377003 );
nor ( n75462 , n396593 , n396599 , n396600 );
buf ( n396602 , n75462 );
buf ( n396603 , n396602 );
xor ( n396604 , n75449 , n396603 );
not ( n75466 , n56275 );
not ( n75467 , n56134 );
nand ( n396607 , n56271 , n75467 );
not ( n396608 , n396607 );
or ( n75470 , n75466 , n396608 );
nor ( n396610 , n376514 , n56278 );
not ( n396611 , n396610 );
nand ( n75473 , n75470 , n396611 );
and ( n396613 , n396610 , n56275 );
nand ( n396614 , n396607 , n396613 );
nand ( n396615 , n75473 , n396614 );
buf ( n396616 , n396615 );
buf ( n396617 , n376990 );
and ( n396618 , n396616 , n396617 );
buf ( n396619 , n396615 );
not ( n396620 , n396619 );
buf ( n396621 , n396620 );
buf ( n396622 , n396621 );
buf ( n396623 , n376997 );
and ( n396624 , n396622 , n396623 );
buf ( n396625 , n377003 );
nor ( n75487 , n396618 , n396624 , n396625 );
buf ( n396627 , n75487 );
buf ( n396628 , n396627 );
buf ( n396629 , n74791 );
not ( n396630 , n396629 );
buf ( n396631 , n396576 );
not ( n75493 , n396631 );
or ( n396633 , n396630 , n75493 );
buf ( n396634 , n75451 );
buf ( n396635 , n376866 );
and ( n396636 , n396634 , n396635 );
buf ( n396637 , n396596 );
buf ( n396638 , n382743 );
and ( n396639 , n396637 , n396638 );
nor ( n396640 , n396636 , n396639 );
buf ( n396641 , n396640 );
buf ( n396642 , n396641 );
buf ( n396643 , n376924 );
or ( n75505 , n396642 , n396643 );
nand ( n396645 , n396633 , n75505 );
buf ( n396646 , n396645 );
buf ( n396647 , n396646 );
and ( n75509 , n396628 , n396647 );
buf ( n396649 , n75509 );
buf ( n396650 , n396649 );
and ( n75512 , n396604 , n396650 );
and ( n75513 , n75449 , n396603 );
or ( n75514 , n75512 , n75513 );
buf ( n396654 , n75514 );
buf ( n396655 , n396654 );
xor ( n75517 , n396568 , n396655 );
buf ( n396657 , n384417 );
not ( n396658 , n396657 );
buf ( n396659 , n378372 );
buf ( n396660 , n394730 );
or ( n396661 , n396659 , n396660 );
buf ( n396662 , n378368 );
buf ( n396663 , n394724 );
or ( n396664 , n396662 , n396663 );
nand ( n396665 , n396661 , n396664 );
buf ( n396666 , n396665 );
buf ( n396667 , n396666 );
not ( n75529 , n396667 );
or ( n396669 , n396658 , n75529 );
buf ( n396670 , n395916 );
buf ( n396671 , n395635 );
or ( n396672 , n396670 , n396671 );
nand ( n396673 , n396669 , n396672 );
buf ( n396674 , n396673 );
buf ( n396675 , n396674 );
and ( n396676 , n75517 , n396675 );
and ( n75538 , n396568 , n396655 );
or ( n396678 , n396676 , n75538 );
buf ( n396679 , n396678 );
buf ( n396680 , n396679 );
and ( n396681 , n396559 , n396680 );
and ( n75543 , n396554 , n396558 );
or ( n75544 , n396681 , n75543 );
buf ( n396684 , n75544 );
buf ( n75546 , n396684 );
xor ( n75547 , n396454 , n75546 );
xor ( n396687 , n395586 , n395592 );
xor ( n396688 , n396687 , n395611 );
xor ( n75550 , n395853 , n395859 );
xor ( n396690 , n396688 , n75550 );
buf ( n396691 , n396690 );
and ( n396692 , n75547 , n396691 );
and ( n75554 , n396454 , n75546 );
or ( n396694 , n396692 , n75554 );
buf ( n396695 , n396694 );
xor ( n75557 , n395745 , n395864 );
xor ( n396697 , n75557 , n74932 );
and ( n75559 , n396695 , n396697 );
xor ( n396699 , n396628 , n396647 );
buf ( n396700 , n396699 );
buf ( n396701 , n74644 );
buf ( n396702 , n57800 );
and ( n396703 , n396701 , n396702 );
buf ( n396704 , n395683 );
buf ( n396705 , n378284 );
and ( n396706 , n396704 , n396705 );
nor ( n75568 , n396703 , n396706 );
buf ( n75569 , n75568 );
buf ( n396709 , n75569 );
buf ( n396710 , n378341 );
or ( n75572 , n396709 , n396710 );
buf ( n396712 , n396507 );
buf ( n396713 , n378424 );
or ( n75575 , n396712 , n396713 );
nand ( n396715 , n75572 , n75575 );
buf ( n396716 , n396715 );
xor ( n75578 , n396700 , n396716 );
buf ( n396718 , n380730 );
not ( n75580 , n396718 );
buf ( n396720 , n396527 );
not ( n396721 , n396720 );
or ( n75583 , n75580 , n396721 );
buf ( n396723 , n63549 );
buf ( n396724 , n380817 );
and ( n396725 , n396723 , n396724 );
buf ( n396726 , n384199 );
buf ( n396727 , n57983 );
and ( n396728 , n396726 , n396727 );
nor ( n75590 , n396725 , n396728 );
buf ( n396730 , n75590 );
buf ( n396731 , n396730 );
buf ( n396732 , n60313 );
or ( n75594 , n396731 , n396732 );
nand ( n75595 , n75583 , n75594 );
buf ( n396735 , n75595 );
and ( n75597 , n75578 , n396735 );
and ( n396737 , n396700 , n396716 );
or ( n75599 , n75597 , n396737 );
buf ( n396739 , n75599 );
not ( n396740 , n396480 );
buf ( n396741 , n57747 );
buf ( n396742 , n394840 );
and ( n396743 , n396741 , n396742 );
buf ( n75605 , n57754 );
buf ( n396745 , n395890 );
and ( n396746 , n75605 , n396745 );
nor ( n396747 , n396743 , n396746 );
buf ( n396748 , n396747 );
not ( n75610 , n396748 );
not ( n396750 , n75610 );
or ( n396751 , n396740 , n396750 );
nand ( n75613 , n75360 , n394832 );
nand ( n396753 , n396751 , n75613 );
buf ( n396754 , n396753 );
xor ( n396755 , n396739 , n396754 );
buf ( n396756 , n384085 );
not ( n396757 , n396756 );
not ( n75619 , n384089 );
not ( n75620 , n380680 );
or ( n396760 , n75619 , n75620 );
or ( n75622 , n380680 , n384089 );
nand ( n396762 , n396760 , n75622 );
buf ( n396763 , n396762 );
not ( n396764 , n396763 );
buf ( n396765 , n396764 );
buf ( n396766 , n396765 );
not ( n396767 , n396766 );
or ( n396768 , n396757 , n396767 );
buf ( n396769 , n396462 );
buf ( n396770 , n384082 );
or ( n75632 , n396769 , n396770 );
nand ( n75633 , n396768 , n75632 );
buf ( n396773 , n75633 );
buf ( n396774 , n396773 );
and ( n75636 , n396755 , n396774 );
and ( n396776 , n396739 , n396754 );
or ( n396777 , n75636 , n396776 );
buf ( n396778 , n396777 );
buf ( n396779 , n396778 );
buf ( n396780 , n61992 );
buf ( n396781 , n382835 );
and ( n396782 , n396780 , n396781 );
buf ( n396783 , n382596 );
buf ( n396784 , n62243 );
and ( n75646 , n396783 , n396784 );
nor ( n75647 , n396782 , n75646 );
buf ( n396787 , n75647 );
buf ( n396788 , n396787 );
buf ( n396789 , n382849 );
or ( n75651 , n396788 , n396789 );
buf ( n396791 , n380838 );
buf ( n396792 , n382835 );
and ( n75654 , n396791 , n396792 );
buf ( n396794 , n380844 );
buf ( n396795 , n62243 );
and ( n75657 , n396794 , n396795 );
nor ( n396797 , n75654 , n75657 );
buf ( n396798 , n396797 );
buf ( n396799 , n396798 );
buf ( n396800 , n384157 );
or ( n396801 , n396799 , n396800 );
nand ( n75663 , n75651 , n396801 );
buf ( n75664 , n75663 );
buf ( n396804 , n75664 );
xor ( n75666 , n75449 , n396603 );
xor ( n75667 , n75666 , n396650 );
buf ( n396807 , n75667 );
buf ( n396808 , n396807 );
xor ( n396809 , n396804 , n396808 );
buf ( n396810 , n384411 );
not ( n396811 , n396810 );
buf ( n396812 , n396666 );
not ( n75674 , n396812 );
or ( n396814 , n396811 , n75674 );
buf ( n396815 , n60089 );
buf ( n396816 , n394724 );
and ( n396817 , n396815 , n396816 );
buf ( n396818 , n60094 );
buf ( n396819 , n394730 );
and ( n396820 , n396818 , n396819 );
nor ( n75682 , n396817 , n396820 );
buf ( n75683 , n75682 );
buf ( n396823 , n75683 );
buf ( n396824 , n384414 );
or ( n396825 , n396823 , n396824 );
nand ( n75687 , n396814 , n396825 );
buf ( n396827 , n75687 );
buf ( n396828 , n396827 );
and ( n75690 , n396809 , n396828 );
and ( n396830 , n396804 , n396808 );
or ( n75692 , n75690 , n396830 );
buf ( n396832 , n75692 );
buf ( n396833 , n396832 );
xor ( n75695 , n396779 , n396833 );
xor ( n396835 , n396471 , n396483 );
xor ( n396836 , n396835 , n396549 );
buf ( n396837 , n396836 );
buf ( n396838 , n396837 );
and ( n75700 , n75695 , n396838 );
and ( n75701 , n396779 , n396833 );
or ( n396841 , n75700 , n75701 );
buf ( n396842 , n396841 );
xor ( n75704 , n396554 , n396558 );
xor ( n396844 , n75704 , n396680 );
buf ( n396845 , n396844 );
xor ( n75707 , n396842 , n396845 );
xor ( n396847 , n395749 , n395766 );
xor ( n396848 , n396847 , n395849 );
buf ( n396849 , n396848 );
buf ( n396850 , n396849 );
xor ( n396851 , n395925 , n395942 );
xor ( n75713 , n396851 , n395954 );
buf ( n396853 , n75713 );
buf ( n396854 , n396853 );
xor ( n75716 , n396850 , n396854 );
or ( n75717 , n396798 , n382849 );
not ( n396857 , n384157 );
nand ( n396858 , n396857 , n74916 );
nand ( n75720 , n75717 , n396858 );
xor ( n396860 , n395775 , n395799 );
xor ( n75722 , n396860 , n395845 );
and ( n75723 , n75720 , n75722 );
xor ( n75724 , n396568 , n396655 );
xor ( n75725 , n75724 , n396675 );
buf ( n75726 , n75725 );
xor ( n396866 , n395775 , n395799 );
xor ( n396867 , n396866 , n395845 );
and ( n75729 , n75726 , n396867 );
and ( n396869 , n75720 , n75726 );
or ( n396870 , n75723 , n75729 , n396869 );
buf ( n396871 , n396870 );
xor ( n75733 , n75716 , n396871 );
buf ( n396873 , n75733 );
and ( n396874 , n75707 , n396873 );
and ( n396875 , n396842 , n396845 );
or ( n75737 , n396874 , n396875 );
buf ( n396877 , n75737 );
xor ( n396878 , n396850 , n396854 );
and ( n75740 , n396878 , n396871 );
and ( n75741 , n396850 , n396854 );
or ( n396881 , n75740 , n75741 );
buf ( n396882 , n396881 );
buf ( n396883 , n396882 );
xor ( n75745 , n396877 , n396883 );
xor ( n396885 , n396454 , n75546 );
xor ( n75747 , n396885 , n396691 );
buf ( n396887 , n75747 );
buf ( n396888 , n396887 );
and ( n396889 , n75745 , n396888 );
and ( n396890 , n396877 , n396883 );
or ( n75752 , n396889 , n396890 );
buf ( n396892 , n75752 );
xor ( n396893 , n395745 , n395864 );
xor ( n396894 , n396893 , n74932 );
and ( n75756 , n396892 , n396894 );
and ( n396896 , n396695 , n396892 );
or ( n396897 , n75559 , n75756 , n396896 );
buf ( n396898 , n396897 );
and ( n75760 , n396449 , n396898 );
not ( n396900 , n396424 );
nor ( n396901 , n396900 , n75326 );
buf ( n396902 , n396901 );
nor ( n75764 , n75760 , n396902 );
buf ( n396904 , n75764 );
buf ( n396905 , n396904 );
not ( n75767 , n396905 );
buf ( n396907 , n75767 );
and ( n75769 , n75302 , n396907 );
and ( n75770 , n396415 , n396396 );
nor ( n75771 , n75769 , n75770 );
buf ( n396911 , n75771 );
not ( n75773 , n396911 );
buf ( n396913 , n75773 );
buf ( n396914 , n396913 );
not ( n396915 , n396914 );
or ( n396916 , n75238 , n396915 );
buf ( n396917 , n75771 );
not ( n396918 , n396917 );
buf ( n396919 , n396352 );
not ( n75781 , n396919 );
or ( n75782 , n396918 , n75781 );
buf ( n396922 , n396389 );
not ( n396923 , n396922 );
buf ( n396924 , n384501 );
not ( n75786 , n396924 );
or ( n396926 , n396923 , n75786 );
buf ( n396927 , n56794 );
buf ( n396928 , n395548 );
nand ( n75790 , n396927 , n396928 );
buf ( n75791 , n75790 );
buf ( n396931 , n75791 );
nand ( n396932 , n396926 , n396931 );
buf ( n396933 , n396932 );
buf ( n396934 , n396933 );
buf ( n396935 , n365242 );
not ( n75797 , n396935 );
buf ( n396937 , n396231 );
not ( n396938 , n396937 );
or ( n75800 , n75797 , n396938 );
buf ( n396940 , n394066 );
not ( n396941 , n396940 );
buf ( n396942 , n394004 );
not ( n75804 , n396942 );
or ( n396944 , n396941 , n75804 );
buf ( n396945 , n351160 );
buf ( n396946 , n394065 );
nand ( n75808 , n396945 , n396946 );
buf ( n396948 , n75808 );
buf ( n396949 , n396948 );
nand ( n75811 , n396944 , n396949 );
buf ( n396951 , n75811 );
buf ( n396952 , n396951 );
buf ( n396953 , n365226 );
nand ( n75815 , n396952 , n396953 );
buf ( n396955 , n75815 );
buf ( n396956 , n396955 );
nand ( n396957 , n75800 , n396956 );
buf ( n396958 , n396957 );
buf ( n396959 , n396958 );
xor ( n396960 , n396934 , n396959 );
xor ( n396961 , n395570 , n395994 );
xor ( n75823 , n396961 , n396030 );
buf ( n396963 , n75823 );
buf ( n396964 , n396963 );
xor ( n396965 , n396960 , n396964 );
buf ( n396966 , n396965 );
buf ( n396967 , n396966 );
nand ( n396968 , n75782 , n396967 );
buf ( n396969 , n396968 );
buf ( n396970 , n396969 );
nand ( n75832 , n396916 , n396970 );
buf ( n75833 , n75832 );
buf ( n396973 , n75833 );
buf ( n396974 , n377782 );
buf ( n396975 , n45592 );
and ( n396976 , n396974 , n396975 );
not ( n396977 , n396974 );
buf ( n396978 , n362420 );
and ( n396979 , n396977 , n396978 );
or ( n396980 , n396976 , n396979 );
buf ( n396981 , n396980 );
buf ( n396982 , n396981 );
buf ( n396983 , n362385 );
or ( n396984 , n396982 , n396983 );
buf ( n396985 , n377757 );
not ( n75847 , n396985 );
buf ( n396987 , n342335 );
not ( n396988 , n396987 );
or ( n396989 , n75847 , n396988 );
buf ( n396990 , n381336 );
buf ( n396991 , n378886 );
nand ( n396992 , n396990 , n396991 );
buf ( n396993 , n396992 );
buf ( n396994 , n396993 );
nand ( n75856 , n396989 , n396994 );
buf ( n396996 , n75856 );
buf ( n396997 , n396996 );
buf ( n396998 , n385243 );
buf ( n396999 , n362385 );
nand ( n397000 , n396997 , n396998 , n396999 );
buf ( n397001 , n397000 );
buf ( n397002 , n397001 );
nand ( n397003 , n396984 , n397002 );
buf ( n397004 , n397003 );
buf ( n397005 , n397004 );
xor ( n75867 , n396973 , n397005 );
buf ( n397007 , n368549 );
not ( n397008 , n397007 );
buf ( n397009 , n73159 );
not ( n75871 , n397009 );
or ( n397011 , n397008 , n75871 );
buf ( n397012 , n45113 );
buf ( n397013 , n380424 );
nand ( n397014 , n397012 , n397013 );
buf ( n397015 , n397014 );
buf ( n397016 , n397015 );
nand ( n75878 , n397011 , n397016 );
buf ( n75879 , n75878 );
buf ( n397019 , n75879 );
not ( n397020 , n397019 );
buf ( n397021 , n397020 );
buf ( n397022 , n397021 );
buf ( n397023 , n368605 );
or ( n397024 , n397022 , n397023 );
buf ( n397025 , n380424 );
buf ( n397026 , n351318 );
and ( n75888 , n397025 , n397026 );
not ( n397028 , n397025 );
buf ( n397029 , n364808 );
and ( n75891 , n397028 , n397029 );
or ( n75892 , n75888 , n75891 );
buf ( n397032 , n75892 );
buf ( n397033 , n397032 );
buf ( n397034 , n368624 );
or ( n75896 , n397033 , n397034 );
nand ( n397036 , n397024 , n75896 );
buf ( n397037 , n397036 );
buf ( n397038 , n397037 );
and ( n75900 , n75867 , n397038 );
and ( n397040 , n396973 , n397005 );
or ( n397041 , n75900 , n397040 );
buf ( n397042 , n397041 );
buf ( n75904 , n397042 );
nand ( n397044 , n396337 , n75904 );
buf ( n397045 , n397044 );
buf ( n397046 , n397045 );
not ( n397047 , n396334 );
buf ( n75909 , n397047 );
not ( n397049 , n75196 );
buf ( n397050 , n397049 );
nand ( n397051 , n75909 , n397050 );
buf ( n397052 , n397051 );
buf ( n397053 , n397052 );
nand ( n397054 , n397046 , n397053 );
buf ( n397055 , n397054 );
buf ( n397056 , n397055 );
nand ( n397057 , n396117 , n397056 );
buf ( n397058 , n397057 );
buf ( n397059 , n397058 );
buf ( n397060 , n396114 );
not ( n397061 , n397060 );
buf ( n397062 , n397061 );
buf ( n397063 , n397062 );
buf ( n397064 , n396079 );
nand ( n397065 , n397063 , n397064 );
buf ( n397066 , n397065 );
buf ( n397067 , n397066 );
nand ( n397068 , n397059 , n397067 );
buf ( n397069 , n397068 );
and ( n397070 , n74389 , n397069 );
and ( n397071 , n395418 , n395421 );
or ( n397072 , n397070 , n397071 );
buf ( n397073 , n397072 );
not ( n397074 , n397073 );
buf ( n397075 , n397074 );
buf ( n397076 , n397075 );
not ( n397077 , n397076 );
xor ( n75939 , n73172 , n394202 );
xor ( n75940 , n75939 , n394211 );
buf ( n397080 , n75940 );
buf ( n397081 , n397080 );
not ( n75943 , n397081 );
buf ( n397083 , n75943 );
buf ( n397084 , n397083 );
not ( n75946 , n397084 );
xor ( n75947 , n394318 , n394355 );
xor ( n397087 , n75947 , n394374 );
buf ( n397088 , n397087 );
buf ( n397089 , n397088 );
not ( n397090 , n397089 );
or ( n397091 , n75946 , n397090 );
buf ( n397092 , n397080 );
not ( n75954 , n397092 );
buf ( n397094 , n397088 );
not ( n397095 , n397094 );
buf ( n397096 , n397095 );
buf ( n397097 , n397096 );
not ( n397098 , n397097 );
or ( n75960 , n75954 , n397098 );
buf ( n397100 , n366317 );
buf ( n397101 , n395476 );
or ( n397102 , n397100 , n397101 );
not ( n75964 , n364744 );
not ( n397104 , n377779 );
and ( n397105 , n75964 , n397104 );
buf ( n397106 , n366329 );
buf ( n397107 , n377779 );
and ( n397108 , n397106 , n397107 );
buf ( n397109 , n397108 );
nor ( n75971 , n397105 , n397109 );
buf ( n75972 , n75971 );
buf ( n75973 , n49692 );
or ( n75974 , n75972 , n75973 );
nand ( n75975 , n397102 , n75974 );
buf ( n75976 , n75975 );
buf ( n397116 , n75976 );
buf ( n397117 , n366751 );
buf ( n397118 , n378098 );
and ( n75980 , n397117 , n397118 );
buf ( n75981 , n75980 );
buf ( n397121 , n75981 );
or ( n75983 , n397116 , n397121 );
xor ( n75984 , n395532 , n396066 );
and ( n75985 , n75984 , n396071 );
and ( n75986 , n395532 , n396066 );
or ( n75987 , n75985 , n75986 );
buf ( n397127 , n75987 );
buf ( n397128 , n397127 );
nand ( n397129 , n75983 , n397128 );
buf ( n397130 , n397129 );
buf ( n397131 , n397130 );
buf ( n397132 , n75976 );
buf ( n397133 , n75981 );
nand ( n397134 , n397132 , n397133 );
buf ( n397135 , n397134 );
buf ( n397136 , n397135 );
nand ( n75998 , n397131 , n397136 );
buf ( n397138 , n75998 );
buf ( n397139 , n397138 );
nand ( n76001 , n75960 , n397139 );
buf ( n397141 , n76001 );
buf ( n397142 , n397141 );
nand ( n76004 , n397091 , n397142 );
buf ( n397144 , n76004 );
buf ( n397145 , n397144 );
not ( n76007 , n397145 );
xor ( n397147 , n384518 , n384543 );
xor ( n76009 , n397147 , n384570 );
buf ( n397149 , n76009 );
not ( n76011 , n397149 );
buf ( n397151 , n365152 );
not ( n76013 , n397151 );
buf ( n397153 , n383680 );
not ( n76015 , n397153 );
or ( n397155 , n76013 , n76015 );
buf ( n397156 , n394178 );
buf ( n397157 , n45015 );
nand ( n397158 , n397156 , n397157 );
buf ( n397159 , n397158 );
buf ( n397160 , n397159 );
nand ( n76022 , n397155 , n397160 );
buf ( n76023 , n76022 );
buf ( n397163 , n76023 );
not ( n397164 , n397163 );
buf ( n397165 , n397164 );
not ( n397166 , n397165 );
and ( n397167 , n76011 , n397166 );
and ( n76029 , n397149 , n397165 );
nor ( n76030 , n397167 , n76029 );
not ( n397170 , n394332 );
not ( n397171 , n47466 );
or ( n76033 , n397170 , n397171 );
buf ( n76034 , n365076 );
or ( n397174 , n383699 , n76034 );
nand ( n397175 , n76033 , n397174 );
not ( n397176 , n397175 );
and ( n397177 , n76030 , n397176 );
not ( n76039 , n76030 );
and ( n76040 , n76039 , n397175 );
nor ( n397180 , n397177 , n76040 );
not ( n76042 , n397180 );
not ( n76043 , n76042 );
buf ( n397183 , n57530 );
not ( n397184 , n397183 );
buf ( n397185 , n393866 );
not ( n397186 , n397185 );
or ( n397187 , n397184 , n397186 );
buf ( n397188 , n395304 );
not ( n76050 , n57147 );
buf ( n397190 , n76050 );
buf ( n397191 , n397190 );
nand ( n76053 , n397188 , n397191 );
buf ( n397193 , n76053 );
buf ( n397194 , n397193 );
nand ( n397195 , n397187 , n397194 );
buf ( n397196 , n397195 );
not ( n397197 , n397196 );
not ( n397198 , n369804 );
not ( n76060 , n395222 );
or ( n397200 , n397198 , n76060 );
buf ( n397201 , n393883 );
buf ( n397202 , n362537 );
and ( n397203 , n397201 , n397202 );
not ( n76065 , n397201 );
buf ( n397205 , n389807 );
and ( n397206 , n76065 , n397205 );
nor ( n397207 , n397203 , n397206 );
buf ( n397208 , n397207 );
or ( n397209 , n397208 , n369813 );
nand ( n76071 , n397200 , n397209 );
not ( n397211 , n76071 );
or ( n397212 , n397197 , n397211 );
or ( n76074 , n76071 , n397196 );
nand ( n76075 , n397212 , n76074 );
not ( n397215 , n76075 );
or ( n397216 , n76043 , n397215 );
or ( n76078 , n76075 , n76042 );
nand ( n397218 , n397216 , n76078 );
buf ( n397219 , n397218 );
not ( n76081 , n397219 );
or ( n76082 , n76007 , n76081 );
buf ( n397222 , n397218 );
buf ( n397223 , n397144 );
or ( n76085 , n397222 , n397223 );
nand ( n397225 , n76082 , n76085 );
buf ( n397226 , n397225 );
buf ( n397227 , n397226 );
not ( n76089 , n397227 );
buf ( n397229 , n57530 );
not ( n397230 , n397229 );
and ( n397231 , n377592 , n352119 );
not ( n397232 , n377592 );
and ( n76094 , n397232 , n32087 );
nor ( n397234 , n397231 , n76094 );
buf ( n397235 , n397234 );
not ( n76097 , n397235 );
or ( n76098 , n397230 , n76097 );
buf ( n397238 , n72861 );
buf ( n397239 , n397190 );
nand ( n76101 , n397238 , n397239 );
buf ( n397241 , n76101 );
buf ( n397242 , n397241 );
nand ( n397243 , n76098 , n397242 );
buf ( n397244 , n397243 );
buf ( n397245 , n397244 );
and ( n76107 , n361625 , n395075 );
not ( n397247 , n361625 );
buf ( n397248 , n377122 );
not ( n76110 , n397248 );
buf ( n397250 , n44717 );
not ( n76112 , n397250 );
or ( n397252 , n76110 , n76112 );
buf ( n397253 , n45908 );
buf ( n397254 , n57463 );
nand ( n397255 , n397253 , n397254 );
buf ( n397256 , n397255 );
buf ( n397257 , n397256 );
nand ( n397258 , n397252 , n397257 );
buf ( n397259 , n397258 );
nand ( n397260 , n397259 , n381426 );
and ( n397261 , n397247 , n397260 );
nor ( n76123 , n76107 , n397261 );
buf ( n397263 , n76123 );
or ( n397264 , n397245 , n397263 );
buf ( n397265 , n396149 );
not ( n76127 , n397265 );
buf ( n397267 , n363429 );
not ( n397268 , n397267 );
or ( n397269 , n76127 , n397268 );
buf ( n397270 , n369374 );
not ( n76132 , n397270 );
buf ( n397272 , n342718 );
not ( n397273 , n397272 );
or ( n76135 , n76132 , n397273 );
buf ( n397275 , n386354 );
buf ( n397276 , n49178 );
nand ( n397277 , n397275 , n397276 );
buf ( n397278 , n397277 );
buf ( n397279 , n397278 );
nand ( n76141 , n76135 , n397279 );
buf ( n397281 , n76141 );
buf ( n397282 , n397281 );
buf ( n397283 , n58231 );
nand ( n397284 , n397282 , n397283 );
buf ( n397285 , n397284 );
buf ( n397286 , n397285 );
nand ( n76148 , n397269 , n397286 );
buf ( n397288 , n76148 );
buf ( n397289 , n397288 );
not ( n76151 , n397289 );
xor ( n76152 , n396200 , n396213 );
and ( n397292 , n76152 , n396239 );
and ( n76154 , n396200 , n396213 );
or ( n76155 , n397292 , n76154 );
buf ( n397295 , n76155 );
buf ( n397296 , n397295 );
xor ( n76158 , n394553 , n395002 );
xor ( n76159 , n76158 , n395028 );
buf ( n397299 , n76159 );
buf ( n397300 , n397299 );
xor ( n76162 , n397296 , n397300 );
buf ( n397302 , n396299 );
not ( n76164 , n397302 );
buf ( n397304 , n366399 );
not ( n76166 , n397304 );
or ( n76167 , n76164 , n76166 );
buf ( n397307 , n395046 );
buf ( n397308 , n377168 );
or ( n397309 , n397307 , n397308 );
buf ( n397310 , n397309 );
buf ( n397311 , n397310 );
nand ( n397312 , n76167 , n397311 );
buf ( n397313 , n397312 );
buf ( n397314 , n397313 );
xnor ( n397315 , n76162 , n397314 );
buf ( n397316 , n397315 );
buf ( n397317 , n397316 );
not ( n397318 , n397317 );
buf ( n397319 , n397318 );
buf ( n397320 , n397319 );
not ( n397321 , n397320 );
or ( n397322 , n76151 , n397321 );
buf ( n397323 , n397288 );
not ( n397324 , n397323 );
buf ( n397325 , n397324 );
buf ( n397326 , n397325 );
not ( n76188 , n397326 );
buf ( n397328 , n397316 );
not ( n76190 , n397328 );
or ( n397330 , n76188 , n76190 );
xor ( n76192 , n396242 , n396267 );
and ( n397332 , n76192 , n396307 );
and ( n76194 , n396242 , n396267 );
or ( n397334 , n397332 , n76194 );
buf ( n397335 , n397334 );
buf ( n397336 , n397335 );
nand ( n397337 , n397330 , n397336 );
buf ( n397338 , n397337 );
buf ( n397339 , n397338 );
nand ( n397340 , n397322 , n397339 );
buf ( n397341 , n397340 );
buf ( n397342 , n397341 );
nand ( n397343 , n397264 , n397342 );
buf ( n397344 , n397343 );
buf ( n397345 , n397344 );
buf ( n397346 , n397244 );
buf ( n397347 , n76123 );
nand ( n76209 , n397346 , n397347 );
buf ( n397349 , n76209 );
buf ( n76211 , n397349 );
nand ( n76212 , n397345 , n76211 );
buf ( n76213 , n76212 );
buf ( n397353 , n76213 );
not ( n76215 , n397353 );
buf ( n397355 , n379274 );
not ( n397356 , n397355 );
buf ( n397357 , n361751 );
not ( n397358 , n397357 );
or ( n397359 , n397356 , n397358 );
buf ( n397360 , n41946 );
buf ( n397361 , n379271 );
nand ( n76223 , n397360 , n397361 );
buf ( n397363 , n76223 );
buf ( n397364 , n397363 );
nand ( n76226 , n397359 , n397364 );
buf ( n397366 , n76226 );
buf ( n397367 , n397366 );
buf ( n397368 , n379263 );
and ( n76230 , n397367 , n397368 );
buf ( n397370 , n379274 );
not ( n76232 , n397370 );
buf ( n397372 , n377961 );
not ( n397373 , n397372 );
or ( n76235 , n76232 , n397373 );
buf ( n397375 , n41528 );
buf ( n397376 , n379271 );
nand ( n76238 , n397375 , n397376 );
buf ( n397378 , n76238 );
buf ( n397379 , n397378 );
nand ( n76241 , n76235 , n397379 );
buf ( n76242 , n76241 );
buf ( n397382 , n76242 );
not ( n76244 , n397382 );
buf ( n397384 , n379296 );
nor ( n397385 , n76244 , n397384 );
buf ( n397386 , n397385 );
buf ( n397387 , n397386 );
nor ( n397388 , n76230 , n397387 );
buf ( n397389 , n397388 );
buf ( n397390 , n397389 );
not ( n397391 , n397390 );
buf ( n397392 , n397391 );
buf ( n397393 , n397392 );
not ( n76255 , n397393 );
or ( n76256 , n76215 , n76255 );
buf ( n397396 , n76213 );
not ( n397397 , n397396 );
buf ( n397398 , n397397 );
buf ( n397399 , n397398 );
not ( n76261 , n397399 );
buf ( n397401 , n397389 );
not ( n76263 , n397401 );
or ( n76264 , n76261 , n76263 );
buf ( n397404 , n394161 );
buf ( n397405 , n365155 );
or ( n76267 , n397404 , n397405 );
buf ( n397407 , n395509 );
buf ( n397408 , n45014 );
nand ( n76270 , n397407 , n397408 );
buf ( n397410 , n76270 );
buf ( n397411 , n397410 );
nand ( n397412 , n76267 , n397411 );
buf ( n397413 , n397412 );
buf ( n397414 , n397413 );
buf ( n397415 , n397281 );
not ( n397416 , n397415 );
buf ( n397417 , n363429 );
not ( n397418 , n397417 );
or ( n397419 , n397416 , n397418 );
buf ( n397420 , n395194 );
buf ( n397421 , n58231 );
nand ( n397422 , n397420 , n397421 );
buf ( n397423 , n397422 );
buf ( n397424 , n397423 );
nand ( n76273 , n397419 , n397424 );
buf ( n397426 , n76273 );
buf ( n397427 , n397426 );
xor ( n397428 , n397414 , n397427 );
buf ( n397429 , n397295 );
not ( n397430 , n397429 );
buf ( n397431 , n397313 );
not ( n397432 , n397431 );
or ( n397433 , n397430 , n397432 );
buf ( n397434 , n397313 );
buf ( n397435 , n397295 );
or ( n397436 , n397434 , n397435 );
buf ( n397437 , n397299 );
nand ( n397438 , n397436 , n397437 );
buf ( n397439 , n397438 );
buf ( n397440 , n397439 );
nand ( n397441 , n397433 , n397440 );
buf ( n397442 , n397441 );
buf ( n397443 , n397442 );
xor ( n397444 , n397428 , n397443 );
buf ( n397445 , n397444 );
buf ( n397446 , n397445 );
buf ( n397447 , n395443 );
not ( n397448 , n397447 );
buf ( n397449 , n397448 );
buf ( n397450 , n397449 );
not ( n397451 , n397450 );
buf ( n397452 , n362027 );
not ( n397453 , n397452 );
or ( n397454 , n397451 , n397453 );
buf ( n397455 , n371063 );
buf ( n397456 , n395246 );
nand ( n397457 , n397455 , n397456 );
buf ( n397458 , n397457 );
buf ( n397459 , n397458 );
nand ( n397460 , n397454 , n397459 );
buf ( n397461 , n397460 );
buf ( n397462 , n397461 );
xor ( n76290 , n397446 , n397462 );
buf ( n76291 , n396322 );
not ( n76292 , n76291 );
buf ( n397466 , n76292 );
buf ( n397467 , n397466 );
not ( n397468 , n397467 );
buf ( n397469 , n361019 );
not ( n76297 , n397469 );
or ( n397471 , n397468 , n76297 );
buf ( n397472 , n361060 );
buf ( n397473 , n395117 );
nand ( n397474 , n397472 , n397473 );
buf ( n397475 , n397474 );
buf ( n397476 , n397475 );
nand ( n76304 , n397471 , n397476 );
buf ( n397478 , n76304 );
buf ( n397479 , n397478 );
and ( n397480 , n76290 , n397479 );
and ( n397481 , n397446 , n397462 );
or ( n76309 , n397480 , n397481 );
buf ( n397483 , n76309 );
buf ( n397484 , n397483 );
nand ( n76312 , n76264 , n397484 );
buf ( n397486 , n76312 );
buf ( n397487 , n397486 );
nand ( n397488 , n76256 , n397487 );
buf ( n397489 , n397488 );
buf ( n397490 , n397489 );
not ( n397491 , n397490 );
buf ( n397492 , n397491 );
buf ( n397493 , n397492 );
not ( n397494 , n397493 );
and ( n397495 , n76089 , n397494 );
buf ( n397496 , n397492 );
buf ( n397497 , n397226 );
and ( n397498 , n397496 , n397497 );
nor ( n76326 , n397495 , n397498 );
buf ( n397500 , n76326 );
buf ( n397501 , n397500 );
not ( n76329 , n397501 );
or ( n397503 , n397077 , n76329 );
xor ( n397504 , n72909 , n393956 );
and ( n76332 , n397504 , n394083 );
not ( n397506 , n397504 );
not ( n397507 , n394083 );
and ( n76335 , n397506 , n397507 );
nor ( n397509 , n76332 , n76335 );
buf ( n397510 , n397509 );
not ( n76338 , n397510 );
buf ( n397512 , n397127 );
buf ( n397513 , n75981 );
xor ( n76341 , n397512 , n397513 );
buf ( n397515 , n75976 );
xnor ( n76343 , n76341 , n397515 );
buf ( n397517 , n76343 );
buf ( n397518 , n397517 );
not ( n76346 , n397518 );
buf ( n76347 , n76346 );
buf ( n397521 , n76347 );
not ( n397522 , n397521 );
or ( n76350 , n76338 , n397522 );
not ( n397524 , n397509 );
not ( n76352 , n397524 );
not ( n397526 , n397517 );
or ( n397527 , n76352 , n397526 );
buf ( n397528 , n387542 );
not ( n397529 , n397528 );
buf ( n397530 , n393934 );
not ( n76358 , n397530 );
or ( n76359 , n397529 , n76358 );
buf ( n397533 , n397032 );
not ( n397534 , n397533 );
buf ( n76362 , n368608 );
nand ( n76363 , n397534 , n76362 );
buf ( n397537 , n76363 );
buf ( n397538 , n397537 );
nand ( n397539 , n76359 , n397538 );
buf ( n397540 , n397539 );
buf ( n397541 , n397540 );
not ( n397542 , n397541 );
buf ( n397543 , n40852 );
not ( n397544 , n397543 );
buf ( n397545 , n44634 );
not ( n76372 , n397545 );
or ( n76373 , n397544 , n76372 );
buf ( n397548 , n378098 );
nand ( n397549 , n76373 , n397548 );
buf ( n397550 , n397549 );
not ( n76377 , n40852 );
nand ( n76378 , n76377 , n45455 );
nand ( n397553 , n397550 , n76378 , n45855 );
buf ( n397554 , n397553 );
not ( n76381 , n397554 );
buf ( n76382 , n76381 );
buf ( n397557 , n76382 );
not ( n76384 , n397557 );
or ( n397559 , n397542 , n76384 );
buf ( n397560 , n397540 );
not ( n397561 , n397560 );
buf ( n397562 , n397561 );
buf ( n397563 , n397562 );
not ( n76390 , n397563 );
buf ( n397565 , n397553 );
not ( n397566 , n397565 );
or ( n76393 , n76390 , n397566 );
xor ( n397568 , n396934 , n396959 );
and ( n397569 , n397568 , n396964 );
and ( n76396 , n396934 , n396959 );
or ( n397571 , n397569 , n76396 );
buf ( n397572 , n397571 );
buf ( n397573 , n397572 );
xor ( n397574 , n395565 , n396035 );
xor ( n397575 , n397574 , n396061 );
buf ( n397576 , n397575 );
buf ( n397577 , n397576 );
xor ( n397578 , n397573 , n397577 );
xor ( n397579 , n394980 , n394983 );
xor ( n76406 , n397579 , n73955 );
xor ( n397581 , n395739 , n395988 );
xor ( n76408 , n76406 , n397581 );
buf ( n397583 , n76408 );
buf ( n397584 , n351345 );
not ( n76411 , n397584 );
buf ( n397586 , n396004 );
not ( n397587 , n397586 );
or ( n397588 , n76411 , n397587 );
buf ( n76415 , n364975 );
buf ( n397590 , n76415 );
buf ( n397591 , n394044 );
nand ( n397592 , n397590 , n397591 );
buf ( n397593 , n397592 );
buf ( n397594 , n397593 );
nand ( n397595 , n397588 , n397594 );
buf ( n397596 , n397595 );
buf ( n397597 , n397596 );
not ( n397598 , n397597 );
buf ( n397599 , n365021 );
not ( n76426 , n397599 );
or ( n397601 , n397598 , n76426 );
buf ( n397602 , n396027 );
buf ( n397603 , n365108 );
nand ( n76430 , n397602 , n397603 );
buf ( n397605 , n76430 );
buf ( n397606 , n397605 );
nand ( n76433 , n397601 , n397606 );
buf ( n76434 , n76433 );
buf ( n397609 , n76434 );
xor ( n76436 , n397583 , n397609 );
buf ( n397611 , n365242 );
not ( n397612 , n397611 );
buf ( n397613 , n396951 );
not ( n76440 , n397613 );
or ( n397615 , n397612 , n76440 );
buf ( n397616 , n45055 );
buf ( n397617 , n75324 );
nand ( n397618 , n397616 , n397617 );
buf ( n397619 , n397618 );
buf ( n397620 , n397619 );
nand ( n76447 , n397615 , n397620 );
buf ( n397622 , n76447 );
buf ( n397623 , n397622 );
and ( n397624 , n76436 , n397623 );
and ( n76451 , n397583 , n397609 );
or ( n397626 , n397624 , n76451 );
buf ( n397627 , n397626 );
buf ( n397628 , n397627 );
buf ( n397629 , n365152 );
not ( n397630 , n397629 );
buf ( n397631 , n396259 );
not ( n76458 , n397631 );
or ( n397633 , n397630 , n76458 );
buf ( n397634 , n396408 );
buf ( n397635 , n45014 );
nand ( n397636 , n397634 , n397635 );
buf ( n397637 , n397636 );
buf ( n397638 , n397637 );
nand ( n397639 , n397633 , n397638 );
buf ( n397640 , n397639 );
buf ( n397641 , n397640 );
xor ( n76468 , n397628 , n397641 );
buf ( n397643 , n368994 );
not ( n76470 , n397643 );
buf ( n397645 , n377279 );
not ( n76472 , n397645 );
or ( n76473 , n76470 , n76472 );
buf ( n397648 , n378135 );
buf ( n397649 , n385238 );
nand ( n76476 , n397648 , n397649 );
buf ( n76477 , n76476 );
buf ( n397652 , n76477 );
nand ( n76479 , n76473 , n397652 );
buf ( n397654 , n76479 );
buf ( n397655 , n397654 );
not ( n397656 , n397655 );
buf ( n397657 , n375896 );
not ( n397658 , n397657 );
or ( n397659 , n397656 , n397658 );
buf ( n397660 , n396048 );
buf ( n397661 , n375920 );
nand ( n397662 , n397660 , n397661 );
buf ( n397663 , n397662 );
buf ( n397664 , n397663 );
nand ( n397665 , n397659 , n397664 );
buf ( n397666 , n397665 );
buf ( n397667 , n397666 );
and ( n397668 , n76468 , n397667 );
and ( n397669 , n397628 , n397641 );
or ( n397670 , n397668 , n397669 );
buf ( n397671 , n397670 );
buf ( n397672 , n397671 );
and ( n397673 , n397578 , n397672 );
and ( n397674 , n397573 , n397577 );
or ( n397675 , n397673 , n397674 );
buf ( n397676 , n397675 );
buf ( n397677 , n397676 );
nand ( n397678 , n76393 , n397677 );
buf ( n397679 , n397678 );
buf ( n397680 , n397679 );
nand ( n397681 , n397559 , n397680 );
buf ( n76482 , n397681 );
nand ( n397683 , n397527 , n76482 );
buf ( n397684 , n397683 );
nand ( n397685 , n76350 , n397684 );
buf ( n397686 , n397685 );
buf ( n397687 , n397686 );
not ( n76488 , n397687 );
buf ( n397689 , n76488 );
buf ( n397690 , n397088 );
buf ( n397691 , n397083 );
and ( n397692 , n397690 , n397691 );
not ( n76493 , n397690 );
buf ( n397694 , n397080 );
and ( n397695 , n76493 , n397694 );
nor ( n76496 , n397692 , n397695 );
buf ( n76497 , n76496 );
and ( n397698 , n76497 , n397138 );
not ( n76499 , n76497 );
buf ( n397700 , n397138 );
not ( n397701 , n397700 );
buf ( n397702 , n397701 );
and ( n397703 , n76499 , n397702 );
nor ( n397704 , n397698 , n397703 );
not ( n397705 , n397704 );
nand ( n76506 , n397689 , n397705 );
buf ( n397707 , n76506 );
not ( n76508 , n397707 );
buf ( n397709 , n76213 );
buf ( n397710 , n397389 );
xor ( n397711 , n397709 , n397710 );
buf ( n397712 , n397483 );
xor ( n397713 , n397711 , n397712 );
buf ( n397714 , n397713 );
buf ( n397715 , n397714 );
not ( n76516 , n397715 );
buf ( n76517 , n76516 );
buf ( n397718 , n76517 );
not ( n76519 , n397718 );
or ( n397720 , n76508 , n76519 );
not ( n397721 , n397689 );
nand ( n76522 , n397721 , n397704 );
buf ( n397723 , n76522 );
nand ( n397724 , n397720 , n397723 );
buf ( n397725 , n397724 );
buf ( n397726 , n397725 );
nand ( n76527 , n397503 , n397726 );
buf ( n397728 , n76527 );
buf ( n397729 , n397728 );
buf ( n397730 , n397500 );
not ( n397731 , n397730 );
buf ( n397732 , n397731 );
buf ( n397733 , n397732 );
buf ( n397734 , n397072 );
nand ( n76535 , n397733 , n397734 );
buf ( n397736 , n76535 );
buf ( n76537 , n397736 );
nand ( n76538 , n397729 , n76537 );
buf ( n76539 , n76538 );
buf ( n76540 , n76539 );
nand ( n76541 , n395394 , n76540 );
buf ( n76542 , n76541 );
buf ( n76543 , n76542 );
buf ( n397744 , n395287 );
buf ( n397745 , n395392 );
nand ( n397746 , n397744 , n397745 );
buf ( n397747 , n397746 );
buf ( n397748 , n397747 );
nand ( n397749 , n76543 , n397748 );
buf ( n397750 , n397749 );
buf ( n397751 , n397750 );
not ( n76552 , n397180 );
or ( n76553 , n397196 , n76071 );
not ( n76554 , n76553 );
or ( n76555 , n76552 , n76554 );
nand ( n397756 , n397196 , n76071 );
nand ( n76557 , n76555 , n397756 );
buf ( n397758 , n76557 );
buf ( n397759 , n379263 );
not ( n397760 , n397759 );
buf ( n397761 , n379274 );
not ( n397762 , n397761 );
buf ( n397763 , n367116 );
not ( n76564 , n397763 );
or ( n397765 , n397762 , n76564 );
buf ( n397766 , n362148 );
buf ( n397767 , n379271 );
nand ( n76568 , n397766 , n397767 );
buf ( n397769 , n76568 );
buf ( n397770 , n397769 );
nand ( n397771 , n397765 , n397770 );
buf ( n397772 , n397771 );
buf ( n397773 , n397772 );
not ( n76574 , n397773 );
or ( n397775 , n397760 , n76574 );
buf ( n397776 , n379274 );
not ( n76577 , n397776 );
buf ( n397778 , n41666 );
not ( n397779 , n397778 );
or ( n76580 , n76577 , n397779 );
buf ( n397781 , n41663 );
buf ( n397782 , n379271 );
nand ( n76583 , n397781 , n397782 );
buf ( n76584 , n76583 );
buf ( n397785 , n76584 );
nand ( n76586 , n76580 , n397785 );
buf ( n397787 , n76586 );
buf ( n397788 , n397787 );
buf ( n397789 , n379299 );
nand ( n76590 , n397788 , n397789 );
buf ( n397791 , n76590 );
buf ( n397792 , n397791 );
nand ( n76593 , n397775 , n397792 );
buf ( n397794 , n76593 );
buf ( n397795 , n397794 );
xor ( n76596 , n397758 , n397795 );
xor ( n76597 , n394312 , n394379 );
and ( n397798 , n76597 , n394405 );
and ( n76599 , n394312 , n394379 );
or ( n397800 , n397798 , n76599 );
buf ( n397801 , n397800 );
buf ( n397802 , n397801 );
xor ( n397803 , n76596 , n397802 );
buf ( n397804 , n397803 );
buf ( n397805 , n397804 );
buf ( n397806 , n76023 );
not ( n397807 , n397806 );
buf ( n397808 , n397175 );
not ( n397809 , n397808 );
or ( n76610 , n397807 , n397809 );
not ( n397811 , n397176 );
not ( n76612 , n397165 );
or ( n397813 , n397811 , n76612 );
nand ( n76614 , n397813 , n397149 );
buf ( n397815 , n76614 );
nand ( n397816 , n76610 , n397815 );
buf ( n397817 , n397816 );
buf ( n397818 , n385223 );
buf ( n397819 , n385245 );
xor ( n397820 , n397818 , n397819 );
buf ( n397821 , n385264 );
xor ( n397822 , n397820 , n397821 );
buf ( n397823 , n397822 );
xor ( n397824 , n397817 , n397823 );
buf ( n397825 , n73364 );
not ( n397826 , n397825 );
buf ( n397827 , n377370 );
not ( n397828 , n397827 );
or ( n397829 , n397826 , n397828 );
buf ( n397830 , n385650 );
buf ( n397831 , n371732 );
nand ( n76632 , n397830 , n397831 );
buf ( n397833 , n76632 );
buf ( n397834 , n397833 );
nand ( n76635 , n397829 , n397834 );
buf ( n397836 , n76635 );
xor ( n76637 , n397824 , n397836 );
buf ( n397838 , n76637 );
buf ( n397839 , n383629 );
not ( n397840 , n397839 );
buf ( n397841 , n359312 );
not ( n397842 , n397841 );
or ( n397843 , n397840 , n397842 );
buf ( n397844 , n359297 );
buf ( n397845 , n378098 );
nand ( n397846 , n397844 , n397845 );
buf ( n397847 , n397846 );
buf ( n397848 , n397847 );
not ( n397849 , n397848 );
buf ( n397850 , n378098 );
not ( n76651 , n397850 );
buf ( n397852 , n57481 );
nand ( n397853 , n76651 , n397852 );
buf ( n397854 , n397853 );
buf ( n397855 , n397854 );
not ( n76656 , n397855 );
or ( n76657 , n397849 , n76656 );
buf ( n397858 , n39205 );
nand ( n397859 , n76657 , n397858 );
buf ( n397860 , n397859 );
buf ( n397861 , n397860 );
buf ( n397862 , n359312 );
or ( n397863 , n397861 , n397862 );
nand ( n397864 , n397843 , n397863 );
buf ( n397865 , n397864 );
buf ( n397866 , n397865 );
buf ( n397867 , n49609 );
not ( n397868 , n397867 );
buf ( n397869 , n383606 );
not ( n397870 , n397869 );
or ( n397871 , n397868 , n397870 );
buf ( n397872 , n397208 );
not ( n397873 , n397872 );
buf ( n397874 , n369804 );
nand ( n397875 , n397873 , n397874 );
buf ( n397876 , n397875 );
buf ( n397877 , n397876 );
nand ( n397878 , n397871 , n397877 );
buf ( n397879 , n397878 );
buf ( n76664 , n397879 );
xor ( n76665 , n397866 , n76664 );
buf ( n397882 , n368608 );
not ( n76667 , n397882 );
not ( n76668 , n380424 );
not ( n76669 , n30912 );
or ( n397886 , n76668 , n76669 );
nand ( n397887 , n368549 , n365328 );
nand ( n76672 , n397886 , n397887 );
buf ( n397889 , n76672 );
not ( n397890 , n397889 );
or ( n76675 , n76667 , n397890 );
buf ( n397892 , n65170 );
buf ( n397893 , n387542 );
nand ( n397894 , n397892 , n397893 );
buf ( n397895 , n397894 );
buf ( n397896 , n397895 );
nand ( n76681 , n76675 , n397896 );
buf ( n397898 , n76681 );
buf ( n397899 , n397898 );
xor ( n76684 , n385707 , n385711 );
xor ( n397901 , n76684 , n385738 );
buf ( n397902 , n397901 );
buf ( n397903 , n397902 );
xor ( n397904 , n397899 , n397903 );
buf ( n397905 , n377353 );
not ( n397906 , n397905 );
buf ( n397907 , n366332 );
not ( n76692 , n397907 );
or ( n397909 , n397906 , n76692 );
buf ( n397910 , n361911 );
buf ( n397911 , n377352 );
nand ( n397912 , n397910 , n397911 );
buf ( n397913 , n397912 );
buf ( n397914 , n397913 );
nand ( n397915 , n397909 , n397914 );
buf ( n397916 , n397915 );
buf ( n397917 , n397916 );
not ( n397918 , n397917 );
buf ( n76696 , n44591 );
not ( n76697 , n76696 );
or ( n76698 , n397918 , n76697 );
buf ( n397922 , n49692 );
not ( n76700 , n397922 );
buf ( n397924 , n385764 );
nand ( n397925 , n76700 , n397924 );
buf ( n397926 , n397925 );
buf ( n397927 , n397926 );
nand ( n397928 , n76698 , n397927 );
buf ( n397929 , n397928 );
buf ( n397930 , n397929 );
and ( n76708 , n397904 , n397930 );
and ( n76709 , n397899 , n397903 );
or ( n397933 , n76708 , n76709 );
buf ( n397934 , n397933 );
buf ( n397935 , n397934 );
xor ( n397936 , n76665 , n397935 );
buf ( n397937 , n397936 );
buf ( n397938 , n397937 );
xor ( n76716 , n397838 , n397938 );
and ( n76717 , n40252 , n379371 );
not ( n397941 , n40252 );
and ( n76719 , n397941 , n379380 );
or ( n397943 , n76717 , n76719 );
and ( n76721 , n397943 , n58923 );
buf ( n397945 , n73255 );
not ( n397946 , n397945 );
buf ( n76724 , n379359 );
nor ( n76725 , n397946 , n76724 );
buf ( n76726 , n76725 );
nor ( n397950 , n76721 , n76726 );
buf ( n397951 , n397950 );
not ( n397952 , n397951 );
buf ( n397953 , n397952 );
buf ( n397954 , n397953 );
xnor ( n76732 , n76716 , n397954 );
buf ( n76733 , n76732 );
buf ( n397957 , n76733 );
not ( n76735 , n397957 );
buf ( n76736 , n76735 );
buf ( n397960 , n76736 );
xor ( n397961 , n397805 , n397960 );
and ( n397962 , n65199 , n385871 );
not ( n76740 , n65199 );
and ( n397964 , n76740 , n385868 );
or ( n76742 , n397962 , n397964 );
xor ( n397966 , n65195 , n76742 );
not ( n397967 , n379912 );
not ( n397968 , n394457 );
or ( n397969 , n397967 , n397968 );
buf ( n397970 , n379841 );
not ( n397971 , n397970 );
buf ( n397972 , n360886 );
not ( n76750 , n397972 );
or ( n397974 , n397971 , n76750 );
buf ( n76752 , n360893 );
buf ( n397976 , n379847 );
nand ( n76754 , n76752 , n397976 );
buf ( n397978 , n76754 );
buf ( n397979 , n397978 );
nand ( n397980 , n397974 , n397979 );
buf ( n397981 , n397980 );
buf ( n397982 , n397981 );
buf ( n397983 , n379890 );
nand ( n397984 , n397982 , n397983 );
buf ( n397985 , n397984 );
nand ( n397986 , n397969 , n397985 );
not ( n397987 , n397986 );
xor ( n76765 , n397966 , n397987 );
buf ( n397989 , n380407 );
not ( n397990 , n397989 );
buf ( n397991 , n394418 );
not ( n76769 , n397991 );
or ( n397993 , n397990 , n76769 );
buf ( n397994 , n380368 );
not ( n397995 , n397994 );
buf ( n397996 , n360308 );
not ( n397997 , n397996 );
or ( n397998 , n397995 , n397997 );
buf ( n397999 , n360930 );
buf ( n398000 , n384667 );
nand ( n398001 , n397999 , n398000 );
buf ( n398002 , n398001 );
buf ( n398003 , n398002 );
nand ( n398004 , n397998 , n398003 );
buf ( n398005 , n398004 );
buf ( n398006 , n398005 );
buf ( n398007 , n380356 );
nand ( n398008 , n398006 , n398007 );
buf ( n398009 , n398008 );
buf ( n398010 , n398009 );
nand ( n398011 , n397993 , n398010 );
buf ( n398012 , n398011 );
xor ( n76790 , n76765 , n398012 );
buf ( n398014 , n76790 );
not ( n398015 , n398014 );
buf ( n398016 , n398015 );
buf ( n398017 , n398016 );
xor ( n398018 , n397961 , n398017 );
buf ( n398019 , n398018 );
buf ( n398020 , n397144 );
not ( n398021 , n398020 );
buf ( n76799 , n397218 );
nand ( n76800 , n398021 , n76799 );
buf ( n398024 , n76800 );
buf ( n398025 , n398024 );
not ( n76803 , n398025 );
buf ( n398027 , n397489 );
not ( n398028 , n398027 );
or ( n398029 , n76803 , n398028 );
buf ( n398030 , n397218 );
not ( n398031 , n398030 );
buf ( n76809 , n397144 );
nand ( n76810 , n398031 , n76809 );
buf ( n398034 , n76810 );
buf ( n398035 , n398034 );
nand ( n76813 , n398029 , n398035 );
buf ( n398037 , n76813 );
buf ( n398038 , n398037 );
xor ( n398039 , n397899 , n397903 );
xor ( n76817 , n398039 , n397930 );
buf ( n76818 , n76817 );
buf ( n398042 , n76818 );
buf ( n398043 , n369444 );
not ( n398044 , n398043 );
buf ( n398045 , n76672 );
not ( n76823 , n398045 );
or ( n398047 , n398044 , n76823 );
buf ( n398048 , n393949 );
buf ( n398049 , n368608 );
nand ( n76827 , n398048 , n398049 );
buf ( n398051 , n76827 );
buf ( n398052 , n398051 );
nand ( n76830 , n398047 , n398052 );
buf ( n76831 , n76830 );
buf ( n398055 , n76831 );
xor ( n398056 , n397414 , n397427 );
and ( n76834 , n398056 , n397443 );
and ( n76835 , n397414 , n397427 );
or ( n398059 , n76834 , n76835 );
buf ( n398060 , n398059 );
buf ( n398061 , n398060 );
xor ( n398062 , n398055 , n398061 );
buf ( n76840 , n75971 );
not ( n398064 , n76840 );
buf ( n398065 , n398064 );
buf ( n398066 , n398065 );
not ( n76842 , n398066 );
buf ( n398068 , n46135 );
not ( n398069 , n398068 );
or ( n76845 , n76842 , n398069 );
buf ( n398071 , n397916 );
buf ( n398072 , n41835 );
nand ( n76848 , n398071 , n398072 );
buf ( n398074 , n76848 );
buf ( n398075 , n398074 );
nand ( n76851 , n76845 , n398075 );
buf ( n398077 , n76851 );
buf ( n398078 , n398077 );
and ( n76854 , n398062 , n398078 );
and ( n398080 , n398055 , n398061 );
or ( n76856 , n76854 , n398080 );
buf ( n398082 , n76856 );
buf ( n398083 , n398082 );
xor ( n76859 , n398042 , n398083 );
buf ( n398085 , n379299 );
not ( n398086 , n398085 );
buf ( n398087 , n397366 );
not ( n398088 , n398087 );
or ( n76864 , n398086 , n398088 );
buf ( n398090 , n397787 );
buf ( n398091 , n379263 );
nand ( n398092 , n398090 , n398091 );
buf ( n398093 , n398092 );
buf ( n398094 , n398093 );
nand ( n398095 , n76864 , n398094 );
buf ( n398096 , n398095 );
buf ( n398097 , n398096 );
xor ( n76873 , n76859 , n398097 );
buf ( n398099 , n76873 );
buf ( n76875 , n398099 );
xor ( n398101 , n398055 , n398061 );
xor ( n76877 , n398101 , n398078 );
buf ( n398103 , n76877 );
buf ( n398104 , n398103 );
not ( n76880 , n398104 );
buf ( n76881 , n76880 );
buf ( n398107 , n76881 );
not ( n398108 , n398107 );
not ( n76884 , n75038 );
not ( n76885 , n59424 );
and ( n398111 , n76884 , n76885 );
and ( n76887 , n394472 , n379890 );
nor ( n76888 , n398111 , n76887 );
buf ( n398114 , n76888 );
not ( n76890 , n398114 );
or ( n76891 , n398108 , n76890 );
buf ( n398117 , n379263 );
not ( n76893 , n398117 );
buf ( n398119 , n76242 );
not ( n76895 , n398119 );
or ( n398121 , n76893 , n76895 );
and ( n76897 , n361712 , n379274 );
not ( n398123 , n361712 );
and ( n398124 , n398123 , n379271 );
or ( n76900 , n76897 , n398124 );
buf ( n398126 , n76900 );
buf ( n398127 , n379299 );
nand ( n76903 , n398126 , n398127 );
buf ( n398129 , n76903 );
buf ( n398130 , n398129 );
nand ( n76906 , n398121 , n398130 );
buf ( n398132 , n76906 );
buf ( n398133 , n44915 );
not ( n76909 , n398133 );
buf ( n398135 , n394528 );
not ( n398136 , n398135 );
or ( n76912 , n76909 , n398136 );
buf ( n398138 , n396171 );
buf ( n398139 , n47466 );
nand ( n398140 , n398138 , n398139 );
buf ( n398141 , n398140 );
buf ( n398142 , n398141 );
nand ( n76918 , n76912 , n398142 );
buf ( n398144 , n76918 );
buf ( n398145 , n398144 );
not ( n398146 , n398145 );
buf ( n398147 , n48502 );
not ( n398148 , n398147 );
buf ( n398149 , n396981 );
not ( n76925 , n398149 );
and ( n398151 , n398148 , n76925 );
buf ( n76927 , n394508 );
buf ( n398153 , n73479 );
nor ( n398154 , n76927 , n398153 );
buf ( n398155 , n398154 );
buf ( n398156 , n398155 );
nor ( n398157 , n398151 , n398156 );
buf ( n398158 , n398157 );
buf ( n398159 , n398158 );
not ( n398160 , n398159 );
buf ( n398161 , n398160 );
buf ( n398162 , n398161 );
not ( n398163 , n398162 );
or ( n398164 , n398146 , n398163 );
buf ( n398165 , n398144 );
not ( n398166 , n398165 );
buf ( n398167 , n398166 );
buf ( n398168 , n398167 );
not ( n398169 , n398168 );
buf ( n398170 , n398158 );
not ( n398171 , n398170 );
or ( n398172 , n398169 , n398171 );
buf ( n398173 , n49609 );
not ( n398174 , n398173 );
buf ( n398175 , n393896 );
not ( n398176 , n398175 );
or ( n398177 , n398174 , n398176 );
buf ( n398178 , n393883 );
not ( n398179 , n398178 );
buf ( n398180 , n366131 );
not ( n76930 , n398180 );
or ( n76931 , n398179 , n76930 );
buf ( n398183 , n351367 );
buf ( n398184 , n369763 );
nand ( n398185 , n398183 , n398184 );
buf ( n398186 , n398185 );
buf ( n398187 , n398186 );
nand ( n76936 , n76931 , n398187 );
buf ( n398189 , n76936 );
buf ( n398190 , n398189 );
buf ( n398191 , n369804 );
nand ( n76940 , n398190 , n398191 );
buf ( n398193 , n76940 );
buf ( n398194 , n398193 );
nand ( n76943 , n398177 , n398194 );
buf ( n398196 , n76943 );
buf ( n398197 , n398196 );
nand ( n76946 , n398172 , n398197 );
buf ( n76947 , n76946 );
buf ( n398200 , n76947 );
nand ( n76949 , n398164 , n398200 );
buf ( n398202 , n76949 );
xor ( n398203 , n398132 , n398202 );
buf ( n398204 , n74024 );
buf ( n398205 , n394538 );
xor ( n76954 , n398204 , n398205 );
buf ( n398207 , n73481 );
xor ( n76956 , n76954 , n398207 );
buf ( n398209 , n76956 );
and ( n76958 , n398203 , n398209 );
and ( n76959 , n398132 , n398202 );
or ( n76960 , n76958 , n76959 );
buf ( n398213 , n76960 );
nand ( n398214 , n76891 , n398213 );
buf ( n398215 , n398214 );
buf ( n398216 , n398215 );
buf ( n398217 , n76888 );
not ( n398218 , n398217 );
buf ( n398219 , n398218 );
buf ( n398220 , n398219 );
buf ( n398221 , n398103 );
nand ( n76970 , n398220 , n398221 );
buf ( n398223 , n76970 );
buf ( n398224 , n398223 );
nand ( n76973 , n398216 , n398224 );
buf ( n398226 , n76973 );
buf ( n398227 , n398226 );
xor ( n76976 , n76875 , n398227 );
not ( n398229 , n395325 );
xor ( n398230 , n395330 , n74329 );
not ( n76979 , n398230 );
not ( n398232 , n76979 );
or ( n76981 , n398229 , n398232 );
not ( n398234 , n395325 );
nand ( n398235 , n398234 , n398230 );
nand ( n398236 , n76981 , n398235 );
buf ( n398237 , n395129 );
not ( n398238 , n398237 );
buf ( n398239 , n395090 );
not ( n76988 , n398239 );
or ( n76989 , n398238 , n76988 );
buf ( n398242 , n395129 );
not ( n398243 , n398242 );
buf ( n398244 , n398243 );
buf ( n398245 , n398244 );
not ( n398246 , n398245 );
buf ( n398247 , n74060 );
not ( n76996 , n398247 );
or ( n398249 , n398246 , n76996 );
buf ( n398250 , n395063 );
nand ( n398251 , n398249 , n398250 );
buf ( n398252 , n398251 );
buf ( n398253 , n398252 );
nand ( n77002 , n76989 , n398253 );
buf ( n398255 , n77002 );
not ( n77004 , n398255 );
xor ( n77005 , n398236 , n77004 );
xor ( n398258 , n395216 , n395233 );
and ( n398259 , n398258 , n395271 );
and ( n77008 , n395216 , n395233 );
or ( n77009 , n398259 , n77008 );
buf ( n398262 , n77009 );
xor ( n398263 , n77005 , n398262 );
buf ( n398264 , n398263 );
and ( n398265 , n76976 , n398264 );
and ( n398266 , n76875 , n398227 );
or ( n77015 , n398265 , n398266 );
buf ( n398268 , n77015 );
buf ( n398269 , n398268 );
xor ( n77018 , n398038 , n398269 );
xor ( n77019 , n398042 , n398083 );
and ( n398272 , n77019 , n398097 );
and ( n77021 , n398042 , n398083 );
or ( n398274 , n398272 , n77021 );
buf ( n398275 , n398274 );
buf ( n398276 , n398275 );
not ( n77025 , n398236 );
not ( n77026 , n77004 );
or ( n77027 , n77025 , n77026 );
nand ( n77028 , n77027 , n398262 );
buf ( n77029 , n77028 );
not ( n398282 , n398236 );
nand ( n77031 , n398282 , n398255 );
buf ( n398284 , n77031 );
nand ( n398285 , n77029 , n398284 );
buf ( n398286 , n398285 );
buf ( n398287 , n398286 );
xor ( n398288 , n398276 , n398287 );
xor ( n77037 , n385743 , n385750 );
xor ( n77038 , n77037 , n385778 );
buf ( n77039 , n77038 );
buf ( n398292 , n77039 );
buf ( n398293 , n386148 );
buf ( n398294 , n385948 );
and ( n77043 , n398293 , n398294 );
not ( n77044 , n398293 );
buf ( n398297 , n385945 );
and ( n398298 , n77044 , n398297 );
nor ( n398299 , n77043 , n398298 );
buf ( n398300 , n398299 );
buf ( n398301 , n398300 );
buf ( n398302 , n385925 );
and ( n77051 , n398301 , n398302 );
not ( n398304 , n398301 );
buf ( n398305 , n385925 );
not ( n77054 , n398305 );
buf ( n77055 , n77054 );
buf ( n398308 , n77055 );
and ( n77057 , n398304 , n398308 );
nor ( n398310 , n77051 , n77057 );
buf ( n398311 , n398310 );
buf ( n398312 , n398311 );
xor ( n398313 , n398292 , n398312 );
not ( n77062 , n394243 );
nor ( n77063 , n77062 , n73142 );
or ( n398316 , n77063 , n394215 );
nand ( n398317 , n73142 , n394240 );
nand ( n77066 , n398316 , n398317 );
buf ( n398319 , n77066 );
xor ( n398320 , n398313 , n398319 );
buf ( n398321 , n398320 );
buf ( n398322 , n398321 );
xor ( n398323 , n398288 , n398322 );
buf ( n398324 , n398323 );
buf ( n398325 , n398324 );
xor ( n77074 , n77018 , n398325 );
buf ( n398327 , n77074 );
xor ( n77076 , n398019 , n398327 );
xor ( n398329 , n76875 , n398227 );
xor ( n398330 , n398329 , n398264 );
buf ( n398331 , n398330 );
buf ( n398332 , n398331 );
buf ( n398333 , n380356 );
not ( n77082 , n398333 );
buf ( n398335 , n74118 );
not ( n77084 , n398335 );
or ( n398337 , n77082 , n77084 );
buf ( n398338 , n380368 );
not ( n77087 , n398338 );
buf ( n398340 , n368474 );
not ( n398341 , n398340 );
or ( n77090 , n77087 , n398341 );
buf ( n398343 , n360893 );
buf ( n398344 , n384667 );
nand ( n77093 , n398343 , n398344 );
buf ( n398346 , n77093 );
buf ( n398347 , n398346 );
nand ( n77096 , n77090 , n398347 );
buf ( n77097 , n77096 );
buf ( n398350 , n77097 );
buf ( n398351 , n380404 );
nand ( n398352 , n398350 , n398351 );
buf ( n398353 , n398352 );
buf ( n398354 , n398353 );
nand ( n77103 , n398337 , n398354 );
buf ( n398356 , n77103 );
buf ( n398357 , n398356 );
buf ( n398358 , n397190 );
not ( n77107 , n398358 );
buf ( n398360 , n397234 );
not ( n77109 , n398360 );
or ( n77110 , n77107 , n77109 );
buf ( n398363 , n377583 );
buf ( n398364 , n398363 );
not ( n398365 , n398364 );
buf ( n398366 , n364771 );
not ( n77115 , n398366 );
or ( n398368 , n398365 , n77115 );
buf ( n398369 , n386390 );
buf ( n398370 , n377592 );
nand ( n398371 , n398369 , n398370 );
buf ( n398372 , n398371 );
buf ( n398373 , n398372 );
nand ( n398374 , n398368 , n398373 );
buf ( n398375 , n398374 );
buf ( n398376 , n398375 );
buf ( n398377 , n57530 );
nand ( n77126 , n398376 , n398377 );
buf ( n398379 , n77126 );
buf ( n398380 , n398379 );
nand ( n77129 , n77110 , n398380 );
buf ( n398382 , n77129 );
buf ( n398383 , n398382 );
buf ( n398384 , n397288 );
buf ( n398385 , n397319 );
xor ( n77134 , n398384 , n398385 );
buf ( n398387 , n397335 );
xor ( n398388 , n77134 , n398387 );
buf ( n398389 , n398388 );
buf ( n398390 , n398389 );
xor ( n398391 , n398383 , n398390 );
buf ( n398392 , n361603 );
buf ( n398393 , n45414 );
not ( n398394 , n398393 );
buf ( n398395 , n379482 );
not ( n77144 , n398395 );
and ( n398397 , n398394 , n77144 );
buf ( n77146 , n361531 );
buf ( n398399 , n379482 );
and ( n398400 , n77146 , n398399 );
nor ( n398401 , n398397 , n398400 );
buf ( n398402 , n398401 );
buf ( n398403 , n398402 );
or ( n77152 , n398392 , n398403 );
buf ( n398405 , n397259 );
not ( n398406 , n398405 );
buf ( n398407 , n398406 );
buf ( n398408 , n398407 );
buf ( n398409 , n364098 );
or ( n398410 , n398408 , n398409 );
nand ( n398411 , n77152 , n398410 );
buf ( n398412 , n398411 );
buf ( n398413 , n398412 );
and ( n398414 , n398391 , n398413 );
and ( n398415 , n398383 , n398390 );
or ( n77164 , n398414 , n398415 );
buf ( n398417 , n77164 );
buf ( n398418 , n398417 );
xor ( n398419 , n398357 , n398418 );
buf ( n398420 , n398144 );
buf ( n398421 , n398196 );
xor ( n398422 , n398420 , n398421 );
buf ( n398423 , n398161 );
xnor ( n398424 , n398422 , n398423 );
buf ( n398425 , n398424 );
buf ( n398426 , n398425 );
not ( n398427 , n398426 );
buf ( n398428 , n398427 );
not ( n77177 , n398428 );
buf ( n398430 , n379263 );
not ( n77179 , n398430 );
buf ( n398432 , n76900 );
not ( n77181 , n398432 );
or ( n398434 , n77179 , n77181 );
buf ( n398435 , n379271 );
buf ( n398436 , n370310 );
and ( n398437 , n398435 , n398436 );
not ( n398438 , n398435 );
buf ( n398439 , n46126 );
and ( n398440 , n398438 , n398439 );
nor ( n398441 , n398437 , n398440 );
buf ( n398442 , n398441 );
buf ( n398443 , n398442 );
not ( n398444 , n398443 );
buf ( n398445 , n379299 );
nand ( n398446 , n398444 , n398445 );
buf ( n398447 , n398446 );
buf ( n398448 , n398447 );
nand ( n398449 , n398434 , n398448 );
buf ( n398450 , n398449 );
not ( n77190 , n398450 );
or ( n77191 , n77177 , n77190 );
not ( n398453 , n398425 );
buf ( n398454 , n398450 );
not ( n77194 , n398454 );
buf ( n398456 , n77194 );
not ( n77196 , n398456 );
or ( n77197 , n398453 , n77196 );
buf ( n398459 , n369804 );
not ( n398460 , n398459 );
buf ( n398461 , n393883 );
not ( n77201 , n398461 );
buf ( n398463 , n31073 );
not ( n398464 , n398463 );
or ( n77204 , n77201 , n398464 );
buf ( n398466 , n351107 );
buf ( n398467 , n369763 );
nand ( n398468 , n398466 , n398467 );
buf ( n398469 , n398468 );
buf ( n398470 , n398469 );
nand ( n398471 , n77204 , n398470 );
buf ( n398472 , n398471 );
buf ( n398473 , n398472 );
not ( n398474 , n398473 );
or ( n398475 , n398460 , n398474 );
buf ( n398476 , n398189 );
buf ( n398477 , n369809 );
nand ( n398478 , n398476 , n398477 );
buf ( n398479 , n398478 );
buf ( n398480 , n398479 );
nand ( n398481 , n398475 , n398480 );
buf ( n398482 , n398481 );
not ( n398483 , n398482 );
buf ( n398484 , n365303 );
buf ( n398485 , n378098 );
nand ( n398486 , n398484 , n398485 );
buf ( n398487 , n398486 );
nand ( n398488 , n398483 , n398487 );
not ( n398489 , n398488 );
buf ( n398490 , n57530 );
not ( n398491 , n398490 );
buf ( n398492 , n398363 );
not ( n398493 , n398492 );
buf ( n398494 , n363041 );
not ( n398495 , n398494 );
or ( n398496 , n398493 , n398495 );
buf ( n398497 , n42891 );
buf ( n398498 , n377592 );
nand ( n398499 , n398497 , n398498 );
buf ( n398500 , n398499 );
buf ( n398501 , n398500 );
nand ( n77213 , n398496 , n398501 );
buf ( n398503 , n77213 );
buf ( n398504 , n398503 );
not ( n77216 , n398504 );
or ( n398506 , n398491 , n77216 );
buf ( n398507 , n398375 );
buf ( n398508 , n397190 );
nand ( n77220 , n398507 , n398508 );
buf ( n77221 , n77220 );
buf ( n398511 , n77221 );
nand ( n77223 , n398506 , n398511 );
buf ( n398513 , n77223 );
not ( n398514 , n398513 );
or ( n398515 , n398489 , n398514 );
buf ( n398516 , n398487 );
not ( n77228 , n398516 );
buf ( n398518 , n398482 );
nand ( n398519 , n77228 , n398518 );
buf ( n398520 , n398519 );
nand ( n77232 , n398515 , n398520 );
nand ( n398522 , n77197 , n77232 );
nand ( n77234 , n77191 , n398522 );
buf ( n398524 , n77234 );
and ( n398525 , n398419 , n398524 );
and ( n77237 , n398357 , n398418 );
or ( n398527 , n398525 , n77237 );
buf ( n398528 , n398527 );
buf ( n398529 , n398528 );
not ( n398530 , n398529 );
buf ( n398531 , n395273 );
buf ( n398532 , n395159 );
xor ( n398533 , n398531 , n398532 );
buf ( n398534 , n395135 );
xor ( n77246 , n398533 , n398534 );
buf ( n398536 , n77246 );
buf ( n77248 , n398536 );
not ( n398538 , n77248 );
buf ( n398539 , n398538 );
buf ( n398540 , n398539 );
not ( n398541 , n398540 );
or ( n77253 , n398530 , n398541 );
buf ( n398543 , n398528 );
not ( n398544 , n398543 );
buf ( n398545 , n398544 );
buf ( n77257 , n398545 );
not ( n77258 , n77257 );
buf ( n398548 , n398536 );
not ( n77260 , n398548 );
or ( n398550 , n77258 , n77260 );
buf ( n398551 , n397341 );
buf ( n398552 , n397244 );
xor ( n398553 , n398551 , n398552 );
buf ( n398554 , n76123 );
xor ( n77266 , n398553 , n398554 );
buf ( n398556 , n77266 );
buf ( n398557 , n398556 );
xor ( n398558 , n397446 , n397462 );
xor ( n77270 , n398558 , n397479 );
buf ( n398560 , n77270 );
buf ( n398561 , n398560 );
xor ( n398562 , n398557 , n398561 );
buf ( n398563 , n58923 );
not ( n77275 , n398563 );
buf ( n398565 , n395408 );
not ( n398566 , n398565 );
or ( n77278 , n77275 , n398566 );
buf ( n398568 , n379371 );
not ( n398569 , n398568 );
buf ( n398570 , n367116 );
not ( n398571 , n398570 );
or ( n77283 , n398569 , n398571 );
buf ( n398573 , n362136 );
buf ( n398574 , n379380 );
nand ( n77286 , n398573 , n398574 );
buf ( n398576 , n77286 );
buf ( n398577 , n398576 );
nand ( n77289 , n77283 , n398577 );
buf ( n77290 , n77289 );
buf ( n398580 , n77290 );
buf ( n398581 , n58871 );
nand ( n398582 , n398580 , n398581 );
buf ( n398583 , n398582 );
buf ( n398584 , n398583 );
nand ( n398585 , n77278 , n398584 );
buf ( n398586 , n398585 );
buf ( n398587 , n398586 );
and ( n398588 , n398562 , n398587 );
and ( n77300 , n398557 , n398561 );
or ( n398590 , n398588 , n77300 );
buf ( n398591 , n398590 );
buf ( n398592 , n398591 );
nand ( n398593 , n398550 , n398592 );
buf ( n398594 , n398593 );
buf ( n398595 , n398594 );
nand ( n398596 , n77253 , n398595 );
buf ( n398597 , n398596 );
buf ( n398598 , n398597 );
xor ( n398599 , n398332 , n398598 );
xor ( n398600 , n395418 , n395421 );
xor ( n77312 , n398600 , n397069 );
buf ( n398602 , n77312 );
buf ( n398603 , n398103 );
buf ( n398604 , n398219 );
xor ( n398605 , n398603 , n398604 );
buf ( n398606 , n76960 );
xnor ( n77318 , n398605 , n398606 );
buf ( n398608 , n77318 );
buf ( n398609 , n398608 );
not ( n77321 , n398609 );
buf ( n398611 , n77321 );
buf ( n398612 , n398611 );
or ( n398613 , n398602 , n398612 );
xor ( n77325 , n398132 , n398202 );
xor ( n77326 , n77325 , n398209 );
buf ( n77327 , n77326 );
xor ( n398617 , n397509 , n76482 );
buf ( n398618 , n398617 );
buf ( n398619 , n76347 );
and ( n398620 , n398618 , n398619 );
not ( n77332 , n398618 );
buf ( n398622 , n397517 );
and ( n398623 , n77332 , n398622 );
nor ( n398624 , n398620 , n398623 );
buf ( n398625 , n398624 );
buf ( n398626 , n398625 );
xor ( n398627 , n77327 , n398626 );
buf ( n398628 , n397562 );
not ( n398629 , n398628 );
buf ( n398630 , n76382 );
not ( n77342 , n398630 );
or ( n398632 , n398629 , n77342 );
buf ( n398633 , n397553 );
buf ( n398634 , n397540 );
nand ( n77346 , n398633 , n398634 );
buf ( n398636 , n77346 );
buf ( n398637 , n398636 );
nand ( n77349 , n398632 , n398637 );
buf ( n398639 , n77349 );
buf ( n398640 , n398639 );
buf ( n398641 , n397676 );
xor ( n398642 , n398640 , n398641 );
buf ( n398643 , n398642 );
buf ( n398644 , n398643 );
xor ( n398645 , n397573 , n397577 );
xor ( n398646 , n398645 , n397672 );
buf ( n398647 , n398646 );
buf ( n398648 , n398647 );
buf ( n398649 , n44915 );
not ( n398650 , n398649 );
buf ( n398651 , n396186 );
not ( n398652 , n398651 );
or ( n398653 , n398650 , n398652 );
xor ( n77365 , n32202 , n380497 );
buf ( n398655 , n77365 );
not ( n398656 , n398655 );
buf ( n398657 , n47466 );
nand ( n77369 , n398656 , n398657 );
buf ( n398659 , n77369 );
buf ( n398660 , n398659 );
nand ( n398661 , n398653 , n398660 );
buf ( n398662 , n398661 );
buf ( n398663 , n398662 );
xor ( n398664 , n397628 , n397641 );
xor ( n77376 , n398664 , n397667 );
buf ( n398666 , n77376 );
buf ( n398667 , n398666 );
xor ( n77379 , n398663 , n398667 );
buf ( n398669 , n43274 );
buf ( n398670 , n377782 );
not ( n398671 , n398670 );
buf ( n398672 , n381286 );
not ( n77384 , n398672 );
or ( n398674 , n398671 , n77384 );
buf ( n398675 , n386354 );
buf ( n398676 , n377779 );
nand ( n77388 , n398675 , n398676 );
buf ( n77389 , n77388 );
buf ( n398679 , n77389 );
nand ( n77391 , n398674 , n398679 );
buf ( n398681 , n77391 );
buf ( n398682 , n398681 );
not ( n77394 , n398682 );
buf ( n398684 , n77394 );
buf ( n398685 , n398684 );
or ( n398686 , n398669 , n398685 );
buf ( n398687 , n396130 );
not ( n398688 , n398687 );
buf ( n398689 , n398688 );
buf ( n398690 , n398689 );
buf ( n398691 , n378183 );
not ( n398692 , n398691 );
buf ( n398693 , n398692 );
buf ( n398694 , n398693 );
or ( n77406 , n398690 , n398694 );
nand ( n398696 , n398686 , n77406 );
buf ( n398697 , n398696 );
buf ( n398698 , n398697 );
and ( n77410 , n77379 , n398698 );
and ( n398700 , n398663 , n398667 );
or ( n77412 , n77410 , n398700 );
buf ( n398702 , n77412 );
buf ( n398703 , n398702 );
xor ( n398704 , n398648 , n398703 );
buf ( n398705 , n361971 );
buf ( n398706 , n377122 );
buf ( n398707 , n367248 );
and ( n398708 , n398706 , n398707 );
not ( n77420 , n398706 );
buf ( n398710 , n364744 );
and ( n398711 , n77420 , n398710 );
nor ( n77423 , n398708 , n398711 );
buf ( n398713 , n77423 );
buf ( n398714 , n398713 );
or ( n398715 , n398705 , n398714 );
buf ( n398716 , n74432 );
buf ( n398717 , n366339 );
or ( n398718 , n398716 , n398717 );
nand ( n398719 , n398715 , n398718 );
buf ( n398720 , n398719 );
buf ( n398721 , n398720 );
and ( n398722 , n398704 , n398721 );
and ( n77434 , n398648 , n398703 );
or ( n77435 , n398722 , n77434 );
buf ( n398725 , n77435 );
buf ( n398726 , n398725 );
xor ( n77438 , n398644 , n398726 );
buf ( n398728 , n396109 );
not ( n77440 , n398728 );
buf ( n398730 , n379890 );
not ( n77442 , n398730 );
or ( n77443 , n77440 , n77442 );
buf ( n398733 , n379838 );
not ( n77445 , n398733 );
buf ( n398735 , n377961 );
not ( n398736 , n398735 );
or ( n398737 , n77445 , n398736 );
buf ( n398738 , n372889 );
buf ( n398739 , n379838 );
not ( n77451 , n398739 );
buf ( n398741 , n77451 );
buf ( n398742 , n398741 );
nand ( n77454 , n398738 , n398742 );
buf ( n398744 , n77454 );
buf ( n398745 , n398744 );
nand ( n398746 , n398737 , n398745 );
buf ( n398747 , n398746 );
buf ( n398748 , n398747 );
buf ( n398749 , n379916 );
nand ( n77461 , n398748 , n398749 );
buf ( n398751 , n77461 );
buf ( n398752 , n398751 );
nand ( n398753 , n77443 , n398752 );
buf ( n398754 , n398753 );
buf ( n398755 , n398754 );
and ( n398756 , n77438 , n398755 );
and ( n77468 , n398644 , n398726 );
or ( n398758 , n398756 , n77468 );
buf ( n398759 , n398758 );
buf ( n398760 , n398759 );
and ( n77472 , n398627 , n398760 );
and ( n398762 , n77327 , n398626 );
or ( n77474 , n77472 , n398762 );
buf ( n398764 , n77474 );
buf ( n77476 , n398764 );
nand ( n398766 , n398613 , n77476 );
buf ( n398767 , n398766 );
buf ( n398768 , n398767 );
buf ( n398769 , n77312 );
buf ( n398770 , n398611 );
nand ( n398771 , n398769 , n398770 );
buf ( n398772 , n398771 );
buf ( n398773 , n398772 );
nand ( n398774 , n398768 , n398773 );
buf ( n398775 , n398774 );
buf ( n398776 , n398775 );
and ( n77488 , n398599 , n398776 );
and ( n398778 , n398332 , n398598 );
or ( n398779 , n77488 , n398778 );
buf ( n398780 , n398779 );
and ( n398781 , n77076 , n398780 );
and ( n398782 , n398019 , n398327 );
or ( n77494 , n398781 , n398782 );
buf ( n398784 , n77494 );
xor ( n398785 , n397751 , n398784 );
buf ( n398786 , n398785 );
buf ( n398787 , n398786 );
xor ( n77499 , n398038 , n398269 );
and ( n398789 , n77499 , n398325 );
and ( n77501 , n398038 , n398269 );
or ( n398791 , n398789 , n77501 );
buf ( n398792 , n398791 );
buf ( n398793 , n398792 );
xor ( n398794 , n385827 , n385900 );
xor ( n77506 , n398794 , n386154 );
buf ( n398796 , n77506 );
buf ( n398797 , n398796 );
xor ( n77509 , n398292 , n398312 );
and ( n398799 , n77509 , n398319 );
and ( n398800 , n398292 , n398312 );
or ( n77512 , n398799 , n398800 );
buf ( n398802 , n77512 );
buf ( n398803 , n398802 );
xor ( n398804 , n398797 , n398803 );
xor ( n77516 , n397758 , n397795 );
and ( n398806 , n77516 , n397802 );
and ( n398807 , n397758 , n397795 );
or ( n77519 , n398806 , n398807 );
buf ( n398809 , n77519 );
buf ( n398810 , n398809 );
xnor ( n398811 , n398804 , n398810 );
buf ( n398812 , n398811 );
buf ( n398813 , n398812 );
buf ( n398814 , n398813 );
buf ( n398815 , n398814 );
buf ( n398816 , n398815 );
not ( n77528 , n398816 );
xor ( n77529 , n398276 , n398287 );
and ( n398819 , n77529 , n398322 );
and ( n77531 , n398276 , n398287 );
or ( n398821 , n398819 , n77531 );
buf ( n398822 , n398821 );
buf ( n77534 , n398822 );
not ( n77535 , n77534 );
buf ( n77536 , n77535 );
buf ( n398826 , n77536 );
not ( n77538 , n398826 );
xor ( n77539 , n395371 , n395380 );
and ( n398829 , n77539 , n395390 );
and ( n398830 , n395371 , n395380 );
or ( n77542 , n398829 , n398830 );
buf ( n398832 , n77542 );
buf ( n398833 , n398832 );
not ( n77545 , n398833 );
or ( n77546 , n77538 , n77545 );
buf ( n398836 , n77536 );
buf ( n398837 , n398832 );
or ( n398838 , n398836 , n398837 );
nand ( n77550 , n77546 , n398838 );
buf ( n398840 , n77550 );
buf ( n398841 , n398840 );
not ( n77553 , n398841 );
or ( n77554 , n77528 , n77553 );
buf ( n398844 , n398840 );
buf ( n398845 , n398815 );
or ( n398846 , n398844 , n398845 );
nand ( n398847 , n77554 , n398846 );
buf ( n398848 , n398847 );
buf ( n398849 , n398848 );
xor ( n398850 , n398793 , n398849 );
xor ( n77562 , n397866 , n76664 );
and ( n77563 , n77562 , n397935 );
and ( n398853 , n397866 , n76664 );
or ( n398854 , n77563 , n398853 );
buf ( n398855 , n398854 );
buf ( n398856 , n398855 );
buf ( n398857 , n379263 );
not ( n398858 , n398857 );
buf ( n398859 , n385806 );
not ( n77571 , n398859 );
or ( n398861 , n398858 , n77571 );
buf ( n398862 , n397772 );
buf ( n398863 , n379299 );
nand ( n77575 , n398862 , n398863 );
buf ( n398865 , n77575 );
buf ( n398866 , n398865 );
nand ( n398867 , n398861 , n398866 );
buf ( n398868 , n398867 );
buf ( n398869 , n398868 );
xor ( n77581 , n398856 , n398869 );
buf ( n398871 , n383728 );
buf ( n398872 , n383612 );
xor ( n77584 , n398871 , n398872 );
buf ( n398874 , n383650 );
xor ( n77586 , n77584 , n398874 );
buf ( n398876 , n77586 );
buf ( n398877 , n398876 );
xnor ( n77589 , n77581 , n398877 );
buf ( n398879 , n77589 );
buf ( n398880 , n398879 );
buf ( n398881 , n397937 );
not ( n77593 , n398881 );
buf ( n398883 , n397953 );
not ( n398884 , n398883 );
or ( n398885 , n77593 , n398884 );
not ( n77597 , n397937 );
not ( n398887 , n77597 );
not ( n398888 , n397950 );
or ( n398889 , n398887 , n398888 );
nand ( n77601 , n398889 , n76637 );
buf ( n77602 , n77601 );
nand ( n77603 , n398885 , n77602 );
buf ( n77604 , n77603 );
buf ( n398894 , n77604 );
and ( n77606 , n398880 , n398894 );
not ( n398896 , n398880 );
buf ( n398897 , n77604 );
not ( n398898 , n398897 );
buf ( n398899 , n398898 );
buf ( n398900 , n398899 );
and ( n398901 , n398896 , n398900 );
nor ( n398902 , n77606 , n398901 );
buf ( n398903 , n398902 );
xor ( n77615 , n395295 , n74279 );
and ( n398905 , n77615 , n395368 );
and ( n398906 , n395295 , n74279 );
or ( n77618 , n398905 , n398906 );
buf ( n398908 , n77618 );
buf ( n398909 , n398908 );
xor ( n77621 , n385662 , n385684 );
xor ( n77622 , n77621 , n385782 );
buf ( n398912 , n77622 );
xor ( n77624 , n398909 , n398912 );
buf ( n398914 , n380356 );
not ( n398915 , n398914 );
buf ( n398916 , n380368 );
not ( n398917 , n398916 );
buf ( n398918 , n359784 );
not ( n398919 , n398918 );
or ( n398920 , n398917 , n398919 );
buf ( n398921 , n359781 );
buf ( n398922 , n380364 );
nand ( n398923 , n398921 , n398922 );
buf ( n398924 , n398923 );
buf ( n398925 , n398924 );
nand ( n398926 , n398920 , n398925 );
buf ( n398927 , n398926 );
buf ( n398928 , n398927 );
not ( n398929 , n398928 );
or ( n77641 , n398915 , n398929 );
buf ( n398931 , n398005 );
buf ( n398932 , n380407 );
nand ( n398933 , n398931 , n398932 );
buf ( n398934 , n398933 );
buf ( n398935 , n398934 );
nand ( n398936 , n77641 , n398935 );
buf ( n398937 , n398936 );
buf ( n398938 , n398937 );
xor ( n398939 , n77624 , n398938 );
buf ( n398940 , n398939 );
buf ( n398941 , n398940 );
not ( n77653 , n398941 );
buf ( n398943 , n77653 );
and ( n77655 , n398903 , n398943 );
not ( n398945 , n398903 );
and ( n77657 , n398945 , n398940 );
nor ( n398947 , n77655 , n77657 );
not ( n77659 , n398947 );
not ( n398949 , n77659 );
not ( n77661 , n398949 );
buf ( n398951 , n76733 );
not ( n398952 , n398951 );
buf ( n398953 , n76790 );
not ( n77665 , n398953 );
or ( n398955 , n398952 , n77665 );
buf ( n398956 , n397804 );
nand ( n77668 , n398955 , n398956 );
buf ( n398958 , n77668 );
buf ( n398959 , n398958 );
buf ( n398960 , n398016 );
buf ( n398961 , n76736 );
nand ( n77673 , n398960 , n398961 );
buf ( n398963 , n77673 );
buf ( n398964 , n398963 );
nand ( n77676 , n398959 , n398964 );
buf ( n398966 , n77676 );
buf ( n398967 , n398966 );
not ( n77679 , n398967 );
buf ( n398969 , n77679 );
buf ( n398970 , n398969 );
not ( n398971 , n398970 );
buf ( n398972 , n384580 );
not ( n398973 , n398972 );
buf ( n398974 , n383940 );
not ( n398975 , n398974 );
or ( n398976 , n398973 , n398975 );
buf ( n398977 , n383912 );
buf ( n398978 , n63935 );
nand ( n398979 , n398977 , n398978 );
buf ( n398980 , n398979 );
buf ( n398981 , n398980 );
nand ( n398982 , n398976 , n398981 );
buf ( n398983 , n398982 );
buf ( n398984 , n398983 );
buf ( n398985 , n63293 );
xor ( n398986 , n398984 , n398985 );
buf ( n398987 , n398986 );
buf ( n398988 , n398987 );
xor ( n77700 , n385325 , n64663 );
xor ( n77701 , n77700 , n385354 );
buf ( n398991 , n77701 );
buf ( n398992 , n398991 );
xor ( n77704 , n398988 , n398992 );
xor ( n77705 , n397817 , n397823 );
and ( n77706 , n77705 , n397836 );
and ( n77707 , n397817 , n397823 );
or ( n77708 , n77706 , n77707 );
buf ( n398998 , n77708 );
xor ( n77710 , n77704 , n398998 );
buf ( n77711 , n77710 );
buf ( n399001 , n77711 );
buf ( n399002 , n379890 );
not ( n77714 , n399002 );
buf ( n399004 , n385504 );
not ( n77716 , n399004 );
or ( n77717 , n77714 , n77716 );
buf ( n399007 , n397981 );
buf ( n77719 , n379916 );
nand ( n77720 , n399007 , n77719 );
buf ( n399010 , n77720 );
buf ( n399011 , n399010 );
nand ( n77723 , n77717 , n399011 );
buf ( n399013 , n77723 );
buf ( n399014 , n399013 );
xor ( n77726 , n383463 , n383500 );
xor ( n77727 , n77726 , n383570 );
buf ( n399017 , n77727 );
buf ( n399018 , n399017 );
xor ( n77730 , n399014 , n399018 );
buf ( n399020 , n58923 );
not ( n77732 , n399020 );
buf ( n399022 , n385475 );
not ( n77734 , n399022 );
or ( n399024 , n77732 , n77734 );
buf ( n399025 , n397943 );
buf ( n399026 , n58871 );
nand ( n399027 , n399025 , n399026 );
buf ( n399028 , n399027 );
buf ( n399029 , n399028 );
nand ( n77741 , n399024 , n399029 );
buf ( n77742 , n77741 );
buf ( n399032 , n77742 );
xor ( n77744 , n77730 , n399032 );
buf ( n399034 , n77744 );
buf ( n77746 , n399034 );
xor ( n77747 , n399001 , n77746 );
not ( n399037 , n398012 );
nand ( n399038 , n399037 , n397987 );
not ( n77750 , n399038 );
not ( n77751 , n397966 );
or ( n77752 , n77750 , n77751 );
buf ( n399042 , n398012 );
buf ( n399043 , n397986 );
nand ( n77755 , n399042 , n399043 );
buf ( n399045 , n77755 );
nand ( n399046 , n77752 , n399045 );
buf ( n399047 , n399046 );
xnor ( n399048 , n77747 , n399047 );
buf ( n399049 , n399048 );
buf ( n399050 , n399049 );
not ( n399051 , n399050 );
buf ( n399052 , n399051 );
buf ( n399053 , n399052 );
not ( n399054 , n399053 );
or ( n77766 , n398971 , n399054 );
buf ( n399056 , n399049 );
not ( n77768 , n399056 );
buf ( n399058 , n77768 );
buf ( n399059 , n399058 );
buf ( n399060 , n398969 );
or ( n399061 , n399059 , n399060 );
nand ( n399062 , n77766 , n399061 );
buf ( n399063 , n399062 );
not ( n399064 , n399063 );
or ( n399065 , n77661 , n399064 );
or ( n77777 , n399063 , n398949 );
nand ( n399067 , n399065 , n77777 );
buf ( n399068 , n399067 );
xor ( n77780 , n398850 , n399068 );
buf ( n399070 , n77780 );
buf ( n399071 , n399070 );
xor ( n77783 , n398787 , n399071 );
buf ( n399073 , n77783 );
xor ( n399074 , n395392 , n76539 );
xnor ( n77786 , n399074 , n395287 );
buf ( n399076 , n77786 );
not ( n399077 , n399076 );
xor ( n77789 , n398019 , n398327 );
xor ( n399079 , n77789 , n398780 );
not ( n399080 , n399079 );
buf ( n399081 , n399080 );
not ( n77793 , n399081 );
or ( n77794 , n399077 , n77793 );
buf ( n399084 , n397714 );
not ( n399085 , n399084 );
and ( n77797 , n397686 , n397704 );
not ( n399087 , n397686 );
and ( n399088 , n399087 , n397705 );
nor ( n77800 , n77797 , n399088 );
buf ( n399090 , n77800 );
not ( n399091 , n399090 );
or ( n77803 , n399085 , n399091 );
buf ( n399093 , n397714 );
buf ( n399094 , n77800 );
or ( n399095 , n399093 , n399094 );
nand ( n399096 , n77803 , n399095 );
buf ( n399097 , n399096 );
buf ( n399098 , n399097 );
not ( n399099 , n398442 );
not ( n77811 , n379445 );
and ( n399101 , n399099 , n77811 );
not ( n77813 , n379274 );
not ( n399103 , n366077 );
or ( n399104 , n77813 , n399103 );
buf ( n399105 , n50871 );
buf ( n399106 , n379271 );
nand ( n399107 , n399105 , n399106 );
buf ( n399108 , n399107 );
nand ( n77819 , n399104 , n399108 );
and ( n399110 , n77819 , n379299 );
nor ( n399111 , n399101 , n399110 );
not ( n77822 , n362063 );
not ( n77823 , n395432 );
and ( n399114 , n77822 , n77823 );
buf ( n399115 , n377094 );
not ( n77826 , n399115 );
buf ( n399117 , n44634 );
not ( n399118 , n399117 );
or ( n399119 , n77826 , n399118 );
buf ( n399120 , n45455 );
buf ( n399121 , n56687 );
nand ( n77832 , n399120 , n399121 );
buf ( n399123 , n77832 );
buf ( n399124 , n399123 );
nand ( n399125 , n399119 , n399124 );
buf ( n399126 , n399125 );
and ( n399127 , n362027 , n399126 );
nor ( n399128 , n399114 , n399127 );
xor ( n77839 , n399111 , n399128 );
buf ( n399130 , n361603 );
not ( n399131 , n399130 );
buf ( n399132 , n378856 );
buf ( n399133 , n44717 );
and ( n77844 , n399132 , n399133 );
not ( n77845 , n399132 );
buf ( n77846 , n366096 );
and ( n399137 , n77845 , n77846 );
nor ( n77848 , n77844 , n399137 );
buf ( n77849 , n77848 );
buf ( n399140 , n77849 );
not ( n77851 , n399140 );
and ( n399142 , n399131 , n77851 );
not ( n399143 , n50987 );
nor ( n77854 , n399143 , n398402 );
buf ( n399145 , n77854 );
nor ( n77856 , n399142 , n399145 );
buf ( n399147 , n77856 );
and ( n77858 , n77839 , n399147 );
and ( n77859 , n399111 , n399128 );
or ( n399150 , n77858 , n77859 );
buf ( n399151 , n399150 );
not ( n399152 , n399151 );
buf ( n399153 , n399152 );
not ( n77864 , n399153 );
buf ( n77865 , n396073 );
buf ( n77866 , n395453 );
xor ( n77867 , n77865 , n77866 );
buf ( n399158 , n395486 );
xnor ( n399159 , n77867 , n399158 );
buf ( n399160 , n399159 );
buf ( n399161 , n399160 );
not ( n399162 , n399161 );
buf ( n399163 , n399162 );
not ( n77874 , n399163 );
or ( n399165 , n77864 , n77874 );
not ( n399166 , n399160 );
not ( n77877 , n399150 );
or ( n399168 , n399166 , n77877 );
xor ( n399169 , n396156 , n396194 );
xor ( n77880 , n399169 , n396310 );
buf ( n399171 , n77880 );
buf ( n399172 , n399171 );
xor ( n77883 , n397583 , n397609 );
xor ( n399174 , n77883 , n397623 );
buf ( n399175 , n399174 );
buf ( n399176 , n399175 );
buf ( n399177 , n369374 );
not ( n77888 , n399177 );
buf ( n399179 , n366659 );
not ( n77890 , n399179 );
or ( n399181 , n77888 , n77890 );
buf ( n77892 , n378135 );
buf ( n77893 , n49178 );
nand ( n77894 , n77892 , n77893 );
buf ( n399185 , n77894 );
buf ( n399186 , n399185 );
nand ( n399187 , n399181 , n399186 );
buf ( n399188 , n399187 );
buf ( n399189 , n399188 );
not ( n399190 , n399189 );
not ( n399191 , n366708 );
buf ( n399192 , n399191 );
not ( n399193 , n399192 );
or ( n399194 , n399190 , n399193 );
buf ( n399195 , n397654 );
buf ( n399196 , n46463 );
nand ( n399197 , n399195 , n399196 );
buf ( n399198 , n399197 );
buf ( n399199 , n399198 );
nand ( n399200 , n399194 , n399199 );
buf ( n399201 , n399200 );
buf ( n399202 , n399201 );
xor ( n399203 , n399176 , n399202 );
buf ( n399204 , n365390 );
not ( n77901 , n399204 );
buf ( n399206 , n396004 );
not ( n77903 , n399206 );
or ( n399208 , n77901 , n77903 );
buf ( n399209 , n76415 );
buf ( n399210 , n365387 );
nand ( n399211 , n399209 , n399210 );
buf ( n399212 , n399211 );
buf ( n399213 , n399212 );
nand ( n77909 , n399208 , n399213 );
buf ( n399215 , n77909 );
buf ( n399216 , n399215 );
not ( n77912 , n399216 );
buf ( n399218 , n365021 );
not ( n77914 , n399218 );
or ( n399220 , n77912 , n77914 );
buf ( n399221 , n397596 );
buf ( n399222 , n365108 );
nand ( n399223 , n399221 , n399222 );
buf ( n399224 , n399223 );
buf ( n399225 , n399224 );
nand ( n399226 , n399220 , n399225 );
buf ( n399227 , n399226 );
buf ( n399228 , n399227 );
buf ( n399229 , n75326 );
buf ( n399230 , n396897 );
buf ( n399231 , n396424 );
xnor ( n399232 , n399230 , n399231 );
buf ( n399233 , n399232 );
buf ( n399234 , n399233 );
xor ( n399235 , n399229 , n399234 );
buf ( n399236 , n399235 );
buf ( n399237 , n399236 );
xor ( n399238 , n399228 , n399237 );
buf ( n399239 , n365152 );
not ( n77935 , n399239 );
buf ( n399241 , n75285 );
not ( n399242 , n399241 );
or ( n77938 , n77935 , n399242 );
buf ( n399244 , n395497 );
not ( n77940 , n399244 );
buf ( n399246 , n381266 );
not ( n399247 , n399246 );
or ( n399248 , n77940 , n399247 );
buf ( n399249 , n351160 );
buf ( n399250 , n45050 );
nand ( n399251 , n399249 , n399250 );
buf ( n399252 , n399251 );
buf ( n399253 , n399252 );
nand ( n399254 , n399248 , n399253 );
buf ( n399255 , n399254 );
buf ( n399256 , n399255 );
buf ( n399257 , n365183 );
nand ( n77953 , n399256 , n399257 );
buf ( n399259 , n77953 );
buf ( n399260 , n399259 );
nand ( n77956 , n77938 , n399260 );
buf ( n77957 , n77956 );
buf ( n399263 , n77957 );
and ( n77959 , n399238 , n399263 );
and ( n399265 , n399228 , n399237 );
or ( n77961 , n77959 , n399265 );
buf ( n399267 , n77961 );
buf ( n399268 , n399267 );
and ( n399269 , n399203 , n399268 );
and ( n77965 , n399176 , n399202 );
or ( n399271 , n399269 , n77965 );
buf ( n399272 , n399271 );
buf ( n399273 , n399272 );
buf ( n399274 , n369444 );
not ( n399275 , n399274 );
buf ( n399276 , n75879 );
not ( n399277 , n399276 );
or ( n77973 , n399275 , n399277 );
buf ( n399279 , n368549 );
not ( n399280 , n399279 );
buf ( n399281 , n365259 );
not ( n77977 , n399281 );
or ( n399283 , n399280 , n77977 );
buf ( n399284 , n352209 );
buf ( n399285 , n380424 );
nand ( n77981 , n399284 , n399285 );
buf ( n399287 , n77981 );
buf ( n399288 , n399287 );
nand ( n77984 , n399283 , n399288 );
buf ( n399290 , n77984 );
buf ( n399291 , n399290 );
buf ( n399292 , n368608 );
nand ( n77988 , n399291 , n399292 );
buf ( n399294 , n77988 );
buf ( n399295 , n399294 );
nand ( n399296 , n77973 , n399295 );
buf ( n399297 , n399296 );
buf ( n399298 , n399297 );
xor ( n77994 , n399273 , n399298 );
buf ( n399300 , n396913 );
not ( n399301 , n399300 );
buf ( n399302 , n396352 );
not ( n399303 , n399302 );
or ( n399304 , n399301 , n399303 );
buf ( n399305 , n396355 );
buf ( n399306 , n75771 );
nand ( n399307 , n399305 , n399306 );
buf ( n399308 , n399307 );
buf ( n399309 , n399308 );
nand ( n399310 , n399304 , n399309 );
buf ( n399311 , n399310 );
xor ( n78007 , n399311 , n396966 );
buf ( n399313 , n78007 );
and ( n399314 , n77994 , n399313 );
and ( n78010 , n399273 , n399298 );
or ( n78011 , n399314 , n78010 );
buf ( n399317 , n78011 );
buf ( n78013 , n399317 );
xor ( n78014 , n399172 , n78013 );
buf ( n399320 , n396904 );
not ( n399321 , n399320 );
buf ( n399322 , n396396 );
not ( n399323 , n399322 );
and ( n399324 , n399321 , n399323 );
buf ( n399325 , n396904 );
buf ( n399326 , n396396 );
and ( n399327 , n399325 , n399326 );
nor ( n399328 , n399324 , n399327 );
buf ( n399329 , n399328 );
buf ( n399330 , n399329 );
buf ( n399331 , n396418 );
and ( n78027 , n399330 , n399331 );
not ( n399333 , n399330 );
buf ( n399334 , n396415 );
and ( n78030 , n399333 , n399334 );
nor ( n399336 , n78027 , n78030 );
buf ( n399337 , n399336 );
not ( n78033 , n399337 );
buf ( n399339 , n377353 );
not ( n399340 , n399339 );
buf ( n399341 , n63905 );
not ( n78037 , n399341 );
or ( n78038 , n399340 , n78037 );
buf ( n399344 , n378956 );
buf ( n399345 , n377352 );
nand ( n78041 , n399344 , n399345 );
buf ( n399347 , n78041 );
buf ( n399348 , n399347 );
nand ( n78044 , n78038 , n399348 );
buf ( n399350 , n78044 );
buf ( n399351 , n399350 );
not ( n399352 , n399351 );
buf ( n399353 , n366399 );
not ( n78049 , n399353 );
or ( n399355 , n399352 , n78049 );
buf ( n399356 , n75222 );
not ( n78052 , n399356 );
buf ( n399358 , n377171 );
nand ( n399359 , n78052 , n399358 );
buf ( n399360 , n399359 );
buf ( n399361 , n399360 );
nand ( n78057 , n399355 , n399361 );
buf ( n399363 , n78057 );
buf ( n399364 , n399363 );
not ( n78060 , n399364 );
buf ( n399366 , n77365 );
not ( n399367 , n399366 );
buf ( n399368 , n365076 );
not ( n78064 , n399368 );
and ( n78065 , n399367 , n78064 );
buf ( n399371 , n380497 );
buf ( n399372 , n31231 );
and ( n399373 , n399371 , n399372 );
not ( n78069 , n399371 );
buf ( n399375 , n382496 );
and ( n78071 , n78069 , n399375 );
nor ( n399377 , n399373 , n78071 );
buf ( n399378 , n399377 );
buf ( n399379 , n399378 );
buf ( n399380 , n44913 );
nor ( n399381 , n399379 , n399380 );
buf ( n399382 , n399381 );
buf ( n399383 , n399382 );
nor ( n399384 , n78065 , n399383 );
buf ( n399385 , n399384 );
buf ( n399386 , n399385 );
nand ( n78082 , n78060 , n399386 );
buf ( n78083 , n78082 );
not ( n399389 , n78083 );
or ( n399390 , n78033 , n399389 );
buf ( n399391 , n399385 );
not ( n399392 , n399391 );
buf ( n399393 , n399363 );
nand ( n78089 , n399392 , n399393 );
buf ( n399395 , n78089 );
nand ( n399396 , n399390 , n399395 );
buf ( n399397 , n399396 );
buf ( n399398 , n48502 );
not ( n78094 , n365915 );
not ( n399400 , n377146 );
and ( n399401 , n78094 , n399400 );
buf ( n399402 , n362423 );
buf ( n399403 , n377146 );
and ( n399404 , n399402 , n399403 );
buf ( n399405 , n399404 );
nor ( n78101 , n399401 , n399405 );
buf ( n399407 , n78101 );
or ( n399408 , n399398 , n399407 );
buf ( n399409 , n396996 );
not ( n78105 , n399409 );
buf ( n399411 , n78105 );
buf ( n399412 , n399411 );
buf ( n399413 , n362385 );
or ( n78109 , n399412 , n399413 );
nand ( n399415 , n399408 , n78109 );
buf ( n399416 , n399415 );
buf ( n399417 , n399416 );
xor ( n78113 , n399397 , n399417 );
buf ( n78114 , n397190 );
not ( n78115 , n78114 );
buf ( n399421 , n398503 );
not ( n399422 , n399421 );
or ( n78118 , n78115 , n399422 );
buf ( n399424 , n398363 );
not ( n399425 , n399424 );
buf ( n399426 , n366131 );
not ( n78122 , n399426 );
or ( n399428 , n399425 , n78122 );
buf ( n399429 , n364858 );
buf ( n399430 , n377592 );
nand ( n78126 , n399429 , n399430 );
buf ( n399432 , n78126 );
buf ( n78128 , n399432 );
nand ( n399434 , n399428 , n78128 );
buf ( n399435 , n399434 );
buf ( n399436 , n399435 );
buf ( n399437 , n57530 );
nand ( n78133 , n399436 , n399437 );
buf ( n399439 , n78133 );
buf ( n399440 , n399439 );
nand ( n78136 , n78118 , n399440 );
buf ( n399442 , n78136 );
buf ( n399443 , n399442 );
and ( n78139 , n78113 , n399443 );
and ( n78140 , n399397 , n399417 );
or ( n78141 , n78139 , n78140 );
buf ( n399447 , n78141 );
buf ( n399448 , n399447 );
and ( n78144 , n78014 , n399448 );
and ( n78145 , n399172 , n78013 );
or ( n78146 , n78144 , n78145 );
buf ( n399452 , n78146 );
nand ( n78148 , n399168 , n399452 );
nand ( n78149 , n399165 , n78148 );
buf ( n399455 , n78149 );
buf ( n399456 , n396079 );
buf ( n399457 , n397062 );
xor ( n399458 , n399456 , n399457 );
buf ( n399459 , n397055 );
xor ( n399460 , n399458 , n399459 );
buf ( n399461 , n399460 );
buf ( n399462 , n399461 );
xor ( n399463 , n399455 , n399462 );
xor ( n78159 , n398383 , n398390 );
xor ( n78160 , n78159 , n398413 );
buf ( n399466 , n78160 );
buf ( n399467 , n399466 );
not ( n399468 , n399467 );
buf ( n399469 , n58923 );
not ( n399470 , n399469 );
buf ( n399471 , n77290 );
not ( n78167 , n399471 );
or ( n78168 , n399470 , n78167 );
buf ( n399474 , n379371 );
not ( n399475 , n399474 );
buf ( n399476 , n369343 );
not ( n399477 , n399476 );
or ( n399478 , n399475 , n399477 );
buf ( n399479 , n367459 );
buf ( n399480 , n379380 );
nand ( n399481 , n399479 , n399480 );
buf ( n399482 , n399481 );
buf ( n399483 , n399482 );
nand ( n399484 , n399478 , n399483 );
buf ( n399485 , n399484 );
buf ( n399486 , n399485 );
buf ( n399487 , n58871 );
nand ( n399488 , n399486 , n399487 );
buf ( n399489 , n399488 );
buf ( n399490 , n399489 );
nand ( n399491 , n78168 , n399490 );
buf ( n399492 , n399491 );
buf ( n399493 , n399492 );
not ( n78189 , n399493 );
or ( n399495 , n399468 , n78189 );
or ( n399496 , n399466 , n399492 );
not ( n78192 , n397049 );
not ( n399498 , n397042 );
not ( n78194 , n399498 );
or ( n399500 , n78192 , n78194 );
nand ( n399501 , n397042 , n75196 );
nand ( n399502 , n399500 , n399501 );
and ( n78198 , n399502 , n396334 );
not ( n399504 , n399502 );
and ( n78200 , n399504 , n397047 );
nor ( n399506 , n78198 , n78200 );
not ( n399507 , n399506 );
nand ( n399508 , n399496 , n399507 );
buf ( n399509 , n399508 );
nand ( n399510 , n399495 , n399509 );
buf ( n399511 , n399510 );
buf ( n399512 , n399511 );
and ( n78208 , n399463 , n399512 );
and ( n399514 , n399455 , n399462 );
or ( n399515 , n78208 , n399514 );
buf ( n399516 , n399515 );
buf ( n399517 , n399516 );
xor ( n399518 , n399098 , n399517 );
xor ( n78214 , n398357 , n398418 );
xor ( n78215 , n78214 , n398524 );
buf ( n399521 , n78215 );
buf ( n399522 , n399521 );
xor ( n78218 , n398557 , n398561 );
xor ( n78219 , n78218 , n398587 );
buf ( n399525 , n78219 );
buf ( n399526 , n399525 );
xor ( n399527 , n399522 , n399526 );
buf ( n399528 , n380407 );
not ( n78224 , n399528 );
buf ( n78225 , n380368 );
not ( n78226 , n78225 );
buf ( n399532 , n363362 );
not ( n399533 , n399532 );
or ( n78229 , n78226 , n399533 );
buf ( n399535 , n42149 );
buf ( n399536 , n380364 );
nand ( n78232 , n399535 , n399536 );
buf ( n399538 , n78232 );
buf ( n399539 , n399538 );
nand ( n399540 , n78229 , n399539 );
buf ( n399541 , n399540 );
buf ( n399542 , n399541 );
not ( n399543 , n399542 );
or ( n399544 , n78224 , n399543 );
buf ( n399545 , n77097 );
buf ( n399546 , n380356 );
nand ( n399547 , n399545 , n399546 );
buf ( n399548 , n399547 );
buf ( n399549 , n399548 );
nand ( n78245 , n399544 , n399549 );
buf ( n399551 , n78245 );
not ( n399552 , n399551 );
buf ( n399553 , n77232 );
buf ( n399554 , n398450 );
xor ( n78250 , n399553 , n399554 );
buf ( n399556 , n398428 );
xor ( n78252 , n78250 , n399556 );
buf ( n399558 , n78252 );
not ( n399559 , n399558 );
or ( n78255 , n399552 , n399559 );
buf ( n399561 , n399551 );
buf ( n399562 , n399558 );
nor ( n399563 , n399561 , n399562 );
buf ( n399564 , n399563 );
xor ( n78260 , n396973 , n397005 );
xor ( n78261 , n78260 , n397038 );
buf ( n399567 , n78261 );
buf ( n399568 , n399567 );
buf ( n399569 , n379916 );
not ( n78265 , n399569 );
buf ( n399571 , n379838 );
not ( n399572 , n399571 );
buf ( n399573 , n42448 );
not ( n78269 , n399573 );
or ( n78270 , n399572 , n78269 );
buf ( n399576 , n361717 );
buf ( n78272 , n379847 );
nand ( n78273 , n399576 , n78272 );
buf ( n399579 , n78273 );
buf ( n399580 , n399579 );
nand ( n78276 , n78270 , n399580 );
buf ( n399582 , n78276 );
buf ( n399583 , n399582 );
not ( n78279 , n399583 );
or ( n78280 , n78265 , n78279 );
buf ( n399586 , n398747 );
buf ( n399587 , n379890 );
nand ( n78283 , n399586 , n399587 );
buf ( n399589 , n78283 );
buf ( n399590 , n399589 );
nand ( n78286 , n78280 , n399590 );
buf ( n399592 , n78286 );
buf ( n399593 , n399592 );
xor ( n399594 , n399568 , n399593 );
buf ( n399595 , n49609 );
not ( n399596 , n399595 );
buf ( n399597 , n398472 );
not ( n78293 , n399597 );
or ( n399599 , n399596 , n78293 );
buf ( n399600 , n393883 );
not ( n78296 , n399600 );
buf ( n399602 , n44638 );
not ( n399603 , n399602 );
or ( n78299 , n78296 , n399603 );
buf ( n399605 , n365561 );
buf ( n399606 , n369763 );
nand ( n78302 , n399605 , n399606 );
buf ( n399608 , n78302 );
buf ( n399609 , n399608 );
nand ( n78305 , n78299 , n399609 );
buf ( n399611 , n78305 );
buf ( n399612 , n399611 );
buf ( n399613 , n369804 );
nand ( n78309 , n399612 , n399613 );
buf ( n399615 , n78309 );
buf ( n399616 , n399615 );
nand ( n399617 , n399599 , n399616 );
buf ( n399618 , n399617 );
buf ( n399619 , n399618 );
buf ( n399620 , n362005 );
not ( n78316 , n399620 );
buf ( n399622 , n366086 );
nand ( n399623 , n78316 , n399622 );
buf ( n399624 , n399623 );
buf ( n399625 , n399624 );
buf ( n399626 , n378098 );
and ( n399627 , n399625 , n399626 );
buf ( n399628 , n362005 );
not ( n399629 , n399628 );
buf ( n399630 , n45908 );
not ( n78326 , n399630 );
or ( n399632 , n399629 , n78326 );
buf ( n399633 , n41892 );
nand ( n78329 , n399632 , n399633 );
buf ( n399635 , n78329 );
buf ( n399636 , n399635 );
nor ( n78332 , n399627 , n399636 );
buf ( n399638 , n78332 );
buf ( n399639 , n399638 );
xor ( n399640 , n399619 , n399639 );
not ( n399641 , n367759 );
buf ( n399642 , n58984 );
not ( n399643 , n399642 );
buf ( n399644 , n41772 );
not ( n78340 , n399644 );
or ( n78341 , n399643 , n78340 );
buf ( n399647 , n47554 );
buf ( n399648 , n379482 );
nand ( n78344 , n399647 , n399648 );
buf ( n399650 , n78344 );
buf ( n399651 , n399650 );
nand ( n399652 , n78341 , n399651 );
buf ( n399653 , n399652 );
not ( n399654 , n399653 );
or ( n78350 , n399641 , n399654 );
or ( n399656 , n398713 , n41836 );
nand ( n78352 , n78350 , n399656 );
buf ( n399658 , n78352 );
and ( n78354 , n399640 , n399658 );
and ( n399660 , n399619 , n399639 );
or ( n399661 , n78354 , n399660 );
buf ( n399662 , n399661 );
buf ( n399663 , n399662 );
and ( n78359 , n399594 , n399663 );
and ( n78360 , n399568 , n399593 );
or ( n78361 , n78359 , n78360 );
buf ( n399667 , n78361 );
buf ( n399668 , n399667 );
not ( n399669 , n399668 );
buf ( n399670 , n399669 );
or ( n399671 , n399564 , n399670 );
nand ( n78367 , n78255 , n399671 );
buf ( n399673 , n78367 );
and ( n78369 , n399527 , n399673 );
and ( n399675 , n399522 , n399526 );
or ( n78371 , n78369 , n399675 );
buf ( n399677 , n78371 );
buf ( n399678 , n399677 );
and ( n78374 , n399518 , n399678 );
and ( n399680 , n399098 , n399517 );
or ( n399681 , n78374 , n399680 );
buf ( n399682 , n399681 );
not ( n399683 , n399682 );
not ( n399684 , n74248 );
nand ( n78380 , n73291 , n73117 );
nand ( n399686 , n78380 , n73295 );
not ( n399687 , n399686 );
and ( n78383 , n399684 , n399687 );
nand ( n399689 , n78380 , n73295 );
and ( n78385 , n74248 , n399689 );
nor ( n78386 , n78383 , n78385 );
not ( n399692 , n73455 );
and ( n399693 , n78386 , n399692 );
not ( n78389 , n78386 );
and ( n399695 , n78389 , n73455 );
nor ( n399696 , n399693 , n399695 );
buf ( n399697 , n399696 );
buf ( n399698 , n397075 );
not ( n399699 , n399698 );
buf ( n399700 , n397732 );
not ( n78396 , n399700 );
or ( n78397 , n399699 , n78396 );
buf ( n399703 , n397500 );
buf ( n78399 , n397072 );
nand ( n78400 , n399703 , n78399 );
buf ( n399706 , n78400 );
buf ( n399707 , n399706 );
nand ( n399708 , n78397 , n399707 );
buf ( n399709 , n399708 );
buf ( n399710 , n399709 );
buf ( n399711 , n397725 );
and ( n399712 , n399710 , n399711 );
not ( n78408 , n399710 );
buf ( n399714 , n397725 );
not ( n399715 , n399714 );
buf ( n399716 , n399715 );
buf ( n399717 , n399716 );
and ( n399718 , n78408 , n399717 );
nor ( n399719 , n399712 , n399718 );
buf ( n399720 , n399719 );
buf ( n399721 , n399720 );
not ( n399722 , n399721 );
buf ( n399723 , n399722 );
buf ( n399724 , n399723 );
nand ( n399725 , n399697 , n399724 );
buf ( n399726 , n399725 );
not ( n78422 , n399726 );
or ( n78423 , n399683 , n78422 );
buf ( n399729 , n399696 );
not ( n399730 , n399729 );
buf ( n399731 , n399730 );
buf ( n399732 , n399731 );
buf ( n399733 , n399720 );
nand ( n399734 , n399732 , n399733 );
buf ( n399735 , n399734 );
nand ( n78431 , n78423 , n399735 );
buf ( n399737 , n78431 );
buf ( n399738 , n399737 );
nand ( n399739 , n77794 , n399738 );
buf ( n399740 , n399739 );
buf ( n399741 , n399740 );
buf ( n399742 , n77786 );
not ( n399743 , n399742 );
buf ( n399744 , n399079 );
nand ( n399745 , n399743 , n399744 );
buf ( n399746 , n399745 );
buf ( n399747 , n399746 );
nand ( n399748 , n399741 , n399747 );
buf ( n399749 , n399748 );
or ( n78445 , n399073 , n399749 );
xor ( n78446 , n64762 , n385447 );
xor ( n78447 , n78446 , n385420 );
buf ( n399753 , n78447 );
and ( n399754 , n385396 , n380356 );
and ( n78450 , n398927 , n380407 );
nor ( n78451 , n399754 , n78450 );
buf ( n399757 , n78451 );
xor ( n399758 , n399753 , n399757 );
buf ( n78454 , n398868 );
not ( n78455 , n78454 );
buf ( n399761 , n78455 );
not ( n399762 , n399761 );
not ( n399763 , n398876 );
and ( n78459 , n399762 , n399763 );
buf ( n399765 , n399761 );
buf ( n399766 , n398876 );
nand ( n399767 , n399765 , n399766 );
buf ( n399768 , n399767 );
and ( n78464 , n399768 , n398855 );
nor ( n399770 , n78459 , n78464 );
buf ( n399771 , n399770 );
xor ( n399772 , n399758 , n399771 );
buf ( n399773 , n399772 );
buf ( n399774 , n399773 );
not ( n399775 , n399774 );
buf ( n399776 , n399775 );
buf ( n399777 , n77604 );
not ( n399778 , n399777 );
not ( n399779 , n398879 );
not ( n78475 , n399779 );
buf ( n399781 , n78475 );
not ( n399782 , n399781 );
or ( n399783 , n399778 , n399782 );
buf ( n399784 , n398940 );
buf ( n399785 , n399779 );
buf ( n399786 , n398899 );
nand ( n78482 , n399785 , n399786 );
buf ( n78483 , n78482 );
buf ( n399789 , n78483 );
nand ( n78485 , n399784 , n399789 );
buf ( n399791 , n78485 );
buf ( n399792 , n399791 );
nand ( n399793 , n399783 , n399792 );
buf ( n399794 , n399793 );
buf ( n399795 , n399794 );
not ( n399796 , n399795 );
buf ( n399797 , n399796 );
xor ( n78493 , n399776 , n399797 );
buf ( n399799 , n77536 );
not ( n78495 , n399799 );
buf ( n399801 , n398812 );
not ( n399802 , n399801 );
or ( n78498 , n78495 , n399802 );
buf ( n399804 , n398832 );
nand ( n78500 , n78498 , n399804 );
buf ( n78501 , n78500 );
buf ( n78502 , n78501 );
buf ( n399808 , n398812 );
not ( n399809 , n399808 );
buf ( n399810 , n398822 );
nand ( n78506 , n399809 , n399810 );
buf ( n399812 , n78506 );
buf ( n399813 , n399812 );
nand ( n78509 , n78502 , n399813 );
buf ( n399815 , n78509 );
xnor ( n78511 , n78493 , n399815 );
buf ( n399817 , n78511 );
xor ( n78513 , n398793 , n398849 );
and ( n399819 , n78513 , n399068 );
and ( n399820 , n398793 , n398849 );
or ( n78516 , n399819 , n399820 );
buf ( n399822 , n78516 );
buf ( n399823 , n399822 );
xor ( n78519 , n399817 , n399823 );
buf ( n399825 , n385511 );
buf ( n78521 , n385523 );
xor ( n78522 , n399825 , n78521 );
buf ( n399828 , n385488 );
xnor ( n399829 , n78522 , n399828 );
buf ( n399830 , n399829 );
not ( n78526 , n399830 );
buf ( n399832 , n385788 );
buf ( n399833 , n385812 );
xor ( n78529 , n399832 , n399833 );
buf ( n399835 , n386158 );
xor ( n399836 , n78529 , n399835 );
buf ( n399837 , n399836 );
not ( n78533 , n399837 );
not ( n399839 , n78533 );
or ( n399840 , n78526 , n399839 );
not ( n78536 , n399830 );
nand ( n78537 , n399837 , n78536 );
nand ( n399843 , n399840 , n78537 );
buf ( n399844 , n399843 );
or ( n78540 , n398809 , n398796 );
nand ( n78541 , n78540 , n398802 );
nand ( n78542 , n398809 , n398796 );
nand ( n399848 , n78541 , n78542 );
buf ( n399849 , n399848 );
xor ( n78545 , n399844 , n399849 );
buf ( n399851 , n78545 );
buf ( n399852 , n399851 );
buf ( n399853 , n398969 );
not ( n399854 , n399853 );
buf ( n399855 , n399854 );
not ( n78551 , n399855 );
not ( n399857 , n77659 );
or ( n399858 , n78551 , n399857 );
not ( n78554 , n398969 );
not ( n399860 , n398947 );
or ( n399861 , n78554 , n399860 );
nand ( n78557 , n399861 , n399058 );
nand ( n399863 , n399858 , n78557 );
buf ( n399864 , n399863 );
xor ( n78560 , n399852 , n399864 );
not ( n78561 , n384584 );
and ( n78562 , n383897 , n63248 );
not ( n78563 , n383897 );
and ( n78564 , n78563 , n383893 );
nor ( n78565 , n78562 , n78564 );
not ( n399871 , n78565 );
or ( n399872 , n78561 , n399871 );
or ( n399873 , n78565 , n384584 );
nand ( n78569 , n399872 , n399873 );
buf ( n399875 , n78569 );
xor ( n399876 , n385285 , n385298 );
xor ( n78572 , n399876 , n385359 );
buf ( n399878 , n78572 );
buf ( n399879 , n399878 );
xor ( n78575 , n399875 , n399879 );
xor ( n399881 , n398988 , n398992 );
and ( n399882 , n399881 , n398998 );
and ( n78578 , n398988 , n398992 );
or ( n78579 , n399882 , n78578 );
buf ( n399885 , n78579 );
buf ( n399886 , n399885 );
xor ( n399887 , n78575 , n399886 );
buf ( n399888 , n399887 );
buf ( n399889 , n399888 );
buf ( n399890 , n399034 );
not ( n78586 , n399890 );
buf ( n399892 , n78586 );
buf ( n399893 , n399892 );
not ( n399894 , n399893 );
buf ( n399895 , n399046 );
not ( n78591 , n399895 );
buf ( n399897 , n78591 );
buf ( n399898 , n399897 );
not ( n78594 , n399898 );
or ( n399900 , n399894 , n78594 );
buf ( n78596 , n77711 );
nand ( n78597 , n399900 , n78596 );
buf ( n78598 , n78597 );
buf ( n78599 , n78598 );
buf ( n399905 , n399892 );
not ( n78601 , n399905 );
buf ( n399907 , n399046 );
nand ( n399908 , n78601 , n399907 );
buf ( n399909 , n399908 );
buf ( n399910 , n399909 );
nand ( n399911 , n78599 , n399910 );
buf ( n399912 , n399911 );
buf ( n399913 , n399912 );
xor ( n78609 , n399889 , n399913 );
xor ( n399915 , n383426 , n383575 );
xor ( n78611 , n399915 , n383740 );
buf ( n399917 , n78611 );
buf ( n78613 , n399917 );
xor ( n399919 , n399014 , n399018 );
and ( n78615 , n399919 , n399032 );
and ( n399921 , n399014 , n399018 );
or ( n399922 , n78615 , n399921 );
buf ( n399923 , n399922 );
buf ( n399924 , n399923 );
xor ( n399925 , n78613 , n399924 );
xor ( n78621 , n398909 , n398912 );
and ( n399927 , n78621 , n398938 );
and ( n78623 , n398909 , n398912 );
or ( n78624 , n399927 , n78623 );
buf ( n399930 , n78624 );
buf ( n399931 , n399930 );
xor ( n78627 , n399925 , n399931 );
buf ( n78628 , n78627 );
buf ( n399934 , n78628 );
xor ( n78630 , n78609 , n399934 );
buf ( n399936 , n78630 );
buf ( n399937 , n399936 );
xor ( n399938 , n78560 , n399937 );
buf ( n399939 , n399938 );
buf ( n399940 , n399939 );
xnor ( n78636 , n78519 , n399940 );
buf ( n399942 , n78636 );
buf ( n399943 , n399070 );
buf ( n399944 , n77494 );
buf ( n399945 , n397750 );
or ( n78641 , n399944 , n399945 );
buf ( n399947 , n78641 );
buf ( n399948 , n399947 );
and ( n399949 , n399943 , n399948 );
and ( n78645 , n397751 , n398784 );
buf ( n399951 , n78645 );
buf ( n78647 , n399951 );
nor ( n78648 , n399949 , n78647 );
buf ( n78649 , n78648 );
nand ( n399955 , n399942 , n78649 );
and ( n399956 , n78445 , n399955 );
not ( n78652 , n399956 );
buf ( n399958 , n398487 );
buf ( n399959 , n398482 );
xor ( n78655 , n399958 , n399959 );
buf ( n399961 , n398513 );
xnor ( n399962 , n78655 , n399961 );
buf ( n399963 , n399962 );
buf ( n399964 , n399963 );
buf ( n399965 , n58871 );
not ( n399966 , n399965 );
buf ( n399967 , n379371 );
not ( n78663 , n399967 );
buf ( n399969 , n41615 );
not ( n399970 , n399969 );
or ( n78666 , n78663 , n399970 );
buf ( n399972 , n361750 );
buf ( n399973 , n379392 );
nand ( n78669 , n399972 , n399973 );
buf ( n78670 , n78669 );
buf ( n399976 , n78670 );
nand ( n78672 , n78666 , n399976 );
buf ( n399978 , n78672 );
buf ( n399979 , n399978 );
not ( n78675 , n399979 );
or ( n399981 , n399966 , n78675 );
buf ( n399982 , n399485 );
buf ( n399983 , n58923 );
nand ( n399984 , n399982 , n399983 );
buf ( n399985 , n399984 );
buf ( n399986 , n399985 );
nand ( n399987 , n399981 , n399986 );
buf ( n399988 , n399987 );
buf ( n399989 , n399988 );
xor ( n78685 , n399964 , n399989 );
and ( n78686 , n368994 , n380923 );
not ( n399992 , n368994 );
and ( n399993 , n399992 , n395541 );
or ( n78689 , n78686 , n399993 );
buf ( n399995 , n78689 );
not ( n78691 , n399995 );
buf ( n399997 , n384501 );
not ( n399998 , n399997 );
or ( n78694 , n78691 , n399998 );
buf ( n400000 , n396369 );
buf ( n400001 , n56794 );
nand ( n400002 , n400000 , n400001 );
buf ( n400003 , n400002 );
buf ( n400004 , n400003 );
nand ( n400005 , n78694 , n400004 );
buf ( n400006 , n400005 );
buf ( n400007 , n400006 );
xor ( n400008 , n395745 , n395864 );
xor ( n400009 , n400008 , n74932 );
xor ( n78705 , n396695 , n396892 );
xor ( n400011 , n400009 , n78705 );
buf ( n400012 , n400011 );
buf ( n400013 , n351345 );
buf ( n400014 , n65349 );
and ( n400015 , n400013 , n400014 );
not ( n78711 , n400013 );
buf ( n400017 , n394065 );
and ( n400018 , n78711 , n400017 );
nor ( n400019 , n400015 , n400018 );
buf ( n400020 , n400019 );
buf ( n400021 , n400020 );
not ( n78717 , n400021 );
buf ( n400023 , n45055 );
not ( n78719 , n400023 );
or ( n400025 , n78717 , n78719 );
buf ( n400026 , n396435 );
not ( n78722 , n400026 );
buf ( n400028 , n365242 );
nand ( n78724 , n78722 , n400028 );
buf ( n400030 , n78724 );
buf ( n400031 , n400030 );
nand ( n78727 , n400025 , n400031 );
buf ( n400033 , n78727 );
buf ( n78729 , n400033 );
xor ( n78730 , n400012 , n78729 );
buf ( n400036 , n395038 );
not ( n400037 , n400036 );
buf ( n400038 , n396004 );
not ( n400039 , n400038 );
or ( n400040 , n400037 , n400039 );
buf ( n400041 , n76415 );
buf ( n78737 , n48458 );
nand ( n78738 , n400041 , n78737 );
buf ( n78739 , n78738 );
buf ( n78740 , n78739 );
nand ( n78741 , n400040 , n78740 );
buf ( n78742 , n78741 );
buf ( n400048 , n78742 );
not ( n400049 , n400048 );
buf ( n400050 , n365021 );
not ( n400051 , n400050 );
or ( n78747 , n400049 , n400051 );
buf ( n400053 , n399215 );
buf ( n400054 , n365108 );
nand ( n400055 , n400053 , n400054 );
buf ( n400056 , n400055 );
buf ( n400057 , n400056 );
nand ( n400058 , n78747 , n400057 );
buf ( n400059 , n400058 );
buf ( n400060 , n400059 );
and ( n78756 , n78730 , n400060 );
and ( n78757 , n400012 , n78729 );
or ( n78758 , n78756 , n78757 );
buf ( n400064 , n78758 );
buf ( n78760 , n400064 );
xor ( n78761 , n400007 , n78760 );
buf ( n400067 , n56970 );
not ( n78763 , n400067 );
buf ( n400069 , n366659 );
not ( n400070 , n400069 );
or ( n78766 , n78763 , n400070 );
buf ( n400072 , n378135 );
buf ( n400073 , n377389 );
nand ( n78769 , n400072 , n400073 );
buf ( n400075 , n78769 );
buf ( n400076 , n400075 );
nand ( n78772 , n78766 , n400076 );
buf ( n400078 , n78772 );
buf ( n400079 , n400078 );
not ( n78775 , n400079 );
buf ( n400081 , n399191 );
not ( n78777 , n400081 );
or ( n78778 , n78775 , n78777 );
buf ( n400084 , n366650 );
not ( n400085 , n400084 );
buf ( n400086 , n399188 );
nand ( n400087 , n400085 , n400086 );
buf ( n400088 , n400087 );
buf ( n400089 , n400088 );
nand ( n78785 , n78778 , n400089 );
buf ( n400091 , n78785 );
buf ( n400092 , n400091 );
and ( n78788 , n78761 , n400092 );
and ( n400094 , n400007 , n78760 );
or ( n78790 , n78788 , n400094 );
buf ( n400096 , n78790 );
buf ( n400097 , n400096 );
buf ( n400098 , n369444 );
not ( n78794 , n400098 );
buf ( n400100 , n399290 );
not ( n400101 , n400100 );
or ( n78797 , n78794 , n400101 );
buf ( n400103 , n380424 );
not ( n400104 , n400103 );
buf ( n400105 , n400104 );
buf ( n400106 , n400105 );
not ( n400107 , n400106 );
buf ( n400108 , n377297 );
not ( n78804 , n400108 );
or ( n400110 , n400107 , n78804 );
buf ( n400111 , n351291 );
buf ( n400112 , n368554 );
nand ( n400113 , n400111 , n400112 );
buf ( n400114 , n400113 );
buf ( n400115 , n400114 );
nand ( n400116 , n400110 , n400115 );
buf ( n400117 , n400116 );
buf ( n400118 , n400117 );
buf ( n400119 , n368608 );
nand ( n78815 , n400118 , n400119 );
buf ( n400121 , n78815 );
buf ( n400122 , n400121 );
nand ( n400123 , n78797 , n400122 );
buf ( n400124 , n400123 );
buf ( n400125 , n400124 );
xor ( n78821 , n400097 , n400125 );
buf ( n400127 , n377757 );
not ( n78823 , n400127 );
buf ( n400129 , n57688 );
not ( n400130 , n400129 );
or ( n78826 , n78823 , n400130 );
buf ( n400132 , n386354 );
buf ( n400133 , n378886 );
nand ( n400134 , n400132 , n400133 );
buf ( n400135 , n400134 );
buf ( n400136 , n400135 );
nand ( n400137 , n78826 , n400136 );
buf ( n400138 , n400137 );
buf ( n400139 , n400138 );
not ( n400140 , n400139 );
buf ( n400141 , n363429 );
not ( n78837 , n400141 );
or ( n400143 , n400140 , n78837 );
buf ( n400144 , n398681 );
buf ( n400145 , n378183 );
nand ( n78841 , n400144 , n400145 );
buf ( n400147 , n78841 );
buf ( n400148 , n400147 );
nand ( n400149 , n400143 , n400148 );
buf ( n400150 , n400149 );
buf ( n400151 , n400150 );
and ( n78847 , n78821 , n400151 );
and ( n400153 , n400097 , n400125 );
or ( n78849 , n78847 , n400153 );
buf ( n400155 , n78849 );
buf ( n78851 , n400155 );
xor ( n78852 , n398663 , n398667 );
xor ( n78853 , n78852 , n398698 );
buf ( n78854 , n78853 );
buf ( n78855 , n78854 );
xor ( n400161 , n78851 , n78855 );
buf ( n400162 , n364852 );
buf ( n400163 , n377068 );
buf ( n400164 , n361534 );
and ( n400165 , n400163 , n400164 );
not ( n400166 , n400163 );
buf ( n400167 , n361531 );
and ( n400168 , n400166 , n400167 );
nor ( n400169 , n400165 , n400168 );
buf ( n400170 , n400169 );
buf ( n400171 , n400170 );
or ( n400172 , n400162 , n400171 );
buf ( n400173 , n77849 );
buf ( n400174 , n361626 );
or ( n400175 , n400173 , n400174 );
nand ( n400176 , n400172 , n400175 );
buf ( n400177 , n400176 );
buf ( n400178 , n400177 );
and ( n400179 , n400161 , n400178 );
and ( n400180 , n78851 , n78855 );
or ( n400181 , n400179 , n400180 );
buf ( n400182 , n400181 );
buf ( n400183 , n400182 );
and ( n400184 , n78685 , n400183 );
and ( n400185 , n399964 , n399989 );
or ( n78858 , n400184 , n400185 );
buf ( n400187 , n78858 );
buf ( n400188 , n400187 );
xor ( n78861 , n398648 , n398703 );
xor ( n400190 , n78861 , n398721 );
buf ( n400191 , n400190 );
buf ( n400192 , n400191 );
buf ( n400193 , n379299 );
not ( n400194 , n400193 );
buf ( n400195 , n379274 );
not ( n400196 , n400195 );
buf ( n400197 , n372201 );
not ( n78870 , n400197 );
or ( n400199 , n400196 , n78870 );
buf ( n400200 , n30912 );
buf ( n400201 , n379271 );
nand ( n78874 , n400200 , n400201 );
buf ( n78875 , n78874 );
buf ( n400204 , n78875 );
nand ( n400205 , n400199 , n400204 );
buf ( n400206 , n400205 );
buf ( n400207 , n400206 );
not ( n78880 , n400207 );
or ( n400209 , n400194 , n78880 );
buf ( n400210 , n379274 );
not ( n78883 , n400210 );
buf ( n400212 , n48496 );
not ( n400213 , n400212 );
or ( n78886 , n78883 , n400213 );
buf ( n400215 , n368700 );
buf ( n400216 , n379271 );
nand ( n400217 , n400215 , n400216 );
buf ( n400218 , n400217 );
buf ( n400219 , n400218 );
nand ( n78892 , n78886 , n400219 );
buf ( n400221 , n78892 );
buf ( n400222 , n400221 );
buf ( n400223 , n379263 );
nand ( n78896 , n400222 , n400223 );
buf ( n400225 , n78896 );
buf ( n400226 , n400225 );
nand ( n400227 , n400209 , n400226 );
buf ( n400228 , n400227 );
not ( n78901 , n400228 );
buf ( n400230 , n371063 );
buf ( n400231 , n378098 );
nand ( n400232 , n400230 , n400231 );
buf ( n400233 , n400232 );
nand ( n400234 , n78901 , n400233 );
not ( n78907 , n400234 );
xor ( n400236 , n399228 , n399237 );
xor ( n78909 , n400236 , n399263 );
buf ( n400238 , n78909 );
buf ( n400239 , n400238 );
buf ( n400240 , n369444 );
not ( n400241 , n400240 );
buf ( n400242 , n400117 );
not ( n78915 , n400242 );
or ( n400244 , n400241 , n78915 );
buf ( n400245 , n400105 );
not ( n78918 , n400245 );
buf ( n400247 , n386837 );
not ( n400248 , n400247 );
or ( n78921 , n78918 , n400248 );
buf ( n400250 , n365440 );
buf ( n400251 , n380424 );
nand ( n78924 , n400250 , n400251 );
buf ( n400253 , n78924 );
buf ( n400254 , n400253 );
nand ( n400255 , n78921 , n400254 );
buf ( n400256 , n400255 );
buf ( n400257 , n400256 );
buf ( n400258 , n368608 );
nand ( n400259 , n400257 , n400258 );
buf ( n400260 , n400259 );
buf ( n400261 , n400260 );
nand ( n400262 , n400244 , n400261 );
buf ( n400263 , n400262 );
buf ( n400264 , n400263 );
xor ( n400265 , n400239 , n400264 );
xor ( n400266 , n400007 , n78760 );
xor ( n400267 , n400266 , n400092 );
buf ( n400268 , n400267 );
buf ( n400269 , n400268 );
and ( n400270 , n400265 , n400269 );
and ( n400271 , n400239 , n400264 );
or ( n400272 , n400270 , n400271 );
buf ( n400273 , n400272 );
not ( n400274 , n400273 );
or ( n400275 , n78907 , n400274 );
buf ( n400276 , n400233 );
not ( n400277 , n400276 );
buf ( n400278 , n400228 );
nand ( n400279 , n400277 , n400278 );
buf ( n400280 , n400279 );
nand ( n78936 , n400275 , n400280 );
buf ( n400282 , n369804 );
not ( n400283 , n400282 );
buf ( n400284 , n393883 );
not ( n78940 , n400284 );
buf ( n400286 , n372382 );
not ( n400287 , n400286 );
or ( n400288 , n78940 , n400287 );
not ( n400289 , n73159 );
buf ( n400290 , n400289 );
buf ( n400291 , n369763 );
nand ( n400292 , n400290 , n400291 );
buf ( n400293 , n400292 );
buf ( n400294 , n400293 );
nand ( n400295 , n400288 , n400294 );
buf ( n400296 , n400295 );
buf ( n400297 , n400296 );
not ( n400298 , n400297 );
or ( n400299 , n400283 , n400298 );
buf ( n400300 , n399611 );
buf ( n400301 , n369809 );
nand ( n400302 , n400300 , n400301 );
buf ( n400303 , n400302 );
buf ( n400304 , n400303 );
nand ( n400305 , n400299 , n400304 );
buf ( n400306 , n400305 );
buf ( n400307 , n400306 );
not ( n400308 , n400307 );
buf ( n400309 , n400308 );
buf ( n400310 , n400309 );
not ( n400311 , n400310 );
buf ( n400312 , n57530 );
not ( n400313 , n400312 );
buf ( n400314 , n398363 );
not ( n400315 , n400314 );
buf ( n400316 , n31073 );
not ( n78950 , n400316 );
or ( n400318 , n400315 , n78950 );
buf ( n400319 , n364827 );
buf ( n400320 , n377592 );
nand ( n400321 , n400319 , n400320 );
buf ( n400322 , n400321 );
buf ( n400323 , n400322 );
nand ( n400324 , n400318 , n400323 );
buf ( n400325 , n400324 );
buf ( n400326 , n400325 );
not ( n78960 , n400326 );
or ( n400328 , n400313 , n78960 );
buf ( n78962 , n399435 );
buf ( n400330 , n397190 );
nand ( n78964 , n78962 , n400330 );
buf ( n400332 , n78964 );
buf ( n400333 , n400332 );
nand ( n78967 , n400328 , n400333 );
buf ( n400335 , n78967 );
buf ( n400336 , n400335 );
not ( n400337 , n400336 );
buf ( n400338 , n400337 );
buf ( n400339 , n400338 );
not ( n400340 , n400339 );
or ( n400341 , n400311 , n400340 );
buf ( n400342 , n399337 );
buf ( n400343 , n399385 );
xor ( n400344 , n400342 , n400343 );
buf ( n400345 , n399363 );
xor ( n400346 , n400344 , n400345 );
buf ( n400347 , n400346 );
buf ( n400348 , n400347 );
not ( n78982 , n400348 );
buf ( n78983 , n78982 );
buf ( n78984 , n78983 );
nand ( n78985 , n400341 , n78984 );
buf ( n78986 , n78985 );
buf ( n78987 , n78986 );
buf ( n400355 , n400335 );
buf ( n400356 , n400306 );
nand ( n400357 , n400355 , n400356 );
buf ( n400358 , n400357 );
buf ( n400359 , n400358 );
nand ( n78993 , n78987 , n400359 );
buf ( n400361 , n78993 );
or ( n78995 , n78936 , n400361 );
xor ( n78996 , n399397 , n399417 );
xor ( n78997 , n78996 , n399443 );
buf ( n400365 , n78997 );
nand ( n78999 , n78995 , n400365 );
buf ( n79000 , n78936 );
buf ( n400368 , n400361 );
nand ( n79002 , n79000 , n400368 );
buf ( n400370 , n79002 );
nand ( n79004 , n78999 , n400370 );
buf ( n400372 , n79004 );
xor ( n400373 , n400192 , n400372 );
not ( n79007 , n379944 );
not ( n400375 , n77819 );
or ( n79009 , n79007 , n400375 );
nand ( n79010 , n400221 , n379299 );
nand ( n400378 , n79009 , n79010 );
buf ( n400379 , n400378 );
buf ( n400380 , n378098 );
not ( n400381 , n400380 );
buf ( n400382 , n365626 );
not ( n79016 , n400382 );
or ( n400384 , n400381 , n79016 );
buf ( n79018 , n45455 );
buf ( n79019 , n379515 );
nand ( n79020 , n79018 , n79019 );
buf ( n79021 , n79020 );
buf ( n79022 , n79021 );
nand ( n79023 , n400384 , n79022 );
buf ( n79024 , n79023 );
buf ( n400392 , n79024 );
not ( n79026 , n400392 );
buf ( n400394 , n364797 );
not ( n79028 , n400394 );
or ( n400396 , n79026 , n79028 );
buf ( n400397 , n41918 );
buf ( n400398 , n399126 );
nand ( n400399 , n400397 , n400398 );
buf ( n400400 , n400399 );
buf ( n400401 , n400400 );
nand ( n400402 , n400396 , n400401 );
buf ( n400403 , n400402 );
buf ( n400404 , n400403 );
xor ( n400405 , n400379 , n400404 );
xor ( n400406 , n399176 , n399202 );
xor ( n79040 , n400406 , n399268 );
buf ( n400408 , n79040 );
buf ( n400409 , n400408 );
buf ( n400410 , n44915 );
not ( n400411 , n400410 );
buf ( n400412 , n399378 );
not ( n79046 , n400412 );
buf ( n400414 , n79046 );
buf ( n400415 , n400414 );
not ( n79049 , n400415 );
or ( n400417 , n400411 , n79049 );
buf ( n400418 , n365041 );
not ( n79052 , n400418 );
buf ( n400420 , n31194 );
not ( n400421 , n400420 );
or ( n79055 , n79052 , n400421 );
buf ( n400423 , n31193 );
buf ( n400424 , n380497 );
nand ( n400425 , n400423 , n400424 );
buf ( n400426 , n400425 );
buf ( n400427 , n400426 );
nand ( n79061 , n79055 , n400427 );
buf ( n400429 , n79061 );
buf ( n400430 , n400429 );
buf ( n400431 , n47466 );
nand ( n400432 , n400430 , n400431 );
buf ( n400433 , n400432 );
buf ( n400434 , n400433 );
nand ( n79068 , n400417 , n400434 );
buf ( n400436 , n79068 );
buf ( n400437 , n400436 );
xor ( n79071 , n396877 , n396883 );
xor ( n400439 , n79071 , n396888 );
buf ( n400440 , n400439 );
buf ( n400441 , n400440 );
xor ( n79075 , n395775 , n395799 );
xor ( n400443 , n79075 , n395845 );
xor ( n400444 , n75720 , n75726 );
xor ( n79078 , n400443 , n400444 );
buf ( n400446 , n73625 );
buf ( n400447 , n380570 );
and ( n79081 , n400446 , n400447 );
buf ( n400449 , n73631 );
buf ( n400450 , n60054 );
and ( n79084 , n400449 , n400450 );
nor ( n79085 , n79081 , n79084 );
buf ( n400453 , n79085 );
buf ( n400454 , n400453 );
buf ( n400455 , n380581 );
or ( n79089 , n400454 , n400455 );
buf ( n400457 , n396492 );
buf ( n400458 , n394774 );
or ( n400459 , n400457 , n400458 );
nand ( n400460 , n79089 , n400459 );
buf ( n400461 , n400460 );
buf ( n400462 , n400461 );
buf ( n400463 , n396615 );
buf ( n400464 , n376866 );
and ( n79098 , n400463 , n400464 );
buf ( n400466 , n396621 );
buf ( n400467 , n382743 );
and ( n400468 , n400466 , n400467 );
nor ( n79102 , n79098 , n400468 );
buf ( n400470 , n79102 );
buf ( n400471 , n400470 );
buf ( n400472 , n376924 );
or ( n400473 , n400471 , n400472 );
buf ( n400474 , n396641 );
buf ( n400475 , n56517 );
or ( n400476 , n400474 , n400475 );
nand ( n400477 , n400473 , n400476 );
buf ( n400478 , n400477 );
buf ( n400479 , n400478 );
nand ( n400480 , n75467 , n56275 );
xnor ( n79114 , n56271 , n400480 );
buf ( n400482 , n79114 );
buf ( n400483 , n376990 );
and ( n79117 , n400482 , n400483 );
buf ( n400485 , n79114 );
not ( n400486 , n400485 );
buf ( n400487 , n400486 );
buf ( n400488 , n400487 );
buf ( n400489 , n376997 );
and ( n79123 , n400488 , n400489 );
buf ( n400491 , n377003 );
nor ( n400492 , n79117 , n79123 , n400491 );
buf ( n400493 , n400492 );
buf ( n400494 , n400493 );
xor ( n400495 , n400479 , n400494 );
not ( n79129 , n376572 );
not ( n79130 , n79129 );
not ( n79131 , n376661 );
or ( n400499 , n79130 , n79131 );
nand ( n400500 , n400499 , n56265 );
not ( n79134 , n376555 );
nand ( n400502 , n79134 , n56268 );
xnor ( n400503 , n400500 , n400502 );
buf ( n400504 , n400503 );
buf ( n400505 , n376990 );
and ( n79139 , n400504 , n400505 );
buf ( n400507 , n400503 );
not ( n400508 , n400507 );
buf ( n400509 , n400508 );
buf ( n400510 , n400509 );
buf ( n400511 , n376997 );
and ( n400512 , n400510 , n400511 );
buf ( n400513 , n377003 );
nor ( n400514 , n79139 , n400512 , n400513 );
buf ( n400515 , n400514 );
buf ( n400516 , n400515 );
buf ( n400517 , n376921 );
not ( n400518 , n400517 );
buf ( n400519 , n79114 );
buf ( n400520 , n376866 );
and ( n79154 , n400519 , n400520 );
buf ( n400522 , n400487 );
buf ( n400523 , n382743 );
and ( n400524 , n400522 , n400523 );
nor ( n79158 , n79154 , n400524 );
buf ( n400526 , n79158 );
buf ( n400527 , n400526 );
not ( n400528 , n400527 );
buf ( n400529 , n400528 );
buf ( n400530 , n400529 );
not ( n79164 , n400530 );
or ( n400532 , n400518 , n79164 );
buf ( n400533 , n400470 );
buf ( n400534 , n56517 );
or ( n400535 , n400533 , n400534 );
nand ( n79169 , n400532 , n400535 );
buf ( n400537 , n79169 );
buf ( n400538 , n400537 );
and ( n79172 , n400516 , n400538 );
buf ( n400540 , n79172 );
buf ( n400541 , n400540 );
and ( n400542 , n400495 , n400541 );
and ( n79176 , n400479 , n400494 );
or ( n79177 , n400542 , n79176 );
buf ( n400545 , n79177 );
buf ( n79179 , n400545 );
xor ( n79180 , n400462 , n79179 );
buf ( n400548 , n382663 );
not ( n400549 , n400548 );
buf ( n400550 , n396787 );
not ( n400551 , n400550 );
buf ( n400552 , n400551 );
buf ( n400553 , n400552 );
not ( n79187 , n400553 );
or ( n400555 , n400549 , n79187 );
buf ( n400556 , n382795 );
buf ( n400557 , n382835 );
and ( n400558 , n400556 , n400557 );
buf ( n400559 , n382803 );
buf ( n400560 , n62243 );
and ( n79194 , n400559 , n400560 );
nor ( n79195 , n400558 , n79194 );
buf ( n400563 , n79195 );
buf ( n400564 , n400563 );
buf ( n400565 , n382849 );
or ( n400566 , n400564 , n400565 );
nand ( n79199 , n400555 , n400566 );
buf ( n400568 , n79199 );
buf ( n400569 , n400568 );
and ( n79202 , n79180 , n400569 );
and ( n400571 , n400462 , n79179 );
or ( n400572 , n79202 , n400571 );
buf ( n400573 , n400572 );
buf ( n400574 , n400573 );
xor ( n400575 , n396497 , n396516 );
xor ( n79205 , n400575 , n396544 );
buf ( n400577 , n79205 );
buf ( n400578 , n400577 );
xor ( n79208 , n400574 , n400578 );
xor ( n79209 , n396804 , n396808 );
xor ( n400581 , n79209 , n396828 );
buf ( n400582 , n400581 );
buf ( n400583 , n400582 );
and ( n79213 , n79208 , n400583 );
and ( n79214 , n400574 , n400578 );
or ( n79215 , n79213 , n79214 );
buf ( n400587 , n79215 );
xor ( n79217 , n79078 , n400587 );
xor ( n79218 , n396779 , n396833 );
xor ( n400590 , n79218 , n396838 );
buf ( n400591 , n400590 );
and ( n79221 , n79217 , n400591 );
and ( n79222 , n79078 , n400587 );
or ( n400594 , n79221 , n79222 );
xor ( n79224 , n396842 , n396845 );
xor ( n79225 , n79224 , n396873 );
and ( n400597 , n400594 , n79225 );
buf ( n400598 , n380838 );
buf ( n400599 , n384343 );
and ( n79229 , n400598 , n400599 );
buf ( n400601 , n380844 );
buf ( n400602 , n384089 );
and ( n79232 , n400601 , n400602 );
nor ( n79233 , n79229 , n79232 );
buf ( n400605 , n79233 );
buf ( n400606 , n400605 );
buf ( n400607 , n384354 );
or ( n79237 , n400606 , n400607 );
buf ( n400609 , n396762 );
buf ( n400610 , n384082 );
or ( n400611 , n400609 , n400610 );
nand ( n79241 , n79237 , n400611 );
buf ( n79242 , n79241 );
xor ( n400614 , n396700 , n396716 );
xor ( n400615 , n400614 , n396735 );
and ( n79245 , n79242 , n400615 );
buf ( n400617 , n63406 );
buf ( n400618 , n382835 );
and ( n79248 , n400617 , n400618 );
buf ( n400620 , n384054 );
buf ( n400621 , n62243 );
and ( n79251 , n400620 , n400621 );
nor ( n400623 , n79248 , n79251 );
buf ( n400624 , n400623 );
buf ( n400625 , n400624 );
buf ( n400626 , n382849 );
or ( n400627 , n400625 , n400626 );
buf ( n400628 , n400563 );
buf ( n400629 , n384157 );
or ( n400630 , n400628 , n400629 );
nand ( n400631 , n400627 , n400630 );
buf ( n400632 , n400631 );
buf ( n400633 , n400632 );
buf ( n400634 , n384380 );
buf ( n400635 , n380817 );
and ( n79265 , n400634 , n400635 );
buf ( n400637 , n384386 );
buf ( n400638 , n57983 );
and ( n79268 , n400637 , n400638 );
nor ( n79269 , n79265 , n79268 );
buf ( n400641 , n79269 );
buf ( n400642 , n400641 );
buf ( n400643 , n60313 );
or ( n400644 , n400642 , n400643 );
buf ( n400645 , n396730 );
buf ( n400646 , n380733 );
or ( n79276 , n400645 , n400646 );
nand ( n79277 , n400644 , n79276 );
buf ( n400649 , n79277 );
buf ( n400650 , n400649 );
xor ( n400651 , n400633 , n400650 );
xor ( n79281 , n400516 , n400538 );
buf ( n400653 , n79281 );
buf ( n400654 , n75451 );
buf ( n400655 , n57800 );
and ( n79285 , n400654 , n400655 );
buf ( n400657 , n396596 );
buf ( n400658 , n376903 );
and ( n79288 , n400657 , n400658 );
nor ( n79289 , n79285 , n79288 );
buf ( n400661 , n79289 );
buf ( n400662 , n400661 );
buf ( n400663 , n378341 );
or ( n400664 , n400662 , n400663 );
buf ( n400665 , n395810 );
buf ( n400666 , n57800 );
and ( n400667 , n400665 , n400666 );
buf ( n400668 , n395816 );
buf ( n400669 , n378284 );
and ( n400670 , n400668 , n400669 );
nor ( n400671 , n400667 , n400670 );
buf ( n400672 , n400671 );
buf ( n400673 , n400672 );
buf ( n400674 , n378424 );
or ( n400675 , n400673 , n400674 );
nand ( n400676 , n400664 , n400675 );
buf ( n400677 , n400676 );
xor ( n400678 , n400653 , n400677 );
buf ( n400679 , n400503 );
buf ( n400680 , n376866 );
and ( n400681 , n400679 , n400680 );
buf ( n400682 , n400509 );
buf ( n400683 , n382743 );
and ( n79299 , n400682 , n400683 );
nor ( n79300 , n400681 , n79299 );
buf ( n400686 , n79300 );
buf ( n400687 , n400686 );
buf ( n400688 , n376924 );
or ( n79304 , n400687 , n400688 );
buf ( n400690 , n400526 );
buf ( n400691 , n56517 );
or ( n79307 , n400690 , n400691 );
nand ( n79308 , n79304 , n79307 );
buf ( n400694 , n79308 );
buf ( n79310 , n400694 );
and ( n400696 , n79129 , n56265 );
xor ( n79312 , n400696 , n376661 );
buf ( n400698 , n79312 );
buf ( n400699 , n376990 );
and ( n400700 , n400698 , n400699 );
buf ( n400701 , n79312 );
not ( n79317 , n400701 );
buf ( n79318 , n79317 );
buf ( n400704 , n79318 );
buf ( n400705 , n376997 );
and ( n400706 , n400704 , n400705 );
buf ( n400707 , n377003 );
nor ( n79323 , n400700 , n400706 , n400707 );
buf ( n79324 , n79323 );
buf ( n400710 , n79324 );
xor ( n79326 , n79310 , n400710 );
buf ( n400712 , n396615 );
buf ( n400713 , n57800 );
and ( n79329 , n400712 , n400713 );
buf ( n400715 , n396621 );
buf ( n400716 , n378284 );
and ( n79332 , n400715 , n400716 );
nor ( n79333 , n79329 , n79332 );
buf ( n400719 , n79333 );
buf ( n400720 , n400719 );
buf ( n400721 , n378341 );
or ( n79337 , n400720 , n400721 );
buf ( n400723 , n400661 );
buf ( n400724 , n378424 );
or ( n79340 , n400723 , n400724 );
nand ( n79341 , n79337 , n79340 );
buf ( n400727 , n79341 );
buf ( n400728 , n400727 );
and ( n400729 , n79326 , n400728 );
and ( n400730 , n79310 , n400710 );
or ( n79346 , n400729 , n400730 );
buf ( n400732 , n79346 );
and ( n400733 , n400678 , n400732 );
and ( n79349 , n400653 , n400677 );
or ( n79350 , n400733 , n79349 );
buf ( n400736 , n79350 );
and ( n400737 , n400651 , n400736 );
and ( n79353 , n400633 , n400650 );
or ( n79354 , n400737 , n79353 );
buf ( n400740 , n79354 );
xor ( n400741 , n396700 , n396716 );
xor ( n400742 , n400741 , n396735 );
and ( n79358 , n400740 , n400742 );
and ( n400744 , n79242 , n400740 );
or ( n79360 , n79245 , n79358 , n400744 );
buf ( n400746 , n79360 );
buf ( n400747 , n73780 );
buf ( n400748 , n380570 );
and ( n400749 , n400747 , n400748 );
buf ( n400750 , n394816 );
buf ( n400751 , n60054 );
and ( n400752 , n400750 , n400751 );
nor ( n400753 , n400749 , n400752 );
buf ( n400754 , n400753 );
buf ( n400755 , n400754 );
buf ( n400756 , n380581 );
or ( n79372 , n400755 , n400756 );
buf ( n400758 , n400453 );
buf ( n400759 , n378453 );
or ( n400760 , n400758 , n400759 );
nand ( n79376 , n79372 , n400760 );
buf ( n79377 , n79376 );
buf ( n400763 , n79377 );
buf ( n400764 , n400672 );
buf ( n400765 , n378341 );
or ( n400766 , n400764 , n400765 );
buf ( n400767 , n75569 );
buf ( n400768 , n378424 );
or ( n79384 , n400767 , n400768 );
nand ( n400770 , n400766 , n79384 );
buf ( n400771 , n400770 );
buf ( n400772 , n400771 );
xor ( n79388 , n400763 , n400772 );
xor ( n400774 , n400479 , n400494 );
xor ( n79390 , n400774 , n400541 );
buf ( n400776 , n79390 );
buf ( n400777 , n400776 );
and ( n400778 , n79388 , n400777 );
and ( n79394 , n400763 , n400772 );
or ( n400780 , n400778 , n79394 );
buf ( n400781 , n400780 );
buf ( n400782 , n400781 );
buf ( n400783 , n378368 );
buf ( n400784 , n394840 );
and ( n79400 , n400783 , n400784 );
buf ( n400786 , n378372 );
buf ( n400787 , n395890 );
and ( n79403 , n400786 , n400787 );
nor ( n400789 , n79400 , n79403 );
buf ( n400790 , n400789 );
buf ( n400791 , n400790 );
buf ( n400792 , n394838 );
or ( n400793 , n400791 , n400792 );
buf ( n400794 , n396748 );
buf ( n400795 , n394835 );
or ( n400796 , n400794 , n400795 );
nand ( n79412 , n400793 , n400796 );
buf ( n400798 , n79412 );
buf ( n400799 , n400798 );
xor ( n79415 , n400782 , n400799 );
buf ( n400801 , n380651 );
buf ( n400802 , n394724 );
and ( n400803 , n400801 , n400802 );
buf ( n400804 , n380657 );
buf ( n400805 , n394730 );
and ( n79421 , n400804 , n400805 );
nor ( n79422 , n400803 , n79421 );
buf ( n400808 , n79422 );
buf ( n400809 , n400808 );
buf ( n400810 , n384414 );
or ( n400811 , n400809 , n400810 );
buf ( n79427 , n75683 );
buf ( n400813 , n395635 );
or ( n400814 , n79427 , n400813 );
nand ( n400815 , n400811 , n400814 );
buf ( n400816 , n400815 );
buf ( n400817 , n400816 );
and ( n79433 , n79415 , n400817 );
and ( n79434 , n400782 , n400799 );
or ( n400820 , n79433 , n79434 );
buf ( n400821 , n400820 );
buf ( n400822 , n400821 );
xor ( n400823 , n400746 , n400822 );
xor ( n400824 , n396739 , n396754 );
xor ( n79440 , n400824 , n396774 );
buf ( n400826 , n79440 );
buf ( n400827 , n400826 );
and ( n79443 , n400823 , n400827 );
and ( n400829 , n400746 , n400822 );
or ( n79445 , n79443 , n400829 );
buf ( n400831 , n79445 );
xor ( n79447 , n79078 , n400587 );
xor ( n79448 , n79447 , n400591 );
and ( n400834 , n400831 , n79448 );
buf ( n400835 , n60089 );
buf ( n400836 , n394840 );
and ( n79452 , n400835 , n400836 );
buf ( n400838 , n60094 );
buf ( n400839 , n395890 );
and ( n400840 , n400838 , n400839 );
nor ( n79456 , n79452 , n400840 );
buf ( n79457 , n79456 );
buf ( n400843 , n79457 );
buf ( n400844 , n394838 );
or ( n400845 , n400843 , n400844 );
buf ( n400846 , n400790 );
buf ( n400847 , n394835 );
or ( n79463 , n400846 , n400847 );
nand ( n400849 , n400845 , n79463 );
buf ( n400850 , n400849 );
buf ( n400851 , n400850 );
buf ( n400852 , n61992 );
buf ( n400853 , n384343 );
and ( n79469 , n400852 , n400853 );
buf ( n400855 , n382596 );
buf ( n400856 , n384089 );
and ( n400857 , n400855 , n400856 );
nor ( n400858 , n79469 , n400857 );
buf ( n400859 , n400858 );
buf ( n400860 , n400859 );
buf ( n400861 , n384354 );
or ( n79477 , n400860 , n400861 );
buf ( n400863 , n400605 );
buf ( n400864 , n384082 );
or ( n400865 , n400863 , n400864 );
nand ( n79481 , n79477 , n400865 );
buf ( n79482 , n79481 );
buf ( n400868 , n79482 );
xor ( n79484 , n400851 , n400868 );
xor ( n400870 , n400763 , n400772 );
xor ( n400871 , n400870 , n400777 );
buf ( n400872 , n400871 );
buf ( n400873 , n400872 );
and ( n79489 , n79484 , n400873 );
and ( n79490 , n400851 , n400868 );
or ( n400876 , n79489 , n79490 );
buf ( n400877 , n400876 );
buf ( n400878 , n400877 );
xor ( n400879 , n400462 , n79179 );
xor ( n400880 , n400879 , n400569 );
buf ( n400881 , n400880 );
buf ( n400882 , n400881 );
xor ( n400883 , n400878 , n400882 );
xor ( n79499 , n400782 , n400799 );
xor ( n79500 , n79499 , n400817 );
buf ( n400886 , n79500 );
buf ( n400887 , n400886 );
and ( n400888 , n400883 , n400887 );
and ( n79504 , n400878 , n400882 );
or ( n79505 , n400888 , n79504 );
buf ( n400891 , n79505 );
xor ( n400892 , n400574 , n400578 );
xor ( n400893 , n400892 , n400583 );
buf ( n400894 , n400893 );
xor ( n79510 , n400891 , n400894 );
xor ( n79511 , n400746 , n400822 );
xor ( n400897 , n79511 , n400827 );
buf ( n400898 , n400897 );
and ( n400899 , n79510 , n400898 );
and ( n79515 , n400891 , n400894 );
or ( n400901 , n400899 , n79515 );
xor ( n79517 , n79078 , n400587 );
xor ( n79518 , n79517 , n400591 );
and ( n400904 , n400901 , n79518 );
and ( n400905 , n400831 , n400901 );
or ( n79521 , n400834 , n400904 , n400905 );
xor ( n400907 , n396842 , n396845 );
xor ( n400908 , n400907 , n396873 );
and ( n79524 , n79521 , n400908 );
and ( n400910 , n400594 , n79521 );
or ( n400911 , n400597 , n79524 , n400910 );
buf ( n400912 , n400911 );
xor ( n400913 , n400441 , n400912 );
buf ( n400914 , n365390 );
not ( n79530 , n400914 );
not ( n400916 , n65349 );
buf ( n400917 , n400916 );
not ( n400918 , n400917 );
or ( n79534 , n79530 , n400918 );
buf ( n400920 , n342879 );
buf ( n400921 , n365387 );
nand ( n79537 , n400920 , n400921 );
buf ( n79538 , n79537 );
buf ( n400924 , n79538 );
nand ( n79540 , n79534 , n400924 );
buf ( n400926 , n79540 );
buf ( n400927 , n400926 );
not ( n400928 , n400927 );
not ( n400929 , n365224 );
buf ( n400930 , n400929 );
not ( n79546 , n400930 );
or ( n79547 , n400928 , n79546 );
buf ( n400933 , n400020 );
buf ( n400934 , n365242 );
nand ( n79550 , n400933 , n400934 );
buf ( n400936 , n79550 );
buf ( n400937 , n400936 );
nand ( n400938 , n79547 , n400937 );
buf ( n400939 , n400938 );
buf ( n400940 , n400939 );
and ( n400941 , n400913 , n400940 );
and ( n400942 , n400441 , n400912 );
or ( n400943 , n400941 , n400942 );
buf ( n400944 , n400943 );
buf ( n400945 , n400944 );
buf ( n400946 , n365152 );
not ( n400947 , n400946 );
buf ( n400948 , n399255 );
not ( n400949 , n400948 );
or ( n400950 , n400947 , n400949 );
buf ( n400951 , n396403 );
not ( n400952 , n400951 );
buf ( n400953 , n364900 );
not ( n400954 , n400953 );
or ( n400955 , n400952 , n400954 );
buf ( n400956 , n75283 );
buf ( n400957 , n352268 );
nand ( n400958 , n400956 , n400957 );
buf ( n400959 , n400958 );
buf ( n400960 , n400959 );
nand ( n400961 , n400955 , n400960 );
buf ( n400962 , n400961 );
buf ( n400963 , n400962 );
buf ( n400964 , n365183 );
nand ( n400965 , n400963 , n400964 );
buf ( n400966 , n400965 );
buf ( n400967 , n400966 );
nand ( n79558 , n400950 , n400967 );
buf ( n400969 , n79558 );
buf ( n400970 , n400969 );
xor ( n79561 , n400945 , n400970 );
buf ( n400972 , n44915 );
not ( n79563 , n400972 );
buf ( n400974 , n400429 );
not ( n400975 , n400974 );
or ( n400976 , n79563 , n400975 );
buf ( n400977 , n365041 );
not ( n400978 , n400977 );
buf ( n400979 , n381220 );
not ( n79570 , n400979 );
or ( n79571 , n400978 , n79570 );
buf ( n79572 , n351195 );
buf ( n400983 , n380497 );
nand ( n79574 , n79572 , n400983 );
buf ( n79575 , n79574 );
buf ( n400986 , n79575 );
nand ( n400987 , n79571 , n400986 );
buf ( n400988 , n400987 );
buf ( n400989 , n400988 );
buf ( n400990 , n47466 );
nand ( n400991 , n400989 , n400990 );
buf ( n400992 , n400991 );
buf ( n400993 , n400992 );
nand ( n400994 , n400976 , n400993 );
buf ( n400995 , n400994 );
buf ( n400996 , n400995 );
and ( n400997 , n79561 , n400996 );
and ( n400998 , n400945 , n400970 );
or ( n400999 , n400997 , n400998 );
buf ( n401000 , n400999 );
buf ( n401001 , n401000 );
xor ( n401002 , n400437 , n401001 );
buf ( n401003 , n50782 );
buf ( n401004 , n378956 );
buf ( n401005 , n377779 );
and ( n401006 , n401004 , n401005 );
buf ( n401007 , n396289 );
buf ( n401008 , n377782 );
and ( n401009 , n401007 , n401008 );
nor ( n79581 , n401006 , n401009 );
buf ( n401011 , n79581 );
buf ( n401012 , n401011 );
or ( n401013 , n401003 , n401012 );
buf ( n79585 , n399350 );
not ( n401015 , n79585 );
buf ( n401016 , n401015 );
buf ( n401017 , n401016 );
buf ( n401018 , n377168 );
or ( n79590 , n401017 , n401018 );
nand ( n401020 , n401013 , n79590 );
buf ( n401021 , n401020 );
buf ( n401022 , n401021 );
and ( n401023 , n401002 , n401022 );
and ( n401024 , n400437 , n401001 );
or ( n79596 , n401023 , n401024 );
buf ( n401026 , n79596 );
buf ( n401027 , n401026 );
xor ( n79599 , n400409 , n401027 );
buf ( n401029 , n42266 );
buf ( n401030 , n377122 );
buf ( n401031 , n365918 );
and ( n401032 , n401030 , n401031 );
not ( n401033 , n401030 );
buf ( n401034 , n365915 );
and ( n401035 , n401033 , n401034 );
nor ( n401036 , n401032 , n401035 );
buf ( n401037 , n401036 );
buf ( n401038 , n401037 );
or ( n401039 , n401029 , n401038 );
buf ( n401040 , n78101 );
buf ( n401041 , n73479 );
or ( n79613 , n401040 , n401041 );
nand ( n79614 , n401039 , n79613 );
buf ( n401044 , n79614 );
buf ( n401045 , n401044 );
and ( n79617 , n79599 , n401045 );
and ( n79618 , n400409 , n401027 );
or ( n79619 , n79617 , n79618 );
buf ( n401049 , n79619 );
buf ( n401050 , n401049 );
and ( n79622 , n400405 , n401050 );
and ( n79623 , n400379 , n400404 );
or ( n79624 , n79622 , n79623 );
buf ( n401054 , n79624 );
buf ( n401055 , n401054 );
and ( n401056 , n400373 , n401055 );
and ( n401057 , n400192 , n400372 );
or ( n79629 , n401056 , n401057 );
buf ( n401059 , n79629 );
buf ( n401060 , n401059 );
xor ( n401061 , n400188 , n401060 );
xor ( n401062 , n398644 , n398726 );
xor ( n401063 , n401062 , n398755 );
buf ( n401064 , n401063 );
buf ( n401065 , n401064 );
and ( n401066 , n401061 , n401065 );
and ( n79638 , n400188 , n401060 );
or ( n79639 , n401066 , n79638 );
buf ( n401069 , n79639 );
buf ( n401070 , n401069 );
xor ( n79642 , n77327 , n398626 );
xor ( n401072 , n79642 , n398760 );
buf ( n401073 , n401072 );
buf ( n401074 , n401073 );
xor ( n79646 , n401070 , n401074 );
xor ( n401076 , n399492 , n399506 );
xor ( n401077 , n401076 , n399466 );
buf ( n401078 , n401077 );
not ( n401079 , n401078 );
buf ( n401080 , n401079 );
not ( n401081 , n401080 );
buf ( n401082 , n399163 );
buf ( n401083 , n399452 );
xor ( n401084 , n401082 , n401083 );
buf ( n401085 , n399153 );
xnor ( n79657 , n401084 , n401085 );
buf ( n401087 , n79657 );
buf ( n401088 , n401087 );
not ( n401089 , n401088 );
buf ( n401090 , n401089 );
not ( n401091 , n401090 );
or ( n79663 , n401081 , n401091 );
not ( n401093 , n401087 );
not ( n401094 , n401077 );
or ( n401095 , n401093 , n401094 );
xor ( n79667 , n399111 , n399128 );
xor ( n79668 , n79667 , n399147 );
buf ( n401098 , n79668 );
not ( n79670 , n401098 );
buf ( n401100 , n79670 );
not ( n401101 , n401100 );
xor ( n79673 , n399172 , n78013 );
xor ( n401103 , n79673 , n399448 );
buf ( n401104 , n401103 );
not ( n401105 , n401104 );
or ( n79677 , n401101 , n401105 );
buf ( n401107 , n401104 );
not ( n79679 , n401107 );
buf ( n79680 , n79679 );
not ( n401110 , n79680 );
not ( n79682 , n79668 );
or ( n401112 , n401110 , n79682 );
xor ( n79684 , n399273 , n399298 );
xor ( n79685 , n79684 , n399313 );
buf ( n401115 , n79685 );
buf ( n401116 , n401115 );
buf ( n401117 , n379890 );
not ( n79689 , n401117 );
buf ( n401119 , n399582 );
not ( n79691 , n401119 );
or ( n79692 , n79689 , n79691 );
buf ( n401122 , n379841 );
not ( n401123 , n401122 );
buf ( n401124 , n362537 );
not ( n401125 , n401124 );
or ( n401126 , n401123 , n401125 );
buf ( n401127 , n362549 );
buf ( n401128 , n398741 );
nand ( n401129 , n401127 , n401128 );
buf ( n401130 , n401129 );
buf ( n401131 , n401130 );
nand ( n401132 , n401126 , n401131 );
buf ( n401133 , n401132 );
buf ( n401134 , n401133 );
buf ( n401135 , n379916 );
nand ( n401136 , n401134 , n401135 );
buf ( n401137 , n401136 );
buf ( n401138 , n401137 );
nand ( n401139 , n79692 , n401138 );
buf ( n401140 , n401139 );
buf ( n401141 , n401140 );
xor ( n79713 , n401116 , n401141 );
xor ( n401143 , n400097 , n400125 );
xor ( n79715 , n401143 , n400151 );
buf ( n401145 , n79715 );
buf ( n401146 , n401145 );
not ( n401147 , n401146 );
buf ( n401148 , n378856 );
not ( n79720 , n401148 );
buf ( n401150 , n367248 );
not ( n401151 , n401150 );
or ( n79723 , n79720 , n401151 );
buf ( n401153 , n364744 );
buf ( n401154 , n378847 );
nand ( n401155 , n401153 , n401154 );
buf ( n401156 , n401155 );
buf ( n401157 , n401156 );
nand ( n401158 , n79723 , n401157 );
buf ( n401159 , n401158 );
buf ( n401160 , n401159 );
not ( n79732 , n401160 );
buf ( n401162 , n367759 );
not ( n401163 , n401162 );
or ( n401164 , n79732 , n401163 );
buf ( n401165 , n399653 );
buf ( n401166 , n41835 );
nand ( n401167 , n401165 , n401166 );
buf ( n401168 , n401167 );
buf ( n401169 , n401168 );
nand ( n79741 , n401164 , n401169 );
buf ( n79742 , n79741 );
buf ( n401172 , n79742 );
not ( n401173 , n401172 );
or ( n79745 , n401147 , n401173 );
buf ( n401175 , n79742 );
buf ( n401176 , n401145 );
or ( n79748 , n401175 , n401176 );
buf ( n401178 , n369374 );
not ( n401179 , n401178 );
buf ( n401180 , n380923 );
not ( n79752 , n401180 );
or ( n401182 , n401179 , n79752 );
buf ( n401183 , n22619 );
buf ( n401184 , n49178 );
nand ( n401185 , n401183 , n401184 );
buf ( n401186 , n401185 );
buf ( n401187 , n401186 );
nand ( n401188 , n401182 , n401187 );
buf ( n401189 , n401188 );
buf ( n401190 , n401189 );
not ( n79762 , n401190 );
buf ( n401192 , n365725 );
not ( n79764 , n401192 );
or ( n79765 , n79762 , n79764 );
buf ( n401195 , n78689 );
buf ( n401196 , n56794 );
nand ( n79768 , n401195 , n401196 );
buf ( n401198 , n79768 );
buf ( n401199 , n401198 );
nand ( n401200 , n79765 , n401199 );
buf ( n401201 , n401200 );
buf ( n401202 , n401201 );
xor ( n401203 , n400012 , n78729 );
xor ( n79775 , n401203 , n400060 );
buf ( n401205 , n79775 );
buf ( n401206 , n401205 );
xor ( n401207 , n401202 , n401206 );
buf ( n401208 , n368994 );
not ( n79780 , n401208 );
buf ( n401210 , n386102 );
not ( n401211 , n401210 );
or ( n79783 , n79780 , n401211 );
buf ( n401213 , n386093 );
buf ( n401214 , n57053 );
nand ( n401215 , n401213 , n401214 );
buf ( n401216 , n401215 );
buf ( n401217 , n401216 );
nand ( n79789 , n79783 , n401217 );
buf ( n401219 , n79789 );
buf ( n401220 , n401219 );
not ( n79792 , n401220 );
buf ( n401222 , n386091 );
not ( n79794 , n401222 );
or ( n401224 , n79792 , n79794 );
buf ( n401225 , n78742 );
buf ( n401226 , n365108 );
nand ( n79798 , n401225 , n401226 );
buf ( n401228 , n79798 );
buf ( n401229 , n401228 );
nand ( n79801 , n401224 , n401229 );
buf ( n401231 , n79801 );
buf ( n401232 , n401231 );
buf ( n401233 , n365149 );
not ( n401234 , n401233 );
buf ( n401235 , n400962 );
not ( n401236 , n401235 );
or ( n401237 , n401234 , n401236 );
buf ( n401238 , n396403 );
not ( n79810 , n401238 );
buf ( n401240 , n60751 );
not ( n79812 , n401240 );
or ( n79813 , n79810 , n79812 );
buf ( n401243 , n396019 );
buf ( n401244 , n342908 );
nand ( n79816 , n401243 , n401244 );
buf ( n401246 , n79816 );
buf ( n401247 , n401246 );
nand ( n401248 , n79813 , n401247 );
buf ( n401249 , n401248 );
buf ( n401250 , n401249 );
buf ( n401251 , n365183 );
nand ( n79823 , n401250 , n401251 );
buf ( n401253 , n79823 );
buf ( n401254 , n401253 );
nand ( n401255 , n401237 , n401254 );
buf ( n401256 , n401255 );
buf ( n401257 , n401256 );
xor ( n401258 , n401232 , n401257 );
xor ( n401259 , n400441 , n400912 );
xor ( n79831 , n401259 , n400940 );
buf ( n401261 , n79831 );
buf ( n401262 , n401261 );
and ( n79834 , n401258 , n401262 );
and ( n79835 , n401232 , n401257 );
or ( n79836 , n79834 , n79835 );
buf ( n401266 , n79836 );
buf ( n401267 , n401266 );
and ( n79839 , n401207 , n401267 );
and ( n79840 , n401202 , n401206 );
or ( n79841 , n79839 , n79840 );
buf ( n401271 , n79841 );
buf ( n401272 , n401271 );
buf ( n401273 , n377143 );
buf ( n401274 , n377683 );
and ( n79846 , n401273 , n401274 );
not ( n79847 , n401273 );
buf ( n401277 , n22769 );
and ( n79849 , n79847 , n401277 );
nor ( n401279 , n79846 , n79849 );
buf ( n401280 , n401279 );
buf ( n401281 , n401280 );
not ( n401282 , n401281 );
buf ( n401283 , n401282 );
buf ( n401284 , n401283 );
not ( n79856 , n401284 );
buf ( n401286 , n363429 );
not ( n401287 , n401286 );
or ( n401288 , n79856 , n401287 );
buf ( n401289 , n400138 );
buf ( n401290 , n43261 );
nand ( n79862 , n401289 , n401290 );
buf ( n401292 , n79862 );
buf ( n401293 , n401292 );
nand ( n79865 , n401288 , n401293 );
buf ( n401295 , n79865 );
buf ( n401296 , n401295 );
xor ( n79868 , n401272 , n401296 );
buf ( n401298 , n377353 );
not ( n79870 , n401298 );
buf ( n401300 , n378138 );
not ( n401301 , n401300 );
or ( n401302 , n79870 , n401301 );
buf ( n401303 , n375901 );
buf ( n401304 , n377352 );
nand ( n79876 , n401303 , n401304 );
buf ( n401306 , n79876 );
buf ( n401307 , n401306 );
nand ( n401308 , n401302 , n401307 );
buf ( n401309 , n401308 );
buf ( n401310 , n401309 );
not ( n401311 , n401310 );
buf ( n401312 , n375896 );
not ( n79884 , n401312 );
or ( n401314 , n401311 , n79884 );
buf ( n401315 , n400078 );
buf ( n401316 , n375920 );
nand ( n79888 , n401315 , n401316 );
buf ( n401318 , n79888 );
buf ( n401319 , n401318 );
nand ( n401320 , n401314 , n401319 );
buf ( n401321 , n401320 );
buf ( n401322 , n401321 );
xor ( n79894 , n400945 , n400970 );
xor ( n401324 , n79894 , n400996 );
buf ( n401325 , n401324 );
buf ( n401326 , n401325 );
xor ( n79898 , n401322 , n401326 );
buf ( n401328 , n50782 );
buf ( n401329 , n377757 );
buf ( n401330 , n396289 );
and ( n79902 , n401329 , n401330 );
not ( n79903 , n401329 );
buf ( n401333 , n56849 );
and ( n401334 , n79903 , n401333 );
nor ( n79906 , n79902 , n401334 );
buf ( n79907 , n79906 );
buf ( n401337 , n79907 );
or ( n401338 , n401328 , n401337 );
buf ( n401339 , n401011 );
buf ( n401340 , n386027 );
or ( n401341 , n401339 , n401340 );
nand ( n401342 , n401338 , n401341 );
buf ( n401343 , n401342 );
buf ( n401344 , n401343 );
and ( n401345 , n79898 , n401344 );
and ( n401346 , n401322 , n401326 );
or ( n79918 , n401345 , n401346 );
buf ( n401348 , n79918 );
buf ( n401349 , n401348 );
and ( n79921 , n79868 , n401349 );
and ( n401351 , n401272 , n401296 );
or ( n401352 , n79921 , n401351 );
buf ( n401353 , n401352 );
buf ( n401354 , n401353 );
nand ( n79926 , n79748 , n401354 );
buf ( n401356 , n79926 );
buf ( n401357 , n401356 );
nand ( n401358 , n79745 , n401357 );
buf ( n401359 , n401358 );
buf ( n401360 , n401359 );
and ( n401361 , n79713 , n401360 );
and ( n79933 , n401116 , n401141 );
or ( n401363 , n401361 , n79933 );
buf ( n401364 , n401363 );
nand ( n79936 , n401112 , n401364 );
nand ( n401366 , n79677 , n79936 );
nand ( n401367 , n401095 , n401366 );
nand ( n79939 , n79663 , n401367 );
buf ( n401369 , n79939 );
xor ( n401370 , n79646 , n401369 );
buf ( n401371 , n401370 );
buf ( n401372 , n401371 );
xor ( n79944 , n400188 , n401060 );
xor ( n79945 , n79944 , n401065 );
buf ( n401375 , n79945 );
xor ( n79947 , n399568 , n399593 );
xor ( n401377 , n79947 , n399663 );
buf ( n401378 , n401377 );
buf ( n401379 , n401378 );
buf ( n401380 , n380356 );
not ( n79952 , n401380 );
buf ( n401382 , n399541 );
not ( n401383 , n401382 );
or ( n79955 , n79952 , n401383 );
buf ( n401385 , n380368 );
not ( n401386 , n401385 );
buf ( n401387 , n362139 );
not ( n79959 , n401387 );
or ( n79960 , n401386 , n79959 );
buf ( n401390 , n362148 );
buf ( n79962 , n384667 );
nand ( n79963 , n401390 , n79962 );
buf ( n401393 , n79963 );
buf ( n401394 , n401393 );
nand ( n401395 , n79960 , n401394 );
buf ( n401396 , n401395 );
buf ( n401397 , n401396 );
buf ( n401398 , n380407 );
nand ( n401399 , n401397 , n401398 );
buf ( n401400 , n401399 );
buf ( n401401 , n401400 );
nand ( n401402 , n79955 , n401401 );
buf ( n401403 , n401402 );
buf ( n401404 , n401403 );
xor ( n401405 , n401379 , n401404 );
buf ( n401406 , n401405 );
buf ( n401407 , n401406 );
xor ( n401408 , n399619 , n399639 );
xor ( n401409 , n401408 , n399658 );
buf ( n401410 , n401409 );
buf ( n401411 , n401410 );
buf ( n401412 , n58923 );
not ( n79984 , n401412 );
buf ( n401414 , n399978 );
not ( n401415 , n401414 );
or ( n79987 , n79984 , n401415 );
buf ( n401417 , n41528 );
not ( n401418 , n401417 );
buf ( n401419 , n379392 );
not ( n401420 , n401419 );
and ( n401421 , n401418 , n401420 );
buf ( n401422 , n361673 );
buf ( n401423 , n379380 );
and ( n79995 , n401422 , n401423 );
nor ( n401425 , n401421 , n79995 );
buf ( n401426 , n401425 );
buf ( n401427 , n401426 );
not ( n79999 , n401427 );
buf ( n401429 , n58871 );
nand ( n80001 , n79999 , n401429 );
buf ( n401431 , n80001 );
buf ( n401432 , n401431 );
nand ( n401433 , n79987 , n401432 );
buf ( n401434 , n401433 );
buf ( n401435 , n401434 );
xor ( n401436 , n401411 , n401435 );
buf ( n401437 , n369809 );
not ( n401438 , n401437 );
buf ( n401439 , n400296 );
not ( n80011 , n401439 );
or ( n80012 , n401438 , n80011 );
buf ( n401442 , n393883 );
not ( n401443 , n401442 );
buf ( n401444 , n365259 );
not ( n80016 , n401444 );
or ( n401446 , n401443 , n80016 );
buf ( n401447 , n352212 );
buf ( n401448 , n369763 );
nand ( n401449 , n401447 , n401448 );
buf ( n401450 , n401449 );
buf ( n401451 , n401450 );
nand ( n401452 , n401446 , n401451 );
buf ( n401453 , n401452 );
buf ( n401454 , n401453 );
buf ( n401455 , n369804 );
nand ( n401456 , n401454 , n401455 );
buf ( n401457 , n401456 );
buf ( n401458 , n401457 );
nand ( n401459 , n80012 , n401458 );
buf ( n401460 , n401459 );
buf ( n401461 , n401460 );
xor ( n401462 , n400437 , n401001 );
xor ( n401463 , n401462 , n401022 );
buf ( n401464 , n401463 );
buf ( n401465 , n401464 );
xor ( n401466 , n401461 , n401465 );
buf ( n401467 , n361531 );
not ( n401468 , n378043 );
not ( n401469 , n41430 );
not ( n401470 , n401469 );
or ( n401471 , n401468 , n401470 );
nand ( n80022 , n401471 , n378098 );
buf ( n401473 , n80022 );
nand ( n401474 , n364744 , n41430 );
buf ( n401475 , n401474 );
and ( n80026 , n401467 , n401473 , n401475 );
buf ( n401477 , n80026 );
buf ( n401478 , n401477 );
and ( n80029 , n401466 , n401478 );
and ( n80030 , n401461 , n401465 );
or ( n80031 , n80029 , n80030 );
buf ( n401482 , n80031 );
buf ( n401483 , n401482 );
not ( n80034 , n401483 );
buf ( n401485 , n361603 );
buf ( n401486 , n56687 );
buf ( n401487 , n363603 );
and ( n80038 , n401486 , n401487 );
not ( n80039 , n401486 );
buf ( n401490 , n361534 );
and ( n80041 , n80039 , n401490 );
nor ( n80042 , n80038 , n80041 );
buf ( n401493 , n80042 );
buf ( n401494 , n401493 );
or ( n80045 , n401485 , n401494 );
buf ( n401496 , n400170 );
buf ( n401497 , n361626 );
or ( n80048 , n401496 , n401497 );
nand ( n80049 , n80045 , n80048 );
buf ( n401500 , n80049 );
buf ( n401501 , n401500 );
not ( n401502 , n401501 );
or ( n80053 , n80034 , n401502 );
buf ( n401504 , n401500 );
buf ( n401505 , n401482 );
or ( n80056 , n401504 , n401505 );
xor ( n401507 , n400409 , n401027 );
xor ( n401508 , n401507 , n401045 );
buf ( n401509 , n401508 );
buf ( n401510 , n401509 );
nand ( n401511 , n80056 , n401510 );
buf ( n401512 , n401511 );
buf ( n401513 , n401512 );
nand ( n80064 , n80053 , n401513 );
buf ( n401515 , n80064 );
buf ( n401516 , n401515 );
and ( n80067 , n401436 , n401516 );
and ( n401518 , n401411 , n401435 );
or ( n401519 , n80067 , n401518 );
buf ( n401520 , n401519 );
buf ( n401521 , n401520 );
xor ( n401522 , n401407 , n401521 );
buf ( n401523 , n401522 );
not ( n80074 , n401523 );
buf ( n401525 , n401364 );
buf ( n401526 , n401104 );
and ( n80077 , n401525 , n401526 );
not ( n401528 , n401525 );
buf ( n401529 , n79680 );
and ( n401530 , n401528 , n401529 );
nor ( n80081 , n80077 , n401530 );
buf ( n401532 , n80081 );
buf ( n401533 , n401532 );
buf ( n401534 , n79668 );
and ( n80085 , n401533 , n401534 );
not ( n401536 , n401533 );
buf ( n401537 , n401100 );
and ( n401538 , n401536 , n401537 );
nor ( n401539 , n80085 , n401538 );
buf ( n401540 , n401539 );
buf ( n401541 , n401540 );
buf ( n401542 , n78983 );
not ( n80093 , n401542 );
buf ( n401544 , n400309 );
not ( n401545 , n401544 );
or ( n80096 , n80093 , n401545 );
buf ( n401547 , n400306 );
buf ( n401548 , n400347 );
nand ( n80099 , n401547 , n401548 );
buf ( n401550 , n80099 );
buf ( n401551 , n401550 );
nand ( n401552 , n80096 , n401551 );
buf ( n401553 , n401552 );
buf ( n401554 , n401553 );
buf ( n401555 , n400338 );
and ( n401556 , n401554 , n401555 );
not ( n80107 , n401554 );
buf ( n401558 , n400335 );
and ( n401559 , n80107 , n401558 );
nor ( n401560 , n401556 , n401559 );
buf ( n401561 , n401560 );
not ( n401562 , n401561 );
buf ( n401563 , n401562 );
not ( n401564 , n401563 );
buf ( n401565 , n400273 );
buf ( n401566 , n400228 );
xor ( n401567 , n401565 , n401566 );
buf ( n401568 , n400233 );
xor ( n401569 , n401567 , n401568 );
buf ( n401570 , n401569 );
buf ( n401571 , n401570 );
not ( n401572 , n401571 );
buf ( n401573 , n401572 );
buf ( n401574 , n401573 );
not ( n401575 , n401574 );
or ( n80126 , n401564 , n401575 );
xor ( n401577 , n400239 , n400264 );
xor ( n401578 , n401577 , n400269 );
buf ( n401579 , n401578 );
buf ( n401580 , n401579 );
buf ( n401581 , n397190 );
not ( n80132 , n401581 );
buf ( n401583 , n400325 );
not ( n401584 , n401583 );
or ( n80135 , n80132 , n401584 );
buf ( n401586 , n398363 );
not ( n401587 , n401586 );
buf ( n401588 , n44638 );
not ( n80139 , n401588 );
or ( n401590 , n401587 , n80139 );
buf ( n401591 , n364804 );
buf ( n401592 , n377592 );
nand ( n80143 , n401591 , n401592 );
buf ( n401594 , n80143 );
buf ( n401595 , n401594 );
nand ( n80146 , n401590 , n401595 );
buf ( n401597 , n80146 );
buf ( n401598 , n401597 );
buf ( n401599 , n57530 );
nand ( n80150 , n401598 , n401599 );
buf ( n401601 , n80150 );
buf ( n401602 , n401601 );
nand ( n401603 , n80135 , n401602 );
buf ( n401604 , n401603 );
buf ( n401605 , n401604 );
xor ( n80156 , n401580 , n401605 );
and ( n401607 , n41772 , n377068 );
not ( n80158 , n41772 );
and ( n80159 , n80158 , n377071 );
or ( n80160 , n401607 , n80159 );
buf ( n401611 , n80160 );
not ( n401612 , n401611 );
buf ( n401613 , n367759 );
not ( n80164 , n401613 );
or ( n401615 , n401612 , n80164 );
buf ( n80166 , n401159 );
buf ( n401617 , n41835 );
nand ( n80168 , n80166 , n401617 );
buf ( n401619 , n80168 );
buf ( n401620 , n401619 );
nand ( n401621 , n401615 , n401620 );
buf ( n401622 , n401621 );
buf ( n401623 , n401622 );
and ( n80174 , n80156 , n401623 );
and ( n80175 , n401580 , n401605 );
or ( n401626 , n80174 , n80175 );
buf ( n401627 , n401626 );
buf ( n401628 , n401627 );
buf ( n401629 , n401570 );
buf ( n401630 , n401561 );
nand ( n80181 , n401629 , n401630 );
buf ( n80182 , n80181 );
buf ( n401633 , n80182 );
nand ( n80184 , n401628 , n401633 );
buf ( n401635 , n80184 );
buf ( n401636 , n401635 );
nand ( n80187 , n80126 , n401636 );
buf ( n401638 , n80187 );
buf ( n401639 , n401638 );
buf ( n401640 , n379916 );
not ( n401641 , n401640 );
buf ( n401642 , n379841 );
not ( n80193 , n401642 );
buf ( n401644 , n52029 );
not ( n401645 , n401644 );
or ( n401646 , n80193 , n401645 );
buf ( n401647 , n50871 );
buf ( n401648 , n398741 );
nand ( n80199 , n401647 , n401648 );
buf ( n401650 , n80199 );
buf ( n401651 , n401650 );
nand ( n80202 , n401646 , n401651 );
buf ( n401653 , n80202 );
buf ( n401654 , n401653 );
not ( n401655 , n401654 );
or ( n401656 , n401641 , n401655 );
buf ( n401657 , n401133 );
buf ( n401658 , n379890 );
nand ( n401659 , n401657 , n401658 );
buf ( n401660 , n401659 );
buf ( n401661 , n401660 );
nand ( n401662 , n401656 , n401661 );
buf ( n401663 , n401662 );
buf ( n401664 , n401663 );
buf ( n401665 , n58984 );
not ( n80216 , n401665 );
buf ( n401667 , n365773 );
not ( n401668 , n401667 );
or ( n80219 , n80216 , n401668 );
buf ( n401670 , n45595 );
buf ( n401671 , n379482 );
nand ( n401672 , n401670 , n401671 );
buf ( n401673 , n401672 );
buf ( n401674 , n401673 );
nand ( n80225 , n80219 , n401674 );
buf ( n401676 , n80225 );
buf ( n401677 , n401676 );
not ( n401678 , n401677 );
buf ( n401679 , n49669 );
not ( n401680 , n401679 );
or ( n401681 , n401678 , n401680 );
buf ( n401682 , n401037 );
not ( n401683 , n401682 );
buf ( n401684 , n48558 );
nand ( n401685 , n401683 , n401684 );
buf ( n401686 , n401685 );
buf ( n401687 , n401686 );
nand ( n80238 , n401681 , n401687 );
buf ( n401689 , n80238 );
not ( n401690 , n401689 );
buf ( n401691 , n379263 );
not ( n401692 , n401691 );
buf ( n401693 , n400206 );
not ( n80244 , n401693 );
or ( n401695 , n401692 , n80244 );
buf ( n401696 , n379271 );
not ( n80247 , n401696 );
buf ( n401698 , n364858 );
not ( n401699 , n401698 );
or ( n80250 , n80247 , n401699 );
buf ( n401701 , n366131 );
buf ( n401702 , n379274 );
nand ( n401703 , n401701 , n401702 );
buf ( n401704 , n401703 );
buf ( n401705 , n401704 );
nand ( n401706 , n80250 , n401705 );
buf ( n401707 , n401706 );
buf ( n401708 , n401707 );
buf ( n401709 , n379299 );
nand ( n401710 , n401708 , n401709 );
buf ( n401711 , n401710 );
buf ( n401712 , n401711 );
nand ( n80263 , n401695 , n401712 );
buf ( n401714 , n80263 );
not ( n80265 , n401714 );
or ( n80266 , n401690 , n80265 );
buf ( n80267 , n401689 );
buf ( n401718 , n401714 );
nor ( n401719 , n80267 , n401718 );
buf ( n401720 , n401719 );
buf ( n401721 , n387542 );
not ( n80272 , n401721 );
buf ( n401723 , n400256 );
not ( n80274 , n401723 );
or ( n401725 , n80272 , n80274 );
buf ( n401726 , n400105 );
not ( n80277 , n401726 );
buf ( n401728 , n382496 );
not ( n80279 , n401728 );
or ( n80280 , n80277 , n80279 );
buf ( n401731 , n378736 );
buf ( n401732 , n380424 );
nand ( n80283 , n401731 , n401732 );
buf ( n401734 , n80283 );
buf ( n401735 , n401734 );
nand ( n80286 , n80280 , n401735 );
buf ( n401737 , n80286 );
buf ( n401738 , n401737 );
buf ( n401739 , n368608 );
nand ( n80290 , n401738 , n401739 );
buf ( n401741 , n80290 );
buf ( n401742 , n401741 );
nand ( n80293 , n401725 , n401742 );
buf ( n401744 , n80293 );
buf ( n401745 , n401744 );
xor ( n401746 , n396842 , n396845 );
xor ( n80297 , n401746 , n396873 );
xor ( n80298 , n400594 , n79521 );
xor ( n80299 , n80297 , n80298 );
buf ( n401750 , n80299 );
buf ( n401751 , n395038 );
not ( n401752 , n401751 );
buf ( n401753 , n394065 );
not ( n401754 , n401753 );
or ( n80305 , n401752 , n401754 );
buf ( n401756 , n394066 );
buf ( n401757 , n48458 );
nand ( n80308 , n401756 , n401757 );
buf ( n401759 , n80308 );
buf ( n401760 , n401759 );
nand ( n401761 , n80305 , n401760 );
buf ( n401762 , n401761 );
buf ( n401763 , n401762 );
not ( n401764 , n401763 );
buf ( n401765 , n45055 );
not ( n80316 , n401765 );
or ( n401767 , n401764 , n80316 );
buf ( n401768 , n400926 );
buf ( n401769 , n365242 );
nand ( n80320 , n401768 , n401769 );
buf ( n401771 , n80320 );
buf ( n401772 , n401771 );
nand ( n401773 , n401767 , n401772 );
buf ( n401774 , n401773 );
buf ( n401775 , n401774 );
xor ( n80326 , n401750 , n401775 );
xor ( n401777 , n79078 , n400587 );
xor ( n401778 , n401777 , n400591 );
xor ( n401779 , n400831 , n400901 );
xor ( n80330 , n401778 , n401779 );
buf ( n401781 , n80330 );
xor ( n80332 , n396700 , n396716 );
xor ( n401783 , n80332 , n396735 );
xor ( n401784 , n79242 , n400740 );
xor ( n401785 , n401783 , n401784 );
buf ( n401786 , n73625 );
buf ( n401787 , n380817 );
and ( n401788 , n401786 , n401787 );
buf ( n401789 , n73631 );
buf ( n401790 , n57983 );
and ( n401791 , n401789 , n401790 );
nor ( n401792 , n401788 , n401791 );
buf ( n401793 , n401792 );
buf ( n401794 , n401793 );
buf ( n401795 , n60313 );
or ( n80346 , n401794 , n401795 );
buf ( n401797 , n400641 );
buf ( n401798 , n380733 );
or ( n80349 , n401797 , n401798 );
nand ( n80350 , n80346 , n80349 );
buf ( n401801 , n80350 );
buf ( n80352 , n401801 );
buf ( n401803 , n74644 );
buf ( n401804 , n380570 );
and ( n401805 , n401803 , n401804 );
buf ( n401806 , n395683 );
buf ( n401807 , n60054 );
and ( n401808 , n401806 , n401807 );
nor ( n80359 , n401805 , n401808 );
buf ( n401810 , n80359 );
buf ( n401811 , n401810 );
buf ( n401812 , n380581 );
or ( n80363 , n401811 , n401812 );
buf ( n401814 , n400754 );
buf ( n401815 , n378453 );
or ( n401816 , n401814 , n401815 );
nand ( n80367 , n80363 , n401816 );
buf ( n401818 , n80367 );
buf ( n401819 , n401818 );
xor ( n80370 , n80352 , n401819 );
buf ( n401821 , n63549 );
buf ( n401822 , n382835 );
and ( n401823 , n401821 , n401822 );
buf ( n401824 , n384199 );
buf ( n401825 , n62243 );
and ( n80376 , n401824 , n401825 );
nor ( n401827 , n401823 , n80376 );
buf ( n401828 , n401827 );
buf ( n401829 , n401828 );
buf ( n401830 , n382849 );
or ( n80381 , n401829 , n401830 );
buf ( n401832 , n400624 );
buf ( n401833 , n384157 );
or ( n401834 , n401832 , n401833 );
nand ( n401835 , n80381 , n401834 );
buf ( n401836 , n401835 );
buf ( n401837 , n401836 );
and ( n401838 , n80370 , n401837 );
and ( n401839 , n80352 , n401819 );
or ( n401840 , n401838 , n401839 );
buf ( n401841 , n401840 );
buf ( n401842 , n401841 );
buf ( n401843 , n380680 );
buf ( n401844 , n394724 );
and ( n80395 , n401843 , n401844 );
buf ( n401846 , n60171 );
buf ( n401847 , n394730 );
and ( n401848 , n401846 , n401847 );
nor ( n80399 , n80395 , n401848 );
buf ( n401850 , n80399 );
buf ( n401851 , n401850 );
buf ( n401852 , n384414 );
or ( n80403 , n401851 , n401852 );
buf ( n401854 , n400808 );
buf ( n401855 , n395635 );
or ( n80406 , n401854 , n401855 );
nand ( n401857 , n80403 , n80406 );
buf ( n401858 , n401857 );
buf ( n401859 , n401858 );
xor ( n401860 , n401842 , n401859 );
xor ( n80411 , n400633 , n400650 );
xor ( n401862 , n80411 , n400736 );
buf ( n401863 , n401862 );
buf ( n401864 , n401863 );
and ( n80415 , n401860 , n401864 );
and ( n401866 , n401842 , n401859 );
or ( n401867 , n80415 , n401866 );
buf ( n401868 , n401867 );
xor ( n401869 , n401785 , n401868 );
xor ( n401870 , n400878 , n400882 );
xor ( n80421 , n401870 , n400887 );
buf ( n401872 , n80421 );
and ( n401873 , n401869 , n401872 );
and ( n80424 , n401785 , n401868 );
or ( n401875 , n401873 , n80424 );
xor ( n401876 , n400891 , n400894 );
xor ( n80427 , n401876 , n400898 );
and ( n80428 , n401875 , n80427 );
buf ( n401879 , n380838 );
buf ( n401880 , n63434 );
not ( n401881 , n401880 );
buf ( n401882 , n401881 );
buf ( n401883 , n401882 );
and ( n80434 , n401879 , n401883 );
buf ( n401885 , n380844 );
buf ( n401886 , n394730 );
and ( n401887 , n401885 , n401886 );
nor ( n80438 , n80434 , n401887 );
buf ( n401889 , n80438 );
buf ( n401890 , n401889 );
buf ( n401891 , n384414 );
or ( n401892 , n401890 , n401891 );
buf ( n401893 , n401850 );
buf ( n401894 , n395635 );
or ( n80445 , n401893 , n401894 );
nand ( n401896 , n401892 , n80445 );
buf ( n401897 , n401896 );
buf ( n401898 , n401897 );
buf ( n401899 , n380651 );
buf ( n401900 , n394840 );
and ( n401901 , n401899 , n401900 );
buf ( n401902 , n380657 );
buf ( n401903 , n395890 );
and ( n401904 , n401902 , n401903 );
nor ( n401905 , n401901 , n401904 );
buf ( n401906 , n401905 );
buf ( n401907 , n401906 );
buf ( n401908 , n394838 );
or ( n401909 , n401907 , n401908 );
buf ( n401910 , n79457 );
buf ( n401911 , n394835 );
or ( n80462 , n401910 , n401911 );
nand ( n80463 , n401909 , n80462 );
buf ( n401914 , n80463 );
buf ( n80465 , n401914 );
xor ( n80466 , n401898 , n80465 );
xor ( n80467 , n376584 , n376586 );
xor ( n80468 , n80467 , n56258 );
buf ( n401919 , n80468 );
not ( n401920 , n401919 );
buf ( n401921 , n401920 );
buf ( n401922 , n401921 );
buf ( n401923 , n376997 );
and ( n401924 , n401922 , n401923 );
buf ( n401925 , n80468 );
buf ( n401926 , n376990 );
and ( n401927 , n401925 , n401926 );
buf ( n401928 , n377003 );
nor ( n401929 , n401924 , n401927 , n401928 );
buf ( n401930 , n401929 );
buf ( n401931 , n401930 );
buf ( n401932 , n376921 );
not ( n80483 , n401932 );
buf ( n401934 , n79312 );
buf ( n401935 , n376866 );
and ( n80486 , n401934 , n401935 );
buf ( n401937 , n79318 );
buf ( n401938 , n382743 );
and ( n401939 , n401937 , n401938 );
nor ( n401940 , n80486 , n401939 );
buf ( n401941 , n401940 );
buf ( n401942 , n401941 );
not ( n80493 , n401942 );
buf ( n80494 , n80493 );
buf ( n401945 , n80494 );
not ( n401946 , n401945 );
or ( n401947 , n80483 , n401946 );
buf ( n401948 , n400686 );
buf ( n401949 , n56517 );
or ( n401950 , n401948 , n401949 );
nand ( n80501 , n401947 , n401950 );
buf ( n401952 , n80501 );
buf ( n401953 , n401952 );
xor ( n401954 , n401931 , n401953 );
buf ( n401955 , n401954 );
buf ( n401956 , n79114 );
buf ( n401957 , n57800 );
and ( n401958 , n401956 , n401957 );
buf ( n401959 , n400487 );
buf ( n401960 , n376903 );
and ( n401961 , n401959 , n401960 );
nor ( n401962 , n401958 , n401961 );
buf ( n401963 , n401962 );
buf ( n80514 , n401963 );
buf ( n80515 , n378341 );
or ( n80516 , n80514 , n80515 );
buf ( n80517 , n400719 );
buf ( n80518 , n378424 );
or ( n80519 , n80517 , n80518 );
nand ( n80520 , n80516 , n80519 );
buf ( n80521 , n80520 );
xor ( n401972 , n401955 , n80521 );
buf ( n401973 , n75451 );
buf ( n401974 , n380570 );
and ( n401975 , n401973 , n401974 );
buf ( n401976 , n396596 );
buf ( n401977 , n60054 );
and ( n80528 , n401976 , n401977 );
nor ( n401979 , n401975 , n80528 );
buf ( n401980 , n401979 );
buf ( n401981 , n401980 );
buf ( n401982 , n380581 );
or ( n80533 , n401981 , n401982 );
buf ( n401984 , n395810 );
buf ( n401985 , n380570 );
and ( n80536 , n401984 , n401985 );
buf ( n401987 , n395816 );
buf ( n401988 , n60054 );
and ( n80539 , n401987 , n401988 );
nor ( n80540 , n80536 , n80539 );
buf ( n401991 , n80540 );
buf ( n401992 , n401991 );
buf ( n401993 , n394774 );
or ( n80544 , n401992 , n401993 );
nand ( n80545 , n80533 , n80544 );
buf ( n401996 , n80545 );
and ( n401997 , n401972 , n401996 );
and ( n80548 , n401955 , n80521 );
or ( n80549 , n401997 , n80548 );
buf ( n402000 , n80549 );
buf ( n402001 , n396499 );
buf ( n402002 , n380817 );
and ( n80553 , n402001 , n402002 );
buf ( n402004 , n394816 );
buf ( n402005 , n57983 );
and ( n402006 , n402004 , n402005 );
nor ( n402007 , n80553 , n402006 );
buf ( n402008 , n402007 );
buf ( n402009 , n402008 );
buf ( n402010 , n60313 );
or ( n402011 , n402009 , n402010 );
buf ( n402012 , n401793 );
buf ( n402013 , n380733 );
or ( n80564 , n402012 , n402013 );
nand ( n80565 , n402011 , n80564 );
buf ( n402016 , n80565 );
buf ( n402017 , n402016 );
xor ( n80568 , n402000 , n402017 );
buf ( n402019 , n63406 );
buf ( n402020 , n384343 );
and ( n402021 , n402019 , n402020 );
buf ( n402022 , n384054 );
buf ( n402023 , n384089 );
and ( n80574 , n402022 , n402023 );
nor ( n402025 , n402021 , n80574 );
buf ( n402026 , n402025 );
buf ( n402027 , n402026 );
buf ( n402028 , n384354 );
or ( n80579 , n402027 , n402028 );
buf ( n402030 , n62202 );
buf ( n402031 , n384343 );
and ( n402032 , n402030 , n402031 );
buf ( n402033 , n382803 );
buf ( n402034 , n384089 );
and ( n80585 , n402033 , n402034 );
nor ( n80586 , n402032 , n80585 );
buf ( n402037 , n80586 );
buf ( n402038 , n402037 );
buf ( n402039 , n384082 );
or ( n402040 , n402038 , n402039 );
nand ( n402041 , n80579 , n402040 );
buf ( n402042 , n402041 );
buf ( n402043 , n402042 );
and ( n402044 , n80568 , n402043 );
and ( n80595 , n402000 , n402017 );
or ( n402046 , n402044 , n80595 );
buf ( n402047 , n402046 );
buf ( n402048 , n402047 );
and ( n402049 , n80466 , n402048 );
and ( n402050 , n401898 , n80465 );
or ( n80601 , n402049 , n402050 );
buf ( n402052 , n80601 );
buf ( n402053 , n402052 );
buf ( n402054 , n401991 );
buf ( n402055 , n380581 );
or ( n80606 , n402054 , n402055 );
buf ( n402057 , n401810 );
buf ( n402058 , n394774 );
or ( n80609 , n402057 , n402058 );
nand ( n402060 , n80606 , n80609 );
buf ( n402061 , n402060 );
buf ( n402062 , n402061 );
and ( n80613 , n401931 , n401953 );
buf ( n402064 , n80613 );
buf ( n402065 , n402064 );
xor ( n80616 , n402062 , n402065 );
xor ( n80617 , n79310 , n400710 );
xor ( n80618 , n80617 , n400728 );
buf ( n402069 , n80618 );
buf ( n402070 , n402069 );
and ( n80621 , n80616 , n402070 );
and ( n402072 , n402062 , n402065 );
or ( n402073 , n80621 , n402072 );
buf ( n402074 , n402073 );
xor ( n402075 , n400653 , n400677 );
xor ( n402076 , n402075 , n400732 );
and ( n80627 , n402074 , n402076 );
buf ( n402078 , n402037 );
buf ( n402079 , n384354 );
or ( n402080 , n402078 , n402079 );
buf ( n402081 , n400859 );
buf ( n402082 , n384082 );
or ( n402083 , n402081 , n402082 );
nand ( n80634 , n402080 , n402083 );
buf ( n402085 , n80634 );
xor ( n80636 , n400653 , n400677 );
xor ( n80637 , n80636 , n400732 );
and ( n402088 , n402085 , n80637 );
and ( n402089 , n402074 , n402085 );
or ( n80640 , n80627 , n402088 , n402089 );
buf ( n402091 , n80640 );
xor ( n402092 , n402053 , n402091 );
xor ( n80643 , n400851 , n400868 );
xor ( n402094 , n80643 , n400873 );
buf ( n402095 , n402094 );
buf ( n402096 , n402095 );
and ( n402097 , n402092 , n402096 );
and ( n80648 , n402053 , n402091 );
or ( n80649 , n402097 , n80648 );
buf ( n402100 , n80649 );
xor ( n402101 , n401785 , n401868 );
xor ( n80652 , n402101 , n401872 );
and ( n402103 , n402100 , n80652 );
buf ( n402104 , n61992 );
buf ( n402105 , n401882 );
and ( n402106 , n402104 , n402105 );
buf ( n402107 , n382596 );
buf ( n402108 , n384421 );
and ( n80659 , n402107 , n402108 );
nor ( n80660 , n402106 , n80659 );
buf ( n402111 , n80660 );
buf ( n402112 , n402111 );
buf ( n402113 , n384414 );
or ( n80664 , n402112 , n402113 );
buf ( n402115 , n401889 );
buf ( n402116 , n395635 );
or ( n402117 , n402115 , n402116 );
nand ( n80668 , n80664 , n402117 );
buf ( n402119 , n80668 );
buf ( n402120 , n384380 );
buf ( n402121 , n382835 );
and ( n402122 , n402120 , n402121 );
buf ( n402123 , n384386 );
buf ( n402124 , n62243 );
and ( n80675 , n402123 , n402124 );
nor ( n402126 , n402122 , n80675 );
buf ( n402127 , n402126 );
buf ( n402128 , n402127 );
buf ( n402129 , n382849 );
or ( n80680 , n402128 , n402129 );
buf ( n402131 , n401828 );
buf ( n402132 , n384157 );
or ( n80683 , n402131 , n402132 );
nand ( n80684 , n80680 , n80683 );
buf ( n402135 , n80684 );
xor ( n402136 , n402119 , n402135 );
xor ( n402137 , n402062 , n402065 );
xor ( n80688 , n402137 , n402070 );
buf ( n402139 , n80688 );
and ( n80690 , n402136 , n402139 );
and ( n402141 , n402119 , n402135 );
or ( n402142 , n80690 , n402141 );
buf ( n402143 , n402142 );
xor ( n80694 , n80352 , n401819 );
xor ( n80695 , n80694 , n401837 );
buf ( n402146 , n80695 );
buf ( n80697 , n402146 );
xor ( n80698 , n402143 , n80697 );
xor ( n80699 , n400653 , n400677 );
xor ( n80700 , n80699 , n400732 );
xor ( n402151 , n402074 , n402085 );
xor ( n402152 , n80700 , n402151 );
buf ( n402153 , n402152 );
and ( n80704 , n80698 , n402153 );
and ( n80705 , n402143 , n80697 );
or ( n402156 , n80704 , n80705 );
buf ( n402157 , n402156 );
xor ( n80708 , n401842 , n401859 );
xor ( n80709 , n80708 , n401864 );
buf ( n402160 , n80709 );
xor ( n80711 , n402157 , n402160 );
xor ( n80712 , n402053 , n402091 );
xor ( n80713 , n80712 , n402096 );
buf ( n402164 , n80713 );
and ( n80715 , n80711 , n402164 );
and ( n80716 , n402157 , n402160 );
or ( n80717 , n80715 , n80716 );
xor ( n80718 , n401785 , n401868 );
xor ( n80719 , n80718 , n401872 );
and ( n80720 , n80717 , n80719 );
and ( n80721 , n402100 , n80717 );
or ( n80722 , n402103 , n80720 , n80721 );
xor ( n80723 , n400891 , n400894 );
xor ( n80724 , n80723 , n400898 );
and ( n80725 , n80722 , n80724 );
and ( n80726 , n401875 , n80722 );
or ( n80727 , n80428 , n80725 , n80726 );
buf ( n402178 , n80727 );
xor ( n80729 , n401781 , n402178 );
buf ( n402180 , n365149 );
not ( n80731 , n402180 );
not ( n80732 , n45050 );
buf ( n402183 , n80732 );
not ( n80734 , n402183 );
not ( n402185 , n31311 );
buf ( n402186 , n402185 );
not ( n402187 , n402186 );
or ( n402188 , n80734 , n402187 );
buf ( n402189 , n351345 );
buf ( n402190 , n22954 );
not ( n402191 , n402190 );
buf ( n402192 , n402191 );
nand ( n402193 , n402189 , n402192 );
buf ( n402194 , n402193 );
buf ( n402195 , n402194 );
nand ( n402196 , n402188 , n402195 );
buf ( n402197 , n402196 );
buf ( n402198 , n402197 );
not ( n402199 , n402198 );
or ( n402200 , n80731 , n402199 );
not ( n402201 , n45010 );
buf ( n402202 , n402201 );
buf ( n402203 , n365384 );
not ( n402204 , n402203 );
buf ( n402205 , n402204 );
buf ( n402206 , n402205 );
not ( n80742 , n402206 );
buf ( n402208 , n402191 );
not ( n402209 , n402208 );
or ( n402210 , n80742 , n402209 );
buf ( n402211 , n80732 );
buf ( n402212 , n365384 );
nand ( n402213 , n402211 , n402212 );
buf ( n402214 , n402213 );
buf ( n402215 , n402214 );
nand ( n402216 , n402210 , n402215 );
buf ( n402217 , n402216 );
buf ( n402218 , n402217 );
nand ( n80754 , n402202 , n402218 );
buf ( n402220 , n80754 );
buf ( n402221 , n402220 );
nand ( n402222 , n402200 , n402221 );
buf ( n402223 , n402222 );
buf ( n402224 , n402223 );
and ( n402225 , n80729 , n402224 );
and ( n80761 , n401781 , n402178 );
or ( n402227 , n402225 , n80761 );
buf ( n402228 , n402227 );
buf ( n402229 , n402228 );
and ( n80765 , n80326 , n402229 );
and ( n402231 , n401750 , n401775 );
or ( n402232 , n80765 , n402231 );
buf ( n402233 , n402232 );
buf ( n402234 , n402233 );
buf ( n402235 , n56970 );
not ( n402236 , n402235 );
buf ( n402237 , n380923 );
not ( n80773 , n402237 );
or ( n402239 , n402236 , n80773 );
buf ( n402240 , n22619 );
buf ( n402241 , n377389 );
nand ( n402242 , n402240 , n402241 );
buf ( n402243 , n402242 );
buf ( n402244 , n402243 );
nand ( n80780 , n402239 , n402244 );
buf ( n402246 , n80780 );
buf ( n402247 , n402246 );
not ( n80783 , n402247 );
buf ( n402249 , n365725 );
not ( n80785 , n402249 );
or ( n80786 , n80783 , n80785 );
buf ( n402252 , n401189 );
buf ( n402253 , n56794 );
nand ( n80789 , n402252 , n402253 );
buf ( n402255 , n80789 );
buf ( n402256 , n402255 );
nand ( n402257 , n80786 , n402256 );
buf ( n402258 , n402257 );
buf ( n402259 , n402258 );
xor ( n80795 , n402234 , n402259 );
buf ( n402261 , n44915 );
not ( n402262 , n402261 );
buf ( n402263 , n400988 );
not ( n402264 , n402263 );
or ( n80800 , n402262 , n402264 );
buf ( n402266 , n365041 );
not ( n402267 , n402266 );
buf ( n402268 , n381266 );
not ( n402269 , n402268 );
or ( n80805 , n402267 , n402269 );
buf ( n402271 , n351160 );
buf ( n402272 , n380497 );
nand ( n80808 , n402271 , n402272 );
buf ( n80809 , n80808 );
buf ( n402275 , n80809 );
nand ( n80811 , n80805 , n402275 );
buf ( n402277 , n80811 );
buf ( n402278 , n402277 );
buf ( n402279 , n47466 );
nand ( n402280 , n402278 , n402279 );
buf ( n402281 , n402280 );
buf ( n402282 , n402281 );
nand ( n80818 , n80800 , n402282 );
buf ( n402284 , n80818 );
buf ( n402285 , n402284 );
and ( n402286 , n80795 , n402285 );
and ( n80822 , n402234 , n402259 );
or ( n402288 , n402286 , n80822 );
buf ( n402289 , n402288 );
buf ( n402290 , n402289 );
xor ( n402291 , n401745 , n402290 );
buf ( n402292 , n369809 );
not ( n80828 , n402292 );
buf ( n402294 , n401453 );
not ( n80830 , n402294 );
or ( n402296 , n80828 , n80830 );
buf ( n402297 , n393883 );
not ( n402298 , n402297 );
not ( n80834 , n377301 );
buf ( n80835 , n80834 );
not ( n80836 , n80835 );
or ( n80837 , n402298 , n80836 );
buf ( n80838 , n31260 );
buf ( n402304 , n369763 );
nand ( n80840 , n80838 , n402304 );
buf ( n402306 , n80840 );
buf ( n402307 , n402306 );
nand ( n80843 , n80837 , n402307 );
buf ( n402309 , n80843 );
buf ( n402310 , n402309 );
buf ( n402311 , n369804 );
nand ( n402312 , n402310 , n402311 );
buf ( n402313 , n402312 );
buf ( n402314 , n402313 );
nand ( n402315 , n402296 , n402314 );
buf ( n402316 , n402315 );
buf ( n402317 , n402316 );
and ( n402318 , n402291 , n402317 );
and ( n402319 , n401745 , n402290 );
or ( n80855 , n402318 , n402319 );
buf ( n402321 , n80855 );
buf ( n402322 , n402321 );
not ( n80858 , n402322 );
buf ( n402324 , n80858 );
or ( n402325 , n401720 , n402324 );
nand ( n80861 , n80266 , n402325 );
buf ( n402327 , n80861 );
xor ( n402328 , n401664 , n402327 );
buf ( n402329 , n361716 );
not ( n402330 , n402329 );
buf ( n402331 , n379380 );
not ( n402332 , n402331 );
and ( n402333 , n402330 , n402332 );
buf ( n402334 , n363547 );
buf ( n402335 , n379392 );
and ( n80871 , n402334 , n402335 );
nor ( n80872 , n402333 , n80871 );
buf ( n402338 , n80872 );
buf ( n402339 , n402338 );
buf ( n402340 , n379359 );
or ( n402341 , n402339 , n402340 );
buf ( n402342 , n401426 );
buf ( n402343 , n381675 );
or ( n80879 , n402342 , n402343 );
nand ( n80880 , n402341 , n80879 );
buf ( n402346 , n80880 );
buf ( n402347 , n402346 );
and ( n80883 , n402328 , n402347 );
and ( n402349 , n401664 , n402327 );
or ( n80885 , n80883 , n402349 );
buf ( n402351 , n80885 );
buf ( n402352 , n402351 );
xor ( n402353 , n401639 , n402352 );
xor ( n80889 , n401116 , n401141 );
xor ( n402355 , n80889 , n401360 );
buf ( n402356 , n402355 );
buf ( n402357 , n402356 );
and ( n402358 , n402353 , n402357 );
and ( n402359 , n401639 , n402352 );
or ( n80895 , n402358 , n402359 );
buf ( n402361 , n80895 );
buf ( n402362 , n402361 );
not ( n80898 , n402362 );
buf ( n80899 , n80898 );
buf ( n402365 , n80899 );
nand ( n80901 , n401541 , n402365 );
buf ( n402367 , n80901 );
not ( n402368 , n402367 );
or ( n402369 , n80074 , n402368 );
buf ( n402370 , n401540 );
not ( n402371 , n402370 );
buf ( n402372 , n402371 );
buf ( n402373 , n402372 );
buf ( n402374 , n402361 );
nand ( n402375 , n402373 , n402374 );
buf ( n402376 , n402375 );
nand ( n80912 , n402369 , n402376 );
xor ( n80913 , n401375 , n80912 );
xor ( n402379 , n401087 , n401366 );
xor ( n402380 , n402379 , n401077 );
and ( n80916 , n80913 , n402380 );
and ( n80917 , n401375 , n80912 );
or ( n80918 , n80916 , n80917 );
buf ( n402384 , n80918 );
xor ( n402385 , n401372 , n402384 );
xor ( n80921 , n399455 , n399462 );
xor ( n80922 , n80921 , n399512 );
buf ( n402388 , n80922 );
buf ( n402389 , n402388 );
xor ( n402390 , n399522 , n399526 );
xor ( n80926 , n402390 , n399673 );
buf ( n402392 , n80926 );
buf ( n402393 , n402392 );
xor ( n402394 , n402389 , n402393 );
buf ( n402395 , n401403 );
buf ( n402396 , n401378 );
or ( n402397 , n402395 , n402396 );
buf ( n402398 , n402397 );
buf ( n402399 , n402398 );
buf ( n402400 , n401520 );
and ( n402401 , n402399 , n402400 );
and ( n402402 , n401379 , n401404 );
buf ( n402403 , n402402 );
buf ( n402404 , n402403 );
nor ( n402405 , n402401 , n402404 );
buf ( n402406 , n402405 );
buf ( n402407 , n402406 );
not ( n402408 , n402407 );
buf ( n402409 , n402408 );
buf ( n402410 , n402409 );
not ( n402411 , n402410 );
buf ( n402412 , n399667 );
buf ( n402413 , n399558 );
xor ( n402414 , n402412 , n402413 );
buf ( n402415 , n399551 );
xnor ( n402416 , n402414 , n402415 );
buf ( n402417 , n402416 );
buf ( n402418 , n402417 );
not ( n402419 , n402418 );
buf ( n402420 , n402419 );
buf ( n402421 , n402420 );
not ( n80932 , n402421 );
or ( n80933 , n402411 , n80932 );
buf ( n402424 , n402406 );
not ( n402425 , n402424 );
buf ( n402426 , n402417 );
not ( n402427 , n402426 );
or ( n80937 , n402425 , n402427 );
xor ( n402429 , n400192 , n400372 );
xor ( n402430 , n402429 , n401055 );
buf ( n402431 , n402430 );
buf ( n402432 , n402431 );
xor ( n402433 , n399964 , n399989 );
xor ( n402434 , n402433 , n400183 );
buf ( n402435 , n402434 );
buf ( n402436 , n402435 );
or ( n80946 , n402432 , n402436 );
xor ( n402438 , n78851 , n78855 );
xor ( n402439 , n402438 , n400178 );
buf ( n402440 , n402439 );
buf ( n402441 , n402440 );
not ( n80951 , n402441 );
buf ( n402443 , n401396 );
buf ( n402444 , n380356 );
and ( n80954 , n402443 , n402444 );
buf ( n402446 , n380368 );
not ( n402447 , n402446 );
buf ( n402448 , n41666 );
not ( n80958 , n402448 );
or ( n80959 , n402447 , n80958 );
buf ( n402451 , n41663 );
buf ( n402452 , n384667 );
nand ( n402453 , n402451 , n402452 );
buf ( n402454 , n402453 );
buf ( n402455 , n402454 );
nand ( n80965 , n80959 , n402455 );
buf ( n402457 , n80965 );
buf ( n402458 , n402457 );
not ( n80968 , n402458 );
buf ( n402460 , n385064 );
nor ( n80970 , n80968 , n402460 );
buf ( n402462 , n80970 );
buf ( n402463 , n402462 );
nor ( n402464 , n80954 , n402463 );
buf ( n402465 , n402464 );
buf ( n402466 , n402465 );
nand ( n402467 , n80951 , n402466 );
buf ( n402468 , n402467 );
buf ( n402469 , n402468 );
xor ( n402470 , n400379 , n400404 );
xor ( n402471 , n402470 , n401050 );
buf ( n402472 , n402471 );
buf ( n402473 , n402472 );
and ( n402474 , n402469 , n402473 );
buf ( n402475 , n402440 );
not ( n402476 , n402475 );
buf ( n402477 , n402465 );
nor ( n402478 , n402476 , n402477 );
buf ( n402479 , n402478 );
buf ( n402480 , n402479 );
nor ( n80990 , n402474 , n402480 );
buf ( n402482 , n80990 );
buf ( n80992 , n402482 );
not ( n402484 , n80992 );
buf ( n402485 , n402484 );
buf ( n402486 , n402485 );
nand ( n402487 , n80946 , n402486 );
buf ( n402488 , n402487 );
buf ( n402489 , n402488 );
buf ( n402490 , n402431 );
buf ( n402491 , n402435 );
nand ( n402492 , n402490 , n402491 );
buf ( n402493 , n402492 );
buf ( n402494 , n402493 );
nand ( n402495 , n402489 , n402494 );
buf ( n402496 , n402495 );
buf ( n402497 , n402496 );
nand ( n81007 , n80937 , n402497 );
buf ( n81008 , n81007 );
buf ( n81009 , n81008 );
nand ( n81010 , n80933 , n81009 );
buf ( n81011 , n81010 );
buf ( n402503 , n81011 );
xor ( n402504 , n402394 , n402503 );
buf ( n402505 , n402504 );
buf ( n402506 , n402505 );
xor ( n81016 , n402385 , n402506 );
buf ( n402508 , n81016 );
buf ( n402509 , n402508 );
not ( n402510 , n402509 );
buf ( n402511 , n402510 );
buf ( n402512 , n402511 );
buf ( n402513 , n402409 );
not ( n402514 , n402513 );
buf ( n402515 , n402417 );
not ( n402516 , n402515 );
or ( n81026 , n402514 , n402516 );
buf ( n402518 , n402420 );
buf ( n402519 , n402406 );
nand ( n81029 , n402518 , n402519 );
buf ( n402521 , n81029 );
buf ( n402522 , n402521 );
nand ( n81032 , n81026 , n402522 );
buf ( n402524 , n81032 );
buf ( n402525 , n402524 );
buf ( n402526 , n402496 );
not ( n402527 , n402526 );
buf ( n402528 , n402527 );
buf ( n402529 , n402528 );
and ( n402530 , n402525 , n402529 );
not ( n81040 , n402525 );
buf ( n402532 , n402496 );
and ( n81042 , n81040 , n402532 );
nor ( n402534 , n402530 , n81042 );
buf ( n402535 , n402534 );
buf ( n402536 , n402535 );
not ( n81046 , n402536 );
buf ( n402538 , n81046 );
buf ( n402539 , n402538 );
not ( n402540 , n402539 );
buf ( n402541 , n78936 );
not ( n402542 , n402541 );
buf ( n402543 , n400365 );
buf ( n402544 , n400361 );
not ( n402545 , n402544 );
buf ( n402546 , n402545 );
buf ( n402547 , n402546 );
and ( n402548 , n402543 , n402547 );
not ( n81058 , n402543 );
buf ( n402550 , n400361 );
and ( n402551 , n81058 , n402550 );
nor ( n402552 , n402548 , n402551 );
buf ( n402553 , n402552 );
buf ( n402554 , n402553 );
not ( n402555 , n402554 );
or ( n81065 , n402542 , n402555 );
buf ( n402557 , n402553 );
buf ( n402558 , n78936 );
or ( n81068 , n402557 , n402558 );
nand ( n81069 , n81065 , n81068 );
buf ( n402561 , n81069 );
buf ( n402562 , n402561 );
xor ( n402563 , n401145 , n401353 );
xnor ( n81073 , n402563 , n79742 );
buf ( n402565 , n81073 );
not ( n81075 , n402565 );
buf ( n402567 , n380404 );
not ( n402568 , n402567 );
and ( n81078 , n380368 , n361751 );
not ( n81079 , n380368 );
and ( n81080 , n81079 , n41616 );
or ( n402572 , n81078 , n81080 );
buf ( n402573 , n402572 );
not ( n81083 , n402573 );
or ( n81084 , n402568 , n81083 );
buf ( n402576 , n402457 );
buf ( n81086 , n380356 );
nand ( n402578 , n402576 , n81086 );
buf ( n402579 , n402578 );
buf ( n402580 , n402579 );
nand ( n402581 , n81084 , n402580 );
buf ( n402582 , n402581 );
buf ( n402583 , n402582 );
not ( n402584 , n402583 );
buf ( n402585 , n402584 );
buf ( n402586 , n402585 );
not ( n402587 , n402586 );
or ( n402588 , n81075 , n402587 );
not ( n402589 , n398693 );
not ( n402590 , n401280 );
and ( n402591 , n402589 , n402590 );
buf ( n402592 , n377122 );
not ( n402593 , n402592 );
buf ( n402594 , n42233 );
not ( n81090 , n402594 );
or ( n402596 , n402593 , n81090 );
buf ( n81092 , n46693 );
buf ( n402598 , n57463 );
nand ( n81094 , n81092 , n402598 );
buf ( n402600 , n81094 );
buf ( n402601 , n402600 );
nand ( n402602 , n402596 , n402601 );
buf ( n402603 , n402602 );
and ( n402604 , n363429 , n402603 );
nor ( n402605 , n402591 , n402604 );
buf ( n402606 , n402605 );
not ( n402607 , n402606 );
buf ( n402608 , n402607 );
not ( n402609 , n402608 );
xor ( n402610 , n401202 , n401206 );
xor ( n402611 , n402610 , n401267 );
buf ( n402612 , n402611 );
not ( n402613 , n402612 );
or ( n402614 , n402609 , n402613 );
buf ( n402615 , n402612 );
not ( n81099 , n402615 );
buf ( n402617 , n81099 );
not ( n402618 , n402617 );
not ( n402619 , n402605 );
or ( n81103 , n402618 , n402619 );
buf ( n402621 , n377782 );
not ( n402622 , n402621 );
buf ( n402623 , n378138 );
not ( n81107 , n402623 );
or ( n81108 , n402622 , n81107 );
buf ( n402626 , n378135 );
buf ( n402627 , n377779 );
nand ( n402628 , n402626 , n402627 );
buf ( n402629 , n402628 );
buf ( n402630 , n402629 );
nand ( n81114 , n81108 , n402630 );
buf ( n402632 , n81114 );
buf ( n402633 , n402632 );
not ( n81117 , n402633 );
buf ( n402635 , n375896 );
not ( n402636 , n402635 );
or ( n402637 , n81117 , n402636 );
buf ( n402638 , n401309 );
buf ( n402639 , n375920 );
nand ( n402640 , n402638 , n402639 );
buf ( n402641 , n402640 );
buf ( n402642 , n402641 );
nand ( n402643 , n402637 , n402642 );
buf ( n402644 , n402643 );
buf ( n402645 , n402644 );
not ( n402646 , n402645 );
buf ( n402647 , n402646 );
buf ( n402648 , n402647 );
not ( n402649 , n402648 );
buf ( n402650 , n401737 );
buf ( n402651 , n387542 );
and ( n402652 , n402650 , n402651 );
buf ( n402653 , n400105 );
not ( n81125 , n402653 );
buf ( n402655 , n351228 );
not ( n402656 , n402655 );
or ( n81128 , n81125 , n402656 );
buf ( n402658 , n57233 );
buf ( n402659 , n380424 );
nand ( n402660 , n402658 , n402659 );
buf ( n402661 , n402660 );
buf ( n402662 , n402661 );
nand ( n81134 , n81128 , n402662 );
buf ( n402664 , n81134 );
buf ( n402665 , n402664 );
not ( n402666 , n402665 );
buf ( n402667 , n368605 );
nor ( n402668 , n402666 , n402667 );
buf ( n402669 , n402668 );
buf ( n402670 , n402669 );
nor ( n402671 , n402652 , n402670 );
buf ( n402672 , n402671 );
buf ( n402673 , n402672 );
not ( n402674 , n402673 );
or ( n402675 , n402649 , n402674 );
xor ( n81147 , n401232 , n401257 );
xor ( n402677 , n81147 , n401262 );
buf ( n402678 , n402677 );
buf ( n402679 , n402678 );
nand ( n81151 , n402675 , n402679 );
buf ( n81152 , n81151 );
buf ( n402682 , n81152 );
buf ( n402683 , n402672 );
not ( n81155 , n402683 );
buf ( n402685 , n402644 );
nand ( n81157 , n81155 , n402685 );
buf ( n402687 , n81157 );
buf ( n402688 , n402687 );
nand ( n81160 , n402682 , n402688 );
buf ( n402690 , n81160 );
nand ( n81162 , n81103 , n402690 );
nand ( n81163 , n402614 , n81162 );
buf ( n402693 , n81163 );
buf ( n402694 , n379838 );
not ( n402695 , n402694 );
buf ( n402696 , n364777 );
not ( n402697 , n402696 );
or ( n81169 , n402695 , n402697 );
buf ( n402699 , n368700 );
buf ( n402700 , n402699 );
buf ( n402701 , n398741 );
nand ( n402702 , n402700 , n402701 );
buf ( n402703 , n402702 );
buf ( n402704 , n402703 );
nand ( n402705 , n81169 , n402704 );
buf ( n402706 , n402705 );
not ( n81178 , n402706 );
not ( n402708 , n379916 );
or ( n402709 , n81178 , n402708 );
buf ( n402710 , n401653 );
not ( n402711 , n402710 );
buf ( n402712 , n402711 );
or ( n81184 , n402712 , n379893 );
nand ( n402714 , n402709 , n81184 );
buf ( n81186 , n402714 );
xor ( n81187 , n402693 , n81186 );
buf ( n402717 , n378856 );
not ( n402718 , n402717 );
buf ( n402719 , n377715 );
not ( n402720 , n402719 );
or ( n402721 , n402718 , n402720 );
buf ( n402722 , n365915 );
buf ( n402723 , n378847 );
nand ( n81195 , n402722 , n402723 );
buf ( n402725 , n81195 );
buf ( n402726 , n402725 );
nand ( n81198 , n402721 , n402726 );
buf ( n402728 , n81198 );
buf ( n402729 , n402728 );
not ( n81201 , n402729 );
buf ( n402731 , n49669 );
not ( n81203 , n402731 );
or ( n402733 , n81201 , n81203 );
buf ( n81205 , n401676 );
buf ( n81206 , n48558 );
nand ( n81207 , n81205 , n81206 );
buf ( n81208 , n81207 );
buf ( n81209 , n81208 );
nand ( n81210 , n402733 , n81209 );
buf ( n81211 , n81210 );
buf ( n402741 , n81211 );
not ( n81213 , n402741 );
buf ( n402743 , n367590 );
buf ( n402744 , n378098 );
nand ( n402745 , n402743 , n402744 );
buf ( n402746 , n402745 );
buf ( n402747 , n402746 );
not ( n402748 , n402747 );
buf ( n402749 , n402748 );
buf ( n402750 , n402749 );
not ( n402751 , n402750 );
or ( n402752 , n81213 , n402751 );
buf ( n402753 , n402746 );
not ( n81225 , n402753 );
buf ( n402755 , n81211 );
not ( n402756 , n402755 );
buf ( n402757 , n402756 );
buf ( n402758 , n402757 );
not ( n402759 , n402758 );
or ( n81231 , n81225 , n402759 );
buf ( n402761 , n365149 );
not ( n81233 , n402761 );
buf ( n402763 , n401249 );
not ( n402764 , n402763 );
or ( n402765 , n81233 , n402764 );
buf ( n402766 , n365183 );
buf ( n402767 , n402197 );
nand ( n81239 , n402766 , n402767 );
buf ( n402769 , n81239 );
buf ( n402770 , n402769 );
nand ( n81242 , n402765 , n402770 );
buf ( n402772 , n81242 );
buf ( n402773 , n402772 );
buf ( n402774 , n369374 );
not ( n402775 , n402774 );
buf ( n402776 , n386102 );
not ( n81248 , n402776 );
or ( n402778 , n402775 , n81248 );
buf ( n402779 , n386093 );
buf ( n402780 , n49178 );
nand ( n81252 , n402779 , n402780 );
buf ( n402782 , n81252 );
buf ( n402783 , n402782 );
nand ( n402784 , n402778 , n402783 );
buf ( n402785 , n402784 );
buf ( n402786 , n402785 );
not ( n402787 , n402786 );
buf ( n402788 , n365024 );
not ( n81260 , n402788 );
or ( n402790 , n402787 , n81260 );
buf ( n402791 , n401219 );
buf ( n402792 , n365108 );
nand ( n402793 , n402791 , n402792 );
buf ( n402794 , n402793 );
buf ( n402795 , n402794 );
nand ( n81267 , n402790 , n402795 );
buf ( n81268 , n81267 );
buf ( n402798 , n81268 );
xor ( n81270 , n402773 , n402798 );
buf ( n402800 , n44915 );
not ( n402801 , n402800 );
buf ( n402802 , n402277 );
not ( n402803 , n402802 );
or ( n81275 , n402801 , n402803 );
buf ( n402805 , n369183 );
buf ( n402806 , n352268 );
and ( n402807 , n402805 , n402806 );
not ( n81279 , n402805 );
buf ( n402809 , n63344 );
and ( n81281 , n81279 , n402809 );
nor ( n402811 , n402807 , n81281 );
buf ( n402812 , n402811 );
buf ( n402813 , n402812 );
not ( n402814 , n402813 );
buf ( n81286 , n47466 );
nand ( n81287 , n402814 , n81286 );
buf ( n81288 , n81287 );
buf ( n402818 , n81288 );
nand ( n81290 , n81275 , n402818 );
buf ( n81291 , n81290 );
buf ( n81292 , n81291 );
and ( n81293 , n81270 , n81292 );
and ( n81294 , n402773 , n402798 );
or ( n81295 , n81293 , n81294 );
buf ( n81296 , n81295 );
buf ( n402826 , n81296 );
xor ( n81298 , n401750 , n401775 );
xor ( n81299 , n81298 , n402229 );
buf ( n81300 , n81299 );
buf ( n81301 , n81300 );
buf ( n81302 , n387542 );
not ( n81303 , n81302 );
buf ( n81304 , n402664 );
not ( n81305 , n81304 );
or ( n81306 , n81303 , n81305 );
buf ( n402836 , n400105 );
not ( n402837 , n402836 );
buf ( n402838 , n378543 );
not ( n402839 , n402838 );
or ( n402840 , n402837 , n402839 );
buf ( n402841 , n381220 );
not ( n402842 , n402841 );
buf ( n81314 , n380424 );
nand ( n81315 , n402842 , n81314 );
buf ( n402845 , n81315 );
buf ( n402846 , n402845 );
nand ( n402847 , n402840 , n402846 );
buf ( n402848 , n402847 );
buf ( n402849 , n402848 );
buf ( n402850 , n368602 );
nand ( n402851 , n402849 , n402850 );
buf ( n402852 , n402851 );
buf ( n402853 , n402852 );
nand ( n402854 , n81306 , n402853 );
buf ( n402855 , n402854 );
buf ( n402856 , n402855 );
xor ( n402857 , n81301 , n402856 );
buf ( n402858 , n402812 );
not ( n402859 , n402858 );
buf ( n402860 , n365076 );
not ( n81332 , n402860 );
and ( n402862 , n402859 , n81332 );
buf ( n402863 , n365041 );
not ( n81335 , n402863 );
buf ( n402865 , n60751 );
not ( n402866 , n402865 );
or ( n81338 , n81335 , n402866 );
buf ( n402868 , n45802 );
buf ( n402869 , n369183 );
nand ( n81341 , n402868 , n402869 );
buf ( n402871 , n81341 );
buf ( n402872 , n402871 );
nand ( n402873 , n81338 , n402872 );
buf ( n402874 , n402873 );
buf ( n402875 , n402874 );
not ( n402876 , n402875 );
buf ( n402877 , n44913 );
nor ( n81349 , n402876 , n402877 );
buf ( n402879 , n81349 );
buf ( n402880 , n402879 );
nor ( n81352 , n402862 , n402880 );
buf ( n81353 , n81352 );
buf ( n81354 , n81353 );
not ( n81355 , n81354 );
buf ( n81356 , n81355 );
buf ( n402886 , n81356 );
buf ( n402887 , n368994 );
not ( n402888 , n402887 );
not ( n81360 , n342879 );
buf ( n402890 , n81360 );
not ( n402891 , n402890 );
or ( n402892 , n402888 , n402891 );
buf ( n402893 , n396441 );
buf ( n402894 , n57053 );
nand ( n402895 , n402893 , n402894 );
buf ( n402896 , n402895 );
buf ( n402897 , n402896 );
nand ( n81369 , n402892 , n402897 );
buf ( n402899 , n81369 );
buf ( n402900 , n402899 );
not ( n81372 , n402900 );
buf ( n402902 , n45055 );
not ( n81374 , n402902 );
or ( n81375 , n81372 , n81374 );
buf ( n402905 , n401762 );
buf ( n402906 , n365242 );
nand ( n402907 , n402905 , n402906 );
buf ( n402908 , n402907 );
buf ( n402909 , n402908 );
nand ( n402910 , n81375 , n402909 );
buf ( n402911 , n402910 );
buf ( n402912 , n402911 );
nand ( n81384 , n402886 , n402912 );
buf ( n402914 , n81384 );
buf ( n402915 , n402914 );
buf ( n402916 , n81356 );
buf ( n402917 , n402911 );
or ( n402918 , n402916 , n402917 );
xor ( n81390 , n401781 , n402178 );
xor ( n81391 , n81390 , n402224 );
buf ( n402921 , n81391 );
buf ( n402922 , n402921 );
nand ( n81394 , n402918 , n402922 );
buf ( n81395 , n81394 );
buf ( n402925 , n81395 );
nand ( n81397 , n402915 , n402925 );
buf ( n81398 , n81397 );
buf ( n402928 , n81398 );
and ( n81400 , n402857 , n402928 );
and ( n402930 , n81301 , n402856 );
or ( n402931 , n81400 , n402930 );
buf ( n402932 , n402931 );
buf ( n402933 , n402932 );
xor ( n402934 , n402826 , n402933 );
buf ( n402935 , n58463 );
buf ( n402936 , n377146 );
and ( n402937 , n402935 , n402936 );
buf ( n402938 , n58471 );
buf ( n402939 , n377143 );
and ( n81408 , n402938 , n402939 );
nor ( n402941 , n402937 , n81408 );
buf ( n402942 , n402941 );
buf ( n402943 , n402942 );
buf ( n402944 , n50782 );
or ( n402945 , n402943 , n402944 );
buf ( n402946 , n79907 );
buf ( n402947 , n377168 );
or ( n402948 , n402946 , n402947 );
nand ( n402949 , n402945 , n402948 );
buf ( n402950 , n402949 );
buf ( n402951 , n402950 );
and ( n402952 , n402934 , n402951 );
and ( n402953 , n402826 , n402933 );
or ( n402954 , n402952 , n402953 );
buf ( n402955 , n402954 );
buf ( n402956 , n402955 );
nand ( n402957 , n81231 , n402956 );
buf ( n402958 , n402957 );
buf ( n402959 , n402958 );
nand ( n402960 , n402752 , n402959 );
buf ( n402961 , n402960 );
buf ( n402962 , n402961 );
and ( n402963 , n81187 , n402962 );
and ( n402964 , n402693 , n81186 );
or ( n402965 , n402963 , n402964 );
buf ( n402966 , n402965 );
buf ( n402967 , n402966 );
nand ( n402968 , n402588 , n402967 );
buf ( n402969 , n402968 );
buf ( n402970 , n402969 );
buf ( n402971 , n81073 );
not ( n402972 , n402971 );
buf ( n402973 , n402582 );
nand ( n81422 , n402972 , n402973 );
buf ( n402975 , n81422 );
buf ( n81424 , n402975 );
nand ( n81425 , n402970 , n81424 );
buf ( n402978 , n81425 );
buf ( n402979 , n402978 );
xor ( n402980 , n402562 , n402979 );
xor ( n402981 , n401411 , n401435 );
xor ( n81430 , n402981 , n401516 );
buf ( n402983 , n81430 );
buf ( n402984 , n402983 );
and ( n402985 , n402980 , n402984 );
and ( n402986 , n402562 , n402979 );
or ( n81435 , n402985 , n402986 );
buf ( n402988 , n81435 );
buf ( n402989 , n402988 );
buf ( n402990 , n402440 );
buf ( n402991 , n402472 );
xor ( n81440 , n402990 , n402991 );
buf ( n402993 , n402465 );
xor ( n402994 , n81440 , n402993 );
buf ( n402995 , n402994 );
buf ( n402996 , n402995 );
not ( n81445 , n402996 );
buf ( n402998 , n81445 );
not ( n402999 , n402998 );
buf ( n403000 , n397190 );
not ( n403001 , n403000 );
buf ( n403002 , n401597 );
not ( n403003 , n403002 );
or ( n403004 , n403001 , n403003 );
not ( n403005 , n398363 );
not ( n403006 , n372382 );
or ( n403007 , n403005 , n403006 );
buf ( n403008 , n375903 );
not ( n403009 , n403008 );
buf ( n403010 , n377592 );
nand ( n403011 , n403009 , n403010 );
buf ( n403012 , n403011 );
nand ( n403013 , n403007 , n403012 );
buf ( n403014 , n403013 );
buf ( n403015 , n57530 );
nand ( n403016 , n403014 , n403015 );
buf ( n403017 , n403016 );
buf ( n403018 , n403017 );
nand ( n403019 , n403004 , n403018 );
buf ( n403020 , n403019 );
buf ( n403021 , n403020 );
xor ( n403022 , n401322 , n401326 );
xor ( n403023 , n403022 , n401344 );
buf ( n403024 , n403023 );
buf ( n403025 , n403024 );
xor ( n403026 , n403021 , n403025 );
not ( n403027 , n401707 );
not ( n403028 , n379263 );
or ( n403029 , n403027 , n403028 );
buf ( n403030 , n351107 );
not ( n81451 , n403030 );
buf ( n403032 , n379271 );
not ( n403033 , n403032 );
and ( n403034 , n81451 , n403033 );
buf ( n403035 , n351107 );
buf ( n403036 , n379271 );
and ( n403037 , n403035 , n403036 );
nor ( n403038 , n403034 , n403037 );
buf ( n403039 , n403038 );
or ( n403040 , n403039 , n379296 );
nand ( n403041 , n403029 , n403040 );
buf ( n403042 , n403041 );
and ( n403043 , n403026 , n403042 );
and ( n81461 , n403021 , n403025 );
or ( n403045 , n403043 , n81461 );
buf ( n403046 , n403045 );
buf ( n403047 , n403046 );
xor ( n81465 , n401461 , n401465 );
xor ( n403049 , n81465 , n401478 );
buf ( n403050 , n403049 );
buf ( n403051 , n403050 );
xor ( n403052 , n403047 , n403051 );
buf ( n403053 , n402338 );
buf ( n403054 , n381675 );
or ( n403055 , n403053 , n403054 );
buf ( n403056 , n379371 );
buf ( n403057 , n362549 );
not ( n403058 , n403057 );
xor ( n403059 , n403056 , n403058 );
buf ( n403060 , n403059 );
buf ( n403061 , n403060 );
not ( n81479 , n403061 );
buf ( n403063 , n58867 );
nand ( n403064 , n81479 , n403063 );
buf ( n403065 , n403064 );
buf ( n403066 , n403065 );
nand ( n403067 , n403055 , n403066 );
buf ( n403068 , n403067 );
buf ( n403069 , n403068 );
and ( n403070 , n403052 , n403069 );
and ( n403071 , n403047 , n403051 );
or ( n81489 , n403070 , n403071 );
buf ( n403073 , n81489 );
buf ( n403074 , n403073 );
not ( n81492 , n403074 );
buf ( n81493 , n81492 );
buf ( n403077 , n81493 );
not ( n81495 , n403077 );
buf ( n403079 , n401482 );
buf ( n403080 , n401509 );
xor ( n403081 , n403079 , n403080 );
buf ( n403082 , n401500 );
xnor ( n403083 , n403081 , n403082 );
buf ( n403084 , n403083 );
buf ( n403085 , n403084 );
not ( n81503 , n403085 );
or ( n403087 , n81495 , n81503 );
xor ( n81505 , n401272 , n401296 );
xor ( n81506 , n81505 , n401349 );
buf ( n403090 , n81506 );
buf ( n403091 , n403090 );
xor ( n81509 , n401745 , n402290 );
xor ( n403093 , n81509 , n402317 );
buf ( n403094 , n403093 );
buf ( n403095 , n403094 );
buf ( n403096 , n379916 );
not ( n403097 , n403096 );
buf ( n403098 , n379838 );
not ( n403099 , n403098 );
buf ( n403100 , n372201 );
not ( n81518 , n403100 );
or ( n403102 , n403099 , n81518 );
buf ( n403103 , n72880 );
buf ( n403104 , n398741 );
nand ( n403105 , n403103 , n403104 );
buf ( n403106 , n403105 );
buf ( n403107 , n403106 );
nand ( n403108 , n403102 , n403107 );
buf ( n403109 , n403108 );
buf ( n403110 , n403109 );
not ( n403111 , n403110 );
or ( n81529 , n403097 , n403111 );
buf ( n403113 , n402706 );
buf ( n403114 , n379890 );
nand ( n403115 , n403113 , n403114 );
buf ( n403116 , n403115 );
buf ( n403117 , n403116 );
nand ( n403118 , n81529 , n403117 );
buf ( n403119 , n403118 );
buf ( n403120 , n403119 );
or ( n403121 , n403095 , n403120 );
buf ( n403122 , n377353 );
not ( n81540 , n403122 );
buf ( n403124 , n380923 );
not ( n403125 , n403124 );
or ( n403126 , n81540 , n403125 );
buf ( n403127 , n22619 );
buf ( n403128 , n377352 );
nand ( n403129 , n403127 , n403128 );
buf ( n403130 , n403129 );
buf ( n403131 , n403130 );
nand ( n403132 , n403126 , n403131 );
buf ( n403133 , n403132 );
buf ( n403134 , n403133 );
not ( n81549 , n403134 );
buf ( n403136 , n365725 );
not ( n403137 , n403136 );
or ( n403138 , n81549 , n403137 );
buf ( n403139 , n402246 );
buf ( n403140 , n56794 );
nand ( n81555 , n403139 , n403140 );
buf ( n403142 , n81555 );
buf ( n403143 , n403142 );
nand ( n81558 , n403138 , n403143 );
buf ( n403145 , n81558 );
buf ( n403146 , n403145 );
buf ( n403147 , n377757 );
not ( n81562 , n403147 );
buf ( n403149 , n378138 );
not ( n403150 , n403149 );
or ( n81565 , n81562 , n403150 );
buf ( n403152 , n375914 );
buf ( n403153 , n378886 );
nand ( n403154 , n403152 , n403153 );
buf ( n403155 , n403154 );
buf ( n403156 , n403155 );
nand ( n403157 , n81565 , n403156 );
buf ( n403158 , n403157 );
buf ( n403159 , n403158 );
not ( n81574 , n403159 );
buf ( n403161 , n375896 );
not ( n403162 , n403161 );
or ( n403163 , n81574 , n403162 );
buf ( n403164 , n402632 );
buf ( n403165 , n375920 );
nand ( n403166 , n403164 , n403165 );
buf ( n403167 , n403166 );
buf ( n403168 , n403167 );
nand ( n403169 , n403163 , n403168 );
buf ( n403170 , n403169 );
buf ( n403171 , n403170 );
xor ( n403172 , n403146 , n403171 );
xor ( n403173 , n402773 , n402798 );
xor ( n403174 , n403173 , n81292 );
buf ( n403175 , n403174 );
buf ( n403176 , n403175 );
and ( n403177 , n403172 , n403176 );
and ( n403178 , n403146 , n403171 );
or ( n403179 , n403177 , n403178 );
buf ( n403180 , n403179 );
buf ( n403181 , n403180 );
not ( n403182 , n403181 );
buf ( n403183 , n369809 );
not ( n403184 , n403183 );
buf ( n403185 , n402309 );
not ( n81579 , n403185 );
or ( n81580 , n403184 , n81579 );
buf ( n403188 , n393883 );
not ( n81582 , n403188 );
buf ( n403190 , n375886 );
not ( n403191 , n403190 );
or ( n403192 , n81582 , n403191 );
buf ( n403193 , n32202 );
buf ( n403194 , n369763 );
nand ( n403195 , n403193 , n403194 );
buf ( n403196 , n403195 );
buf ( n403197 , n403196 );
nand ( n403198 , n403192 , n403197 );
buf ( n403199 , n403198 );
buf ( n403200 , n403199 );
buf ( n403201 , n369804 );
nand ( n403202 , n403200 , n403201 );
buf ( n403203 , n403202 );
buf ( n403204 , n403203 );
nand ( n403205 , n81580 , n403204 );
buf ( n403206 , n403205 );
buf ( n403207 , n403206 );
not ( n403208 , n403207 );
or ( n403209 , n403182 , n403208 );
buf ( n403210 , n403180 );
buf ( n403211 , n403206 );
or ( n403212 , n403210 , n403211 );
xor ( n403213 , n402234 , n402259 );
xor ( n403214 , n403213 , n402285 );
buf ( n403215 , n403214 );
buf ( n403216 , n403215 );
nand ( n403217 , n403212 , n403216 );
buf ( n403218 , n403217 );
buf ( n403219 , n403218 );
nand ( n81586 , n403209 , n403219 );
buf ( n403221 , n81586 );
buf ( n403222 , n403221 );
nand ( n81587 , n403121 , n403222 );
buf ( n403224 , n81587 );
buf ( n403225 , n403224 );
buf ( n403226 , n403119 );
buf ( n81591 , n403094 );
nand ( n81592 , n403226 , n81591 );
buf ( n403229 , n81592 );
buf ( n403230 , n403229 );
nand ( n81595 , n403225 , n403230 );
buf ( n403232 , n81595 );
buf ( n403233 , n403232 );
xor ( n403234 , n403091 , n403233 );
buf ( n403235 , n361603 );
buf ( n403236 , n378098 );
buf ( n403237 , n363603 );
and ( n403238 , n403236 , n403237 );
not ( n81603 , n403236 );
buf ( n403240 , n361534 );
and ( n403241 , n81603 , n403240 );
or ( n81606 , n403238 , n403241 );
buf ( n81607 , n81606 );
buf ( n403244 , n81607 );
or ( n81609 , n403235 , n403244 );
buf ( n403246 , n401493 );
buf ( n403247 , n364098 );
or ( n403248 , n403246 , n403247 );
nand ( n403249 , n81609 , n403248 );
buf ( n403250 , n403249 );
buf ( n403251 , n403250 );
and ( n403252 , n403234 , n403251 );
and ( n81617 , n403091 , n403233 );
or ( n81618 , n403252 , n81617 );
buf ( n403255 , n81618 );
buf ( n403256 , n403255 );
nand ( n403257 , n403087 , n403256 );
buf ( n403258 , n403257 );
buf ( n403259 , n403258 );
buf ( n403260 , n403084 );
not ( n81625 , n403260 );
buf ( n403262 , n81625 );
buf ( n403263 , n403262 );
buf ( n403264 , n403073 );
nand ( n81629 , n403263 , n403264 );
buf ( n403266 , n81629 );
buf ( n403267 , n403266 );
and ( n403268 , n403259 , n403267 );
buf ( n403269 , n403268 );
buf ( n403270 , n403269 );
not ( n403271 , n403270 );
buf ( n403272 , n403271 );
not ( n81637 , n403272 );
or ( n81638 , n402999 , n81637 );
not ( n403275 , n403269 );
not ( n403276 , n402995 );
or ( n81641 , n403275 , n403276 );
xor ( n403278 , n401639 , n402352 );
xor ( n403279 , n403278 , n402357 );
buf ( n403280 , n403279 );
nand ( n81645 , n81641 , n403280 );
nand ( n403282 , n81638 , n81645 );
buf ( n403283 , n403282 );
xor ( n403284 , n402989 , n403283 );
buf ( n403285 , n402431 );
not ( n81650 , n403285 );
xor ( n403287 , n402482 , n402435 );
buf ( n403288 , n403287 );
not ( n81653 , n403288 );
or ( n403290 , n81650 , n81653 );
buf ( n403291 , n403287 );
buf ( n403292 , n402431 );
or ( n403293 , n403291 , n403292 );
nand ( n403294 , n403290 , n403293 );
buf ( n403295 , n403294 );
buf ( n403296 , n403295 );
and ( n403297 , n403284 , n403296 );
and ( n81662 , n402989 , n403283 );
or ( n403299 , n403297 , n81662 );
buf ( n403300 , n403299 );
buf ( n403301 , n403300 );
not ( n81666 , n403301 );
or ( n403303 , n402540 , n81666 );
not ( n403304 , n402535 );
buf ( n403305 , n403300 );
not ( n81670 , n403305 );
buf ( n81671 , n81670 );
not ( n403308 , n81671 );
or ( n81673 , n403304 , n403308 );
xor ( n403310 , n401375 , n80912 );
xor ( n403311 , n403310 , n402380 );
nand ( n81676 , n81673 , n403311 );
buf ( n403313 , n81676 );
nand ( n403314 , n403303 , n403313 );
buf ( n403315 , n403314 );
buf ( n403316 , n403315 );
not ( n81681 , n403316 );
buf ( n403318 , n81681 );
buf ( n403319 , n403318 );
nand ( n403320 , n402512 , n403319 );
buf ( n403321 , n403320 );
buf ( n403322 , n403321 );
xor ( n403323 , n402989 , n403283 );
xor ( n81688 , n403323 , n403296 );
buf ( n403325 , n81688 );
not ( n403326 , n403325 );
buf ( n403327 , n401523 );
not ( n403328 , n403327 );
buf ( n403329 , n402372 );
buf ( n403330 , n402361 );
and ( n81695 , n403329 , n403330 );
not ( n403332 , n403329 );
buf ( n403333 , n80899 );
and ( n403334 , n403332 , n403333 );
nor ( n81699 , n81695 , n403334 );
buf ( n403336 , n81699 );
buf ( n403337 , n403336 );
not ( n81702 , n403337 );
buf ( n403339 , n81702 );
buf ( n403340 , n403339 );
not ( n403341 , n403340 );
or ( n403342 , n403328 , n403341 );
buf ( n403343 , n401523 );
not ( n81708 , n403343 );
buf ( n403345 , n403336 );
nand ( n403346 , n81708 , n403345 );
buf ( n403347 , n403346 );
buf ( n403348 , n403347 );
nand ( n81713 , n403342 , n403348 );
buf ( n403350 , n81713 );
buf ( n403351 , n403350 );
buf ( n403352 , n401570 );
not ( n81717 , n401561 );
buf ( n403354 , n81717 );
and ( n403355 , n403352 , n403354 );
not ( n403356 , n403352 );
buf ( n403357 , n401561 );
and ( n403358 , n403356 , n403357 );
nor ( n403359 , n403355 , n403358 );
buf ( n403360 , n403359 );
xnor ( n81725 , n401627 , n403360 );
buf ( n403362 , n81725 );
xor ( n403363 , n401664 , n402327 );
xor ( n81728 , n403363 , n402347 );
buf ( n403365 , n81728 );
buf ( n81730 , n403365 );
xor ( n81731 , n403362 , n81730 );
and ( n403368 , n401714 , n402324 );
not ( n403369 , n401714 );
and ( n81734 , n403369 , n402321 );
or ( n403371 , n403368 , n81734 );
xor ( n403372 , n401689 , n403371 );
buf ( n403373 , n403372 );
xor ( n81738 , n401580 , n401605 );
xor ( n403375 , n81738 , n401623 );
buf ( n403376 , n403375 );
buf ( n403377 , n403376 );
xor ( n403378 , n403373 , n403377 );
and ( n81743 , n81152 , n402687 );
and ( n403380 , n402612 , n81743 );
not ( n403381 , n402612 );
and ( n81746 , n403381 , n402690 );
or ( n81747 , n403380 , n81746 );
buf ( n403384 , n81747 );
buf ( n403385 , n402605 );
and ( n403386 , n403384 , n403385 );
not ( n81751 , n403384 );
buf ( n403388 , n402608 );
and ( n81753 , n81751 , n403388 );
nor ( n403390 , n403386 , n81753 );
buf ( n403391 , n403390 );
buf ( n403392 , n403391 );
not ( n81757 , n403392 );
buf ( n403394 , n81757 );
buf ( n403395 , n403394 );
not ( n81760 , n403395 );
buf ( n403397 , n377094 );
not ( n81762 , n403397 );
buf ( n403399 , n41772 );
not ( n81764 , n403399 );
or ( n403401 , n81762 , n81764 );
buf ( n403402 , n366329 );
buf ( n403403 , n56687 );
nand ( n81768 , n403402 , n403403 );
buf ( n403405 , n81768 );
buf ( n403406 , n403405 );
nand ( n81771 , n403401 , n403406 );
buf ( n403408 , n81771 );
buf ( n403409 , n403408 );
not ( n403410 , n403409 );
buf ( n403411 , n41830 );
not ( n81776 , n403411 );
or ( n403413 , n403410 , n81776 );
buf ( n403414 , n80160 );
buf ( n403415 , n41835 );
nand ( n81780 , n403414 , n403415 );
buf ( n81781 , n81780 );
buf ( n403418 , n81781 );
nand ( n403419 , n403413 , n403418 );
buf ( n403420 , n403419 );
buf ( n403421 , n403420 );
not ( n403422 , n403421 );
or ( n403423 , n81760 , n403422 );
buf ( n403424 , n403420 );
buf ( n403425 , n403394 );
or ( n403426 , n403424 , n403425 );
buf ( n403427 , n361955 );
not ( n403428 , n403427 );
buf ( n403429 , n342335 );
not ( n403430 , n403429 );
or ( n403431 , n403428 , n403430 );
buf ( n403432 , n378098 );
nand ( n81797 , n403431 , n403432 );
buf ( n81798 , n81797 );
buf ( n81799 , n81798 );
buf ( n403436 , n365319 );
buf ( n403437 , n361955 );
not ( n403438 , n403437 );
buf ( n81803 , n381336 );
nand ( n81804 , n403438 , n81803 );
buf ( n403441 , n81804 );
buf ( n403442 , n403441 );
and ( n81807 , n81799 , n403436 , n403442 );
buf ( n403444 , n81807 );
buf ( n403445 , n403444 );
not ( n403446 , n403445 );
buf ( n403447 , n403446 );
buf ( n403448 , n403447 );
not ( n403449 , n403448 );
buf ( n403450 , n58984 );
not ( n81815 , n403450 );
buf ( n403452 , n342718 );
not ( n403453 , n403452 );
or ( n81818 , n81815 , n403453 );
buf ( n403455 , n386354 );
buf ( n403456 , n379482 );
nand ( n403457 , n403455 , n403456 );
buf ( n403458 , n403457 );
buf ( n81823 , n403458 );
nand ( n403460 , n81818 , n81823 );
buf ( n403461 , n403460 );
buf ( n403462 , n403461 );
not ( n403463 , n403462 );
buf ( n403464 , n363429 );
not ( n81829 , n403464 );
or ( n81830 , n403463 , n81829 );
buf ( n403467 , n402603 );
buf ( n403468 , n378183 );
nand ( n81833 , n403467 , n403468 );
buf ( n403470 , n81833 );
buf ( n403471 , n403470 );
nand ( n403472 , n81830 , n403471 );
buf ( n403473 , n403472 );
buf ( n403474 , n403473 );
not ( n81839 , n403474 );
buf ( n403476 , n81839 );
buf ( n403477 , n403476 );
not ( n81842 , n403477 );
or ( n81843 , n403449 , n81842 );
buf ( n403480 , n369809 );
not ( n403481 , n403480 );
buf ( n403482 , n403199 );
not ( n81847 , n403482 );
or ( n81848 , n403481 , n81847 );
and ( n81849 , n375873 , n393883 );
not ( n403486 , n375873 );
and ( n81851 , n403486 , n369763 );
or ( n81852 , n81849 , n81851 );
buf ( n403489 , n81852 );
buf ( n403490 , n369804 );
nand ( n81855 , n403489 , n403490 );
buf ( n403492 , n81855 );
buf ( n403493 , n403492 );
nand ( n81858 , n81848 , n403493 );
buf ( n403495 , n81858 );
buf ( n403496 , n403495 );
xor ( n81861 , n400891 , n400894 );
xor ( n81862 , n81861 , n400898 );
xor ( n81863 , n401875 , n80722 );
xor ( n81864 , n81862 , n81863 );
buf ( n403501 , n81864 );
buf ( n403502 , n368656 );
not ( n81867 , n396401 );
buf ( n403504 , n81867 );
and ( n403505 , n403502 , n403504 );
not ( n403506 , n403502 );
not ( n81871 , n81867 );
buf ( n403508 , n81871 );
and ( n81873 , n403506 , n403508 );
nor ( n403510 , n403505 , n81873 );
buf ( n403511 , n403510 );
buf ( n403512 , n403511 );
not ( n403513 , n403512 );
buf ( n403514 , n45012 );
not ( n81879 , n403514 );
or ( n403516 , n403513 , n81879 );
buf ( n403517 , n402217 );
buf ( n403518 , n365149 );
nand ( n403519 , n403517 , n403518 );
buf ( n403520 , n403519 );
buf ( n403521 , n403520 );
nand ( n403522 , n403516 , n403521 );
buf ( n403523 , n403522 );
buf ( n403524 , n403523 );
xor ( n403525 , n403501 , n403524 );
xor ( n403526 , n401785 , n401868 );
xor ( n81891 , n403526 , n401872 );
xor ( n403528 , n402100 , n80717 );
xor ( n403529 , n81891 , n403528 );
buf ( n403530 , n403529 );
xor ( n403531 , n401898 , n80465 );
xor ( n403532 , n403531 , n402048 );
buf ( n403533 , n403532 );
buf ( n403534 , n380680 );
buf ( n403535 , n394840 );
and ( n403536 , n403534 , n403535 );
buf ( n403537 , n60171 );
buf ( n403538 , n395890 );
and ( n81903 , n403537 , n403538 );
nor ( n403540 , n403536 , n81903 );
buf ( n403541 , n403540 );
buf ( n403542 , n403541 );
buf ( n403543 , n394838 );
or ( n403544 , n403542 , n403543 );
buf ( n403545 , n401906 );
buf ( n403546 , n394835 );
or ( n81911 , n403545 , n403546 );
nand ( n81912 , n403544 , n81911 );
buf ( n403549 , n81912 );
buf ( n403550 , n403549 );
buf ( n403551 , n74644 );
buf ( n403552 , n380817 );
and ( n403553 , n403551 , n403552 );
buf ( n403554 , n395683 );
buf ( n403555 , n63664 );
and ( n403556 , n403554 , n403555 );
nor ( n81921 , n403553 , n403556 );
buf ( n81922 , n81921 );
buf ( n403559 , n81922 );
buf ( n403560 , n60313 );
or ( n403561 , n403559 , n403560 );
buf ( n403562 , n402008 );
buf ( n403563 , n380733 );
or ( n403564 , n403562 , n403563 );
nand ( n81929 , n403561 , n403564 );
buf ( n403566 , n81929 );
buf ( n403567 , n403566 );
buf ( n403568 , n80468 );
buf ( n403569 , n376866 );
and ( n81934 , n403568 , n403569 );
buf ( n403571 , n401921 );
buf ( n403572 , n382743 );
and ( n403573 , n403571 , n403572 );
nor ( n81938 , n81934 , n403573 );
buf ( n81939 , n81938 );
buf ( n403576 , n81939 );
buf ( n403577 , n376924 );
or ( n81942 , n403576 , n403577 );
buf ( n403579 , n401941 );
buf ( n403580 , n56517 );
or ( n403581 , n403579 , n403580 );
nand ( n81946 , n81942 , n403581 );
buf ( n403583 , n81946 );
buf ( n403584 , n403583 );
and ( n81949 , n56198 , n376657 );
xor ( n81950 , n81949 , n376654 );
buf ( n403587 , n81950 );
not ( n81952 , n403587 );
buf ( n403589 , n81952 );
buf ( n403590 , n403589 );
buf ( n403591 , n376997 );
and ( n403592 , n403590 , n403591 );
buf ( n403593 , n81950 );
buf ( n403594 , n376990 );
and ( n81959 , n403593 , n403594 );
buf ( n403596 , n377003 );
nor ( n403597 , n403592 , n81959 , n403596 );
buf ( n403598 , n403597 );
buf ( n403599 , n403598 );
xor ( n403600 , n403584 , n403599 );
buf ( n403601 , n400503 );
buf ( n403602 , n57800 );
and ( n403603 , n403601 , n403602 );
buf ( n403604 , n400509 );
buf ( n403605 , n376903 );
and ( n403606 , n403604 , n403605 );
nor ( n403607 , n403603 , n403606 );
buf ( n403608 , n403607 );
buf ( n403609 , n403608 );
buf ( n403610 , n378341 );
or ( n403611 , n403609 , n403610 );
buf ( n403612 , n401963 );
buf ( n403613 , n378424 );
or ( n81967 , n403612 , n403613 );
nand ( n403615 , n403611 , n81967 );
buf ( n403616 , n403615 );
buf ( n403617 , n403616 );
and ( n403618 , n403600 , n403617 );
and ( n403619 , n403584 , n403599 );
or ( n81973 , n403618 , n403619 );
buf ( n403621 , n81973 );
buf ( n403622 , n403621 );
xor ( n403623 , n403567 , n403622 );
buf ( n403624 , n396615 );
buf ( n403625 , n57789 );
and ( n403626 , n403624 , n403625 );
buf ( n403627 , n396621 );
buf ( n403628 , n60054 );
and ( n403629 , n403627 , n403628 );
nor ( n81983 , n403626 , n403629 );
buf ( n403631 , n81983 );
buf ( n403632 , n403631 );
buf ( n403633 , n380581 );
or ( n81987 , n403632 , n403633 );
buf ( n403635 , n401980 );
buf ( n403636 , n394774 );
or ( n403637 , n403635 , n403636 );
nand ( n81991 , n81987 , n403637 );
buf ( n403639 , n81991 );
buf ( n403640 , n403639 );
and ( n403641 , n376612 , n376653 );
xor ( n81995 , n403641 , n376650 );
buf ( n403643 , n81995 );
not ( n81997 , n403643 );
buf ( n403645 , n81997 );
buf ( n403646 , n403645 );
buf ( n403647 , n376997 );
and ( n82001 , n403646 , n403647 );
buf ( n403649 , n81995 );
buf ( n403650 , n376990 );
and ( n403651 , n403649 , n403650 );
buf ( n403652 , n377003 );
nor ( n403653 , n82001 , n403651 , n403652 );
buf ( n403654 , n403653 );
buf ( n403655 , n403654 );
buf ( n403656 , n376866 );
buf ( n403657 , n81950 );
and ( n403658 , n403656 , n403657 );
not ( n403659 , n403656 );
buf ( n403660 , n403589 );
and ( n403661 , n403659 , n403660 );
nor ( n403662 , n403658 , n403661 );
buf ( n403663 , n403662 );
buf ( n403664 , n403663 );
buf ( n403665 , n376924 );
or ( n82005 , n403664 , n403665 );
buf ( n403667 , n81939 );
buf ( n403668 , n56517 );
or ( n403669 , n403667 , n403668 );
nand ( n403670 , n82005 , n403669 );
buf ( n403671 , n403670 );
buf ( n403672 , n403671 );
and ( n82012 , n403655 , n403672 );
buf ( n403674 , n82012 );
buf ( n403675 , n403674 );
xor ( n82015 , n403640 , n403675 );
xor ( n403677 , n403584 , n403599 );
xor ( n403678 , n403677 , n403617 );
buf ( n403679 , n403678 );
buf ( n403680 , n403679 );
and ( n82020 , n82015 , n403680 );
and ( n82021 , n403640 , n403675 );
or ( n403683 , n82020 , n82021 );
buf ( n403684 , n403683 );
buf ( n403685 , n403684 );
and ( n82025 , n403623 , n403685 );
and ( n403687 , n403567 , n403622 );
or ( n403688 , n82025 , n403687 );
buf ( n403689 , n403688 );
buf ( n403690 , n403689 );
xor ( n403691 , n403550 , n403690 );
buf ( n403692 , n73625 );
buf ( n403693 , n382835 );
and ( n403694 , n403692 , n403693 );
buf ( n82034 , n73631 );
buf ( n403696 , n62243 );
and ( n403697 , n82034 , n403696 );
nor ( n403698 , n403694 , n403697 );
buf ( n403699 , n403698 );
buf ( n403700 , n403699 );
buf ( n403701 , n382849 );
or ( n403702 , n403700 , n403701 );
buf ( n403703 , n402127 );
buf ( n403704 , n384157 );
or ( n403705 , n403703 , n403704 );
nand ( n82045 , n403702 , n403705 );
buf ( n403707 , n82045 );
xor ( n82047 , n401955 , n80521 );
xor ( n82048 , n82047 , n401996 );
and ( n403710 , n403707 , n82048 );
buf ( n403711 , n63549 );
buf ( n403712 , n384343 );
and ( n403713 , n403711 , n403712 );
buf ( n403714 , n384199 );
buf ( n403715 , n384089 );
and ( n403716 , n403714 , n403715 );
nor ( n403717 , n403713 , n403716 );
buf ( n403718 , n403717 );
buf ( n403719 , n403718 );
buf ( n403720 , n384354 );
or ( n82060 , n403719 , n403720 );
buf ( n403722 , n402026 );
buf ( n403723 , n384082 );
or ( n82063 , n403722 , n403723 );
nand ( n403725 , n82060 , n82063 );
buf ( n403726 , n403725 );
xor ( n82066 , n401955 , n80521 );
xor ( n403728 , n82066 , n401996 );
and ( n403729 , n403726 , n403728 );
and ( n82069 , n403707 , n403726 );
or ( n403731 , n403710 , n403729 , n82069 );
buf ( n403732 , n403731 );
and ( n82072 , n403691 , n403732 );
and ( n403734 , n403550 , n403690 );
or ( n403735 , n82072 , n403734 );
buf ( n403736 , n403735 );
xor ( n82076 , n403533 , n403736 );
xor ( n82077 , n402143 , n80697 );
xor ( n403739 , n82077 , n402153 );
buf ( n403740 , n403739 );
and ( n82080 , n82076 , n403740 );
and ( n82081 , n403533 , n403736 );
or ( n403743 , n82080 , n82081 );
xor ( n403744 , n402157 , n402160 );
xor ( n82084 , n403744 , n402164 );
and ( n403746 , n403743 , n82084 );
xor ( n403747 , n402000 , n402017 );
xor ( n82087 , n403747 , n402043 );
buf ( n403749 , n82087 );
xor ( n403750 , n402119 , n402135 );
xor ( n403751 , n403750 , n402139 );
and ( n403752 , n403749 , n403751 );
buf ( n403753 , n376924 );
buf ( n403754 , n81995 );
buf ( n403755 , n376866 );
and ( n82095 , n403754 , n403755 );
buf ( n403757 , n403645 );
buf ( n403758 , n377030 );
and ( n403759 , n403757 , n403758 );
nor ( n403760 , n82095 , n403759 );
buf ( n403761 , n403760 );
buf ( n403762 , n403761 );
or ( n403763 , n403753 , n403762 );
buf ( n403764 , n403663 );
buf ( n403765 , n56517 );
or ( n82105 , n403764 , n403765 );
nand ( n403767 , n403763 , n82105 );
buf ( n403768 , n403767 );
buf ( n403769 , n403768 );
not ( n82109 , n376647 );
nand ( n403771 , n82109 , n56249 );
xor ( n403772 , n56242 , n403771 );
buf ( n403773 , n403772 );
not ( n403774 , n403773 );
buf ( n403775 , n403774 );
buf ( n403776 , n403775 );
buf ( n403777 , n376997 );
and ( n403778 , n403776 , n403777 );
buf ( n403779 , n403772 );
buf ( n403780 , n376990 );
and ( n403781 , n403779 , n403780 );
buf ( n403782 , n377003 );
nor ( n82122 , n403778 , n403781 , n403782 );
buf ( n403784 , n82122 );
buf ( n403785 , n403784 );
xor ( n82125 , n403769 , n403785 );
buf ( n403787 , n376997 );
and ( n403788 , n56237 , n376640 );
not ( n403789 , n403788 );
not ( n82129 , n56226 );
nor ( n403791 , n82129 , n56216 );
not ( n403792 , n403791 );
or ( n403793 , n403789 , n403792 );
or ( n82133 , n403791 , n403788 );
nand ( n403795 , n403793 , n82133 );
buf ( n403796 , n403795 );
not ( n82136 , n403796 );
buf ( n403798 , n82136 );
buf ( n403799 , n403798 );
and ( n403800 , n403787 , n403799 );
buf ( n403801 , n376990 );
buf ( n403802 , n403795 );
and ( n403803 , n403801 , n403802 );
buf ( n403804 , n377003 );
nor ( n82144 , n403800 , n403803 , n403804 );
buf ( n82145 , n82144 );
buf ( n82146 , n82145 );
buf ( n403808 , n376924 );
buf ( n403809 , n376866 );
buf ( n403810 , n403772 );
and ( n403811 , n403809 , n403810 );
buf ( n403812 , n377030 );
buf ( n403813 , n403775 );
and ( n403814 , n403812 , n403813 );
nor ( n403815 , n403811 , n403814 );
buf ( n403816 , n403815 );
buf ( n403817 , n403816 );
or ( n82157 , n403808 , n403817 );
buf ( n403819 , n403761 );
buf ( n403820 , n56517 );
or ( n82160 , n403819 , n403820 );
nand ( n82161 , n82157 , n82160 );
buf ( n403823 , n82161 );
buf ( n403824 , n403823 );
and ( n82164 , n82146 , n403824 );
buf ( n403826 , n82164 );
buf ( n403827 , n403826 );
and ( n82167 , n82125 , n403827 );
and ( n82168 , n403769 , n403785 );
or ( n403830 , n82167 , n82168 );
buf ( n403831 , n403830 );
buf ( n403832 , n403831 );
buf ( n403833 , n79312 );
buf ( n403834 , n57800 );
and ( n403835 , n403833 , n403834 );
buf ( n403836 , n79318 );
buf ( n403837 , n378284 );
and ( n82177 , n403836 , n403837 );
nor ( n82178 , n403835 , n82177 );
buf ( n403840 , n82178 );
buf ( n403841 , n403840 );
buf ( n403842 , n378341 );
or ( n82182 , n403841 , n403842 );
buf ( n403844 , n403608 );
buf ( n403845 , n378424 );
or ( n403846 , n403844 , n403845 );
nand ( n82186 , n82182 , n403846 );
buf ( n403848 , n82186 );
buf ( n403849 , n403848 );
xor ( n403850 , n403832 , n403849 );
xor ( n82190 , n403655 , n403672 );
buf ( n403852 , n82190 );
buf ( n403853 , n403852 );
and ( n82193 , n403850 , n403853 );
and ( n403855 , n403832 , n403849 );
or ( n82195 , n82193 , n403855 );
buf ( n403857 , n82195 );
buf ( n403858 , n395810 );
buf ( n403859 , n380817 );
and ( n403860 , n403858 , n403859 );
buf ( n403861 , n395816 );
not ( n82201 , n57982 );
buf ( n403863 , n82201 );
and ( n403864 , n403861 , n403863 );
nor ( n82204 , n403860 , n403864 );
buf ( n82205 , n82204 );
buf ( n403867 , n82205 );
buf ( n403868 , n60313 );
or ( n82208 , n403867 , n403868 );
buf ( n403870 , n81922 );
buf ( n403871 , n380733 );
or ( n82211 , n403870 , n403871 );
nand ( n403873 , n82208 , n82211 );
buf ( n403874 , n403873 );
xor ( n82214 , n403857 , n403874 );
buf ( n403876 , n396499 );
buf ( n403877 , n382835 );
and ( n82217 , n403876 , n403877 );
buf ( n403879 , n394816 );
buf ( n403880 , n62243 );
and ( n403881 , n403879 , n403880 );
nor ( n403882 , n82217 , n403881 );
buf ( n403883 , n403882 );
buf ( n403884 , n403883 );
buf ( n403885 , n382849 );
or ( n403886 , n403884 , n403885 );
buf ( n403887 , n403699 );
buf ( n403888 , n384157 );
or ( n82228 , n403887 , n403888 );
nand ( n82229 , n403886 , n82228 );
buf ( n403891 , n82229 );
and ( n403892 , n82214 , n403891 );
and ( n82232 , n403857 , n403874 );
or ( n82233 , n403892 , n82232 );
buf ( n403895 , n82233 );
buf ( n403896 , n382795 );
buf ( n403897 , n401882 );
and ( n403898 , n403896 , n403897 );
buf ( n403899 , n382803 );
buf ( n403900 , n384421 );
and ( n82240 , n403899 , n403900 );
nor ( n82241 , n403898 , n82240 );
buf ( n403903 , n82241 );
buf ( n403904 , n403903 );
buf ( n403905 , n384414 );
or ( n82245 , n403904 , n403905 );
buf ( n403907 , n402111 );
buf ( n403908 , n395635 );
or ( n403909 , n403907 , n403908 );
nand ( n82249 , n82245 , n403909 );
buf ( n82250 , n82249 );
buf ( n403912 , n82250 );
xor ( n82252 , n403895 , n403912 );
xor ( n403914 , n403567 , n403622 );
xor ( n403915 , n403914 , n403685 );
buf ( n403916 , n403915 );
buf ( n403917 , n403916 );
and ( n403918 , n82252 , n403917 );
and ( n403919 , n403895 , n403912 );
or ( n82259 , n403918 , n403919 );
buf ( n403921 , n82259 );
xor ( n403922 , n402119 , n402135 );
xor ( n82262 , n403922 , n402139 );
and ( n403924 , n403921 , n82262 );
and ( n403925 , n403749 , n403921 );
or ( n82265 , n403752 , n403924 , n403925 );
xor ( n403927 , n403533 , n403736 );
xor ( n403928 , n403927 , n403740 );
and ( n82268 , n82265 , n403928 );
xor ( n82269 , n403640 , n403675 );
xor ( n82270 , n82269 , n403680 );
buf ( n403932 , n82270 );
buf ( n403933 , n403932 );
buf ( n403934 , n75451 );
buf ( n403935 , n380817 );
and ( n82275 , n403934 , n403935 );
buf ( n403937 , n396596 );
buf ( n403938 , n82201 );
and ( n403939 , n403937 , n403938 );
nor ( n82279 , n82275 , n403939 );
buf ( n82280 , n82279 );
buf ( n403942 , n82280 );
buf ( n403943 , n60313 );
or ( n82283 , n403942 , n403943 );
buf ( n403945 , n82205 );
buf ( n403946 , n380733 );
or ( n82286 , n403945 , n403946 );
nand ( n403948 , n82283 , n82286 );
buf ( n403949 , n403948 );
buf ( n403950 , n403949 );
buf ( n403951 , n79114 );
buf ( n403952 , n57789 );
and ( n403953 , n403951 , n403952 );
buf ( n403954 , n400487 );
buf ( n403955 , n60054 );
and ( n82295 , n403954 , n403955 );
nor ( n82296 , n403953 , n82295 );
buf ( n403958 , n82296 );
buf ( n403959 , n403958 );
buf ( n403960 , n380581 );
or ( n82300 , n403959 , n403960 );
buf ( n403962 , n403631 );
buf ( n403963 , n394774 );
or ( n82303 , n403962 , n403963 );
nand ( n403965 , n82300 , n82303 );
buf ( n403966 , n403965 );
buf ( n403967 , n403966 );
xor ( n403968 , n403950 , n403967 );
buf ( n403969 , n400503 );
buf ( n403970 , n57789 );
and ( n82310 , n403969 , n403970 );
buf ( n403972 , n400509 );
buf ( n403973 , n60054 );
and ( n82313 , n403972 , n403973 );
nor ( n403975 , n82310 , n82313 );
buf ( n403976 , n403975 );
buf ( n403977 , n403976 );
buf ( n403978 , n380581 );
or ( n403979 , n403977 , n403978 );
buf ( n403980 , n403958 );
buf ( n403981 , n394774 );
or ( n403982 , n403980 , n403981 );
nand ( n82322 , n403979 , n403982 );
buf ( n403984 , n82322 );
buf ( n403985 , n403984 );
buf ( n403986 , n80468 );
buf ( n403987 , n57800 );
and ( n403988 , n403986 , n403987 );
buf ( n403989 , n401921 );
buf ( n403990 , n378284 );
and ( n403991 , n403989 , n403990 );
nor ( n82331 , n403988 , n403991 );
buf ( n82332 , n82331 );
buf ( n403994 , n82332 );
buf ( n403995 , n378341 );
or ( n403996 , n403994 , n403995 );
buf ( n403997 , n403840 );
buf ( n403998 , n378424 );
or ( n403999 , n403997 , n403998 );
nand ( n404000 , n403996 , n403999 );
buf ( n404001 , n404000 );
buf ( n404002 , n404001 );
xor ( n82342 , n403985 , n404002 );
xor ( n404004 , n403769 , n403785 );
xor ( n82344 , n404004 , n403827 );
buf ( n404006 , n82344 );
buf ( n82346 , n404006 );
and ( n82347 , n82342 , n82346 );
and ( n82348 , n403985 , n404002 );
or ( n82349 , n82347 , n82348 );
buf ( n82350 , n82349 );
buf ( n404012 , n82350 );
and ( n82352 , n403968 , n404012 );
and ( n82353 , n403950 , n403967 );
or ( n82354 , n82352 , n82353 );
buf ( n404016 , n82354 );
buf ( n404017 , n404016 );
xor ( n404018 , n403933 , n404017 );
buf ( n404019 , n63406 );
buf ( n404020 , n401882 );
and ( n404021 , n404019 , n404020 );
buf ( n404022 , n384054 );
buf ( n404023 , n394730 );
and ( n404024 , n404022 , n404023 );
nor ( n82364 , n404021 , n404024 );
buf ( n82365 , n82364 );
buf ( n404027 , n82365 );
buf ( n404028 , n384414 );
or ( n404029 , n404027 , n404028 );
buf ( n404030 , n403903 );
buf ( n404031 , n395635 );
or ( n82371 , n404030 , n404031 );
nand ( n82372 , n404029 , n82371 );
buf ( n404034 , n82372 );
buf ( n404035 , n404034 );
and ( n82375 , n404018 , n404035 );
and ( n82376 , n403933 , n404017 );
or ( n82377 , n82375 , n82376 );
buf ( n404039 , n82377 );
buf ( n404040 , n404039 );
buf ( n404041 , n380838 );
buf ( n404042 , n394840 );
and ( n82382 , n404041 , n404042 );
buf ( n404044 , n380844 );
buf ( n404045 , n395890 );
and ( n82385 , n404044 , n404045 );
nor ( n82386 , n82382 , n82385 );
buf ( n404048 , n82386 );
buf ( n404049 , n404048 );
buf ( n404050 , n394838 );
or ( n404051 , n404049 , n404050 );
buf ( n404052 , n403541 );
buf ( n404053 , n394835 );
or ( n82393 , n404052 , n404053 );
nand ( n82394 , n404051 , n82393 );
buf ( n404056 , n82394 );
buf ( n404057 , n404056 );
xor ( n404058 , n404040 , n404057 );
xor ( n404059 , n401955 , n80521 );
xor ( n404060 , n404059 , n401996 );
xor ( n82398 , n403707 , n403726 );
xor ( n82399 , n404060 , n82398 );
buf ( n404063 , n82399 );
and ( n404064 , n404058 , n404063 );
and ( n404065 , n404040 , n404057 );
or ( n82403 , n404064 , n404065 );
buf ( n404067 , n82403 );
xor ( n82405 , n403550 , n403690 );
xor ( n404069 , n82405 , n403732 );
buf ( n404070 , n404069 );
xor ( n404071 , n404067 , n404070 );
xor ( n404072 , n402119 , n402135 );
xor ( n82410 , n404072 , n402139 );
xor ( n404074 , n403749 , n403921 );
xor ( n82412 , n82410 , n404074 );
and ( n404076 , n404071 , n82412 );
and ( n82414 , n404067 , n404070 );
or ( n404078 , n404076 , n82414 );
xor ( n82416 , n403533 , n403736 );
xor ( n404080 , n82416 , n403740 );
and ( n404081 , n404078 , n404080 );
and ( n82419 , n82265 , n404078 );
or ( n404083 , n82268 , n404081 , n82419 );
xor ( n82421 , n402157 , n402160 );
xor ( n82422 , n82421 , n402164 );
and ( n404086 , n404083 , n82422 );
and ( n404087 , n403743 , n404083 );
or ( n82425 , n403746 , n404086 , n404087 );
buf ( n404089 , n82425 );
xor ( n404090 , n403530 , n404089 );
buf ( n404091 , n44915 );
not ( n82429 , n404091 );
buf ( n404093 , n365041 );
not ( n404094 , n404093 );
buf ( n404095 , n402185 );
not ( n82433 , n404095 );
or ( n404097 , n404094 , n82433 );
nand ( n82435 , n351345 , n369183 );
buf ( n404099 , n82435 );
nand ( n404100 , n404097 , n404099 );
buf ( n404101 , n404100 );
buf ( n404102 , n404101 );
not ( n82440 , n404102 );
or ( n404104 , n82429 , n82440 );
buf ( n404105 , n365041 );
not ( n82443 , n404105 );
buf ( n404107 , n365384 );
not ( n404108 , n404107 );
or ( n404109 , n82443 , n404108 );
nand ( n82447 , n402205 , n369183 );
buf ( n404111 , n82447 );
nand ( n404112 , n404109 , n404111 );
buf ( n404113 , n404112 );
buf ( n404114 , n404113 );
not ( n404115 , n44912 );
buf ( n404116 , n404115 );
nand ( n82454 , n404114 , n404116 );
buf ( n404118 , n82454 );
buf ( n404119 , n404118 );
nand ( n404120 , n404104 , n404119 );
buf ( n404121 , n404120 );
buf ( n404122 , n404121 );
and ( n404123 , n404090 , n404122 );
and ( n404124 , n403530 , n404089 );
or ( n404125 , n404123 , n404124 );
buf ( n404126 , n404125 );
buf ( n404127 , n404126 );
and ( n404128 , n403525 , n404127 );
and ( n404129 , n403501 , n403524 );
or ( n404130 , n404128 , n404129 );
buf ( n404131 , n404130 );
buf ( n404132 , n404131 );
and ( n404133 , n56970 , n364978 );
not ( n404134 , n56970 );
and ( n404135 , n404134 , n62340 );
or ( n82461 , n404133 , n404135 );
not ( n404137 , n82461 );
not ( n404138 , n365024 );
or ( n82464 , n404137 , n404138 );
buf ( n404140 , n402785 );
buf ( n404141 , n365108 );
nand ( n404142 , n404140 , n404141 );
buf ( n404143 , n404142 );
nand ( n82469 , n82464 , n404143 );
buf ( n404145 , n82469 );
xor ( n82470 , n404132 , n404145 );
and ( n404147 , n22619 , n377782 );
not ( n404148 , n22619 );
and ( n404149 , n404148 , n377779 );
nor ( n82473 , n404147 , n404149 );
buf ( n404151 , n82473 );
not ( n82475 , n404151 );
buf ( n404153 , n365725 );
not ( n82477 , n404153 );
or ( n82478 , n82475 , n82477 );
buf ( n404156 , n403133 );
buf ( n404157 , n56794 );
nand ( n82481 , n404156 , n404157 );
buf ( n404159 , n82481 );
buf ( n404160 , n404159 );
nand ( n404161 , n82478 , n404160 );
buf ( n404162 , n404161 );
buf ( n404163 , n404162 );
and ( n404164 , n82470 , n404163 );
and ( n404165 , n404132 , n404145 );
or ( n404166 , n404164 , n404165 );
buf ( n404167 , n404166 );
buf ( n404168 , n404167 );
xor ( n404169 , n403496 , n404168 );
buf ( n404170 , n377122 );
buf ( n404171 , n58471 );
and ( n404172 , n404170 , n404171 );
not ( n404173 , n404170 );
buf ( n404174 , n386807 );
and ( n404175 , n404173 , n404174 );
nor ( n82486 , n404172 , n404175 );
buf ( n404177 , n82486 );
buf ( n404178 , n404177 );
buf ( n404179 , n50782 );
or ( n82490 , n404178 , n404179 );
buf ( n404181 , n402942 );
buf ( n404182 , n377168 );
or ( n82493 , n404181 , n404182 );
nand ( n404184 , n82490 , n82493 );
buf ( n404185 , n404184 );
buf ( n404186 , n404185 );
and ( n82497 , n404169 , n404186 );
and ( n82498 , n403496 , n404168 );
or ( n82499 , n82497 , n82498 );
buf ( n404190 , n82499 );
buf ( n404191 , n404190 );
nand ( n82502 , n81843 , n404191 );
buf ( n82503 , n82502 );
buf ( n404194 , n82503 );
buf ( n404195 , n403444 );
buf ( n404196 , n403473 );
nand ( n404197 , n404195 , n404196 );
buf ( n404198 , n404197 );
buf ( n404199 , n404198 );
nand ( n404200 , n404194 , n404199 );
buf ( n404201 , n404200 );
buf ( n404202 , n404201 );
nand ( n404203 , n403426 , n404202 );
buf ( n404204 , n404203 );
buf ( n404205 , n404204 );
nand ( n404206 , n403423 , n404205 );
buf ( n404207 , n404206 );
buf ( n404208 , n404207 );
and ( n404209 , n403378 , n404208 );
and ( n404210 , n403373 , n403377 );
or ( n404211 , n404209 , n404210 );
buf ( n404212 , n404211 );
buf ( n404213 , n404212 );
and ( n404214 , n81731 , n404213 );
and ( n404215 , n403362 , n81730 );
or ( n404216 , n404214 , n404215 );
buf ( n404217 , n404216 );
buf ( n404218 , n404217 );
xor ( n404219 , n402562 , n402979 );
xor ( n404220 , n404219 , n402984 );
buf ( n404221 , n404220 );
buf ( n404222 , n404221 );
xor ( n82510 , n404218 , n404222 );
buf ( n404224 , n380356 );
not ( n404225 , n404224 );
buf ( n404226 , n402572 );
not ( n82514 , n404226 );
or ( n82515 , n404225 , n82514 );
buf ( n404229 , n380368 );
not ( n404230 , n404229 );
buf ( n404231 , n374547 );
not ( n404232 , n404231 );
or ( n82520 , n404230 , n404232 );
buf ( n82521 , n361673 );
buf ( n404235 , n380364 );
nand ( n404236 , n82521 , n404235 );
buf ( n404237 , n404236 );
buf ( n404238 , n404237 );
nand ( n404239 , n82520 , n404238 );
buf ( n404240 , n404239 );
buf ( n404241 , n404240 );
buf ( n404242 , n380404 );
nand ( n404243 , n404241 , n404242 );
buf ( n404244 , n404243 );
buf ( n404245 , n404244 );
nand ( n82533 , n82515 , n404245 );
buf ( n404247 , n82533 );
buf ( n404248 , n404247 );
not ( n82536 , n404248 );
buf ( n404250 , n403060 );
not ( n82538 , n404250 );
buf ( n404252 , n381675 );
not ( n82540 , n404252 );
and ( n404254 , n82538 , n82540 );
buf ( n404255 , n379371 );
not ( n82543 , n404255 );
buf ( n404257 , n352119 );
not ( n404258 , n404257 );
or ( n82546 , n82543 , n404258 );
buf ( n404260 , n42355 );
buf ( n404261 , n379392 );
nand ( n82549 , n404260 , n404261 );
buf ( n404263 , n82549 );
buf ( n404264 , n404263 );
nand ( n404265 , n82546 , n404264 );
buf ( n404266 , n404265 );
buf ( n404267 , n404266 );
buf ( n404268 , n58867 );
and ( n404269 , n404267 , n404268 );
nor ( n404270 , n404254 , n404269 );
buf ( n404271 , n404270 );
buf ( n404272 , n404271 );
not ( n404273 , n404272 );
buf ( n404274 , n377068 );
not ( n404275 , n404274 );
buf ( n404276 , n377715 );
not ( n404277 , n404276 );
or ( n404278 , n404275 , n404277 );
buf ( n404279 , n45595 );
buf ( n404280 , n377071 );
nand ( n404281 , n404279 , n404280 );
buf ( n404282 , n404281 );
buf ( n404283 , n404282 );
nand ( n404284 , n404278 , n404283 );
buf ( n404285 , n404284 );
buf ( n404286 , n404285 );
not ( n404287 , n404286 );
buf ( n404288 , n42263 );
not ( n404289 , n404288 );
or ( n404290 , n404287 , n404289 );
buf ( n404291 , n402728 );
buf ( n404292 , n48490 );
nand ( n404293 , n404291 , n404292 );
buf ( n404294 , n404293 );
buf ( n404295 , n404294 );
nand ( n404296 , n404290 , n404295 );
buf ( n404297 , n404296 );
buf ( n404298 , n404297 );
not ( n82561 , n404298 );
and ( n82562 , n398363 , n365259 );
not ( n404301 , n398363 );
and ( n404302 , n404301 , n352212 );
or ( n82565 , n82562 , n404302 );
not ( n404304 , n82565 );
not ( n82566 , n404304 );
not ( n404306 , n377618 );
and ( n404307 , n82566 , n404306 );
and ( n82569 , n403013 , n397190 );
nor ( n82570 , n404307 , n82569 );
buf ( n404310 , n82570 );
not ( n404311 , n404310 );
buf ( n404312 , n404311 );
buf ( n404313 , n404312 );
not ( n404314 , n404313 );
or ( n404315 , n82561 , n404314 );
buf ( n404316 , n404297 );
buf ( n404317 , n404312 );
or ( n404318 , n404316 , n404317 );
buf ( n404319 , n402678 );
buf ( n404320 , n402644 );
xor ( n404321 , n404319 , n404320 );
buf ( n404322 , n402672 );
not ( n404323 , n404322 );
xor ( n404324 , n404321 , n404323 );
buf ( n404325 , n404324 );
buf ( n404326 , n404325 );
nand ( n404327 , n404318 , n404326 );
buf ( n404328 , n404327 );
buf ( n404329 , n404328 );
nand ( n404330 , n404315 , n404329 );
buf ( n82573 , n404330 );
not ( n404332 , n82573 );
buf ( n404333 , n404332 );
not ( n82575 , n404333 );
or ( n82576 , n404273 , n82575 );
xor ( n404336 , n403021 , n403025 );
xor ( n404337 , n404336 , n403042 );
buf ( n404338 , n404337 );
buf ( n404339 , n404338 );
nand ( n82581 , n82576 , n404339 );
buf ( n404341 , n82581 );
buf ( n404342 , n404341 );
buf ( n404343 , n82573 );
not ( n82585 , n404271 );
buf ( n404345 , n82585 );
nand ( n404346 , n404343 , n404345 );
buf ( n404347 , n404346 );
buf ( n404348 , n404347 );
and ( n82590 , n404342 , n404348 );
buf ( n404350 , n82590 );
buf ( n404351 , n404350 );
not ( n82593 , n404351 );
buf ( n82594 , n82593 );
buf ( n404354 , n82594 );
not ( n82596 , n404354 );
or ( n82597 , n82536 , n82596 );
xor ( n82598 , n403091 , n403233 );
xor ( n404358 , n82598 , n403251 );
buf ( n404359 , n404358 );
buf ( n404360 , n404359 );
buf ( n404361 , n404247 );
not ( n82603 , n404361 );
buf ( n404363 , n404350 );
nand ( n404364 , n82603 , n404363 );
buf ( n404365 , n404364 );
buf ( n404366 , n404365 );
nand ( n404367 , n404360 , n404366 );
buf ( n404368 , n404367 );
buf ( n404369 , n404368 );
nand ( n404370 , n82597 , n404369 );
buf ( n404371 , n404370 );
buf ( n404372 , n404371 );
buf ( n404373 , n402966 );
not ( n404374 , n404373 );
buf ( n404375 , n402585 );
not ( n404376 , n404375 );
or ( n82618 , n404374 , n404376 );
buf ( n404378 , n402585 );
buf ( n404379 , n402966 );
or ( n404380 , n404378 , n404379 );
nand ( n82622 , n82618 , n404380 );
buf ( n82623 , n82622 );
xnor ( n404383 , n81073 , n82623 );
buf ( n404384 , n404383 );
xor ( n404385 , n404372 , n404384 );
buf ( n404386 , n81493 );
not ( n82628 , n404386 );
buf ( n404388 , n403255 );
not ( n404389 , n404388 );
or ( n82631 , n82628 , n404389 );
buf ( n82632 , n81493 );
buf ( n82633 , n403255 );
or ( n82634 , n82632 , n82633 );
nand ( n82635 , n82631 , n82634 );
buf ( n82636 , n82635 );
xnor ( n404396 , n403084 , n82636 );
buf ( n404397 , n404396 );
and ( n82639 , n404385 , n404397 );
and ( n404399 , n404372 , n404384 );
or ( n404400 , n82639 , n404399 );
buf ( n404401 , n404400 );
buf ( n404402 , n404401 );
and ( n404403 , n82510 , n404402 );
and ( n404404 , n404218 , n404222 );
or ( n404405 , n404403 , n404404 );
buf ( n404406 , n404405 );
buf ( n404407 , n404406 );
or ( n82649 , n403351 , n404407 );
buf ( n404409 , n82649 );
not ( n404410 , n404409 );
or ( n82652 , n403326 , n404410 );
buf ( n404412 , n404406 );
buf ( n404413 , n403350 );
nand ( n404414 , n404412 , n404413 );
buf ( n404415 , n404414 );
nand ( n404416 , n82652 , n404415 );
not ( n404417 , n404416 );
buf ( n404418 , n81671 );
buf ( n404419 , n402535 );
and ( n404420 , n404418 , n404419 );
not ( n404421 , n404418 );
buf ( n404422 , n402538 );
and ( n404423 , n404421 , n404422 );
nor ( n404424 , n404420 , n404423 );
buf ( n404425 , n404424 );
buf ( n404426 , n404425 );
buf ( n404427 , n403311 );
not ( n404428 , n404427 );
buf ( n404429 , n404428 );
buf ( n404430 , n404429 );
and ( n82672 , n404426 , n404430 );
not ( n404432 , n404426 );
buf ( n404433 , n403311 );
and ( n82675 , n404432 , n404433 );
nor ( n404435 , n82672 , n82675 );
buf ( n404436 , n404435 );
nand ( n82678 , n404417 , n404436 );
buf ( n404438 , n82678 );
and ( n404439 , n403322 , n404438 );
buf ( n404440 , n404439 );
buf ( n404441 , n404440 );
xor ( n82683 , n402389 , n402393 );
and ( n404443 , n82683 , n402503 );
and ( n82685 , n402389 , n402393 );
or ( n82686 , n404443 , n82685 );
buf ( n404446 , n82686 );
buf ( n404447 , n404446 );
xor ( n404448 , n399098 , n399517 );
xor ( n82690 , n404448 , n399678 );
buf ( n404450 , n82690 );
buf ( n404451 , n404450 );
and ( n404452 , n404447 , n404451 );
not ( n404453 , n404447 );
buf ( n404454 , n404450 );
not ( n82696 , n404454 );
buf ( n404456 , n82696 );
buf ( n404457 , n404456 );
and ( n82699 , n404453 , n404457 );
nor ( n82700 , n404452 , n82699 );
buf ( n82701 , n82700 );
buf ( n404461 , n398528 );
buf ( n404462 , n398591 );
xor ( n82704 , n404461 , n404462 );
buf ( n404464 , n398539 );
xnor ( n404465 , n82704 , n404464 );
buf ( n404466 , n404465 );
not ( n82708 , n404466 );
and ( n404468 , n77312 , n398611 );
not ( n82710 , n77312 );
and ( n82711 , n82710 , n398608 );
nor ( n404471 , n404468 , n82711 );
buf ( n404472 , n398764 );
not ( n82714 , n404472 );
buf ( n404474 , n82714 );
and ( n404475 , n404471 , n404474 );
not ( n82717 , n404471 );
and ( n82718 , n82717 , n398764 );
nor ( n404478 , n404475 , n82718 );
not ( n404479 , n404478 );
not ( n82721 , n404479 );
or ( n82722 , n82708 , n82721 );
or ( n82723 , n404466 , n404479 );
nand ( n404483 , n82722 , n82723 );
buf ( n404484 , n404483 );
not ( n82726 , n404484 );
xor ( n82727 , n401070 , n401074 );
and ( n82728 , n82727 , n401369 );
and ( n404488 , n401070 , n401074 );
or ( n82730 , n82728 , n404488 );
buf ( n404490 , n82730 );
buf ( n404491 , n404490 );
not ( n82733 , n404491 );
buf ( n404493 , n82733 );
buf ( n404494 , n404493 );
not ( n82736 , n404494 );
and ( n82737 , n82726 , n82736 );
buf ( n404497 , n404493 );
buf ( n404498 , n404483 );
and ( n82740 , n404497 , n404498 );
nor ( n404500 , n82737 , n82740 );
buf ( n404501 , n404500 );
and ( n404502 , n82701 , n404501 );
not ( n82744 , n82701 );
buf ( n404504 , n404501 );
not ( n82746 , n404504 );
buf ( n404506 , n82746 );
and ( n82748 , n82744 , n404506 );
nor ( n82749 , n404502 , n82748 );
xor ( n404509 , n401372 , n402384 );
and ( n82751 , n404509 , n402506 );
and ( n82752 , n401372 , n402384 );
or ( n404512 , n82751 , n82752 );
buf ( n404513 , n404512 );
not ( n82755 , n404513 );
nand ( n82756 , n82749 , n82755 );
buf ( n404516 , n82756 );
and ( n82758 , n404441 , n404516 );
buf ( n82759 , n82758 );
xor ( n404519 , n404218 , n404222 );
xor ( n82761 , n404519 , n404402 );
buf ( n404521 , n82761 );
xor ( n404522 , n402693 , n81186 );
xor ( n404523 , n404522 , n402962 );
buf ( n404524 , n404523 );
buf ( n404525 , n404524 );
xor ( n404526 , n403047 , n403051 );
xor ( n404527 , n404526 , n403069 );
buf ( n404528 , n404527 );
buf ( n404529 , n404528 );
xor ( n404530 , n404525 , n404529 );
xor ( n82772 , n402826 , n402933 );
xor ( n82773 , n82772 , n402951 );
buf ( n404533 , n82773 );
buf ( n404534 , n404533 );
buf ( n404535 , n379890 );
not ( n82777 , n404535 );
buf ( n404537 , n403109 );
not ( n404538 , n404537 );
or ( n404539 , n82777 , n404538 );
buf ( n404540 , n379838 );
not ( n404541 , n404540 );
buf ( n404542 , n364870 );
not ( n404543 , n404542 );
or ( n404544 , n404541 , n404543 );
buf ( n404545 , n364858 );
buf ( n404546 , n398741 );
nand ( n404547 , n404545 , n404546 );
buf ( n404548 , n404547 );
buf ( n404549 , n404548 );
nand ( n404550 , n404544 , n404549 );
buf ( n404551 , n404550 );
buf ( n404552 , n404551 );
buf ( n404553 , n379916 );
nand ( n404554 , n404552 , n404553 );
buf ( n404555 , n404554 );
buf ( n404556 , n404555 );
nand ( n404557 , n404539 , n404556 );
buf ( n82780 , n404557 );
buf ( n82781 , n82780 );
xor ( n82782 , n404534 , n82781 );
buf ( n82783 , n379263 );
not ( n82784 , n82783 );
buf ( n82785 , n403039 );
not ( n82786 , n82785 );
buf ( n82787 , n82786 );
buf ( n82788 , n82787 );
not ( n82789 , n82788 );
or ( n82790 , n82784 , n82789 );
buf ( n404569 , n379274 );
not ( n404570 , n404569 );
buf ( n404571 , n351318 );
not ( n404572 , n404571 );
or ( n404573 , n404570 , n404572 );
buf ( n404574 , n365561 );
buf ( n404575 , n379271 );
nand ( n404576 , n404574 , n404575 );
buf ( n404577 , n404576 );
buf ( n404578 , n404577 );
nand ( n82801 , n404573 , n404578 );
buf ( n404580 , n82801 );
buf ( n404581 , n404580 );
buf ( n404582 , n379299 );
nand ( n404583 , n404581 , n404582 );
buf ( n404584 , n404583 );
buf ( n404585 , n404584 );
nand ( n404586 , n82790 , n404585 );
buf ( n404587 , n404586 );
buf ( n404588 , n404587 );
and ( n404589 , n82782 , n404588 );
and ( n404590 , n404534 , n82781 );
or ( n82813 , n404589 , n404590 );
buf ( n404592 , n82813 );
buf ( n82815 , n404592 );
buf ( n404594 , n380404 );
not ( n82817 , n404594 );
buf ( n404596 , n380368 );
not ( n404597 , n404596 );
buf ( n404598 , n43377 );
not ( n404599 , n404598 );
or ( n404600 , n404597 , n404599 );
buf ( n404601 , n361717 );
buf ( n404602 , n384667 );
nand ( n82824 , n404601 , n404602 );
buf ( n404604 , n82824 );
buf ( n404605 , n404604 );
nand ( n404606 , n404600 , n404605 );
buf ( n404607 , n404606 );
buf ( n82829 , n404607 );
not ( n82830 , n82829 );
or ( n82831 , n82817 , n82830 );
buf ( n82832 , n404240 );
buf ( n404612 , n380356 );
nand ( n82834 , n82832 , n404612 );
buf ( n404614 , n82834 );
buf ( n404615 , n404614 );
nand ( n404616 , n82831 , n404615 );
buf ( n404617 , n404616 );
buf ( n404618 , n404617 );
xor ( n404619 , n82815 , n404618 );
buf ( n404620 , n402955 );
buf ( n404621 , n402749 );
xor ( n404622 , n404620 , n404621 );
buf ( n404623 , n81211 );
xor ( n404624 , n404622 , n404623 );
buf ( n404625 , n404624 );
buf ( n404626 , n404625 );
and ( n404627 , n404619 , n404626 );
and ( n404628 , n82815 , n404618 );
or ( n404629 , n404627 , n404628 );
buf ( n404630 , n404629 );
buf ( n404631 , n404630 );
and ( n404632 , n404530 , n404631 );
and ( n404633 , n404525 , n404529 );
or ( n82855 , n404632 , n404633 );
buf ( n404635 , n82855 );
buf ( n404636 , n404635 );
not ( n82858 , n404636 );
xor ( n404638 , n403362 , n81730 );
xor ( n404639 , n404638 , n404213 );
buf ( n404640 , n404639 );
buf ( n404641 , n404640 );
not ( n82863 , n404641 );
or ( n404643 , n82858 , n82863 );
buf ( n404644 , n404640 );
buf ( n404645 , n404635 );
or ( n404646 , n404644 , n404645 );
not ( n404647 , n82585 );
not ( n82869 , n404332 );
or ( n404649 , n404647 , n82869 );
nand ( n404650 , n82573 , n404271 );
nand ( n82872 , n404649 , n404650 );
buf ( n404652 , n404338 );
not ( n404653 , n404652 );
buf ( n404654 , n404653 );
and ( n404655 , n82872 , n404654 );
not ( n82877 , n82872 );
and ( n404657 , n82877 , n404338 );
nor ( n404658 , n404655 , n404657 );
not ( n82880 , n404658 );
not ( n404660 , n82880 );
buf ( n404661 , n403444 );
buf ( n404662 , n403473 );
and ( n404663 , n404661 , n404662 );
not ( n82885 , n404661 );
buf ( n404665 , n403476 );
and ( n82887 , n82885 , n404665 );
nor ( n82888 , n404663 , n82887 );
buf ( n404668 , n82888 );
buf ( n404669 , n404668 );
buf ( n404670 , n404190 );
xnor ( n404671 , n404669 , n404670 );
buf ( n404672 , n404671 );
buf ( n404673 , n404672 );
xor ( n404674 , n82570 , n404325 );
xor ( n404675 , n404297 , n404674 );
buf ( n404676 , n404675 );
nand ( n404677 , n404673 , n404676 );
buf ( n404678 , n404677 );
buf ( n404679 , n404678 );
xor ( n404680 , n403146 , n403171 );
xor ( n404681 , n404680 , n403176 );
buf ( n404682 , n404681 );
buf ( n404683 , n404682 );
buf ( n404684 , n379299 );
not ( n82906 , n404684 );
buf ( n404686 , n379274 );
not ( n404687 , n404686 );
buf ( n404688 , n32160 );
not ( n82910 , n404688 );
or ( n404690 , n404687 , n82910 );
buf ( n404691 , n400289 );
buf ( n404692 , n379271 );
nand ( n404693 , n404691 , n404692 );
buf ( n404694 , n404693 );
buf ( n404695 , n404694 );
nand ( n82917 , n404690 , n404695 );
buf ( n404697 , n82917 );
buf ( n404698 , n404697 );
not ( n404699 , n404698 );
or ( n404700 , n82906 , n404699 );
buf ( n82922 , n404580 );
buf ( n82923 , n379263 );
nand ( n82924 , n82922 , n82923 );
buf ( n82925 , n82924 );
buf ( n404705 , n82925 );
nand ( n82927 , n404700 , n404705 );
buf ( n82928 , n82927 );
buf ( n404708 , n82928 );
xor ( n82930 , n404683 , n404708 );
xor ( n82931 , n404132 , n404145 );
xor ( n82932 , n82931 , n404163 );
buf ( n404712 , n82932 );
buf ( n404713 , n404712 );
buf ( n404714 , n397190 );
not ( n82936 , n404714 );
buf ( n404716 , n398363 );
not ( n404717 , n404716 );
buf ( n404718 , n377297 );
not ( n82940 , n404718 );
or ( n404720 , n404717 , n82940 );
buf ( n404721 , n31260 );
buf ( n404722 , n377592 );
nand ( n404723 , n404721 , n404722 );
buf ( n404724 , n404723 );
buf ( n404725 , n404724 );
nand ( n404726 , n404720 , n404725 );
buf ( n404727 , n404726 );
buf ( n404728 , n404727 );
not ( n404729 , n404728 );
or ( n404730 , n82936 , n404729 );
buf ( n404731 , n398363 );
not ( n404732 , n404731 );
buf ( n404733 , n386837 );
not ( n404734 , n404733 );
or ( n404735 , n404732 , n404734 );
buf ( n404736 , n32202 );
buf ( n404737 , n377592 );
nand ( n404738 , n404736 , n404737 );
buf ( n404739 , n404738 );
buf ( n404740 , n404739 );
nand ( n82950 , n404735 , n404740 );
buf ( n404742 , n82950 );
buf ( n82952 , n404742 );
buf ( n404744 , n57530 );
nand ( n82954 , n82952 , n404744 );
buf ( n404746 , n82954 );
buf ( n404747 , n404746 );
nand ( n404748 , n404730 , n404747 );
buf ( n404749 , n404748 );
buf ( n404750 , n404749 );
xor ( n404751 , n404713 , n404750 );
buf ( n404752 , n50782 );
buf ( n404753 , n58463 );
buf ( n404754 , n379482 );
and ( n82964 , n404753 , n404754 );
buf ( n404756 , n396289 );
buf ( n404757 , n58984 );
and ( n82967 , n404756 , n404757 );
nor ( n404759 , n82964 , n82967 );
buf ( n404760 , n404759 );
buf ( n404761 , n404760 );
or ( n404762 , n404752 , n404761 );
buf ( n404763 , n404177 );
buf ( n404764 , n386027 );
or ( n404765 , n404763 , n404764 );
nand ( n404766 , n404762 , n404765 );
buf ( n404767 , n404766 );
buf ( n404768 , n404767 );
and ( n404769 , n404751 , n404768 );
and ( n404770 , n404713 , n404750 );
or ( n404771 , n404769 , n404770 );
buf ( n404772 , n404771 );
buf ( n404773 , n404772 );
and ( n404774 , n82930 , n404773 );
and ( n404775 , n404683 , n404708 );
or ( n404776 , n404774 , n404775 );
buf ( n404777 , n404776 );
buf ( n404778 , n404777 );
and ( n404779 , n404679 , n404778 );
buf ( n404780 , n404675 );
buf ( n404781 , n404672 );
nor ( n404782 , n404780 , n404781 );
buf ( n404783 , n404782 );
buf ( n404784 , n404783 );
nor ( n404785 , n404779 , n404784 );
buf ( n404786 , n404785 );
buf ( n404787 , n404786 );
not ( n404788 , n404787 );
buf ( n404789 , n404788 );
not ( n404790 , n404789 );
or ( n404791 , n404660 , n404790 );
buf ( n404792 , n404786 );
not ( n404793 , n404792 );
buf ( n404794 , n404658 );
not ( n404795 , n404794 );
or ( n82982 , n404793 , n404795 );
buf ( n404797 , n378098 );
buf ( n404798 , n366329 );
and ( n82985 , n404797 , n404798 );
not ( n404800 , n404797 );
buf ( n404801 , n41772 );
and ( n82988 , n404800 , n404801 );
nor ( n404803 , n82985 , n82988 );
buf ( n404804 , n404803 );
buf ( n404805 , n404804 );
not ( n404806 , n404805 );
buf ( n82993 , n367759 );
not ( n82994 , n82993 );
or ( n82995 , n404806 , n82994 );
buf ( n82996 , n403408 );
buf ( n404811 , n41835 );
nand ( n82998 , n82996 , n404811 );
buf ( n404813 , n82998 );
buf ( n404814 , n404813 );
nand ( n83001 , n82995 , n404814 );
buf ( n404816 , n83001 );
not ( n404817 , n404816 );
buf ( n404818 , n58923 );
not ( n404819 , n404818 );
buf ( n404820 , n404266 );
not ( n83007 , n404820 );
or ( n404822 , n404819 , n83007 );
buf ( n404823 , n379371 );
not ( n83010 , n404823 );
buf ( n404825 , n364771 );
not ( n404826 , n404825 );
or ( n83013 , n83010 , n404826 );
buf ( n404828 , n49988 );
not ( n404829 , n404828 );
buf ( n404830 , n379392 );
nand ( n404831 , n404829 , n404830 );
buf ( n404832 , n404831 );
buf ( n404833 , n404832 );
nand ( n404834 , n83013 , n404833 );
buf ( n404835 , n404834 );
buf ( n404836 , n404835 );
buf ( n404837 , n58867 );
nand ( n83023 , n404836 , n404837 );
buf ( n404839 , n83023 );
buf ( n404840 , n404839 );
nand ( n404841 , n404822 , n404840 );
buf ( n404842 , n404841 );
buf ( n404843 , n404842 );
not ( n404844 , n404843 );
buf ( n404845 , n404844 );
nand ( n83031 , n404817 , n404845 );
not ( n404847 , n83031 );
xor ( n404848 , n403496 , n404168 );
xor ( n83034 , n404848 , n404186 );
buf ( n404850 , n83034 );
buf ( n404851 , n404850 );
buf ( n404852 , n377757 );
not ( n404853 , n404852 );
buf ( n404854 , n61903 );
not ( n83040 , n404854 );
or ( n404856 , n404853 , n83040 );
buf ( n404857 , n22619 );
buf ( n404858 , n378886 );
nand ( n404859 , n404857 , n404858 );
buf ( n404860 , n404859 );
buf ( n404861 , n404860 );
nand ( n404862 , n404856 , n404861 );
buf ( n404863 , n404862 );
buf ( n404864 , n404863 );
not ( n83050 , n404864 );
buf ( n404866 , n365725 );
not ( n404867 , n404866 );
or ( n404868 , n83050 , n404867 );
buf ( n404869 , n82473 );
buf ( n404870 , n56794 );
nand ( n83056 , n404869 , n404870 );
buf ( n404872 , n83056 );
buf ( n404873 , n404872 );
nand ( n404874 , n404868 , n404873 );
buf ( n404875 , n404874 );
buf ( n404876 , n404875 );
buf ( n404877 , n369809 );
not ( n404878 , n404877 );
buf ( n404879 , n393883 );
not ( n404880 , n404879 );
buf ( n404881 , n351228 );
not ( n404882 , n404881 );
or ( n83068 , n404880 , n404882 );
not ( n83069 , n351228 );
buf ( n83070 , n83069 );
buf ( n83071 , n369763 );
nand ( n83072 , n83070 , n83071 );
buf ( n83073 , n83072 );
buf ( n83074 , n83073 );
nand ( n83075 , n83068 , n83074 );
buf ( n83076 , n83075 );
buf ( n404892 , n83076 );
not ( n83078 , n404892 );
or ( n404894 , n404878 , n83078 );
buf ( n404895 , n393883 );
not ( n83081 , n404895 );
buf ( n404897 , n378543 );
not ( n404898 , n404897 );
or ( n83084 , n83081 , n404898 );
buf ( n404900 , n378543 );
not ( n404901 , n404900 );
buf ( n404902 , n404901 );
buf ( n404903 , n404902 );
buf ( n83089 , n369763 );
nand ( n83090 , n404903 , n83089 );
buf ( n404906 , n83090 );
buf ( n404907 , n404906 );
nand ( n83093 , n83084 , n404907 );
buf ( n404909 , n83093 );
buf ( n404910 , n404909 );
buf ( n404911 , n369804 );
nand ( n83097 , n404910 , n404911 );
buf ( n404913 , n83097 );
buf ( n404914 , n404913 );
nand ( n404915 , n404894 , n404914 );
buf ( n404916 , n404915 );
buf ( n404917 , n404916 );
xor ( n404918 , n404876 , n404917 );
buf ( n404919 , n377782 );
not ( n404920 , n404919 );
buf ( n404921 , n396004 );
not ( n404922 , n404921 );
or ( n404923 , n404920 , n404922 );
buf ( n404924 , n386093 );
buf ( n404925 , n377779 );
nand ( n404926 , n404924 , n404925 );
buf ( n404927 , n404926 );
buf ( n404928 , n404927 );
nand ( n404929 , n404923 , n404928 );
buf ( n404930 , n404929 );
buf ( n404931 , n404930 );
not ( n83104 , n404931 );
buf ( n404933 , n365024 );
not ( n404934 , n404933 );
or ( n83107 , n83104 , n404934 );
buf ( n404936 , n377352 );
buf ( n404937 , n386102 );
and ( n404938 , n404936 , n404937 );
not ( n83111 , n404936 );
buf ( n404940 , n76415 );
and ( n404941 , n83111 , n404940 );
nor ( n404942 , n404938 , n404941 );
buf ( n404943 , n404942 );
buf ( n404944 , n404943 );
buf ( n404945 , n365108 );
nand ( n404946 , n404944 , n404945 );
buf ( n404947 , n404946 );
buf ( n404948 , n404947 );
nand ( n404949 , n83107 , n404948 );
buf ( n404950 , n404949 );
buf ( n404951 , n404950 );
buf ( n404952 , n368621 );
not ( n404953 , n404952 );
buf ( n404954 , n400105 );
not ( n83113 , n404954 );
buf ( n404956 , n63344 );
not ( n404957 , n404956 );
or ( n83116 , n83113 , n404957 );
buf ( n404959 , n63345 );
buf ( n404960 , n380424 );
nand ( n404961 , n404959 , n404960 );
buf ( n404962 , n404961 );
buf ( n404963 , n404962 );
nand ( n83122 , n83116 , n404963 );
buf ( n404965 , n83122 );
buf ( n404966 , n404965 );
not ( n83125 , n404966 );
or ( n404968 , n404953 , n83125 );
buf ( n404969 , n400105 );
not ( n404970 , n404969 );
buf ( n404971 , n60751 );
not ( n404972 , n404971 );
or ( n404973 , n404970 , n404972 );
buf ( n404974 , n45802 );
buf ( n404975 , n380424 );
nand ( n83134 , n404974 , n404975 );
buf ( n404977 , n83134 );
buf ( n404978 , n404977 );
nand ( n404979 , n404973 , n404978 );
buf ( n404980 , n404979 );
buf ( n404981 , n404980 );
buf ( n404982 , n368602 );
nand ( n83141 , n404981 , n404982 );
buf ( n83142 , n83141 );
buf ( n404985 , n83142 );
nand ( n404986 , n404968 , n404985 );
buf ( n404987 , n404986 );
buf ( n404988 , n404987 );
or ( n404989 , n404951 , n404988 );
xor ( n83148 , n403530 , n404089 );
xor ( n404991 , n83148 , n404122 );
buf ( n404992 , n404991 );
buf ( n404993 , n404992 );
nand ( n83152 , n404989 , n404993 );
buf ( n83153 , n83152 );
buf ( n404996 , n83153 );
buf ( n404997 , n404950 );
buf ( n404998 , n404987 );
nand ( n404999 , n404997 , n404998 );
buf ( n405000 , n404999 );
buf ( n405001 , n405000 );
nand ( n405002 , n404996 , n405001 );
buf ( n405003 , n405002 );
buf ( n405004 , n405003 );
and ( n405005 , n404918 , n405004 );
and ( n405006 , n404876 , n404917 );
or ( n405007 , n405005 , n405006 );
buf ( n405008 , n405007 );
buf ( n405009 , n405008 );
not ( n405010 , n405009 );
buf ( n405011 , n405010 );
buf ( n405012 , n405011 );
not ( n405013 , n405012 );
nand ( n405014 , n22769 , n342019 );
not ( n405015 , n342718 );
not ( n83160 , n42254 );
or ( n83161 , n405015 , n83160 );
nand ( n405018 , n83161 , n378098 );
nand ( n405019 , n405014 , n405018 , n45595 );
buf ( n405020 , n405019 );
not ( n83165 , n405020 );
or ( n405022 , n405013 , n83165 );
buf ( n405023 , n44915 );
not ( n83168 , n405023 );
buf ( n405025 , n402874 );
not ( n405026 , n405025 );
or ( n83171 , n83168 , n405026 );
buf ( n405028 , n404101 );
buf ( n405029 , n404115 );
nand ( n83174 , n405028 , n405029 );
buf ( n405031 , n83174 );
buf ( n405032 , n405031 );
nand ( n83177 , n83171 , n405032 );
buf ( n405034 , n83177 );
buf ( n405035 , n405034 );
and ( n405036 , n369374 , n386040 );
not ( n83181 , n369374 );
and ( n83182 , n83181 , n396441 );
or ( n83183 , n405036 , n83182 );
buf ( n405040 , n83183 );
not ( n405041 , n405040 );
buf ( n405042 , n45055 );
not ( n405043 , n405042 );
or ( n83188 , n405041 , n405043 );
buf ( n405045 , n402899 );
buf ( n405046 , n365242 );
nand ( n405047 , n405045 , n405046 );
buf ( n405048 , n405047 );
buf ( n83193 , n405048 );
nand ( n83194 , n83188 , n83193 );
buf ( n83195 , n83194 );
buf ( n405052 , n83195 );
xor ( n83197 , n405035 , n405052 );
buf ( n405054 , n404943 );
not ( n405055 , n405054 );
buf ( n405056 , n405055 );
or ( n405057 , n44862 , n405056 );
not ( n83202 , n44946 );
nand ( n405059 , n83202 , n82461 );
nand ( n405060 , n405057 , n405059 );
buf ( n405061 , n405060 );
and ( n83206 , n83197 , n405061 );
and ( n405063 , n405035 , n405052 );
or ( n405064 , n83206 , n405063 );
buf ( n405065 , n405064 );
xor ( n83210 , n402921 , n402911 );
xor ( n405067 , n83210 , n81353 );
not ( n405068 , n387542 );
not ( n83213 , n402848 );
or ( n83214 , n405068 , n83213 );
buf ( n405071 , n400105 );
not ( n405072 , n405071 );
buf ( n405073 , n394004 );
not ( n405074 , n405073 );
or ( n405075 , n405072 , n405074 );
buf ( n405076 , n351160 );
buf ( n405077 , n380424 );
nand ( n405078 , n405076 , n405077 );
buf ( n405079 , n405078 );
buf ( n405080 , n405079 );
nand ( n83225 , n405075 , n405080 );
buf ( n83226 , n83225 );
buf ( n405083 , n83226 );
buf ( n405084 , n368602 );
nand ( n405085 , n405083 , n405084 );
buf ( n405086 , n405085 );
nand ( n83231 , n83214 , n405086 );
not ( n83232 , n83231 );
and ( n405089 , n405067 , n83232 );
not ( n405090 , n405067 );
and ( n83235 , n405090 , n83231 );
nor ( n83236 , n405089 , n83235 );
xor ( n83237 , n405065 , n83236 );
buf ( n405094 , n83237 );
nand ( n83239 , n405022 , n405094 );
buf ( n405096 , n83239 );
buf ( n405097 , n405096 );
buf ( n405098 , n405019 );
not ( n405099 , n405098 );
buf ( n405100 , n405008 );
nand ( n405101 , n405099 , n405100 );
buf ( n405102 , n405101 );
buf ( n405103 , n405102 );
nand ( n405104 , n405097 , n405103 );
buf ( n405105 , n405104 );
buf ( n405106 , n405105 );
xor ( n83251 , n404851 , n405106 );
buf ( n405108 , n404285 );
not ( n405109 , n405108 );
buf ( n405110 , n42242 );
not ( n405111 , n405110 );
or ( n405112 , n405109 , n405111 );
buf ( n405113 , n42266 );
buf ( n405114 , n365915 );
buf ( n405115 , n56687 );
and ( n405116 , n405114 , n405115 );
buf ( n405117 , n377715 );
buf ( n405118 , n377094 );
and ( n83263 , n405117 , n405118 );
nor ( n405120 , n405116 , n83263 );
buf ( n405121 , n405120 );
buf ( n405122 , n405121 );
or ( n405123 , n405113 , n405122 );
nand ( n83268 , n405112 , n405123 );
buf ( n83269 , n83268 );
buf ( n405126 , n83269 );
and ( n83271 , n83251 , n405126 );
and ( n405128 , n404851 , n405106 );
or ( n405129 , n83271 , n405128 );
buf ( n405130 , n405129 );
not ( n83275 , n405130 );
or ( n83276 , n404847 , n83275 );
buf ( n405133 , n404842 );
buf ( n405134 , n404816 );
nand ( n83279 , n405133 , n405134 );
buf ( n405136 , n83279 );
nand ( n83281 , n83276 , n405136 );
buf ( n405138 , n83281 );
nand ( n83283 , n82982 , n405138 );
buf ( n405140 , n83283 );
nand ( n83285 , n404791 , n405140 );
not ( n83286 , n83285 );
xor ( n83287 , n403373 , n403377 );
xor ( n83288 , n83287 , n404208 );
buf ( n405145 , n83288 );
buf ( n405146 , n405145 );
not ( n83291 , n405146 );
buf ( n405148 , n365311 );
buf ( n405149 , n378098 );
nand ( n83294 , n405148 , n405149 );
buf ( n405151 , n83294 );
not ( n83296 , n405151 );
xor ( n405153 , n81301 , n402856 );
xor ( n405154 , n405153 , n402928 );
buf ( n405155 , n405154 );
buf ( n405156 , n405155 );
not ( n83301 , n405156 );
buf ( n405158 , n83301 );
not ( n83303 , n405158 );
and ( n405160 , n83296 , n83303 );
buf ( n405161 , n405151 );
buf ( n405162 , n405158 );
nand ( n83307 , n405161 , n405162 );
buf ( n405164 , n83307 );
buf ( n405165 , n83231 );
buf ( n405166 , n405065 );
or ( n405167 , n405165 , n405166 );
buf ( n405168 , n405067 );
not ( n83313 , n405168 );
buf ( n405170 , n83313 );
buf ( n405171 , n405170 );
nand ( n83316 , n405167 , n405171 );
buf ( n405173 , n83316 );
buf ( n405174 , n405173 );
buf ( n405175 , n83231 );
buf ( n405176 , n405065 );
nand ( n405177 , n405175 , n405176 );
buf ( n405178 , n405177 );
buf ( n405179 , n405178 );
nand ( n83324 , n405174 , n405179 );
buf ( n405181 , n83324 );
and ( n83326 , n405164 , n405181 );
nor ( n405183 , n405160 , n83326 );
buf ( n83328 , n405183 );
buf ( n405185 , n403215 );
buf ( n405186 , n403180 );
xor ( n83331 , n405185 , n405186 );
buf ( n405188 , n403206 );
xnor ( n405189 , n83331 , n405188 );
buf ( n405190 , n405189 );
buf ( n405191 , n405190 );
xor ( n83336 , n83328 , n405191 );
buf ( n405193 , n397190 );
not ( n405194 , n405193 );
buf ( n405195 , n82565 );
not ( n83340 , n405195 );
or ( n405197 , n405194 , n83340 );
buf ( n405198 , n404727 );
buf ( n405199 , n57530 );
nand ( n83344 , n405198 , n405199 );
buf ( n405201 , n83344 );
buf ( n405202 , n405201 );
nand ( n405203 , n405197 , n405202 );
buf ( n405204 , n405203 );
buf ( n405205 , n405204 );
not ( n405206 , n405205 );
not ( n405207 , n363429 );
buf ( n405208 , n405207 );
not ( n405209 , n405208 );
buf ( n405210 , n378847 );
buf ( n405211 , n22768 );
and ( n405212 , n405210 , n405211 );
not ( n405213 , n405210 );
buf ( n405214 , n362377 );
and ( n405215 , n405213 , n405214 );
or ( n83360 , n405212 , n405215 );
buf ( n405217 , n83360 );
buf ( n405218 , n405217 );
not ( n405219 , n405218 );
and ( n83364 , n405209 , n405219 );
buf ( n405221 , n403461 );
not ( n405222 , n405221 );
buf ( n405223 , n398693 );
nor ( n405224 , n405222 , n405223 );
buf ( n405225 , n405224 );
buf ( n405226 , n405225 );
nor ( n83371 , n83364 , n405226 );
buf ( n405228 , n83371 );
buf ( n405229 , n405228 );
nand ( n83374 , n405206 , n405229 );
buf ( n405231 , n83374 );
buf ( n405232 , n405231 );
buf ( n405233 , n377143 );
not ( n83378 , n405233 );
buf ( n405235 , n388576 );
not ( n405236 , n405235 );
or ( n83381 , n83378 , n405236 );
buf ( n405238 , n378135 );
buf ( n405239 , n377153 );
nand ( n83384 , n405238 , n405239 );
buf ( n405241 , n83384 );
buf ( n405242 , n405241 );
nand ( n83387 , n83381 , n405242 );
buf ( n405244 , n83387 );
buf ( n405245 , n405244 );
not ( n405246 , n405245 );
buf ( n405247 , n375896 );
not ( n405248 , n405247 );
or ( n405249 , n405246 , n405248 );
buf ( n405250 , n403158 );
buf ( n405251 , n375920 );
nand ( n405252 , n405250 , n405251 );
buf ( n405253 , n405252 );
buf ( n405254 , n405253 );
nand ( n405255 , n405249 , n405254 );
buf ( n405256 , n405255 );
buf ( n405257 , n405256 );
not ( n405258 , n405257 );
buf ( n405259 , n405258 );
buf ( n405260 , n405259 );
not ( n405261 , n405260 );
buf ( n405262 , n369809 );
not ( n405263 , n405262 );
buf ( n405264 , n81852 );
not ( n405265 , n405264 );
or ( n405266 , n405263 , n405265 );
buf ( n405267 , n83076 );
buf ( n405268 , n369804 );
nand ( n405269 , n405267 , n405268 );
buf ( n405270 , n405269 );
buf ( n405271 , n405270 );
nand ( n405272 , n405266 , n405271 );
buf ( n405273 , n405272 );
buf ( n405274 , n405273 );
not ( n83391 , n405274 );
buf ( n405276 , n83391 );
buf ( n405277 , n405276 );
not ( n83392 , n405277 );
or ( n405279 , n405261 , n83392 );
xor ( n405280 , n403501 , n403524 );
xor ( n83395 , n405280 , n404127 );
buf ( n405282 , n83395 );
not ( n83397 , n405282 );
buf ( n405284 , n387542 );
not ( n83399 , n405284 );
buf ( n405286 , n83226 );
not ( n83401 , n405286 );
or ( n83402 , n83399 , n83401 );
buf ( n83403 , n404965 );
buf ( n405290 , n368602 );
nand ( n83405 , n83403 , n405290 );
buf ( n405292 , n83405 );
buf ( n405293 , n405292 );
nand ( n83408 , n83402 , n405293 );
buf ( n405295 , n83408 );
not ( n405296 , n405295 );
or ( n405297 , n83397 , n405296 );
or ( n405298 , n405282 , n405295 );
buf ( n405299 , n45012 );
not ( n405300 , n405299 );
buf ( n405301 , n368994 );
not ( n405302 , n405301 );
buf ( n405303 , n342908 );
not ( n405304 , n405303 );
or ( n405305 , n405302 , n405304 );
buf ( n405306 , n81867 );
buf ( n405307 , n57053 );
nand ( n405308 , n405306 , n405307 );
buf ( n405309 , n405308 );
buf ( n405310 , n405309 );
nand ( n405311 , n405305 , n405310 );
buf ( n405312 , n405311 );
buf ( n405313 , n405312 );
not ( n405314 , n405313 );
or ( n405315 , n405300 , n405314 );
buf ( n405316 , n403511 );
buf ( n405317 , n365149 );
nand ( n405318 , n405316 , n405317 );
buf ( n405319 , n405318 );
buf ( n405320 , n405319 );
nand ( n83414 , n405315 , n405320 );
buf ( n405322 , n83414 );
not ( n405323 , n405322 );
buf ( n405324 , n56970 );
not ( n405325 , n405324 );
buf ( n405326 , n400916 );
not ( n83420 , n405326 );
or ( n405328 , n405325 , n83420 );
buf ( n405329 , n396441 );
buf ( n405330 , n377389 );
nand ( n405331 , n405329 , n405330 );
buf ( n405332 , n405331 );
buf ( n405333 , n405332 );
nand ( n405334 , n405328 , n405333 );
buf ( n405335 , n405334 );
not ( n83429 , n405335 );
not ( n83430 , n45055 );
or ( n83431 , n83429 , n83430 );
nand ( n405339 , n83183 , n365242 );
nand ( n405340 , n83431 , n405339 );
not ( n83434 , n405340 );
or ( n405342 , n405323 , n83434 );
or ( n405343 , n405340 , n405322 );
xor ( n83437 , n402157 , n402160 );
xor ( n405345 , n83437 , n402164 );
xor ( n405346 , n403743 , n404083 );
xor ( n83440 , n405345 , n405346 );
buf ( n405348 , n83440 );
buf ( n405349 , n44915 );
not ( n405350 , n405349 );
buf ( n405351 , n404113 );
not ( n405352 , n405351 );
or ( n405353 , n405350 , n405352 );
buf ( n405354 , n404115 );
buf ( n405355 , n365136 );
not ( n405356 , n405355 );
buf ( n405357 , n405356 );
and ( n83451 , n405357 , n48458 );
not ( n83452 , n405357 );
and ( n405360 , n83452 , n368656 );
or ( n405361 , n83451 , n405360 );
buf ( n405362 , n405361 );
nand ( n405363 , n405354 , n405362 );
buf ( n405364 , n405363 );
buf ( n405365 , n405364 );
nand ( n83459 , n405353 , n405365 );
buf ( n405367 , n83459 );
buf ( n405368 , n405367 );
xor ( n405369 , n405348 , n405368 );
buf ( n405370 , n49172 );
buf ( n405371 , n405370 );
not ( n405372 , n405371 );
buf ( n405373 , n75283 );
not ( n405374 , n405373 );
or ( n83468 , n405372 , n405374 );
buf ( n405376 , n81867 );
buf ( n405377 , n405370 );
not ( n405378 , n405377 );
buf ( n405379 , n405378 );
buf ( n405380 , n405379 );
nand ( n405381 , n405376 , n405380 );
buf ( n405382 , n405381 );
buf ( n405383 , n405382 );
nand ( n405384 , n83468 , n405383 );
buf ( n405385 , n405384 );
buf ( n405386 , n405385 );
not ( n83480 , n405386 );
buf ( n405388 , n45012 );
not ( n405389 , n405388 );
or ( n405390 , n83480 , n405389 );
buf ( n405391 , n405312 );
buf ( n405392 , n365149 );
nand ( n405393 , n405391 , n405392 );
buf ( n405394 , n405393 );
buf ( n405395 , n405394 );
nand ( n405396 , n405390 , n405395 );
buf ( n405397 , n405396 );
buf ( n405398 , n405397 );
and ( n405399 , n405369 , n405398 );
and ( n405400 , n405348 , n405368 );
or ( n405401 , n405399 , n405400 );
buf ( n405402 , n405401 );
nand ( n405403 , n405343 , n405402 );
nand ( n405404 , n405342 , n405403 );
nand ( n405405 , n405298 , n405404 );
nand ( n405406 , n405297 , n405405 );
buf ( n405407 , n405406 );
nand ( n405408 , n405279 , n405407 );
buf ( n405409 , n405408 );
buf ( n405410 , n405409 );
buf ( n405411 , n405273 );
buf ( n405412 , n405256 );
nand ( n405413 , n405411 , n405412 );
buf ( n405414 , n405413 );
buf ( n405415 , n405414 );
nand ( n405416 , n405410 , n405415 );
buf ( n405417 , n405416 );
buf ( n405418 , n405417 );
and ( n405419 , n405232 , n405418 );
buf ( n405420 , n405204 );
not ( n405421 , n405420 );
buf ( n405422 , n405228 );
nor ( n405423 , n405421 , n405422 );
buf ( n83486 , n405423 );
buf ( n405425 , n83486 );
nor ( n83488 , n405419 , n405425 );
buf ( n405427 , n83488 );
buf ( n405428 , n405427 );
and ( n405429 , n83336 , n405428 );
and ( n83492 , n83328 , n405191 );
or ( n405431 , n405429 , n83492 );
buf ( n405432 , n405431 );
buf ( n405433 , n405432 );
buf ( n405434 , n403094 );
buf ( n405435 , n403221 );
xor ( n405436 , n405434 , n405435 );
buf ( n405437 , n403119 );
xnor ( n405438 , n405436 , n405437 );
buf ( n405439 , n405438 );
buf ( n405440 , n405439 );
xor ( n83503 , n405433 , n405440 );
xor ( n405442 , n404201 , n403391 );
xor ( n405443 , n405442 , n403420 );
buf ( n405444 , n405443 );
and ( n405445 , n83503 , n405444 );
and ( n405446 , n405433 , n405440 );
or ( n83509 , n405445 , n405446 );
buf ( n405448 , n83509 );
buf ( n405449 , n405448 );
nand ( n83512 , n83291 , n405449 );
buf ( n405451 , n83512 );
not ( n405452 , n405451 );
or ( n83515 , n83286 , n405452 );
buf ( n405454 , n405448 );
not ( n405455 , n405454 );
buf ( n405456 , n405145 );
nand ( n83519 , n405455 , n405456 );
buf ( n405458 , n83519 );
nand ( n83521 , n83515 , n405458 );
buf ( n405460 , n83521 );
nand ( n83523 , n404646 , n405460 );
buf ( n405462 , n83523 );
buf ( n405463 , n405462 );
nand ( n405464 , n404643 , n405463 );
buf ( n405465 , n405464 );
buf ( n405466 , n405465 );
buf ( n405467 , n403280 );
buf ( n405468 , n403269 );
and ( n405469 , n405467 , n405468 );
not ( n83532 , n405467 );
buf ( n405471 , n403272 );
and ( n83534 , n83532 , n405471 );
nor ( n83535 , n405469 , n83534 );
buf ( n405474 , n83535 );
buf ( n405475 , n405474 );
buf ( n405476 , n402995 );
and ( n405477 , n405475 , n405476 );
not ( n83540 , n405475 );
buf ( n405479 , n402998 );
and ( n405480 , n83540 , n405479 );
nor ( n405481 , n405477 , n405480 );
buf ( n405482 , n405481 );
buf ( n405483 , n405482 );
not ( n405484 , n405483 );
buf ( n405485 , n405484 );
buf ( n405486 , n405485 );
and ( n405487 , n405466 , n405486 );
not ( n405488 , n405466 );
buf ( n405489 , n405482 );
and ( n405490 , n405488 , n405489 );
nor ( n405491 , n405487 , n405490 );
buf ( n405492 , n405491 );
xnor ( n405493 , n404521 , n405492 );
buf ( n405494 , n404635 );
buf ( n405495 , n404640 );
xor ( n83555 , n405494 , n405495 );
buf ( n405497 , n83521 );
xnor ( n405498 , n83555 , n405497 );
buf ( n405499 , n405498 );
buf ( n405500 , n405499 );
not ( n405501 , n405500 );
buf ( n405502 , n405501 );
not ( n405503 , n405502 );
xor ( n405504 , n404372 , n404384 );
xor ( n83564 , n405504 , n404397 );
buf ( n405506 , n83564 );
not ( n405507 , n405506 );
or ( n405508 , n405503 , n405507 );
buf ( n405509 , n405506 );
not ( n83569 , n405509 );
buf ( n405511 , n83569 );
not ( n405512 , n405511 );
not ( n83572 , n405499 );
or ( n83573 , n405512 , n83572 );
buf ( n405515 , n404247 );
buf ( n83575 , n404350 );
xor ( n83576 , n405515 , n83575 );
buf ( n405518 , n404359 );
xnor ( n405519 , n83576 , n405518 );
buf ( n405520 , n405519 );
buf ( n405521 , n405520 );
xor ( n405522 , n405433 , n405440 );
xor ( n83582 , n405522 , n405444 );
buf ( n405524 , n83582 );
buf ( n405525 , n405524 );
not ( n405526 , n405525 );
buf ( n405527 , n405526 );
buf ( n405528 , n405527 );
not ( n405529 , n405528 );
xor ( n405530 , n82815 , n404618 );
xor ( n83590 , n405530 , n404626 );
buf ( n405532 , n83590 );
buf ( n405533 , n405532 );
not ( n405534 , n405533 );
or ( n405535 , n405529 , n405534 );
buf ( n405536 , n405524 );
not ( n83596 , n405536 );
buf ( n405538 , n405532 );
not ( n405539 , n405538 );
buf ( n405540 , n405539 );
buf ( n405541 , n405540 );
not ( n405542 , n405541 );
or ( n83602 , n83596 , n405542 );
xor ( n405544 , n83328 , n405191 );
xor ( n405545 , n405544 , n405428 );
buf ( n405546 , n405545 );
buf ( n405547 , n405546 );
not ( n405548 , n405547 );
buf ( n405549 , n384667 );
buf ( n405550 , n373764 );
and ( n405551 , n405549 , n405550 );
not ( n83611 , n405549 );
buf ( n405553 , n362549 );
and ( n405554 , n83611 , n405553 );
or ( n405555 , n405551 , n405554 );
buf ( n405556 , n405555 );
not ( n405557 , n405556 );
not ( n83617 , n385064 );
and ( n405559 , n405557 , n83617 );
and ( n405560 , n404607 , n380356 );
nor ( n83620 , n405559 , n405560 );
buf ( n405562 , n83620 );
not ( n405563 , n405562 );
or ( n83623 , n405548 , n405563 );
and ( n405565 , n405181 , n405158 );
not ( n405566 , n405181 );
and ( n83626 , n405566 , n405155 );
or ( n83627 , n405565 , n83626 );
xnor ( n83628 , n83627 , n405151 );
buf ( n405570 , n83628 );
buf ( n405571 , n379916 );
not ( n83631 , n405571 );
buf ( n405573 , n379838 );
not ( n83633 , n405573 );
buf ( n405575 , n31073 );
not ( n405576 , n405575 );
or ( n83636 , n83633 , n405576 );
buf ( n405578 , n351107 );
buf ( n405579 , n398741 );
nand ( n83639 , n405578 , n405579 );
buf ( n405581 , n83639 );
buf ( n405582 , n405581 );
nand ( n83642 , n83636 , n405582 );
buf ( n83643 , n83642 );
buf ( n405585 , n83643 );
not ( n83645 , n405585 );
or ( n405587 , n83631 , n83645 );
buf ( n405588 , n404551 );
buf ( n405589 , n379890 );
nand ( n405590 , n405588 , n405589 );
buf ( n405591 , n405590 );
buf ( n405592 , n405591 );
nand ( n405593 , n405587 , n405592 );
buf ( n405594 , n405593 );
buf ( n405595 , n405594 );
xor ( n405596 , n405570 , n405595 );
buf ( n405597 , n58867 );
not ( n83657 , n405597 );
buf ( n405599 , n379368 );
not ( n83659 , n405599 );
buf ( n405601 , n45152 );
not ( n405602 , n405601 );
or ( n83662 , n83659 , n405602 );
buf ( n405604 , n30912 );
buf ( n405605 , n379392 );
nand ( n83665 , n405604 , n405605 );
buf ( n405607 , n83665 );
buf ( n405608 , n405607 );
nand ( n83668 , n83662 , n405608 );
buf ( n405610 , n83668 );
buf ( n405611 , n405610 );
not ( n405612 , n405611 );
or ( n83672 , n83657 , n405612 );
buf ( n405614 , n404835 );
buf ( n405615 , n58923 );
nand ( n405616 , n405614 , n405615 );
buf ( n405617 , n405616 );
buf ( n405618 , n405617 );
nand ( n405619 , n83672 , n405618 );
buf ( n405620 , n405619 );
buf ( n405621 , n405620 );
and ( n405622 , n405596 , n405621 );
and ( n405623 , n405570 , n405595 );
or ( n405624 , n405622 , n405623 );
buf ( n405625 , n405624 );
buf ( n405626 , n405625 );
nand ( n405627 , n83623 , n405626 );
buf ( n405628 , n405627 );
buf ( n405629 , n405628 );
buf ( n405630 , n83620 );
not ( n405631 , n405630 );
buf ( n405632 , n405631 );
buf ( n405633 , n405632 );
buf ( n405634 , n405546 );
not ( n405635 , n405634 );
buf ( n405636 , n405635 );
buf ( n405637 , n405636 );
nand ( n405638 , n405633 , n405637 );
buf ( n405639 , n405638 );
buf ( n405640 , n405639 );
nand ( n83678 , n405629 , n405640 );
buf ( n405642 , n83678 );
buf ( n405643 , n405642 );
nand ( n83681 , n83602 , n405643 );
buf ( n405645 , n83681 );
buf ( n405646 , n405645 );
nand ( n83684 , n405535 , n405646 );
buf ( n83685 , n83684 );
buf ( n405649 , n83685 );
xor ( n83687 , n405521 , n405649 );
xor ( n83688 , n404525 , n404529 );
xor ( n83689 , n83688 , n404631 );
buf ( n405653 , n83689 );
buf ( n405654 , n405653 );
and ( n83692 , n83687 , n405654 );
and ( n405656 , n405521 , n405649 );
or ( n83694 , n83692 , n405656 );
buf ( n405658 , n83694 );
nand ( n405659 , n83573 , n405658 );
nand ( n405660 , n405508 , n405659 );
or ( n405661 , n405493 , n405660 );
buf ( n405662 , n405661 );
buf ( n405663 , n403350 );
buf ( n405664 , n404406 );
xor ( n405665 , n405663 , n405664 );
buf ( n405666 , n403325 );
xnor ( n405667 , n405665 , n405666 );
buf ( n405668 , n405667 );
buf ( n405669 , n405668 );
buf ( n405670 , n404521 );
not ( n83706 , n405670 );
buf ( n405672 , n83706 );
not ( n83708 , n405672 );
not ( n83709 , n405485 );
and ( n405675 , n83708 , n83709 );
buf ( n405676 , n405482 );
not ( n405677 , n405676 );
buf ( n405678 , n405672 );
nand ( n405679 , n405677 , n405678 );
buf ( n405680 , n405679 );
and ( n405681 , n405680 , n405465 );
nor ( n405682 , n405675 , n405681 );
buf ( n405683 , n405682 );
nand ( n405684 , n405669 , n405683 );
buf ( n405685 , n405684 );
buf ( n405686 , n405685 );
and ( n405687 , n405662 , n405686 );
buf ( n405688 , n405687 );
buf ( n405689 , n405688 );
not ( n405690 , n405689 );
buf ( n405691 , n379890 );
not ( n83727 , n405691 );
and ( n405693 , n370652 , n379838 );
not ( n405694 , n370652 );
and ( n405695 , n405694 , n398741 );
or ( n83731 , n405693 , n405695 );
buf ( n405697 , n83731 );
not ( n405698 , n405697 );
or ( n83732 , n83727 , n405698 );
buf ( n405700 , n379838 );
not ( n405701 , n405700 );
buf ( n405702 , n372382 );
not ( n405703 , n405702 );
or ( n405704 , n405701 , n405703 );
buf ( n405705 , n391133 );
buf ( n405706 , n398741 );
nand ( n405707 , n405705 , n405706 );
buf ( n405708 , n405707 );
buf ( n405709 , n405708 );
nand ( n405710 , n405704 , n405709 );
buf ( n405711 , n405710 );
buf ( n405712 , n405711 );
buf ( n405713 , n379916 );
nand ( n405714 , n405712 , n405713 );
buf ( n405715 , n405714 );
buf ( n405716 , n405715 );
nand ( n405717 , n83732 , n405716 );
buf ( n405718 , n405717 );
buf ( n405719 , n405718 );
xor ( n405720 , n403895 , n403912 );
xor ( n405721 , n405720 , n403917 );
buf ( n405722 , n405721 );
buf ( n405723 , n384380 );
buf ( n405724 , n384343 );
and ( n405725 , n405723 , n405724 );
buf ( n405726 , n384386 );
buf ( n405727 , n384089 );
and ( n405728 , n405726 , n405727 );
nor ( n405729 , n405725 , n405728 );
buf ( n405730 , n405729 );
buf ( n405731 , n405730 );
buf ( n405732 , n384354 );
or ( n83744 , n405731 , n405732 );
buf ( n405734 , n403718 );
buf ( n405735 , n384082 );
or ( n405736 , n405734 , n405735 );
nand ( n405737 , n83744 , n405736 );
buf ( n405738 , n405737 );
xor ( n405739 , n403857 , n403874 );
xor ( n405740 , n405739 , n403891 );
and ( n405741 , n405738 , n405740 );
buf ( n405742 , n61992 );
buf ( n405743 , n394840 );
and ( n405744 , n405742 , n405743 );
buf ( n405745 , n382596 );
buf ( n405746 , n395890 );
and ( n405747 , n405745 , n405746 );
nor ( n405748 , n405744 , n405747 );
buf ( n405749 , n405748 );
buf ( n405750 , n405749 );
buf ( n405751 , n394838 );
or ( n405752 , n405750 , n405751 );
buf ( n405753 , n404048 );
buf ( n405754 , n394835 );
or ( n405755 , n405753 , n405754 );
nand ( n405756 , n405752 , n405755 );
buf ( n83750 , n405756 );
xor ( n405758 , n403857 , n403874 );
xor ( n405759 , n405758 , n403891 );
and ( n405760 , n83750 , n405759 );
and ( n405761 , n405738 , n83750 );
or ( n83753 , n405741 , n405760 , n405761 );
xor ( n405763 , n405722 , n83753 );
xor ( n405764 , n404040 , n404057 );
xor ( n83756 , n405764 , n404063 );
buf ( n405766 , n83756 );
and ( n405767 , n405763 , n405766 );
and ( n83759 , n405722 , n83753 );
or ( n405769 , n405767 , n83759 );
xor ( n405770 , n404067 , n404070 );
xor ( n405771 , n405770 , n82412 );
and ( n405772 , n405769 , n405771 );
xor ( n405773 , n82146 , n403824 );
buf ( n405774 , n405773 );
buf ( n405775 , n405774 );
buf ( n405776 , n378341 );
buf ( n405777 , n81950 );
buf ( n405778 , n57800 );
and ( n83766 , n405777 , n405778 );
buf ( n405780 , n403589 );
buf ( n405781 , n378284 );
and ( n405782 , n405780 , n405781 );
nor ( n83770 , n83766 , n405782 );
buf ( n83771 , n83770 );
buf ( n405785 , n83771 );
or ( n83773 , n405776 , n405785 );
buf ( n405787 , n82332 );
buf ( n405788 , n378262 );
or ( n405789 , n405787 , n405788 );
nand ( n405790 , n83773 , n405789 );
buf ( n405791 , n405790 );
buf ( n405792 , n405791 );
xor ( n405793 , n405775 , n405792 );
buf ( n405794 , n376924 );
buf ( n405795 , n376866 );
buf ( n405796 , n403795 );
and ( n405797 , n405795 , n405796 );
buf ( n405798 , n377030 );
buf ( n405799 , n403798 );
and ( n83787 , n405798 , n405799 );
nor ( n405801 , n405797 , n83787 );
buf ( n405802 , n405801 );
buf ( n405803 , n405802 );
or ( n405804 , n405794 , n405803 );
buf ( n405805 , n403816 );
buf ( n405806 , n56517 );
or ( n405807 , n405805 , n405806 );
nand ( n405808 , n405804 , n405807 );
buf ( n405809 , n405808 );
buf ( n405810 , n405809 );
buf ( n405811 , n376997 );
xor ( n405812 , n376618 , n56216 );
xnor ( n405813 , n405812 , n56225 );
buf ( n405814 , n405813 );
not ( n405815 , n405814 );
buf ( n405816 , n405815 );
buf ( n405817 , n405816 );
and ( n405818 , n405811 , n405817 );
buf ( n405819 , n376990 );
buf ( n405820 , n405813 );
and ( n405821 , n405819 , n405820 );
buf ( n405822 , n377003 );
nor ( n83794 , n405818 , n405821 , n405822 );
buf ( n405824 , n83794 );
buf ( n405825 , n405824 );
xor ( n405826 , n405810 , n405825 );
buf ( n405827 , n378291 );
not ( n83799 , n405827 );
buf ( n405829 , n83771 );
not ( n405830 , n405829 );
buf ( n405831 , n405830 );
buf ( n405832 , n405831 );
not ( n405833 , n405832 );
or ( n405834 , n83799 , n405833 );
buf ( n405835 , n378341 );
buf ( n405836 , n57800 );
buf ( n405837 , n81995 );
and ( n405838 , n405836 , n405837 );
buf ( n405839 , n403645 );
buf ( n405840 , n378284 );
and ( n405841 , n405839 , n405840 );
nor ( n83808 , n405838 , n405841 );
buf ( n405843 , n83808 );
buf ( n405844 , n405843 );
or ( n83810 , n405835 , n405844 );
nand ( n83811 , n405834 , n83810 );
buf ( n405847 , n83811 );
buf ( n405848 , n405847 );
and ( n405849 , n405826 , n405848 );
and ( n83813 , n405810 , n405825 );
or ( n405851 , n405849 , n83813 );
buf ( n405852 , n405851 );
buf ( n405853 , n405852 );
and ( n83816 , n405793 , n405853 );
and ( n83817 , n405775 , n405792 );
or ( n83818 , n83816 , n83817 );
buf ( n405857 , n83818 );
buf ( n405858 , n405857 );
buf ( n405859 , n396615 );
buf ( n405860 , n380817 );
and ( n405861 , n405859 , n405860 );
buf ( n405862 , n396621 );
buf ( n405863 , n82201 );
and ( n405864 , n405862 , n405863 );
nor ( n405865 , n405861 , n405864 );
buf ( n405866 , n405865 );
buf ( n405867 , n405866 );
buf ( n405868 , n60313 );
or ( n405869 , n405867 , n405868 );
buf ( n405870 , n82280 );
buf ( n405871 , n380733 );
or ( n405872 , n405870 , n405871 );
nand ( n405873 , n405869 , n405872 );
buf ( n405874 , n405873 );
buf ( n405875 , n405874 );
xor ( n405876 , n405858 , n405875 );
buf ( n405877 , n382655 );
not ( n405878 , n405877 );
buf ( n405879 , n395810 );
buf ( n405880 , n382835 );
and ( n405881 , n405879 , n405880 );
buf ( n405882 , n395816 );
buf ( n405883 , n62243 );
and ( n83827 , n405882 , n405883 );
nor ( n83828 , n405881 , n83827 );
buf ( n405886 , n83828 );
buf ( n405887 , n405886 );
not ( n83831 , n405887 );
buf ( n405889 , n83831 );
buf ( n405890 , n405889 );
not ( n83834 , n405890 );
or ( n83835 , n405878 , n83834 );
buf ( n405893 , n74644 );
buf ( n405894 , n382835 );
and ( n405895 , n405893 , n405894 );
buf ( n405896 , n395683 );
buf ( n405897 , n62243 );
and ( n83840 , n405896 , n405897 );
nor ( n405899 , n405895 , n83840 );
buf ( n405900 , n405899 );
buf ( n405901 , n405900 );
buf ( n405902 , n384157 );
or ( n83845 , n405901 , n405902 );
nand ( n83846 , n83835 , n83845 );
buf ( n405905 , n83846 );
buf ( n405906 , n405905 );
and ( n83849 , n405876 , n405906 );
and ( n83850 , n405858 , n405875 );
or ( n83851 , n83849 , n83850 );
buf ( n405910 , n83851 );
buf ( n405911 , n405910 );
buf ( n405912 , n73625 );
buf ( n405913 , n384343 );
and ( n405914 , n405912 , n405913 );
buf ( n405915 , n73631 );
buf ( n405916 , n384089 );
and ( n405917 , n405915 , n405916 );
nor ( n405918 , n405914 , n405917 );
buf ( n405919 , n405918 );
buf ( n405920 , n405919 );
buf ( n405921 , n384354 );
or ( n405922 , n405920 , n405921 );
buf ( n405923 , n405730 );
buf ( n405924 , n384082 );
or ( n405925 , n405923 , n405924 );
nand ( n405926 , n405922 , n405925 );
buf ( n405927 , n405926 );
buf ( n405928 , n405927 );
xor ( n405929 , n405911 , n405928 );
xor ( n405930 , n403950 , n403967 );
xor ( n405931 , n405930 , n404012 );
buf ( n405932 , n405931 );
buf ( n405933 , n405932 );
and ( n405934 , n405929 , n405933 );
and ( n83858 , n405911 , n405928 );
or ( n83859 , n405934 , n83858 );
buf ( n405937 , n83859 );
buf ( n405938 , n405937 );
buf ( n405939 , n405900 );
buf ( n405940 , n382849 );
or ( n405941 , n405939 , n405940 );
buf ( n405942 , n403883 );
buf ( n405943 , n384157 );
or ( n405944 , n405942 , n405943 );
nand ( n405945 , n405941 , n405944 );
buf ( n405946 , n405945 );
buf ( n405947 , n405946 );
xor ( n405948 , n403832 , n403849 );
xor ( n83872 , n405948 , n403853 );
buf ( n405950 , n83872 );
buf ( n405951 , n405950 );
xor ( n405952 , n405947 , n405951 );
buf ( n405953 , n63549 );
buf ( n405954 , n394724 );
and ( n405955 , n405953 , n405954 );
buf ( n405956 , n384199 );
buf ( n405957 , n394730 );
and ( n405958 , n405956 , n405957 );
nor ( n405959 , n405955 , n405958 );
buf ( n405960 , n405959 );
buf ( n405961 , n405960 );
buf ( n405962 , n384414 );
or ( n405963 , n405961 , n405962 );
buf ( n405964 , n82365 );
buf ( n405965 , n395635 );
or ( n405966 , n405964 , n405965 );
nand ( n405967 , n405963 , n405966 );
buf ( n405968 , n405967 );
buf ( n405969 , n405968 );
and ( n405970 , n405952 , n405969 );
and ( n405971 , n405947 , n405951 );
or ( n405972 , n405970 , n405971 );
buf ( n405973 , n405972 );
buf ( n405974 , n405973 );
xor ( n405975 , n405938 , n405974 );
xor ( n405976 , n403933 , n404017 );
xor ( n405977 , n405976 , n404035 );
buf ( n405978 , n405977 );
buf ( n405979 , n405978 );
and ( n83892 , n405975 , n405979 );
and ( n405981 , n405938 , n405974 );
or ( n405982 , n83892 , n405981 );
buf ( n405983 , n405982 );
xor ( n405984 , n405722 , n83753 );
xor ( n405985 , n405984 , n405766 );
and ( n83896 , n405983 , n405985 );
buf ( n405987 , n79114 );
buf ( n405988 , n380817 );
and ( n83899 , n405987 , n405988 );
buf ( n83900 , n400487 );
buf ( n83901 , n82201 );
and ( n83902 , n83900 , n83901 );
nor ( n83903 , n83899 , n83902 );
buf ( n83904 , n83903 );
buf ( n405995 , n83904 );
buf ( n405996 , n60313 );
or ( n83907 , n405995 , n405996 );
buf ( n405998 , n405866 );
buf ( n405999 , n380733 );
or ( n406000 , n405998 , n405999 );
nand ( n83908 , n83907 , n406000 );
buf ( n83909 , n83908 );
buf ( n406003 , n79312 );
buf ( n406004 , n57789 );
and ( n406005 , n406003 , n406004 );
buf ( n406006 , n79318 );
buf ( n406007 , n60054 );
and ( n406008 , n406006 , n406007 );
nor ( n406009 , n406005 , n406008 );
buf ( n406010 , n406009 );
buf ( n406011 , n406010 );
buf ( n406012 , n380581 );
or ( n406013 , n406011 , n406012 );
buf ( n406014 , n403976 );
buf ( n406015 , n394774 );
or ( n406016 , n406014 , n406015 );
nand ( n406017 , n406013 , n406016 );
buf ( n406018 , n406017 );
xor ( n406019 , n83909 , n406018 );
xor ( n406020 , n405775 , n405792 );
xor ( n406021 , n406020 , n405853 );
buf ( n406022 , n406021 );
and ( n83913 , n406019 , n406022 );
and ( n83914 , n83909 , n406018 );
or ( n406025 , n83913 , n83914 );
xor ( n406026 , n403985 , n404002 );
xor ( n83917 , n406026 , n82346 );
buf ( n406028 , n83917 );
xor ( n83919 , n406025 , n406028 );
buf ( n406030 , n73780 );
buf ( n406031 , n384343 );
and ( n83922 , n406030 , n406031 );
buf ( n406033 , n394816 );
buf ( n406034 , n384089 );
and ( n406035 , n406033 , n406034 );
nor ( n406036 , n83922 , n406035 );
buf ( n406037 , n406036 );
buf ( n406038 , n406037 );
buf ( n406039 , n384354 );
or ( n406040 , n406038 , n406039 );
buf ( n406041 , n405919 );
buf ( n406042 , n384082 );
or ( n83932 , n406041 , n406042 );
nand ( n83933 , n406040 , n83932 );
buf ( n406045 , n83933 );
and ( n406046 , n83919 , n406045 );
and ( n83936 , n406025 , n406028 );
or ( n406048 , n406046 , n83936 );
buf ( n406049 , n406048 );
buf ( n406050 , n62202 );
buf ( n406051 , n394840 );
and ( n406052 , n406050 , n406051 );
buf ( n406053 , n382803 );
buf ( n406054 , n395890 );
and ( n83940 , n406053 , n406054 );
nor ( n83941 , n406052 , n83940 );
buf ( n83942 , n83941 );
buf ( n406058 , n83942 );
buf ( n406059 , n394838 );
or ( n406060 , n406058 , n406059 );
buf ( n406061 , n405749 );
buf ( n406062 , n394835 );
or ( n83948 , n406061 , n406062 );
nand ( n406064 , n406060 , n83948 );
buf ( n406065 , n406064 );
buf ( n406066 , n406065 );
xor ( n406067 , n406049 , n406066 );
xor ( n406068 , n405947 , n405951 );
xor ( n83954 , n406068 , n405969 );
buf ( n406070 , n83954 );
buf ( n83956 , n406070 );
and ( n83957 , n406067 , n83956 );
and ( n406073 , n406049 , n406066 );
or ( n83958 , n83957 , n406073 );
buf ( n83959 , n83958 );
xor ( n406076 , n403857 , n403874 );
xor ( n406077 , n406076 , n403891 );
xor ( n406078 , n405738 , n83750 );
xor ( n406079 , n406077 , n406078 );
xor ( n406080 , n83959 , n406079 );
xor ( n406081 , n405938 , n405974 );
xor ( n406082 , n406081 , n405979 );
buf ( n406083 , n406082 );
and ( n406084 , n406080 , n406083 );
and ( n406085 , n83959 , n406079 );
or ( n406086 , n406084 , n406085 );
xor ( n406087 , n405722 , n83753 );
xor ( n406088 , n406087 , n405766 );
and ( n406089 , n406086 , n406088 );
and ( n406090 , n405983 , n406086 );
or ( n406091 , n83896 , n406089 , n406090 );
xor ( n406092 , n404067 , n404070 );
xor ( n406093 , n406092 , n82412 );
and ( n406094 , n406091 , n406093 );
and ( n406095 , n405769 , n406091 );
or ( n406096 , n405772 , n406094 , n406095 );
buf ( n406097 , n406096 );
xor ( n406098 , n403533 , n403736 );
xor ( n406099 , n406098 , n403740 );
xor ( n406100 , n82265 , n404078 );
xor ( n406101 , n406099 , n406100 );
buf ( n406102 , n406101 );
xor ( n406103 , n406097 , n406102 );
buf ( n406104 , n48792 );
not ( n406105 , n406104 );
buf ( n406106 , n369183 );
not ( n406107 , n406106 );
or ( n406108 , n406105 , n406107 );
buf ( n406109 , n405357 );
buf ( n406110 , n48791 );
nand ( n406111 , n406109 , n406110 );
buf ( n406112 , n406111 );
buf ( n406113 , n406112 );
nand ( n406114 , n406108 , n406113 );
buf ( n406115 , n406114 );
buf ( n406116 , n406115 );
not ( n406117 , n406116 );
buf ( n406118 , n404115 );
not ( n83965 , n406118 );
or ( n83966 , n406117 , n83965 );
buf ( n406121 , n405361 );
buf ( n406122 , n44915 );
nand ( n406123 , n406121 , n406122 );
buf ( n406124 , n406123 );
buf ( n406125 , n406124 );
nand ( n83972 , n83966 , n406125 );
buf ( n406127 , n83972 );
buf ( n406128 , n406127 );
and ( n406129 , n406103 , n406128 );
and ( n406130 , n406097 , n406102 );
or ( n406131 , n406129 , n406130 );
buf ( n406132 , n406131 );
buf ( n406133 , n406132 );
buf ( n406134 , n368621 );
not ( n406135 , n406134 );
buf ( n406136 , n404980 );
not ( n406137 , n406136 );
or ( n406138 , n406135 , n406137 );
buf ( n406139 , n380424 );
buf ( n406140 , n394044 );
not ( n406141 , n406140 );
xor ( n406142 , n406139 , n406141 );
buf ( n406143 , n406142 );
buf ( n406144 , n406143 );
not ( n406145 , n406144 );
buf ( n406146 , n368602 );
nand ( n406147 , n406145 , n406146 );
buf ( n406148 , n406147 );
buf ( n406149 , n406148 );
nand ( n406150 , n406138 , n406149 );
buf ( n406151 , n406150 );
buf ( n406152 , n406151 );
xor ( n406153 , n406133 , n406152 );
buf ( n406154 , n377353 );
buf ( n406155 , n396441 );
and ( n406156 , n406154 , n406155 );
not ( n406157 , n406154 );
buf ( n406158 , n81360 );
and ( n406159 , n406157 , n406158 );
nor ( n406160 , n406156 , n406159 );
buf ( n406161 , n406160 );
buf ( n406162 , n406161 );
not ( n406163 , n406162 );
buf ( n406164 , n45055 );
not ( n406165 , n406164 );
or ( n406166 , n406163 , n406165 );
buf ( n406167 , n405335 );
buf ( n406168 , n365242 );
nand ( n406169 , n406167 , n406168 );
buf ( n406170 , n406169 );
buf ( n406171 , n406170 );
nand ( n406172 , n406166 , n406171 );
buf ( n406173 , n406172 );
buf ( n406174 , n406173 );
and ( n406175 , n406153 , n406174 );
and ( n406176 , n406133 , n406152 );
or ( n406177 , n406175 , n406176 );
buf ( n406178 , n406177 );
buf ( n406179 , n406178 );
buf ( n406180 , n377143 );
not ( n406181 , n406180 );
buf ( n406182 , n380923 );
not ( n406183 , n406182 );
or ( n406184 , n406181 , n406183 );
buf ( n406185 , n22619 );
buf ( n406186 , n377153 );
nand ( n406187 , n406185 , n406186 );
buf ( n406188 , n406187 );
buf ( n406189 , n406188 );
nand ( n406190 , n406184 , n406189 );
buf ( n406191 , n406190 );
buf ( n406192 , n406191 );
not ( n406193 , n406192 );
buf ( n406194 , n384501 );
not ( n406195 , n406194 );
or ( n406196 , n406193 , n406195 );
buf ( n406197 , n404863 );
buf ( n406198 , n56794 );
nand ( n406199 , n406197 , n406198 );
buf ( n406200 , n406199 );
buf ( n406201 , n406200 );
nand ( n406202 , n406196 , n406201 );
buf ( n406203 , n406202 );
buf ( n406204 , n406203 );
xor ( n406205 , n406179 , n406204 );
buf ( n406206 , n369809 );
not ( n406207 , n406206 );
buf ( n406208 , n404909 );
not ( n83992 , n406208 );
or ( n406210 , n406207 , n83992 );
buf ( n406211 , n393883 );
not ( n406212 , n406211 );
buf ( n406213 , n394004 );
not ( n406214 , n406213 );
or ( n406215 , n406212 , n406214 );
buf ( n406216 , n351160 );
buf ( n406217 , n369763 );
nand ( n406218 , n406216 , n406217 );
buf ( n406219 , n406218 );
buf ( n406220 , n406219 );
nand ( n406221 , n406215 , n406220 );
buf ( n406222 , n406221 );
buf ( n406223 , n406222 );
buf ( n406224 , n369804 );
nand ( n406225 , n406223 , n406224 );
buf ( n406226 , n406225 );
buf ( n406227 , n406226 );
nand ( n406228 , n406210 , n406227 );
buf ( n406229 , n406228 );
buf ( n406230 , n406229 );
xor ( n406231 , n406205 , n406230 );
buf ( n406232 , n406231 );
buf ( n406233 , n406232 );
xor ( n406234 , n404067 , n404070 );
xor ( n406235 , n406234 , n82412 );
xor ( n406236 , n405769 , n406091 );
xor ( n406237 , n406235 , n406236 );
buf ( n406238 , n406237 );
buf ( n406239 , n405370 );
not ( n406240 , n406239 );
buf ( n406241 , n369183 );
not ( n406242 , n406241 );
or ( n406243 , n406240 , n406242 );
buf ( n406244 , n342965 );
not ( n406245 , n406244 );
buf ( n406246 , n406245 );
buf ( n406247 , n406246 );
not ( n406248 , n406247 );
buf ( n406249 , n406248 );
buf ( n406250 , n406249 );
buf ( n406251 , n405379 );
nand ( n406252 , n406250 , n406251 );
buf ( n406253 , n406252 );
buf ( n406254 , n406253 );
nand ( n84018 , n406243 , n406254 );
buf ( n406256 , n84018 );
buf ( n406257 , n406256 );
not ( n406258 , n406257 );
not ( n84022 , n44912 );
buf ( n406260 , n84022 );
buf ( n406261 , n406260 );
not ( n84025 , n406261 );
or ( n406263 , n406258 , n84025 );
buf ( n406264 , n406115 );
buf ( n406265 , n44915 );
nand ( n406266 , n406264 , n406265 );
buf ( n406267 , n406266 );
buf ( n406268 , n406267 );
nand ( n406269 , n406263 , n406268 );
buf ( n406270 , n406269 );
buf ( n84034 , n406270 );
xor ( n84035 , n406238 , n84034 );
not ( n406273 , n369444 );
not ( n84037 , n368549 );
not ( n84038 , n365384 );
or ( n406276 , n84037 , n84038 );
buf ( n406277 , n351062 );
buf ( n84041 , n406277 );
buf ( n84042 , n84041 );
buf ( n406280 , n84042 );
buf ( n406281 , n380424 );
nand ( n406282 , n406280 , n406281 );
buf ( n406283 , n406282 );
nand ( n84047 , n406276 , n406283 );
not ( n406285 , n84047 );
or ( n406286 , n406273 , n406285 );
buf ( n406287 , n368549 );
not ( n406288 , n406287 );
buf ( n406289 , n48458 );
not ( n84053 , n406289 );
or ( n406291 , n406288 , n84053 );
buf ( n406292 , n368656 );
buf ( n406293 , n380424 );
nand ( n406294 , n406292 , n406293 );
buf ( n406295 , n406294 );
buf ( n406296 , n406295 );
nand ( n406297 , n406291 , n406296 );
buf ( n406298 , n406297 );
nand ( n406299 , n406298 , n368602 );
nand ( n406300 , n406286 , n406299 );
buf ( n406301 , n406300 );
and ( n406302 , n84035 , n406301 );
and ( n406303 , n406238 , n84034 );
or ( n406304 , n406302 , n406303 );
buf ( n406305 , n406304 );
buf ( n406306 , n406305 );
buf ( n406307 , n369809 );
not ( n406308 , n406307 );
buf ( n406309 , n393883 );
not ( n406310 , n406309 );
buf ( n406311 , n364900 );
not ( n406312 , n406311 );
or ( n406313 , n406310 , n406312 );
buf ( n406314 , n63345 );
buf ( n406315 , n369763 );
nand ( n406316 , n406314 , n406315 );
buf ( n406317 , n406316 );
buf ( n406318 , n406317 );
nand ( n406319 , n406313 , n406318 );
buf ( n406320 , n406319 );
buf ( n406321 , n406320 );
not ( n406322 , n406321 );
or ( n406323 , n406308 , n406322 );
buf ( n406324 , n393883 );
not ( n84071 , n406324 );
buf ( n406326 , n74977 );
not ( n84073 , n406326 );
or ( n406328 , n84071 , n84073 );
nand ( n84075 , n369763 , n45802 );
buf ( n406330 , n84075 );
nand ( n406331 , n406328 , n406330 );
buf ( n406332 , n406331 );
buf ( n406333 , n406332 );
buf ( n406334 , n369804 );
nand ( n406335 , n406333 , n406334 );
buf ( n406336 , n406335 );
buf ( n406337 , n406336 );
nand ( n84084 , n406323 , n406337 );
buf ( n406339 , n84084 );
buf ( n406340 , n406339 );
xor ( n84087 , n406306 , n406340 );
buf ( n406342 , n394065 );
not ( n406343 , n406342 );
buf ( n84090 , n377779 );
not ( n406345 , n84090 );
buf ( n406346 , n406345 );
buf ( n406347 , n406346 );
not ( n406348 , n406347 );
or ( n84095 , n406343 , n406348 );
buf ( n406350 , n394066 );
buf ( n406351 , n377779 );
nand ( n406352 , n406350 , n406351 );
buf ( n406353 , n406352 );
buf ( n406354 , n406353 );
nand ( n84101 , n84095 , n406354 );
buf ( n406356 , n84101 );
buf ( n406357 , n406356 );
not ( n406358 , n406357 );
buf ( n406359 , n45055 );
not ( n84106 , n406359 );
or ( n406361 , n406358 , n84106 );
buf ( n406362 , n365242 );
buf ( n406363 , n406161 );
nand ( n406364 , n406362 , n406363 );
buf ( n406365 , n406364 );
buf ( n406366 , n406365 );
nand ( n406367 , n406361 , n406366 );
buf ( n406368 , n406367 );
buf ( n406369 , n406368 );
and ( n84116 , n84087 , n406369 );
and ( n406371 , n406306 , n406340 );
or ( n406372 , n84116 , n406371 );
buf ( n406373 , n406372 );
buf ( n406374 , n406373 );
and ( n84121 , n377122 , n22619 );
not ( n406376 , n377122 );
and ( n84123 , n406376 , n380923 );
nor ( n406378 , n84121 , n84123 );
buf ( n406379 , n406378 );
not ( n84126 , n406379 );
buf ( n406381 , n384501 );
not ( n406382 , n406381 );
or ( n406383 , n84126 , n406382 );
buf ( n406384 , n406191 );
buf ( n406385 , n56794 );
nand ( n406386 , n406384 , n406385 );
buf ( n84129 , n406386 );
buf ( n406388 , n84129 );
nand ( n84131 , n406383 , n406388 );
buf ( n84132 , n84131 );
buf ( n84133 , n84132 );
xor ( n84134 , n406374 , n84133 );
buf ( n406393 , n45012 );
not ( n84136 , n406393 );
and ( n84137 , n377353 , n81867 );
not ( n406396 , n377353 );
and ( n84139 , n406396 , n402191 );
nor ( n406398 , n84137 , n84139 );
buf ( n406399 , n406398 );
not ( n406400 , n406399 );
or ( n84143 , n84136 , n406400 );
buf ( n406402 , n56970 );
not ( n406403 , n406402 );
buf ( n406404 , n81871 );
not ( n406405 , n406404 );
or ( n84148 , n406403 , n406405 );
buf ( n406407 , n81867 );
buf ( n406408 , n377389 );
nand ( n406409 , n406407 , n406408 );
buf ( n406410 , n406409 );
buf ( n406411 , n406410 );
nand ( n406412 , n84148 , n406411 );
buf ( n406413 , n406412 );
buf ( n406414 , n406413 );
buf ( n406415 , n365149 );
nand ( n406416 , n406414 , n406415 );
buf ( n406417 , n406416 );
buf ( n406418 , n406417 );
nand ( n406419 , n84143 , n406418 );
buf ( n406420 , n406419 );
buf ( n406421 , n406420 );
xor ( n406422 , n405911 , n405928 );
xor ( n406423 , n406422 , n405933 );
buf ( n406424 , n406423 );
buf ( n406425 , n384380 );
buf ( n406426 , n394724 );
and ( n406427 , n406425 , n406426 );
buf ( n406428 , n384386 );
buf ( n406429 , n394730 );
and ( n84154 , n406428 , n406429 );
nor ( n406431 , n406427 , n84154 );
buf ( n406432 , n406431 );
buf ( n406433 , n406432 );
buf ( n406434 , n384414 );
or ( n84159 , n406433 , n406434 );
buf ( n406436 , n405960 );
buf ( n406437 , n395635 );
or ( n84162 , n406436 , n406437 );
nand ( n406439 , n84159 , n84162 );
buf ( n406440 , n406439 );
xor ( n84165 , n405858 , n405875 );
xor ( n84166 , n84165 , n405906 );
buf ( n406443 , n84166 );
xor ( n406444 , n406440 , n406443 );
buf ( n406445 , n63406 );
buf ( n406446 , n394840 );
and ( n406447 , n406445 , n406446 );
buf ( n406448 , n384054 );
buf ( n406449 , n395890 );
and ( n84174 , n406448 , n406449 );
nor ( n406451 , n406447 , n84174 );
buf ( n406452 , n406451 );
buf ( n406453 , n406452 );
buf ( n406454 , n394838 );
or ( n406455 , n406453 , n406454 );
buf ( n406456 , n83942 );
buf ( n406457 , n394835 );
or ( n406458 , n406456 , n406457 );
nand ( n84182 , n406455 , n406458 );
buf ( n84183 , n84182 );
and ( n406461 , n406444 , n84183 );
and ( n84185 , n406440 , n406443 );
or ( n406463 , n406461 , n84185 );
xor ( n406464 , n406424 , n406463 );
buf ( n406465 , n75451 );
buf ( n406466 , n382835 );
and ( n406467 , n406465 , n406466 );
buf ( n406468 , n396596 );
buf ( n406469 , n62243 );
and ( n84193 , n406468 , n406469 );
nor ( n84194 , n406467 , n84193 );
buf ( n406472 , n84194 );
buf ( n406473 , n406472 );
buf ( n406474 , n382849 );
or ( n84198 , n406473 , n406474 );
buf ( n406476 , n405886 );
buf ( n406477 , n384157 );
or ( n84201 , n406476 , n406477 );
nand ( n406479 , n84198 , n84201 );
buf ( n406480 , n406479 );
buf ( n406481 , n406480 );
buf ( n406482 , n80468 );
buf ( n406483 , n57789 );
and ( n406484 , n406482 , n406483 );
buf ( n406485 , n401921 );
buf ( n406486 , n378470 );
and ( n84210 , n406485 , n406486 );
nor ( n84211 , n406484 , n84210 );
buf ( n406489 , n84211 );
buf ( n406490 , n406489 );
buf ( n406491 , n380581 );
or ( n406492 , n406490 , n406491 );
buf ( n84216 , n406010 );
buf ( n406494 , n378476 );
or ( n406495 , n84216 , n406494 );
nand ( n406496 , n406492 , n406495 );
buf ( n406497 , n406496 );
buf ( n406498 , n406497 );
buf ( n406499 , n376924 );
buf ( n406500 , n376866 );
buf ( n406501 , n405813 );
and ( n406502 , n406500 , n406501 );
buf ( n406503 , n377030 );
buf ( n406504 , n405816 );
and ( n84226 , n406503 , n406504 );
nor ( n406506 , n406502 , n84226 );
buf ( n406507 , n406506 );
buf ( n406508 , n406507 );
or ( n84230 , n406499 , n406508 );
buf ( n406510 , n405802 );
buf ( n406511 , n56517 );
or ( n406512 , n406510 , n406511 );
nand ( n406513 , n84230 , n406512 );
buf ( n406514 , n406513 );
buf ( n406515 , n406514 );
buf ( n406516 , n57800 );
buf ( n406517 , n403772 );
and ( n84239 , n406516 , n406517 );
buf ( n406519 , n378284 );
buf ( n406520 , n403775 );
and ( n406521 , n406519 , n406520 );
nor ( n406522 , n84239 , n406521 );
buf ( n406523 , n406522 );
buf ( n406524 , n406523 );
not ( n406525 , n406524 );
buf ( n406526 , n406525 );
buf ( n406527 , n406526 );
not ( n84249 , n406527 );
buf ( n406529 , n378280 );
not ( n406530 , n406529 );
or ( n84252 , n84249 , n406530 );
buf ( n406532 , n378262 );
buf ( n406533 , n405843 );
or ( n84255 , n406532 , n406533 );
nand ( n406535 , n84252 , n84255 );
buf ( n406536 , n406535 );
buf ( n84258 , n406536 );
and ( n84259 , n406515 , n84258 );
buf ( n406539 , n84259 );
buf ( n406540 , n406539 );
xor ( n406541 , n406498 , n406540 );
xor ( n84263 , n405810 , n405825 );
xor ( n406543 , n84263 , n405848 );
buf ( n406544 , n406543 );
buf ( n406545 , n406544 );
and ( n406546 , n406541 , n406545 );
and ( n406547 , n406498 , n406540 );
or ( n84269 , n406546 , n406547 );
buf ( n406549 , n84269 );
buf ( n406550 , n406549 );
xor ( n406551 , n406481 , n406550 );
buf ( n406552 , n81950 );
buf ( n406553 , n57789 );
and ( n406554 , n406552 , n406553 );
buf ( n84276 , n403589 );
buf ( n406556 , n378470 );
and ( n406557 , n84276 , n406556 );
nor ( n84279 , n406554 , n406557 );
buf ( n406559 , n84279 );
buf ( n406560 , n406559 );
buf ( n406561 , n380581 );
or ( n84283 , n406560 , n406561 );
buf ( n406563 , n406489 );
buf ( n406564 , n378453 );
or ( n84286 , n406563 , n406564 );
nand ( n84287 , n84283 , n84286 );
buf ( n406567 , n84287 );
buf ( n406568 , n376997 );
xor ( n406569 , n376615 , n56214 );
buf ( n406570 , n406569 );
not ( n406571 , n406570 );
buf ( n406572 , n406571 );
buf ( n406573 , n406572 );
and ( n84295 , n406568 , n406573 );
buf ( n406575 , n376990 );
buf ( n406576 , n406569 );
and ( n84298 , n406575 , n406576 );
buf ( n406578 , n377003 );
nor ( n84300 , n84295 , n84298 , n406578 );
buf ( n406580 , n84300 );
xor ( n84302 , n406567 , n406580 );
xor ( n406582 , n406515 , n84258 );
buf ( n406583 , n406582 );
and ( n406584 , n84302 , n406583 );
and ( n84306 , n406567 , n406580 );
or ( n406586 , n406584 , n84306 );
buf ( n406587 , n400503 );
not ( n406588 , n57983 );
buf ( n406589 , n406588 );
and ( n84311 , n406587 , n406589 );
buf ( n406591 , n400509 );
buf ( n406592 , n63664 );
and ( n406593 , n406591 , n406592 );
nor ( n84315 , n84311 , n406593 );
buf ( n406595 , n84315 );
buf ( n406596 , n406595 );
buf ( n406597 , n60313 );
or ( n406598 , n406596 , n406597 );
buf ( n406599 , n83904 );
buf ( n406600 , n380733 );
or ( n84322 , n406599 , n406600 );
nand ( n406602 , n406598 , n84322 );
buf ( n406603 , n406602 );
xor ( n84325 , n406586 , n406603 );
buf ( n406605 , n382835 );
buf ( n406606 , n396615 );
and ( n406607 , n406605 , n406606 );
not ( n406608 , n406605 );
buf ( n406609 , n396621 );
and ( n84331 , n406608 , n406609 );
nor ( n84332 , n406607 , n84331 );
buf ( n406612 , n84332 );
buf ( n406613 , n406612 );
buf ( n406614 , n382849 );
or ( n84336 , n406613 , n406614 );
buf ( n406616 , n406472 );
buf ( n406617 , n384157 );
or ( n84339 , n406616 , n406617 );
nand ( n84340 , n84336 , n84339 );
buf ( n406620 , n84340 );
and ( n84342 , n84325 , n406620 );
and ( n84343 , n406586 , n406603 );
or ( n406623 , n84342 , n84343 );
buf ( n406624 , n406623 );
and ( n84346 , n406551 , n406624 );
and ( n84347 , n406481 , n406550 );
or ( n84348 , n84346 , n84347 );
buf ( n406628 , n84348 );
xor ( n406629 , n406025 , n406028 );
xor ( n406630 , n406629 , n406045 );
and ( n84352 , n406628 , n406630 );
buf ( n406632 , n74644 );
buf ( n406633 , n384343 );
and ( n406634 , n406632 , n406633 );
buf ( n406635 , n395683 );
buf ( n406636 , n384089 );
and ( n84358 , n406635 , n406636 );
nor ( n406638 , n406634 , n84358 );
buf ( n406639 , n406638 );
buf ( n406640 , n406639 );
buf ( n406641 , n384354 );
or ( n84363 , n406640 , n406641 );
buf ( n406643 , n406037 );
buf ( n406644 , n384082 );
or ( n406645 , n406643 , n406644 );
nand ( n84367 , n84363 , n406645 );
buf ( n406647 , n84367 );
xor ( n406648 , n83909 , n406018 );
xor ( n406649 , n406648 , n406022 );
and ( n84371 , n406647 , n406649 );
buf ( n406651 , n63549 );
buf ( n406652 , n394840 );
and ( n84374 , n406651 , n406652 );
buf ( n84375 , n384199 );
buf ( n406655 , n395890 );
and ( n406656 , n84375 , n406655 );
nor ( n406657 , n84374 , n406656 );
buf ( n406658 , n406657 );
buf ( n406659 , n406658 );
buf ( n406660 , n394838 );
or ( n406661 , n406659 , n406660 );
buf ( n406662 , n406452 );
buf ( n406663 , n394835 );
or ( n406664 , n406662 , n406663 );
nand ( n406665 , n406661 , n406664 );
buf ( n406666 , n406665 );
xor ( n406667 , n83909 , n406018 );
xor ( n84389 , n406667 , n406022 );
and ( n84390 , n406666 , n84389 );
and ( n406670 , n406647 , n406666 );
or ( n84392 , n84371 , n84390 , n406670 );
xor ( n84393 , n406025 , n406028 );
xor ( n84394 , n84393 , n406045 );
and ( n84395 , n84392 , n84394 );
and ( n406675 , n406628 , n84392 );
or ( n406676 , n84352 , n84395 , n406675 );
and ( n84398 , n406464 , n406676 );
and ( n406678 , n406424 , n406463 );
or ( n84400 , n84398 , n406678 );
xor ( n406680 , n83959 , n406079 );
xor ( n84402 , n406680 , n406083 );
and ( n84403 , n84400 , n84402 );
xor ( n406683 , n406049 , n406066 );
xor ( n406684 , n406683 , n83956 );
buf ( n406685 , n406684 );
xor ( n84407 , n406424 , n406463 );
xor ( n406687 , n84407 , n406676 );
and ( n84409 , n406685 , n406687 );
buf ( n406689 , n73625 );
buf ( n406690 , n394724 );
and ( n406691 , n406689 , n406690 );
buf ( n406692 , n73631 );
buf ( n406693 , n63434 );
and ( n406694 , n406692 , n406693 );
nor ( n406695 , n406691 , n406694 );
buf ( n406696 , n406695 );
buf ( n84418 , n406696 );
buf ( n406698 , n384414 );
or ( n84420 , n84418 , n406698 );
buf ( n406700 , n406432 );
buf ( n406701 , n395635 );
or ( n84423 , n406700 , n406701 );
nand ( n84424 , n84420 , n84423 );
buf ( n406704 , n84424 );
buf ( n406705 , n406704 );
buf ( n406706 , n395810 );
buf ( n406707 , n384343 );
and ( n84429 , n406706 , n406707 );
buf ( n406709 , n395816 );
buf ( n406710 , n384089 );
and ( n84432 , n406709 , n406710 );
nor ( n84433 , n84429 , n84432 );
buf ( n406713 , n84433 );
buf ( n406714 , n406713 );
buf ( n406715 , n384354 );
or ( n84437 , n406714 , n406715 );
buf ( n406717 , n406639 );
buf ( n406718 , n384082 );
or ( n406719 , n406717 , n406718 );
nand ( n84440 , n84437 , n406719 );
buf ( n406721 , n84440 );
buf ( n406722 , n406721 );
xor ( n406723 , n406498 , n406540 );
xor ( n84444 , n406723 , n406545 );
buf ( n406725 , n84444 );
buf ( n406726 , n406725 );
xor ( n84447 , n406722 , n406726 );
buf ( n406728 , n376924 );
buf ( n406729 , n376866 );
buf ( n406730 , n406569 );
and ( n84451 , n406729 , n406730 );
buf ( n406732 , n377030 );
buf ( n406733 , n406572 );
and ( n84454 , n406732 , n406733 );
nor ( n406735 , n84451 , n84454 );
buf ( n406736 , n406735 );
buf ( n406737 , n406736 );
or ( n84458 , n406728 , n406737 );
buf ( n406739 , n406507 );
buf ( n406740 , n56517 );
or ( n84461 , n406739 , n406740 );
nand ( n406742 , n84458 , n84461 );
buf ( n406743 , n406742 );
buf ( n406744 , n406743 );
buf ( n406745 , n376997 );
and ( n406746 , n376615 , n622 );
buf ( n406747 , n406746 );
not ( n406748 , n406747 );
buf ( n406749 , n406748 );
buf ( n406750 , n406749 );
and ( n406751 , n406745 , n406750 );
buf ( n406752 , n376990 );
buf ( n406753 , n406746 );
and ( n406754 , n406752 , n406753 );
buf ( n406755 , n377003 );
nor ( n84476 , n406751 , n406754 , n406755 );
buf ( n84477 , n84476 );
buf ( n406758 , n84477 );
xor ( n84479 , n406744 , n406758 );
buf ( n406760 , n378341 );
buf ( n406761 , n57800 );
buf ( n406762 , n403795 );
and ( n84483 , n406761 , n406762 );
buf ( n406764 , n378284 );
buf ( n406765 , n403798 );
and ( n84486 , n406764 , n406765 );
nor ( n406767 , n84483 , n84486 );
buf ( n406768 , n406767 );
buf ( n406769 , n406768 );
or ( n84490 , n406760 , n406769 );
buf ( n406771 , n378262 );
buf ( n406772 , n406523 );
or ( n84493 , n406771 , n406772 );
nand ( n406774 , n84490 , n84493 );
buf ( n406775 , n406774 );
buf ( n406776 , n406775 );
and ( n406777 , n84479 , n406776 );
and ( n406778 , n406744 , n406758 );
or ( n84499 , n406777 , n406778 );
buf ( n406780 , n84499 );
buf ( n406781 , n406780 );
buf ( n406782 , n79312 );
buf ( n406783 , n406588 );
and ( n406784 , n406782 , n406783 );
buf ( n406785 , n79318 );
buf ( n406786 , n82201 );
and ( n406787 , n406785 , n406786 );
nor ( n406788 , n406784 , n406787 );
buf ( n406789 , n406788 );
buf ( n406790 , n406789 );
buf ( n406791 , n60313 );
or ( n406792 , n406790 , n406791 );
buf ( n406793 , n406595 );
buf ( n406794 , n380733 );
or ( n406795 , n406793 , n406794 );
nand ( n406796 , n406792 , n406795 );
buf ( n406797 , n406796 );
buf ( n406798 , n406797 );
xor ( n406799 , n406781 , n406798 );
buf ( n406800 , n382663 );
not ( n406801 , n406800 );
buf ( n406802 , n406612 );
not ( n406803 , n406802 );
buf ( n406804 , n406803 );
buf ( n406805 , n406804 );
not ( n406806 , n406805 );
or ( n406807 , n406801 , n406806 );
buf ( n406808 , n79114 );
buf ( n406809 , n382835 );
and ( n84507 , n406808 , n406809 );
buf ( n406811 , n400487 );
buf ( n406812 , n62243 );
and ( n406813 , n406811 , n406812 );
nor ( n406814 , n84507 , n406813 );
buf ( n406815 , n406814 );
buf ( n406816 , n406815 );
buf ( n406817 , n382849 );
or ( n406818 , n406816 , n406817 );
nand ( n406819 , n406807 , n406818 );
buf ( n406820 , n406819 );
buf ( n406821 , n406820 );
and ( n406822 , n406799 , n406821 );
and ( n84514 , n406781 , n406798 );
or ( n406824 , n406822 , n84514 );
buf ( n406825 , n406824 );
buf ( n406826 , n406825 );
and ( n84518 , n84447 , n406826 );
and ( n84519 , n406722 , n406726 );
or ( n84520 , n84518 , n84519 );
buf ( n406830 , n84520 );
buf ( n406831 , n406830 );
xor ( n406832 , n406705 , n406831 );
xor ( n84524 , n406481 , n406550 );
xor ( n406834 , n84524 , n406624 );
buf ( n406835 , n406834 );
buf ( n406836 , n406835 );
and ( n406837 , n406832 , n406836 );
and ( n84529 , n406705 , n406831 );
or ( n406839 , n406837 , n84529 );
buf ( n406840 , n406839 );
xor ( n84532 , n406440 , n406443 );
xor ( n406842 , n84532 , n84183 );
and ( n406843 , n406840 , n406842 );
xor ( n84535 , n406025 , n406028 );
xor ( n84536 , n84535 , n406045 );
xor ( n406846 , n406628 , n84392 );
xor ( n84537 , n84536 , n406846 );
xor ( n406848 , n406440 , n406443 );
xor ( n84539 , n406848 , n84183 );
and ( n84540 , n84537 , n84539 );
and ( n84541 , n406840 , n84537 );
or ( n84542 , n406843 , n84540 , n84541 );
xor ( n84543 , n406424 , n406463 );
xor ( n84544 , n84543 , n406676 );
and ( n84545 , n84542 , n84544 );
and ( n84546 , n406685 , n84542 );
or ( n84547 , n84409 , n84545 , n84546 );
xor ( n84548 , n83959 , n406079 );
xor ( n406859 , n84548 , n406083 );
and ( n84550 , n84547 , n406859 );
and ( n406861 , n84400 , n84547 );
or ( n84552 , n84403 , n84550 , n406861 );
buf ( n406863 , n84552 );
xor ( n84554 , n405722 , n83753 );
xor ( n84555 , n84554 , n405766 );
xor ( n406866 , n405983 , n406086 );
xor ( n406867 , n84555 , n406866 );
buf ( n406868 , n406867 );
xor ( n406869 , n406863 , n406868 );
buf ( n406870 , n377379 );
not ( n84561 , n406870 );
buf ( n406872 , n406246 );
not ( n406873 , n406872 );
or ( n84564 , n84561 , n406873 );
buf ( n406875 , n369183 );
buf ( n406876 , n377379 );
or ( n406877 , n406875 , n406876 );
buf ( n406878 , n406877 );
buf ( n406879 , n406878 );
nand ( n406880 , n84564 , n406879 );
buf ( n406881 , n406880 );
buf ( n406882 , n406881 );
not ( n84573 , n406882 );
buf ( n406884 , n406260 );
not ( n84575 , n406884 );
or ( n84576 , n84573 , n84575 );
buf ( n406887 , n365076 );
not ( n406888 , n406887 );
buf ( n84579 , n406256 );
nand ( n84580 , n406888 , n84579 );
buf ( n84581 , n84580 );
buf ( n406892 , n84581 );
nand ( n84583 , n84576 , n406892 );
buf ( n406894 , n84583 );
buf ( n406895 , n406894 );
and ( n84586 , n406869 , n406895 );
and ( n406897 , n406863 , n406868 );
or ( n84588 , n84586 , n406897 );
buf ( n406899 , n84588 );
buf ( n406900 , n406899 );
xor ( n84591 , n406421 , n406900 );
buf ( n406902 , n369444 );
not ( n84593 , n406902 );
buf ( n406904 , n406298 );
not ( n406905 , n406904 );
or ( n406906 , n84593 , n406905 );
and ( n84597 , n48791 , n368549 );
not ( n406908 , n48791 );
and ( n406909 , n406908 , n44906 );
or ( n84600 , n84597 , n406909 );
buf ( n406911 , n84600 );
buf ( n406912 , n368602 );
nand ( n406913 , n406911 , n406912 );
buf ( n406914 , n406913 );
buf ( n406915 , n406914 );
nand ( n406916 , n406906 , n406915 );
buf ( n406917 , n406916 );
buf ( n406918 , n406917 );
nand ( n84609 , n84600 , n48418 );
xor ( n84610 , n83959 , n406079 );
xor ( n84611 , n84610 , n406083 );
xor ( n84612 , n84400 , n84547 );
xor ( n84613 , n84611 , n84612 );
not ( n84614 , n84613 );
buf ( n84615 , n368599 );
buf ( n406926 , n84615 );
buf ( n406927 , n23037 );
buf ( n406928 , n352353 );
not ( n84619 , n406928 );
buf ( n406930 , n84619 );
buf ( n406931 , n406930 );
not ( n84622 , n406931 );
buf ( n406933 , n84622 );
buf ( n406934 , n406933 );
and ( n84625 , n406927 , n406934 );
not ( n84626 , n406927 );
buf ( n406937 , n369372 );
and ( n406938 , n84626 , n406937 );
nor ( n84629 , n84625 , n406938 );
buf ( n406940 , n84629 );
buf ( n406941 , n406940 );
nand ( n84632 , n406926 , n406941 );
buf ( n84633 , n84632 );
nand ( n84634 , n84609 , n84614 , n84633 );
not ( n84635 , n84634 );
buf ( n406946 , n377353 );
not ( n406947 , n406946 );
buf ( n406948 , n342964 );
buf ( n84639 , n406948 );
buf ( n406950 , n84639 );
buf ( n406951 , n406950 );
not ( n406952 , n406951 );
buf ( n406953 , n406952 );
buf ( n406954 , n406953 );
not ( n84645 , n406954 );
or ( n406956 , n406947 , n84645 );
buf ( n406957 , n406950 );
buf ( n406958 , n377352 );
nand ( n406959 , n406957 , n406958 );
buf ( n406960 , n406959 );
buf ( n406961 , n406960 );
nand ( n406962 , n406956 , n406961 );
buf ( n406963 , n406962 );
buf ( n406964 , n406963 );
not ( n406965 , n406964 );
buf ( n406966 , n406260 );
not ( n406967 , n406966 );
or ( n84658 , n406965 , n406967 );
buf ( n84659 , n406881 );
buf ( n84660 , n44915 );
nand ( n84661 , n84659 , n84660 );
buf ( n84662 , n84661 );
buf ( n84663 , n84662 );
nand ( n84664 , n84658 , n84663 );
buf ( n84665 , n84664 );
not ( n406976 , n84665 );
or ( n84667 , n84635 , n406976 );
nand ( n406978 , n84609 , n84633 );
nand ( n406979 , n406978 , n84613 );
nand ( n84670 , n84667 , n406979 );
buf ( n406981 , n84670 );
xor ( n84672 , n406918 , n406981 );
xor ( n84673 , n406863 , n406868 );
xor ( n406984 , n84673 , n406895 );
buf ( n406985 , n406984 );
buf ( n406986 , n406985 );
and ( n84677 , n84672 , n406986 );
and ( n84678 , n406918 , n406981 );
or ( n406989 , n84677 , n84678 );
buf ( n406990 , n406989 );
buf ( n406991 , n406990 );
and ( n406992 , n84591 , n406991 );
and ( n406993 , n406421 , n406900 );
or ( n84684 , n406992 , n406993 );
buf ( n406995 , n84684 );
buf ( n84686 , n406995 );
buf ( n406997 , n406413 );
not ( n406998 , n406997 );
buf ( n406999 , n45012 );
not ( n84690 , n406999 );
or ( n407001 , n406998 , n84690 );
buf ( n84692 , n405385 );
buf ( n407003 , n365149 );
nand ( n407004 , n84692 , n407003 );
buf ( n407005 , n407004 );
buf ( n407006 , n407005 );
nand ( n407007 , n407001 , n407006 );
buf ( n407008 , n407007 );
buf ( n407009 , n407008 );
xor ( n84700 , n406097 , n406102 );
xor ( n84701 , n84700 , n406128 );
buf ( n407012 , n84701 );
buf ( n407013 , n407012 );
xor ( n84704 , n407009 , n407013 );
buf ( n407015 , n406143 );
buf ( n407016 , n368624 );
or ( n407017 , n407015 , n407016 );
buf ( n407018 , n84047 );
buf ( n407019 , n368602 );
nand ( n407020 , n407018 , n407019 );
buf ( n407021 , n407020 );
buf ( n407022 , n407021 );
nand ( n407023 , n407017 , n407022 );
buf ( n407024 , n407023 );
buf ( n407025 , n407024 );
xor ( n407026 , n84704 , n407025 );
buf ( n407027 , n407026 );
buf ( n407028 , n407027 );
xor ( n84719 , n84686 , n407028 );
buf ( n407030 , n377143 );
buf ( n407031 , n386093 );
and ( n407032 , n407030 , n407031 );
not ( n84723 , n407030 );
buf ( n407034 , n386102 );
and ( n84725 , n84723 , n407034 );
nor ( n407036 , n407032 , n84725 );
buf ( n407037 , n407036 );
buf ( n407038 , n407037 );
not ( n407039 , n407038 );
buf ( n407040 , n365024 );
not ( n407041 , n407040 );
or ( n84732 , n407039 , n407041 );
buf ( n407043 , n377757 );
not ( n407044 , n407043 );
buf ( n407045 , n364978 );
not ( n84736 , n407045 );
or ( n407047 , n407044 , n84736 );
buf ( n407048 , n386093 );
buf ( n407049 , n378886 );
nand ( n407050 , n407048 , n407049 );
buf ( n407051 , n407050 );
buf ( n407052 , n407051 );
nand ( n84743 , n407047 , n407052 );
buf ( n84744 , n84743 );
buf ( n407055 , n84744 );
buf ( n407056 , n365108 );
nand ( n407057 , n407055 , n407056 );
buf ( n407058 , n407057 );
buf ( n407059 , n407058 );
nand ( n407060 , n84732 , n407059 );
buf ( n407061 , n407060 );
buf ( n407062 , n407061 );
and ( n84753 , n84719 , n407062 );
and ( n84754 , n84686 , n407028 );
or ( n84755 , n84753 , n84754 );
buf ( n407066 , n84755 );
buf ( n407067 , n407066 );
and ( n84758 , n84134 , n407067 );
and ( n84759 , n406374 , n84133 );
or ( n84760 , n84758 , n84759 );
buf ( n407071 , n84760 );
buf ( n407072 , n407071 );
xor ( n84763 , n406233 , n407072 );
xor ( n84764 , n405348 , n405368 );
xor ( n84765 , n84764 , n405398 );
buf ( n407076 , n84765 );
buf ( n407077 , n407076 );
xor ( n84768 , n407009 , n407013 );
and ( n407079 , n84768 , n407025 );
and ( n407080 , n407009 , n407013 );
or ( n84771 , n407079 , n407080 );
buf ( n407082 , n84771 );
buf ( n407083 , n407082 );
xor ( n84774 , n407077 , n407083 );
buf ( n407085 , n84744 );
not ( n407086 , n407085 );
buf ( n407087 , n365024 );
not ( n84778 , n407087 );
or ( n407089 , n407086 , n84778 );
buf ( n407090 , n404930 );
buf ( n407091 , n365108 );
nand ( n407092 , n407090 , n407091 );
buf ( n407093 , n407092 );
buf ( n407094 , n407093 );
nand ( n407095 , n407089 , n407094 );
buf ( n407096 , n407095 );
buf ( n407097 , n407096 );
xor ( n407098 , n84774 , n407097 );
buf ( n407099 , n407098 );
buf ( n407100 , n407099 );
buf ( n407101 , n363416 );
buf ( n407102 , n379515 );
nor ( n407103 , n407101 , n407102 );
buf ( n407104 , n407103 );
buf ( n407105 , n407104 );
xor ( n407106 , n407100 , n407105 );
buf ( n84781 , n378843 );
buf ( n84782 , n375914 );
and ( n84783 , n84781 , n84782 );
not ( n84784 , n84781 );
buf ( n84785 , n377279 );
and ( n84786 , n84784 , n84785 );
nor ( n84787 , n84783 , n84786 );
buf ( n84788 , n84787 );
buf ( n407115 , n84788 );
not ( n84790 , n407115 );
buf ( n407117 , n399191 );
not ( n407118 , n407117 );
or ( n84793 , n84790 , n407118 );
buf ( n407120 , n58984 );
buf ( n407121 , n375901 );
and ( n84796 , n407120 , n407121 );
not ( n407123 , n407120 );
buf ( n407124 , n377279 );
and ( n84799 , n407123 , n407124 );
nor ( n407126 , n84796 , n84799 );
buf ( n407127 , n407126 );
buf ( n407128 , n407127 );
buf ( n407129 , n375920 );
nand ( n407130 , n407128 , n407129 );
buf ( n407131 , n407130 );
buf ( n407132 , n407131 );
nand ( n407133 , n84793 , n407132 );
buf ( n407134 , n407133 );
buf ( n407135 , n407134 );
and ( n407136 , n407106 , n407135 );
and ( n84811 , n407100 , n407105 );
or ( n407138 , n407136 , n84811 );
buf ( n407139 , n407138 );
buf ( n407140 , n407139 );
and ( n84815 , n84763 , n407140 );
and ( n84816 , n406233 , n407072 );
or ( n407143 , n84815 , n84816 );
buf ( n407144 , n407143 );
buf ( n407145 , n407144 );
xor ( n407146 , n405719 , n407145 );
buf ( n407147 , n58867 );
not ( n84822 , n407147 );
buf ( n407149 , n379371 );
not ( n407150 , n407149 );
buf ( n407151 , n31073 );
not ( n84826 , n407151 );
or ( n407153 , n407150 , n84826 );
buf ( n407154 , n351107 );
buf ( n407155 , n379392 );
nand ( n407156 , n407154 , n407155 );
buf ( n407157 , n407156 );
buf ( n407158 , n407157 );
nand ( n407159 , n407153 , n407158 );
buf ( n407160 , n407159 );
buf ( n407161 , n407160 );
not ( n84836 , n407161 );
or ( n84837 , n84822 , n84836 );
buf ( n407164 , n379368 );
not ( n407165 , n407164 );
buf ( n407166 , n45459 );
not ( n84841 , n407166 );
or ( n84842 , n407165 , n84841 );
buf ( n407169 , n364858 );
buf ( n407170 , n379392 );
nand ( n84845 , n407169 , n407170 );
buf ( n407172 , n84845 );
buf ( n407173 , n407172 );
nand ( n84848 , n84842 , n407173 );
buf ( n407175 , n84848 );
buf ( n407176 , n407175 );
buf ( n407177 , n58923 );
nand ( n84852 , n407176 , n407177 );
buf ( n407179 , n84852 );
buf ( n407180 , n407179 );
nand ( n407181 , n84837 , n407180 );
buf ( n407182 , n407181 );
buf ( n407183 , n407182 );
xor ( n407184 , n407146 , n407183 );
buf ( n407185 , n407184 );
xor ( n407186 , n406233 , n407072 );
xor ( n84861 , n407186 , n407140 );
buf ( n407188 , n84861 );
buf ( n84863 , n407188 );
buf ( n407190 , n380356 );
not ( n84865 , n407190 );
buf ( n407192 , n380368 );
buf ( n407193 , n42891 );
and ( n84868 , n407192 , n407193 );
not ( n407195 , n407192 );
buf ( n407196 , n42898 );
and ( n84871 , n407195 , n407196 );
nor ( n407198 , n84868 , n84871 );
buf ( n407199 , n407198 );
buf ( n407200 , n407199 );
not ( n407201 , n407200 );
or ( n407202 , n84865 , n407201 );
buf ( n407203 , n380368 );
buf ( n407204 , n364858 );
and ( n84879 , n407203 , n407204 );
not ( n407206 , n407203 );
buf ( n407207 , n45459 );
and ( n407208 , n407206 , n407207 );
nor ( n84883 , n84879 , n407208 );
buf ( n407210 , n84883 );
buf ( n84885 , n407210 );
buf ( n84886 , n380404 );
nand ( n84887 , n84885 , n84886 );
buf ( n84888 , n84887 );
buf ( n84889 , n84888 );
nand ( n84890 , n407202 , n84889 );
buf ( n84891 , n84890 );
buf ( n407218 , n84891 );
xor ( n84893 , n84863 , n407218 );
buf ( n407220 , n379371 );
not ( n407221 , n407220 );
buf ( n407222 , n351318 );
not ( n84897 , n407222 );
or ( n407224 , n407221 , n84897 );
buf ( n407225 , n364808 );
buf ( n407226 , n379368 );
not ( n407227 , n407226 );
buf ( n407228 , n407227 );
buf ( n407229 , n407228 );
nand ( n407230 , n407225 , n407229 );
buf ( n407231 , n407230 );
buf ( n407232 , n407231 );
nand ( n407233 , n407224 , n407232 );
buf ( n407234 , n407233 );
not ( n84909 , n407234 );
not ( n407236 , n58867 );
or ( n84911 , n84909 , n407236 );
buf ( n407238 , n407160 );
not ( n407239 , n407238 );
buf ( n407240 , n407239 );
or ( n407241 , n407240 , n381675 );
nand ( n407242 , n84911 , n407241 );
buf ( n407243 , n407242 );
and ( n407244 , n84893 , n407243 );
and ( n407245 , n84863 , n407218 );
or ( n84914 , n407244 , n407245 );
buf ( n407247 , n84914 );
xor ( n84916 , n407185 , n407247 );
buf ( n84917 , n405322 );
buf ( n407250 , n405340 );
xor ( n407251 , n84917 , n407250 );
buf ( n407252 , n405402 );
xnor ( n84921 , n407251 , n407252 );
buf ( n407254 , n84921 );
buf ( n407255 , n407254 );
not ( n84924 , n407255 );
buf ( n407257 , n84924 );
not ( n84926 , n407257 );
buf ( n407259 , n404992 );
buf ( n407260 , n404987 );
xor ( n84929 , n407259 , n407260 );
buf ( n407262 , n404950 );
xnor ( n407263 , n84929 , n407262 );
buf ( n407264 , n407263 );
buf ( n407265 , n407264 );
not ( n84934 , n407265 );
buf ( n407267 , n84934 );
not ( n84936 , n407267 );
or ( n84937 , n84926 , n84936 );
not ( n84938 , n407254 );
not ( n84939 , n407264 );
or ( n84940 , n84938 , n84939 );
xor ( n84941 , n407077 , n407083 );
and ( n407274 , n84941 , n407097 );
and ( n84943 , n407077 , n407083 );
or ( n407276 , n407274 , n84943 );
buf ( n407277 , n407276 );
nand ( n407278 , n84940 , n407277 );
nand ( n407279 , n84937 , n407278 );
buf ( n407280 , n407279 );
buf ( n407281 , n48490 );
buf ( n407282 , n378098 );
and ( n84951 , n407281 , n407282 );
buf ( n407284 , n84951 );
buf ( n84953 , n407284 );
xor ( n84954 , n407280 , n84953 );
xor ( n407287 , n404876 , n404917 );
xor ( n407288 , n407287 , n405004 );
buf ( n407289 , n407288 );
buf ( n407290 , n407289 );
xor ( n84959 , n84954 , n407290 );
buf ( n407292 , n84959 );
buf ( n407293 , n407292 );
buf ( n407294 , n380404 );
not ( n84963 , n407294 );
buf ( n407296 , n407199 );
not ( n84965 , n407296 );
or ( n407298 , n84963 , n84965 );
buf ( n407299 , n380368 );
not ( n407300 , n407299 );
buf ( n407301 , n364771 );
not ( n84970 , n407301 );
or ( n84971 , n407300 , n84970 );
buf ( n407304 , n42911 );
buf ( n407305 , n384667 );
nand ( n407306 , n407304 , n407305 );
buf ( n407307 , n407306 );
buf ( n407308 , n407307 );
nand ( n407309 , n84971 , n407308 );
buf ( n407310 , n407309 );
buf ( n407311 , n407310 );
buf ( n407312 , n380356 );
nand ( n84981 , n407311 , n407312 );
buf ( n407314 , n84981 );
buf ( n407315 , n407314 );
nand ( n407316 , n407298 , n407315 );
buf ( n407317 , n407316 );
buf ( n407318 , n407317 );
xor ( n407319 , n407293 , n407318 );
buf ( n407320 , n379274 );
not ( n84989 , n407320 );
buf ( n407322 , n365259 );
not ( n84991 , n407322 );
or ( n407324 , n84989 , n84991 );
buf ( n407325 , n352209 );
buf ( n407326 , n379271 );
nand ( n407327 , n407325 , n407326 );
buf ( n407328 , n407327 );
buf ( n407329 , n407328 );
nand ( n407330 , n407324 , n407329 );
buf ( n407331 , n407330 );
buf ( n407332 , n407331 );
buf ( n407333 , n379263 );
and ( n407334 , n407332 , n407333 );
buf ( n407335 , n379274 );
not ( n407336 , n407335 );
buf ( n407337 , n365474 );
not ( n85004 , n407337 );
or ( n407339 , n407336 , n85004 );
buf ( n407340 , n66894 );
buf ( n407341 , n379271 );
nand ( n407342 , n407340 , n407341 );
buf ( n407343 , n407342 );
buf ( n407344 , n407343 );
nand ( n407345 , n407339 , n407344 );
buf ( n85009 , n407345 );
buf ( n407347 , n85009 );
not ( n85011 , n407347 );
buf ( n407349 , n379296 );
nor ( n407350 , n85011 , n407349 );
buf ( n407351 , n407350 );
buf ( n407352 , n407351 );
nor ( n407353 , n407334 , n407352 );
buf ( n407354 , n407353 );
buf ( n407355 , n407354 );
buf ( n407356 , n398363 );
not ( n407357 , n407356 );
buf ( n407358 , n365344 );
not ( n407359 , n407358 );
or ( n407360 , n407357 , n407359 );
buf ( n407361 , n378736 );
buf ( n407362 , n377592 );
nand ( n407363 , n407361 , n407362 );
buf ( n85022 , n407363 );
buf ( n407365 , n85022 );
nand ( n85024 , n407360 , n407365 );
buf ( n85025 , n85024 );
buf ( n407368 , n85025 );
buf ( n407369 , n397190 );
and ( n407370 , n407368 , n407369 );
buf ( n407371 , n377585 );
not ( n85030 , n407371 );
buf ( n407373 , n31194 );
not ( n85032 , n407373 );
or ( n85033 , n85030 , n85032 );
buf ( n407376 , n83069 );
buf ( n407377 , n377592 );
nand ( n407378 , n407376 , n407377 );
buf ( n407379 , n407378 );
buf ( n407380 , n407379 );
nand ( n85039 , n85033 , n407380 );
buf ( n407382 , n85039 );
buf ( n407383 , n407382 );
not ( n85042 , n407383 );
buf ( n407385 , n377618 );
nor ( n407386 , n85042 , n407385 );
buf ( n407387 , n407386 );
buf ( n407388 , n407387 );
nor ( n407389 , n407370 , n407388 );
buf ( n407390 , n407389 );
buf ( n407391 , n407390 );
not ( n407392 , n407391 );
buf ( n407393 , n407392 );
buf ( n407394 , n407393 );
not ( n407395 , n407394 );
buf ( n407396 , n362377 );
buf ( n407397 , n363411 );
not ( n407398 , n407397 );
buf ( n407399 , n63905 );
not ( n85058 , n407399 );
or ( n407401 , n407398 , n85058 );
buf ( n407402 , n378098 );
nand ( n407403 , n407401 , n407402 );
buf ( n407404 , n407403 );
buf ( n407405 , n407404 );
buf ( n407406 , n363411 );
not ( n85065 , n407406 );
buf ( n407408 , n342656 );
nand ( n407409 , n85065 , n407408 );
buf ( n407410 , n407409 );
buf ( n407411 , n407410 );
nand ( n407412 , n407396 , n407405 , n407411 );
buf ( n407413 , n407412 );
buf ( n407414 , n407413 );
not ( n407415 , n407414 );
buf ( n407416 , n407415 );
buf ( n407417 , n407416 );
not ( n407418 , n407417 );
or ( n85077 , n407395 , n407418 );
buf ( n407420 , n407413 );
not ( n407421 , n407420 );
buf ( n407422 , n407390 );
not ( n407423 , n407422 );
or ( n85082 , n407421 , n407423 );
buf ( n407425 , n407127 );
not ( n85084 , n407425 );
buf ( n407427 , n375896 );
not ( n85086 , n407427 );
or ( n85087 , n85084 , n85086 );
buf ( n407430 , n377122 );
not ( n407431 , n407430 );
buf ( n407432 , n388576 );
not ( n407433 , n407432 );
or ( n407434 , n407431 , n407433 );
buf ( n407435 , n375901 );
buf ( n407436 , n57463 );
nand ( n407437 , n407435 , n407436 );
buf ( n407438 , n407437 );
buf ( n407439 , n407438 );
nand ( n407440 , n407434 , n407439 );
buf ( n407441 , n407440 );
buf ( n407442 , n407441 );
buf ( n407443 , n375920 );
nand ( n407444 , n407442 , n407443 );
buf ( n407445 , n407444 );
buf ( n407446 , n407445 );
nand ( n85105 , n85087 , n407446 );
buf ( n85106 , n85105 );
buf ( n407449 , n85106 );
nand ( n85108 , n85082 , n407449 );
buf ( n407451 , n85108 );
buf ( n407452 , n407451 );
nand ( n85111 , n85077 , n407452 );
buf ( n407454 , n85111 );
buf ( n407455 , n407454 );
not ( n85114 , n407455 );
buf ( n407457 , n85114 );
buf ( n407458 , n407457 );
and ( n407459 , n407355 , n407458 );
not ( n407460 , n407355 );
buf ( n407461 , n407454 );
and ( n407462 , n407460 , n407461 );
nor ( n407463 , n407459 , n407462 );
buf ( n407464 , n407463 );
buf ( n407465 , n407464 );
xor ( n407466 , n405035 , n405052 );
xor ( n407467 , n407466 , n405061 );
buf ( n407468 , n407467 );
buf ( n407469 , n407468 );
buf ( n407470 , n407441 );
not ( n407471 , n407470 );
buf ( n407472 , n375896 );
not ( n407473 , n407472 );
or ( n407474 , n407471 , n407473 );
buf ( n407475 , n405244 );
buf ( n407476 , n46463 );
nand ( n407477 , n407475 , n407476 );
buf ( n407478 , n407477 );
buf ( n407479 , n407478 );
nand ( n407480 , n407474 , n407479 );
buf ( n407481 , n407480 );
buf ( n407482 , n407481 );
xor ( n407483 , n407469 , n407482 );
buf ( n407484 , n50782 );
or ( n85120 , n396289 , n58378 );
nand ( n85121 , n22707 , n58378 );
nand ( n85122 , n85120 , n85121 );
buf ( n407488 , n85122 );
or ( n85124 , n407484 , n407488 );
buf ( n407490 , n377168 );
buf ( n407491 , n404760 );
or ( n85127 , n407490 , n407491 );
nand ( n407493 , n85124 , n85127 );
buf ( n407494 , n407493 );
buf ( n407495 , n407494 );
xor ( n85131 , n407483 , n407495 );
buf ( n407497 , n85131 );
buf ( n407498 , n407497 );
and ( n407499 , n407465 , n407498 );
not ( n85135 , n407465 );
buf ( n407501 , n407497 );
not ( n407502 , n407501 );
buf ( n407503 , n407502 );
buf ( n407504 , n407503 );
and ( n407505 , n85135 , n407504 );
nor ( n85141 , n407499 , n407505 );
buf ( n407507 , n85141 );
buf ( n407508 , n407507 );
xor ( n407509 , n407319 , n407508 );
buf ( n407510 , n407509 );
xor ( n85146 , n84916 , n407510 );
buf ( n407512 , n85146 );
xor ( n85148 , n84863 , n407218 );
xor ( n85149 , n85148 , n407243 );
buf ( n407515 , n85149 );
buf ( n407516 , n407515 );
buf ( n407517 , n369809 );
not ( n407518 , n407517 );
buf ( n407519 , n406222 );
not ( n407520 , n407519 );
or ( n407521 , n407518 , n407520 );
buf ( n407522 , n406320 );
buf ( n407523 , n369804 );
nand ( n407524 , n407522 , n407523 );
buf ( n407525 , n407524 );
buf ( n407526 , n407525 );
nand ( n407527 , n407521 , n407526 );
buf ( n407528 , n407527 );
buf ( n407529 , n407528 );
xor ( n407530 , n406133 , n406152 );
xor ( n407531 , n407530 , n406174 );
buf ( n407532 , n407531 );
buf ( n407533 , n407532 );
xor ( n407534 , n407529 , n407533 );
buf ( n407535 , n397190 );
not ( n407536 , n407535 );
buf ( n407537 , n407382 );
not ( n85163 , n407537 );
or ( n407539 , n407536 , n85163 );
buf ( n407540 , n377585 );
not ( n407541 , n407540 );
buf ( n407542 , n45336 );
not ( n85168 , n407542 );
or ( n407544 , n407541 , n85168 );
buf ( n407545 , n404902 );
buf ( n407546 , n377592 );
nand ( n407547 , n407545 , n407546 );
buf ( n407548 , n407547 );
buf ( n407549 , n407548 );
nand ( n407550 , n407544 , n407549 );
buf ( n407551 , n407550 );
buf ( n407552 , n407551 );
not ( n407553 , n57170 );
buf ( n85179 , n407553 );
buf ( n407555 , n85179 );
nand ( n407556 , n407552 , n407555 );
buf ( n407557 , n407556 );
buf ( n407558 , n407557 );
nand ( n85184 , n407539 , n407558 );
buf ( n407560 , n85184 );
buf ( n407561 , n407560 );
xor ( n85187 , n407534 , n407561 );
buf ( n407563 , n85187 );
buf ( n407564 , n407563 );
xor ( n85190 , n406374 , n84133 );
xor ( n407566 , n85190 , n407067 );
buf ( n407567 , n407566 );
buf ( n407568 , n407567 );
xor ( n407569 , n407564 , n407568 );
buf ( n407570 , n379890 );
not ( n85196 , n407570 );
buf ( n407572 , n379838 );
not ( n407573 , n407572 );
buf ( n407574 , n386359 );
not ( n85200 , n407574 );
or ( n407576 , n407573 , n85200 );
buf ( n407577 , n352212 );
buf ( n407578 , n398741 );
nand ( n85204 , n407577 , n407578 );
buf ( n407580 , n85204 );
buf ( n407581 , n407580 );
nand ( n85207 , n407576 , n407581 );
buf ( n407583 , n85207 );
buf ( n407584 , n407583 );
not ( n85210 , n407584 );
or ( n85211 , n85196 , n85210 );
buf ( n407587 , n379838 );
not ( n85213 , n407587 );
buf ( n407589 , n351292 );
not ( n85215 , n407589 );
or ( n85216 , n85213 , n85215 );
buf ( n407592 , n66894 );
buf ( n407593 , n398741 );
nand ( n85219 , n407592 , n407593 );
buf ( n407595 , n85219 );
buf ( n407596 , n407595 );
nand ( n407597 , n85216 , n407596 );
buf ( n407598 , n407597 );
buf ( n407599 , n407598 );
buf ( n407600 , n379916 );
nand ( n85226 , n407599 , n407600 );
buf ( n407602 , n85226 );
buf ( n407603 , n407602 );
nand ( n85229 , n85211 , n407603 );
buf ( n407605 , n85229 );
buf ( n407606 , n407605 );
and ( n85232 , n407569 , n407606 );
and ( n407608 , n407564 , n407568 );
or ( n85234 , n85232 , n407608 );
buf ( n407610 , n85234 );
buf ( n407611 , n407610 );
buf ( n407612 , n58984 );
buf ( n407613 , n395541 );
and ( n407614 , n407612 , n407613 );
not ( n85240 , n407612 );
buf ( n407616 , n380923 );
and ( n407617 , n85240 , n407616 );
nor ( n85243 , n407614 , n407617 );
buf ( n85244 , n85243 );
buf ( n407620 , n85244 );
not ( n407621 , n407620 );
buf ( n407622 , n384501 );
not ( n407623 , n407622 );
or ( n407624 , n407621 , n407623 );
buf ( n407625 , n406378 );
buf ( n407626 , n56794 );
nand ( n85252 , n407625 , n407626 );
buf ( n407628 , n85252 );
buf ( n407629 , n407628 );
nand ( n407630 , n407624 , n407629 );
buf ( n407631 , n407630 );
buf ( n407632 , n407631 );
buf ( n407633 , n397190 );
not ( n85259 , n407633 );
buf ( n407635 , n407551 );
not ( n407636 , n407635 );
or ( n85262 , n85259 , n407636 );
buf ( n85263 , n377585 );
not ( n85264 , n85263 );
buf ( n85265 , n381266 );
not ( n85266 , n85265 );
or ( n85267 , n85264 , n85266 );
buf ( n85268 , n351160 );
buf ( n85269 , n377592 );
nand ( n85270 , n85268 , n85269 );
buf ( n85271 , n85270 );
buf ( n85272 , n85271 );
nand ( n85273 , n85267 , n85272 );
buf ( n85274 , n85273 );
buf ( n407650 , n85274 );
buf ( n407651 , n85179 );
nand ( n85277 , n407650 , n407651 );
buf ( n407653 , n85277 );
buf ( n407654 , n407653 );
nand ( n85280 , n85262 , n407654 );
buf ( n85281 , n85280 );
buf ( n407657 , n85281 );
xor ( n85283 , n407632 , n407657 );
buf ( n407659 , n377068 );
not ( n85285 , n407659 );
buf ( n407661 , n388576 );
not ( n85287 , n407661 );
or ( n407663 , n85285 , n85287 );
buf ( n407664 , n378135 );
buf ( n407665 , n377071 );
nand ( n407666 , n407664 , n407665 );
buf ( n407667 , n407666 );
buf ( n407668 , n407667 );
nand ( n407669 , n407663 , n407668 );
buf ( n407670 , n407669 );
buf ( n407671 , n407670 );
not ( n407672 , n407671 );
buf ( n407673 , n375896 );
not ( n85299 , n407673 );
or ( n85300 , n407672 , n85299 );
buf ( n407676 , n84788 );
buf ( n85302 , n375920 );
nand ( n85303 , n407676 , n85302 );
buf ( n407679 , n85303 );
buf ( n407680 , n407679 );
nand ( n85306 , n85300 , n407680 );
buf ( n407682 , n85306 );
buf ( n407683 , n407682 );
and ( n407684 , n85283 , n407683 );
and ( n85310 , n407632 , n407657 );
or ( n407686 , n407684 , n85310 );
buf ( n407687 , n407686 );
buf ( n407688 , n407687 );
xor ( n85314 , n84686 , n407028 );
xor ( n85315 , n85314 , n407062 );
buf ( n407691 , n85315 );
buf ( n407692 , n407691 );
buf ( n407693 , n406346 );
not ( n407694 , n407693 );
buf ( n407695 , n396401 );
not ( n407696 , n407695 );
or ( n85322 , n407694 , n407696 );
buf ( n407698 , n80732 );
buf ( n407699 , n377779 );
nand ( n85325 , n407698 , n407699 );
buf ( n407701 , n85325 );
buf ( n407702 , n407701 );
nand ( n85328 , n85322 , n407702 );
buf ( n407704 , n85328 );
buf ( n407705 , n407704 );
not ( n85331 , n407705 );
buf ( n407707 , n365181 );
not ( n407708 , n407707 );
or ( n85334 , n85331 , n407708 );
buf ( n407710 , n406398 );
buf ( n407711 , n365146 );
not ( n407712 , n407711 );
buf ( n407713 , n407712 );
buf ( n407714 , n407713 );
nand ( n407715 , n407710 , n407714 );
buf ( n407716 , n407715 );
buf ( n407717 , n407716 );
nand ( n407718 , n85334 , n407717 );
buf ( n407719 , n407718 );
buf ( n407720 , n407719 );
buf ( n407721 , n369809 );
not ( n85347 , n407721 );
buf ( n407723 , n393883 );
not ( n407724 , n407723 );
buf ( n407725 , n402185 );
not ( n85351 , n407725 );
or ( n85352 , n407724 , n85351 );
buf ( n407728 , n351345 );
buf ( n407729 , n369763 );
nand ( n85355 , n407728 , n407729 );
buf ( n407731 , n85355 );
buf ( n407732 , n407731 );
nand ( n407733 , n85352 , n407732 );
buf ( n407734 , n407733 );
buf ( n407735 , n407734 );
not ( n407736 , n407735 );
or ( n85362 , n85347 , n407736 );
buf ( n407738 , n393883 );
not ( n407739 , n407738 );
buf ( n407740 , n365384 );
not ( n85366 , n407740 );
or ( n85367 , n407739 , n85366 );
buf ( n407743 , n402205 );
buf ( n407744 , n369763 );
nand ( n85370 , n407743 , n407744 );
buf ( n85371 , n85370 );
buf ( n407747 , n85371 );
nand ( n85373 , n85367 , n407747 );
buf ( n407749 , n85373 );
buf ( n407750 , n407749 );
buf ( n407751 , n369804 );
nand ( n407752 , n407750 , n407751 );
buf ( n407753 , n407752 );
buf ( n407754 , n407753 );
nand ( n407755 , n85362 , n407754 );
buf ( n407756 , n407755 );
buf ( n407757 , n407756 );
xor ( n407758 , n407720 , n407757 );
xor ( n407759 , n406424 , n406463 );
xor ( n407760 , n407759 , n406676 );
xor ( n85386 , n406685 , n84542 );
xor ( n407762 , n407760 , n85386 );
buf ( n407763 , n407762 );
xor ( n85389 , n406440 , n406443 );
xor ( n407765 , n85389 , n84183 );
xor ( n407766 , n406840 , n84537 );
xor ( n85392 , n407765 , n407766 );
buf ( n407768 , n85392 );
xor ( n407769 , n83909 , n406018 );
xor ( n85395 , n407769 , n406022 );
xor ( n407771 , n406647 , n406666 );
xor ( n85397 , n85395 , n407771 );
buf ( n407773 , n396499 );
buf ( n407774 , n394724 );
and ( n85400 , n407773 , n407774 );
buf ( n407776 , n394816 );
buf ( n407777 , n394730 );
and ( n85403 , n407776 , n407777 );
nor ( n85404 , n85400 , n85403 );
buf ( n407780 , n85404 );
buf ( n407781 , n407780 );
buf ( n407782 , n384414 );
or ( n85408 , n407781 , n407782 );
buf ( n407784 , n406696 );
buf ( n407785 , n395635 );
or ( n407786 , n407784 , n407785 );
nand ( n85412 , n85408 , n407786 );
buf ( n407788 , n85412 );
xor ( n85414 , n406586 , n406603 );
xor ( n85415 , n85414 , n406620 );
and ( n85416 , n407788 , n85415 );
buf ( n407792 , n384380 );
buf ( n407793 , n394840 );
and ( n85419 , n407792 , n407793 );
buf ( n407795 , n384386 );
buf ( n407796 , n395890 );
and ( n407797 , n407795 , n407796 );
nor ( n85423 , n85419 , n407797 );
buf ( n407799 , n85423 );
buf ( n407800 , n407799 );
buf ( n407801 , n394838 );
or ( n85427 , n407800 , n407801 );
buf ( n407803 , n406658 );
buf ( n407804 , n394835 );
or ( n407805 , n407803 , n407804 );
nand ( n85431 , n85427 , n407805 );
buf ( n407807 , n85431 );
xor ( n407808 , n406586 , n406603 );
xor ( n407809 , n407808 , n406620 );
and ( n85435 , n407807 , n407809 );
and ( n407811 , n407788 , n407807 );
or ( n85437 , n85416 , n85435 , n407811 );
xor ( n85438 , n85397 , n85437 );
xor ( n407814 , n406781 , n406798 );
xor ( n407815 , n407814 , n406821 );
buf ( n407816 , n407815 );
buf ( n407817 , n75451 );
buf ( n407818 , n384343 );
and ( n85444 , n407817 , n407818 );
buf ( n407820 , n396596 );
buf ( n407821 , n384089 );
and ( n85447 , n407820 , n407821 );
nor ( n85448 , n85444 , n85447 );
buf ( n407824 , n85448 );
buf ( n407825 , n407824 );
buf ( n407826 , n384354 );
or ( n85452 , n407825 , n407826 );
buf ( n407828 , n406713 );
buf ( n407829 , n384082 );
or ( n85455 , n407828 , n407829 );
nand ( n85456 , n85452 , n85455 );
buf ( n407832 , n85456 );
xor ( n85458 , n407816 , n407832 );
buf ( n407834 , n74644 );
buf ( n407835 , n394724 );
and ( n85461 , n407834 , n407835 );
buf ( n407837 , n395683 );
buf ( n407838 , n63434 );
and ( n407839 , n407837 , n407838 );
nor ( n407840 , n85461 , n407839 );
buf ( n407841 , n407840 );
buf ( n407842 , n407841 );
buf ( n407843 , n384414 );
or ( n407844 , n407842 , n407843 );
buf ( n407845 , n407780 );
buf ( n407846 , n395635 );
or ( n407847 , n407845 , n407846 );
nand ( n407848 , n407844 , n407847 );
buf ( n407849 , n407848 );
and ( n407850 , n85458 , n407849 );
and ( n407851 , n407816 , n407832 );
or ( n407852 , n407850 , n407851 );
buf ( n407853 , n407852 );
buf ( n407854 , n80468 );
buf ( n407855 , n406588 );
and ( n407856 , n407854 , n407855 );
buf ( n407857 , n401921 );
buf ( n407858 , n82201 );
and ( n407859 , n407857 , n407858 );
nor ( n407860 , n407856 , n407859 );
buf ( n85464 , n407860 );
buf ( n407862 , n85464 );
buf ( n407863 , n60313 );
or ( n85467 , n407862 , n407863 );
buf ( n407865 , n406789 );
buf ( n407866 , n380733 );
or ( n85470 , n407865 , n407866 );
nand ( n85471 , n85467 , n85470 );
buf ( n407869 , n85471 );
buf ( n407870 , n407869 );
buf ( n407871 , n380581 );
buf ( n407872 , n57789 );
buf ( n407873 , n81995 );
and ( n85477 , n407872 , n407873 );
buf ( n407875 , n403645 );
buf ( n407876 , n378470 );
and ( n407877 , n407875 , n407876 );
nor ( n85481 , n85477 , n407877 );
buf ( n407879 , n85481 );
buf ( n407880 , n407879 );
or ( n85484 , n407871 , n407880 );
buf ( n407882 , n406559 );
buf ( n407883 , n378476 );
or ( n407884 , n407882 , n407883 );
nand ( n85488 , n85484 , n407884 );
buf ( n85489 , n85488 );
buf ( n407887 , n85489 );
xor ( n85491 , n407870 , n407887 );
buf ( n407889 , n380581 );
buf ( n407890 , n57789 );
buf ( n407891 , n403772 );
and ( n407892 , n407890 , n407891 );
buf ( n407893 , n378470 );
buf ( n407894 , n403775 );
and ( n85498 , n407893 , n407894 );
nor ( n85499 , n407892 , n85498 );
buf ( n407897 , n85499 );
buf ( n407898 , n407897 );
or ( n407899 , n407889 , n407898 );
buf ( n407900 , n407879 );
buf ( n407901 , n378476 );
or ( n407902 , n407900 , n407901 );
nand ( n407903 , n407899 , n407902 );
buf ( n407904 , n407903 );
buf ( n407905 , n377030 );
buf ( n85509 , n376997 );
buf ( n407907 , n623 );
nor ( n407908 , n407905 , n85509 , n407907 );
buf ( n407909 , n407908 );
xor ( n85513 , n407904 , n407909 );
buf ( n407911 , n57800 );
buf ( n407912 , n405813 );
and ( n85516 , n407911 , n407912 );
buf ( n407914 , n378284 );
buf ( n407915 , n405816 );
and ( n407916 , n407914 , n407915 );
nor ( n85520 , n85516 , n407916 );
buf ( n85521 , n85520 );
buf ( n407919 , n85521 );
not ( n85523 , n407919 );
buf ( n85524 , n85523 );
buf ( n407922 , n85524 );
not ( n85526 , n407922 );
buf ( n407924 , n378280 );
not ( n85528 , n407924 );
or ( n407926 , n85526 , n85528 );
buf ( n407927 , n378262 );
buf ( n407928 , n406768 );
or ( n407929 , n407927 , n407928 );
nand ( n85533 , n407926 , n407929 );
buf ( n407931 , n85533 );
and ( n407932 , n85513 , n407931 );
and ( n407933 , n407904 , n407909 );
or ( n85537 , n407932 , n407933 );
buf ( n407935 , n85537 );
and ( n407936 , n85491 , n407935 );
and ( n85540 , n407870 , n407887 );
or ( n407938 , n407936 , n85540 );
buf ( n407939 , n407938 );
xor ( n85543 , n406567 , n406580 );
xor ( n407941 , n85543 , n406583 );
and ( n407942 , n407939 , n407941 );
buf ( n407943 , n400503 );
buf ( n407944 , n382835 );
and ( n85548 , n407943 , n407944 );
buf ( n407946 , n400509 );
buf ( n407947 , n62243 );
and ( n85551 , n407946 , n407947 );
nor ( n407949 , n85548 , n85551 );
buf ( n407950 , n407949 );
buf ( n407951 , n407950 );
buf ( n407952 , n382849 );
or ( n407953 , n407951 , n407952 );
buf ( n407954 , n406815 );
buf ( n407955 , n384157 );
or ( n407956 , n407954 , n407955 );
nand ( n407957 , n407953 , n407956 );
buf ( n407958 , n407957 );
buf ( n407959 , n407958 );
xor ( n407960 , n406744 , n406758 );
xor ( n85564 , n407960 , n406776 );
buf ( n407962 , n85564 );
buf ( n407963 , n407962 );
xor ( n407964 , n407959 , n407963 );
buf ( n407965 , n376924 );
buf ( n407966 , n376866 );
buf ( n407967 , n406746 );
and ( n85571 , n407966 , n407967 );
buf ( n407969 , n377030 );
buf ( n407970 , n406749 );
and ( n85574 , n407969 , n407970 );
nor ( n407972 , n85571 , n85574 );
buf ( n407973 , n407972 );
buf ( n407974 , n407973 );
or ( n407975 , n407965 , n407974 );
buf ( n407976 , n406736 );
buf ( n407977 , n56517 );
or ( n85581 , n407976 , n407977 );
nand ( n407979 , n407975 , n85581 );
buf ( n407980 , n407979 );
buf ( n407981 , n407980 );
buf ( n407982 , n56639 );
xor ( n407983 , n407981 , n407982 );
buf ( n407984 , n377003 );
buf ( n407985 , n623 );
not ( n85589 , n407985 );
buf ( n85590 , n85589 );
buf ( n407988 , n85590 );
nor ( n85592 , n407984 , n407988 );
buf ( n407990 , n85592 );
buf ( n85594 , n407990 );
buf ( n407992 , n380581 );
buf ( n407993 , n57789 );
buf ( n407994 , n403795 );
and ( n407995 , n407993 , n407994 );
buf ( n407996 , n378470 );
buf ( n407997 , n403798 );
and ( n407998 , n407996 , n407997 );
nor ( n407999 , n407995 , n407998 );
buf ( n408000 , n407999 );
buf ( n408001 , n408000 );
or ( n408002 , n407992 , n408001 );
buf ( n408003 , n407897 );
buf ( n408004 , n394774 );
or ( n408005 , n408003 , n408004 );
nand ( n408006 , n408002 , n408005 );
buf ( n408007 , n408006 );
buf ( n408008 , n408007 );
and ( n408009 , n85594 , n408008 );
buf ( n408010 , n408009 );
buf ( n408011 , n408010 );
and ( n85597 , n407983 , n408011 );
and ( n408013 , n407981 , n407982 );
or ( n408014 , n85597 , n408013 );
buf ( n408015 , n408014 );
buf ( n408016 , n408015 );
and ( n408017 , n407964 , n408016 );
and ( n408018 , n407959 , n407963 );
or ( n85602 , n408017 , n408018 );
buf ( n408020 , n85602 );
xor ( n408021 , n406567 , n406580 );
xor ( n85605 , n408021 , n406583 );
and ( n85606 , n408020 , n85605 );
and ( n85607 , n407939 , n408020 );
or ( n85608 , n407942 , n85606 , n85607 );
buf ( n408026 , n85608 );
xor ( n85610 , n407853 , n408026 );
xor ( n85611 , n406722 , n406726 );
xor ( n85612 , n85611 , n406826 );
buf ( n408030 , n85612 );
buf ( n408031 , n408030 );
and ( n85615 , n85610 , n408031 );
and ( n85616 , n407853 , n408026 );
or ( n85617 , n85615 , n85616 );
buf ( n408035 , n85617 );
and ( n85619 , n85438 , n408035 );
and ( n408037 , n85397 , n85437 );
or ( n85621 , n85619 , n408037 );
buf ( n408039 , n85621 );
xor ( n85623 , n407768 , n408039 );
xor ( n85624 , n406705 , n406831 );
xor ( n85625 , n85624 , n406836 );
buf ( n408043 , n85625 );
xor ( n408044 , n85397 , n85437 );
xor ( n85628 , n408044 , n408035 );
and ( n408046 , n408043 , n85628 );
buf ( n408047 , n73625 );
buf ( n408048 , n394840 );
and ( n85632 , n408047 , n408048 );
buf ( n408050 , n73631 );
buf ( n408051 , n395890 );
and ( n408052 , n408050 , n408051 );
nor ( n85636 , n85632 , n408052 );
buf ( n408054 , n85636 );
buf ( n408055 , n408054 );
buf ( n408056 , n394838 );
or ( n408057 , n408055 , n408056 );
buf ( n408058 , n407799 );
buf ( n408059 , n394835 );
or ( n85642 , n408058 , n408059 );
nand ( n85643 , n408057 , n85642 );
buf ( n408062 , n85643 );
buf ( n408063 , n408062 );
buf ( n408064 , n81950 );
buf ( n408065 , n406588 );
and ( n408066 , n408064 , n408065 );
buf ( n408067 , n403589 );
buf ( n408068 , n57983 );
and ( n85651 , n408067 , n408068 );
nor ( n85652 , n408066 , n85651 );
buf ( n408071 , n85652 );
buf ( n408072 , n408071 );
buf ( n408073 , n60313 );
or ( n408074 , n408072 , n408073 );
buf ( n408075 , n85464 );
buf ( n408076 , n380733 );
or ( n408077 , n408075 , n408076 );
nand ( n85660 , n408074 , n408077 );
buf ( n85661 , n85660 );
xor ( n408080 , n407904 , n407909 );
xor ( n85663 , n408080 , n407931 );
and ( n85664 , n85661 , n85663 );
buf ( n408083 , n407973 );
buf ( n408084 , n56517 );
or ( n408085 , n408083 , n408084 );
buf ( n408086 , n56623 );
nand ( n85669 , n408085 , n408086 );
buf ( n85670 , n85669 );
buf ( n408089 , n85670 );
buf ( n408090 , n378341 );
buf ( n408091 , n57800 );
buf ( n408092 , n406569 );
and ( n85675 , n408091 , n408092 );
buf ( n408094 , n378284 );
buf ( n408095 , n406572 );
and ( n85678 , n408094 , n408095 );
nor ( n85679 , n85675 , n85678 );
buf ( n408098 , n85679 );
buf ( n408099 , n408098 );
or ( n408100 , n408090 , n408099 );
buf ( n408101 , n378262 );
buf ( n408102 , n85521 );
or ( n85685 , n408101 , n408102 );
nand ( n85686 , n408100 , n85685 );
buf ( n408105 , n85686 );
buf ( n408106 , n408105 );
xor ( n408107 , n408089 , n408106 );
buf ( n408108 , n60313 );
buf ( n408109 , n406588 );
buf ( n408110 , n81995 );
and ( n85693 , n408109 , n408110 );
buf ( n408112 , n403645 );
buf ( n408113 , n63664 );
and ( n408114 , n408112 , n408113 );
nor ( n408115 , n85693 , n408114 );
buf ( n408116 , n408115 );
buf ( n408117 , n408116 );
or ( n408118 , n408108 , n408117 );
buf ( n408119 , n408071 );
buf ( n408120 , n380733 );
or ( n85703 , n408119 , n408120 );
nand ( n408122 , n408118 , n85703 );
buf ( n408123 , n408122 );
buf ( n408124 , n408123 );
and ( n408125 , n408107 , n408124 );
and ( n85708 , n408089 , n408106 );
or ( n85709 , n408125 , n85708 );
buf ( n408128 , n85709 );
xor ( n85711 , n407904 , n407909 );
xor ( n85712 , n85711 , n407931 );
and ( n85713 , n408128 , n85712 );
and ( n408132 , n85661 , n408128 );
or ( n85715 , n85664 , n85713 , n408132 );
buf ( n408134 , n85715 );
buf ( n408135 , n396615 );
buf ( n408136 , n384343 );
and ( n85719 , n408135 , n408136 );
buf ( n408138 , n396621 );
buf ( n408139 , n384089 );
and ( n85722 , n408138 , n408139 );
nor ( n85723 , n85719 , n85722 );
buf ( n408142 , n85723 );
buf ( n408143 , n408142 );
buf ( n408144 , n384354 );
or ( n85727 , n408143 , n408144 );
buf ( n408146 , n407824 );
buf ( n408147 , n384082 );
or ( n85730 , n408146 , n408147 );
nand ( n408149 , n85727 , n85730 );
buf ( n408150 , n408149 );
buf ( n408151 , n408150 );
xor ( n408152 , n408134 , n408151 );
xor ( n408153 , n407870 , n407887 );
xor ( n85736 , n408153 , n407935 );
buf ( n408155 , n85736 );
buf ( n408156 , n408155 );
and ( n408157 , n408152 , n408156 );
and ( n408158 , n408134 , n408151 );
or ( n85741 , n408157 , n408158 );
buf ( n408160 , n85741 );
buf ( n408161 , n408160 );
xor ( n85744 , n408063 , n408161 );
xor ( n85745 , n406567 , n406580 );
xor ( n85746 , n85745 , n406583 );
xor ( n85747 , n407939 , n408020 );
xor ( n85748 , n85746 , n85747 );
buf ( n408167 , n85748 );
and ( n85750 , n85744 , n408167 );
and ( n85751 , n408063 , n408161 );
or ( n408170 , n85750 , n85751 );
buf ( n408171 , n408170 );
xor ( n408172 , n406586 , n406603 );
xor ( n408173 , n408172 , n406620 );
xor ( n408174 , n407788 , n407807 );
xor ( n408175 , n408173 , n408174 );
xor ( n408176 , n408171 , n408175 );
xor ( n408177 , n407853 , n408026 );
xor ( n408178 , n408177 , n408031 );
buf ( n408179 , n408178 );
and ( n408180 , n408176 , n408179 );
and ( n408181 , n408171 , n408175 );
or ( n408182 , n408180 , n408181 );
xor ( n408183 , n85397 , n85437 );
xor ( n408184 , n408183 , n408035 );
and ( n408185 , n408182 , n408184 );
and ( n408186 , n408043 , n408182 );
or ( n408187 , n408046 , n408185 , n408186 );
buf ( n408188 , n408187 );
and ( n408189 , n85623 , n408188 );
and ( n408190 , n407768 , n408039 );
or ( n408191 , n408189 , n408190 );
buf ( n408192 , n408191 );
buf ( n408193 , n408192 );
xor ( n408194 , n407763 , n408193 );
buf ( n408195 , n377379 );
not ( n85755 , n408195 );
buf ( n85756 , n343001 );
buf ( n408198 , n85756 );
not ( n85758 , n408198 );
or ( n85759 , n85755 , n85758 );
not ( n408201 , n377379 );
buf ( n408202 , n408201 );
buf ( n408203 , n23037 );
nand ( n408204 , n408202 , n408203 );
buf ( n408205 , n408204 );
buf ( n408206 , n408205 );
nand ( n408207 , n85759 , n408206 );
buf ( n408208 , n408207 );
buf ( n408209 , n408208 );
not ( n408210 , n408209 );
buf ( n408211 , n368599 );
not ( n408212 , n408211 );
or ( n408213 , n408210 , n408212 );
buf ( n408214 , n406940 );
buf ( n408215 , n369444 );
nand ( n408216 , n408214 , n408215 );
buf ( n408217 , n408216 );
buf ( n408218 , n408217 );
nand ( n408219 , n408213 , n408218 );
buf ( n408220 , n408219 );
buf ( n408221 , n408220 );
and ( n85778 , n408194 , n408221 );
and ( n408223 , n407763 , n408193 );
or ( n408224 , n85778 , n408223 );
buf ( n408225 , n408224 );
buf ( n408226 , n408225 );
buf ( n408227 , n369809 );
not ( n85784 , n408227 );
buf ( n408229 , n407749 );
not ( n408230 , n408229 );
or ( n85787 , n85784 , n408230 );
buf ( n408232 , n393883 );
not ( n408233 , n408232 );
buf ( n408234 , n352314 );
not ( n408235 , n408234 );
buf ( n408236 , n408235 );
buf ( n408237 , n408236 );
not ( n408238 , n408237 );
or ( n85795 , n408233 , n408238 );
buf ( n408240 , n368656 );
buf ( n408241 , n369763 );
nand ( n85798 , n408240 , n408241 );
buf ( n85799 , n85798 );
buf ( n408244 , n85799 );
nand ( n85801 , n85795 , n408244 );
buf ( n408246 , n85801 );
buf ( n408247 , n408246 );
buf ( n408248 , n369804 );
nand ( n408249 , n408247 , n408248 );
buf ( n408250 , n408249 );
buf ( n408251 , n408250 );
nand ( n85808 , n85787 , n408251 );
buf ( n408253 , n85808 );
buf ( n408254 , n408253 );
xor ( n408255 , n408226 , n408254 );
buf ( n408256 , n369809 );
not ( n408257 , n408256 );
buf ( n408258 , n408246 );
not ( n85815 , n408258 );
or ( n408260 , n408257 , n85815 );
not ( n408261 , n393883 );
not ( n85818 , n48791 );
or ( n408263 , n408261 , n85818 );
buf ( n408264 , n48792 );
buf ( n408265 , n369763 );
nand ( n408266 , n408264 , n408265 );
buf ( n408267 , n408266 );
nand ( n408268 , n408263 , n408267 );
buf ( n408269 , n408268 );
buf ( n408270 , n369804 );
nand ( n85827 , n408269 , n408270 );
buf ( n408272 , n85827 );
buf ( n408273 , n408272 );
nand ( n408274 , n408260 , n408273 );
buf ( n408275 , n408274 );
buf ( n408276 , n408275 );
xor ( n85833 , n407763 , n408193 );
xor ( n408278 , n85833 , n408221 );
buf ( n408279 , n408278 );
buf ( n408280 , n408279 );
xor ( n408281 , n408276 , n408280 );
buf ( n408282 , n406346 );
not ( n85839 , n408282 );
buf ( n408284 , n406953 );
not ( n85841 , n408284 );
or ( n408286 , n85839 , n85841 );
buf ( n408287 , n405357 );
buf ( n408288 , n377779 );
nand ( n408289 , n408287 , n408288 );
buf ( n408290 , n408289 );
buf ( n408291 , n408290 );
nand ( n408292 , n408286 , n408291 );
buf ( n408293 , n408292 );
buf ( n408294 , n408293 );
not ( n408295 , n408294 );
buf ( n408296 , n406260 );
not ( n408297 , n408296 );
or ( n408298 , n408295 , n408297 );
buf ( n408299 , n406963 );
buf ( n408300 , n44915 );
nand ( n85846 , n408299 , n408300 );
buf ( n408302 , n85846 );
buf ( n408303 , n408302 );
nand ( n408304 , n408298 , n408303 );
buf ( n408305 , n408304 );
buf ( n408306 , n408305 );
and ( n408307 , n408281 , n408306 );
and ( n85853 , n408276 , n408280 );
or ( n85854 , n408307 , n85853 );
buf ( n408310 , n85854 );
buf ( n408311 , n408310 );
and ( n408312 , n408255 , n408311 );
and ( n85858 , n408226 , n408254 );
or ( n408314 , n408312 , n85858 );
buf ( n408315 , n408314 );
buf ( n408316 , n408315 );
and ( n408317 , n407758 , n408316 );
and ( n408318 , n407720 , n407757 );
or ( n85864 , n408317 , n408318 );
buf ( n408320 , n85864 );
buf ( n408321 , n408320 );
xor ( n408322 , n406421 , n406900 );
xor ( n408323 , n408322 , n406991 );
buf ( n408324 , n408323 );
buf ( n408325 , n408324 );
xor ( n85871 , n408321 , n408325 );
buf ( n408327 , n377122 );
not ( n408328 , n408327 );
buf ( n408329 , n396004 );
not ( n85875 , n408329 );
or ( n408331 , n408328 , n85875 );
buf ( n408332 , n76415 );
buf ( n408333 , n57463 );
nand ( n408334 , n408332 , n408333 );
buf ( n408335 , n408334 );
buf ( n408336 , n408335 );
nand ( n85882 , n408331 , n408336 );
buf ( n408338 , n85882 );
buf ( n408339 , n408338 );
not ( n85885 , n408339 );
buf ( n408341 , n365024 );
not ( n85887 , n408341 );
or ( n85888 , n85885 , n85887 );
buf ( n408344 , n407037 );
buf ( n408345 , n365108 );
nand ( n85891 , n408344 , n408345 );
buf ( n408347 , n85891 );
buf ( n408348 , n408347 );
nand ( n85894 , n85888 , n408348 );
buf ( n408350 , n85894 );
buf ( n408351 , n408350 );
and ( n85897 , n85871 , n408351 );
and ( n408353 , n408321 , n408325 );
or ( n85899 , n85897 , n408353 );
buf ( n408355 , n85899 );
buf ( n408356 , n408355 );
xor ( n408357 , n407692 , n408356 );
buf ( n408358 , n379260 );
not ( n408359 , n408358 );
buf ( n408360 , n379274 );
not ( n408361 , n408360 );
buf ( n408362 , n365344 );
not ( n408363 , n408362 );
or ( n408364 , n408361 , n408363 );
buf ( n408365 , n378736 );
buf ( n408366 , n379271 );
nand ( n408367 , n408365 , n408366 );
buf ( n408368 , n408367 );
buf ( n408369 , n408368 );
nand ( n408370 , n408364 , n408369 );
buf ( n408371 , n408370 );
buf ( n408372 , n408371 );
not ( n408373 , n408372 );
or ( n408374 , n408359 , n408373 );
buf ( n408375 , n379274 );
not ( n408376 , n408375 );
buf ( n408377 , n31194 );
not ( n408378 , n408377 );
or ( n408379 , n408376 , n408378 );
buf ( n408380 , n57233 );
buf ( n408381 , n379271 );
nand ( n408382 , n408380 , n408381 );
buf ( n408383 , n408382 );
buf ( n408384 , n408383 );
nand ( n408385 , n408379 , n408384 );
buf ( n408386 , n408385 );
buf ( n408387 , n408386 );
buf ( n408388 , n379962 );
nand ( n408389 , n408387 , n408388 );
buf ( n408390 , n408389 );
buf ( n408391 , n408390 );
nand ( n408392 , n408374 , n408391 );
buf ( n408393 , n408392 );
buf ( n408394 , n408393 );
and ( n408395 , n408357 , n408394 );
and ( n408396 , n407692 , n408356 );
or ( n85917 , n408395 , n408396 );
buf ( n408398 , n85917 );
buf ( n408399 , n408398 );
xor ( n85920 , n407688 , n408399 );
xor ( n85921 , n406238 , n84034 );
xor ( n408402 , n85921 , n406301 );
buf ( n408403 , n408402 );
buf ( n408404 , n408403 );
buf ( n408405 , n369809 );
not ( n408406 , n408405 );
buf ( n408407 , n406332 );
not ( n408408 , n408407 );
or ( n408409 , n408406 , n408408 );
buf ( n408410 , n407734 );
buf ( n408411 , n369804 );
nand ( n408412 , n408410 , n408411 );
buf ( n408413 , n408412 );
buf ( n408414 , n408413 );
nand ( n85933 , n408409 , n408414 );
buf ( n408416 , n85933 );
buf ( n408417 , n408416 );
xor ( n408418 , n408404 , n408417 );
and ( n85936 , n377757 , n394065 );
not ( n408420 , n377757 );
not ( n85938 , n400916 );
and ( n85939 , n408420 , n85938 );
or ( n408423 , n85936 , n85939 );
buf ( n408424 , n408423 );
not ( n408425 , n408424 );
buf ( n408426 , n45055 );
not ( n85944 , n408426 );
or ( n85945 , n408425 , n85944 );
buf ( n408429 , n365242 );
buf ( n408430 , n406356 );
nand ( n85948 , n408429 , n408430 );
buf ( n408432 , n85948 );
buf ( n408433 , n408432 );
nand ( n85951 , n85945 , n408433 );
buf ( n408435 , n85951 );
buf ( n408436 , n408435 );
xor ( n85954 , n408418 , n408436 );
buf ( n85955 , n85954 );
buf ( n408439 , n85955 );
buf ( n408440 , n397190 );
not ( n408441 , n408440 );
buf ( n408442 , n85274 );
not ( n408443 , n408442 );
or ( n85961 , n408441 , n408443 );
not ( n85962 , n377592 );
not ( n85963 , n364901 );
or ( n85964 , n85962 , n85963 );
nand ( n85965 , n364900 , n398363 );
nand ( n85966 , n85964 , n85965 );
buf ( n408450 , n85966 );
buf ( n408451 , n85179 );
nand ( n85969 , n408450 , n408451 );
buf ( n408453 , n85969 );
buf ( n408454 , n408453 );
nand ( n408455 , n85961 , n408454 );
buf ( n408456 , n408455 );
buf ( n408457 , n408456 );
xor ( n408458 , n408439 , n408457 );
buf ( n408459 , n377168 );
buf ( n408460 , n379515 );
nor ( n85978 , n408459 , n408460 );
buf ( n85979 , n85978 );
buf ( n408463 , n85979 );
and ( n408464 , n408458 , n408463 );
and ( n85982 , n408439 , n408457 );
or ( n408466 , n408464 , n85982 );
buf ( n408467 , n408466 );
buf ( n408468 , n408467 );
buf ( n85986 , n22619 );
buf ( n85987 , n58378 );
nand ( n85988 , n85986 , n85987 );
buf ( n85989 , n85988 );
nand ( n408473 , n380923 , n378843 );
nand ( n85991 , n85989 , n408473 );
buf ( n408475 , n85991 );
not ( n408476 , n408475 );
buf ( n408477 , n365725 );
not ( n85995 , n408477 );
or ( n85996 , n408476 , n85995 );
buf ( n408480 , n85244 );
buf ( n408481 , n56794 );
nand ( n85999 , n408480 , n408481 );
buf ( n408483 , n85999 );
buf ( n408484 , n408483 );
nand ( n86002 , n85996 , n408484 );
buf ( n408486 , n86002 );
buf ( n86004 , n408486 );
xor ( n86005 , n406918 , n406981 );
xor ( n408489 , n86005 , n406986 );
buf ( n408490 , n408489 );
buf ( n408491 , n408490 );
and ( n86009 , n377143 , n394065 );
not ( n408493 , n377143 );
and ( n86011 , n408493 , n65351 );
or ( n86012 , n86009 , n86011 );
buf ( n408496 , n86012 );
not ( n86014 , n408496 );
buf ( n408498 , n45055 );
not ( n408499 , n408498 );
or ( n86017 , n86014 , n408499 );
buf ( n408501 , n408423 );
buf ( n408502 , n365242 );
nand ( n86020 , n408501 , n408502 );
buf ( n408504 , n86020 );
buf ( n408505 , n408504 );
nand ( n408506 , n86017 , n408505 );
buf ( n408507 , n408506 );
buf ( n408508 , n408507 );
xor ( n408509 , n408491 , n408508 );
buf ( n408510 , n397190 );
not ( n408511 , n408510 );
buf ( n408512 , n85966 );
not ( n86027 , n408512 );
or ( n86028 , n408511 , n86027 );
buf ( n408515 , n377585 );
not ( n408516 , n408515 );
buf ( n408517 , n60751 );
not ( n86031 , n408517 );
or ( n86032 , n408516 , n86031 );
buf ( n408520 , n45802 );
buf ( n408521 , n377592 );
nand ( n86035 , n408520 , n408521 );
buf ( n408523 , n86035 );
buf ( n408524 , n408523 );
nand ( n86038 , n86032 , n408524 );
buf ( n408526 , n86038 );
buf ( n408527 , n408526 );
buf ( n408528 , n85179 );
nand ( n408529 , n408527 , n408528 );
buf ( n408530 , n408529 );
buf ( n408531 , n408530 );
nand ( n408532 , n86028 , n408531 );
buf ( n408533 , n408532 );
buf ( n408534 , n408533 );
and ( n86048 , n408509 , n408534 );
and ( n408536 , n408491 , n408508 );
or ( n86050 , n86048 , n408536 );
buf ( n408538 , n86050 );
buf ( n408539 , n408538 );
xor ( n86053 , n86004 , n408539 );
buf ( n408541 , n379260 );
not ( n408542 , n408541 );
buf ( n408543 , n408386 );
not ( n408544 , n408543 );
or ( n86058 , n408542 , n408544 );
buf ( n408546 , n379274 );
not ( n86060 , n408546 );
buf ( n408548 , n378543 );
not ( n408549 , n408548 );
or ( n86063 , n86060 , n408549 );
buf ( n408551 , n365490 );
buf ( n408552 , n379271 );
nand ( n86066 , n408551 , n408552 );
buf ( n408554 , n86066 );
buf ( n408555 , n408554 );
nand ( n408556 , n86063 , n408555 );
buf ( n408557 , n408556 );
buf ( n408558 , n408557 );
buf ( n408559 , n379962 );
nand ( n408560 , n408558 , n408559 );
buf ( n408561 , n408560 );
buf ( n408562 , n408561 );
nand ( n408563 , n86058 , n408562 );
buf ( n408564 , n408563 );
buf ( n408565 , n408564 );
and ( n86079 , n86053 , n408565 );
and ( n408567 , n86004 , n408539 );
or ( n86081 , n86079 , n408567 );
buf ( n408569 , n86081 );
buf ( n408570 , n408569 );
xor ( n86084 , n408468 , n408570 );
buf ( n408572 , n50782 );
buf ( n408573 , n378098 );
buf ( n408574 , n65993 );
and ( n86088 , n408573 , n408574 );
not ( n86089 , n408573 );
buf ( n408577 , n342656 );
and ( n86091 , n86089 , n408577 );
nor ( n86092 , n86088 , n86091 );
buf ( n408580 , n86092 );
buf ( n408581 , n408580 );
or ( n408582 , n408572 , n408581 );
buf ( n408583 , n56849 );
buf ( n408584 , n56687 );
nor ( n408585 , n408583 , n408584 );
buf ( n408586 , n408585 );
buf ( n408587 , n408586 );
buf ( n408588 , n386807 );
buf ( n408589 , n56687 );
and ( n86099 , n408588 , n408589 );
buf ( n408591 , n86099 );
buf ( n408592 , n408591 );
nor ( n408593 , n408587 , n408592 );
buf ( n408594 , n408593 );
buf ( n408595 , n408594 );
buf ( n408596 , n377268 );
or ( n408597 , n408595 , n408596 );
nand ( n408598 , n408582 , n408597 );
buf ( n408599 , n408598 );
buf ( n408600 , n408599 );
and ( n408601 , n86084 , n408600 );
and ( n408602 , n408468 , n408570 );
or ( n408603 , n408601 , n408602 );
buf ( n408604 , n408603 );
buf ( n408605 , n408604 );
and ( n408606 , n85920 , n408605 );
and ( n86102 , n407688 , n408399 );
or ( n408608 , n408606 , n86102 );
buf ( n408609 , n408608 );
buf ( n408610 , n408609 );
xor ( n408611 , n407611 , n408610 );
buf ( n408612 , n407267 );
not ( n408613 , n408612 );
buf ( n408614 , n407277 );
buf ( n408615 , n407254 );
and ( n408616 , n408614 , n408615 );
not ( n86112 , n408614 );
buf ( n408618 , n407257 );
and ( n408619 , n86112 , n408618 );
nor ( n408620 , n408616 , n408619 );
buf ( n408621 , n408620 );
buf ( n408622 , n408621 );
not ( n408623 , n408622 );
or ( n86119 , n408613 , n408623 );
buf ( n408625 , n408621 );
buf ( n408626 , n407267 );
or ( n408627 , n408625 , n408626 );
nand ( n86123 , n86119 , n408627 );
buf ( n408629 , n86123 );
buf ( n408630 , n408629 );
buf ( n408631 , n378098 );
buf ( n408632 , n46693 );
and ( n86128 , n408631 , n408632 );
not ( n408634 , n408631 );
buf ( n408635 , n364953 );
and ( n86131 , n408634 , n408635 );
nor ( n408637 , n86128 , n86131 );
buf ( n408638 , n408637 );
buf ( n408639 , n408638 );
not ( n408640 , n408639 );
buf ( n408641 , n363429 );
not ( n408642 , n408641 );
or ( n408643 , n408640 , n408642 );
buf ( n408644 , n377094 );
not ( n408645 , n408644 );
buf ( n408646 , n342718 );
not ( n408647 , n408646 );
or ( n86137 , n408645 , n408647 );
buf ( n408649 , n369497 );
buf ( n408650 , n56687 );
nand ( n86140 , n408649 , n408650 );
buf ( n408652 , n86140 );
buf ( n408653 , n408652 );
nand ( n86143 , n86137 , n408653 );
buf ( n408655 , n86143 );
buf ( n408656 , n408655 );
buf ( n408657 , n43261 );
nand ( n86147 , n408656 , n408657 );
buf ( n408659 , n86147 );
buf ( n408660 , n408659 );
nand ( n408661 , n408643 , n408660 );
buf ( n408662 , n408661 );
buf ( n408663 , n408662 );
xor ( n408664 , n408630 , n408663 );
buf ( n408665 , n85106 );
buf ( n408666 , n407393 );
and ( n86156 , n408665 , n408666 );
not ( n86157 , n408665 );
buf ( n408669 , n407390 );
and ( n408670 , n86157 , n408669 );
nor ( n86160 , n86156 , n408670 );
buf ( n86161 , n86160 );
buf ( n408673 , n86161 );
buf ( n408674 , n407416 );
and ( n408675 , n408673 , n408674 );
not ( n408676 , n408673 );
buf ( n408677 , n407413 );
and ( n408678 , n408676 , n408677 );
nor ( n408679 , n408675 , n408678 );
buf ( n408680 , n408679 );
buf ( n408681 , n408680 );
xor ( n408682 , n408664 , n408681 );
buf ( n408683 , n408682 );
buf ( n408684 , n408683 );
xor ( n86172 , n408611 , n408684 );
buf ( n408686 , n86172 );
buf ( n408687 , n408686 );
xor ( n408688 , n407516 , n408687 );
buf ( n408689 , n377094 );
not ( n86177 , n408689 );
buf ( n408691 , n388576 );
not ( n86179 , n408691 );
or ( n408693 , n86177 , n86179 );
buf ( n408694 , n378135 );
buf ( n408695 , n56687 );
nand ( n86183 , n408694 , n408695 );
buf ( n408697 , n86183 );
buf ( n408698 , n408697 );
nand ( n86186 , n408693 , n408698 );
buf ( n408700 , n86186 );
buf ( n408701 , n408700 );
not ( n408702 , n408701 );
buf ( n408703 , n399191 );
not ( n86191 , n408703 );
or ( n86192 , n408702 , n86191 );
buf ( n408706 , n407670 );
buf ( n408707 , n375920 );
nand ( n408708 , n408706 , n408707 );
buf ( n408709 , n408708 );
buf ( n408710 , n408709 );
nand ( n408711 , n86192 , n408710 );
buf ( n408712 , n408711 );
buf ( n408713 , n408712 );
buf ( n408714 , n58984 );
not ( n86202 , n408714 );
buf ( n408716 , n386102 );
not ( n408717 , n408716 );
or ( n86205 , n86202 , n408717 );
buf ( n408719 , n386093 );
buf ( n408720 , n58984 );
not ( n408721 , n408720 );
buf ( n408722 , n408721 );
buf ( n408723 , n408722 );
nand ( n408724 , n408719 , n408723 );
buf ( n408725 , n408724 );
buf ( n408726 , n408725 );
nand ( n408727 , n86205 , n408726 );
buf ( n408728 , n408727 );
buf ( n408729 , n408728 );
not ( n86217 , n408729 );
buf ( n408731 , n365024 );
not ( n408732 , n408731 );
or ( n408733 , n86217 , n408732 );
buf ( n408734 , n408338 );
buf ( n408735 , n365108 );
nand ( n86223 , n408734 , n408735 );
buf ( n408737 , n86223 );
buf ( n408738 , n408737 );
nand ( n86226 , n408733 , n408738 );
buf ( n408740 , n86226 );
buf ( n408741 , n408740 );
xor ( n408742 , n407720 , n407757 );
xor ( n408743 , n408742 , n408316 );
buf ( n408744 , n408743 );
buf ( n408745 , n408744 );
xor ( n86233 , n408741 , n408745 );
buf ( n408747 , n378135 );
buf ( n408748 , n380923 );
not ( n86236 , n408748 );
buf ( n408750 , n366646 );
not ( n408751 , n408750 );
or ( n86239 , n86236 , n408751 );
buf ( n408753 , n378098 );
nand ( n408754 , n86239 , n408753 );
buf ( n408755 , n408754 );
buf ( n408756 , n408755 );
buf ( n86244 , n22619 );
buf ( n408758 , n342590 );
nand ( n408759 , n86244 , n408758 );
buf ( n408760 , n408759 );
buf ( n408761 , n408760 );
and ( n408762 , n408747 , n408756 , n408761 );
buf ( n408763 , n408762 );
buf ( n408764 , n408763 );
and ( n408765 , n86233 , n408764 );
and ( n408766 , n408741 , n408745 );
or ( n86254 , n408765 , n408766 );
buf ( n408768 , n86254 );
buf ( n86256 , n408768 );
xor ( n86257 , n408713 , n86256 );
xor ( n408771 , n408321 , n408325 );
xor ( n86259 , n408771 , n408351 );
buf ( n408773 , n86259 );
buf ( n86261 , n408773 );
and ( n86262 , n86257 , n86261 );
and ( n86263 , n408713 , n86256 );
or ( n86264 , n86262 , n86263 );
buf ( n86265 , n86264 );
buf ( n408779 , n86265 );
xor ( n86267 , n407692 , n408356 );
xor ( n408781 , n86267 , n408394 );
buf ( n408782 , n408781 );
buf ( n408783 , n408782 );
xor ( n86271 , n408779 , n408783 );
xor ( n408785 , n408468 , n408570 );
xor ( n86273 , n408785 , n408600 );
buf ( n408787 , n86273 );
buf ( n408788 , n408787 );
and ( n408789 , n86271 , n408788 );
and ( n86277 , n408779 , n408783 );
or ( n408791 , n408789 , n86277 );
buf ( n408792 , n408791 );
buf ( n408793 , n408792 );
xor ( n408794 , n407688 , n408399 );
xor ( n408795 , n408794 , n408605 );
buf ( n408796 , n408795 );
buf ( n408797 , n408796 );
xor ( n408798 , n408793 , n408797 );
buf ( n408799 , n380356 );
not ( n86287 , n408799 );
and ( n86288 , n380368 , n31073 );
not ( n86289 , n380368 );
and ( n86290 , n86289 , n367576 );
or ( n408804 , n86288 , n86290 );
buf ( n408805 , n408804 );
not ( n86293 , n408805 );
or ( n408807 , n86287 , n86293 );
buf ( n408808 , n380368 );
not ( n86296 , n408808 );
buf ( n408810 , n351318 );
not ( n86298 , n408810 );
or ( n408812 , n86296 , n86298 );
buf ( n408813 , n364804 );
buf ( n408814 , n380364 );
nand ( n86302 , n408813 , n408814 );
buf ( n408816 , n86302 );
buf ( n408817 , n408816 );
nand ( n408818 , n408812 , n408817 );
buf ( n408819 , n408818 );
buf ( n408820 , n408819 );
buf ( n408821 , n380404 );
nand ( n408822 , n408820 , n408821 );
buf ( n408823 , n408822 );
buf ( n408824 , n408823 );
nand ( n408825 , n408807 , n408824 );
buf ( n408826 , n408825 );
buf ( n408827 , n408826 );
buf ( n408828 , n58923 );
not ( n86316 , n408828 );
buf ( n408830 , n379371 );
not ( n408831 , n408830 );
buf ( n408832 , n45125 );
not ( n86320 , n408832 );
or ( n408834 , n408831 , n86320 );
buf ( n408835 , n45113 );
buf ( n408836 , n407228 );
nand ( n86324 , n408835 , n408836 );
buf ( n408838 , n86324 );
buf ( n86326 , n408838 );
nand ( n86327 , n408834 , n86326 );
buf ( n86328 , n86327 );
buf ( n408842 , n86328 );
not ( n86330 , n408842 );
or ( n408844 , n86316 , n86330 );
buf ( n408845 , n379368 );
buf ( n408846 , n352212 );
and ( n408847 , n408845 , n408846 );
not ( n408848 , n408845 );
buf ( n408849 , n386359 );
and ( n408850 , n408848 , n408849 );
nor ( n408851 , n408847 , n408850 );
buf ( n408852 , n408851 );
buf ( n86340 , n408852 );
buf ( n86341 , n58867 );
nand ( n86342 , n86340 , n86341 );
buf ( n86343 , n86342 );
buf ( n408857 , n86343 );
nand ( n86345 , n408844 , n408857 );
buf ( n408859 , n86345 );
buf ( n408860 , n408859 );
xor ( n408861 , n408827 , n408860 );
not ( n86349 , n379890 );
buf ( n408863 , n379838 );
not ( n86351 , n408863 );
buf ( n408865 , n386837 );
not ( n408866 , n408865 );
or ( n86354 , n86351 , n408866 );
buf ( n408868 , n32202 );
buf ( n86356 , n398741 );
nand ( n408870 , n408868 , n86356 );
buf ( n408871 , n408870 );
buf ( n408872 , n408871 );
nand ( n408873 , n86354 , n408872 );
buf ( n408874 , n408873 );
not ( n86362 , n408874 );
or ( n408876 , n86349 , n86362 );
buf ( n408877 , n379838 );
not ( n86365 , n408877 );
buf ( n408879 , n382496 );
not ( n408880 , n408879 );
or ( n408881 , n86365 , n408880 );
buf ( n408882 , n378736 );
buf ( n408883 , n398741 );
nand ( n408884 , n408882 , n408883 );
buf ( n408885 , n408884 );
buf ( n408886 , n408885 );
nand ( n408887 , n408881 , n408886 );
buf ( n408888 , n408887 );
buf ( n408889 , n408888 );
buf ( n408890 , n379916 );
nand ( n408891 , n408889 , n408890 );
buf ( n408892 , n408891 );
nand ( n86380 , n408876 , n408892 );
nand ( n408894 , n84665 , n406978 , n84613 );
not ( n408895 , n84634 );
nand ( n86383 , n408895 , n84665 );
not ( n86384 , n84665 );
nor ( n86385 , n406978 , n84614 );
nand ( n86386 , n86384 , n86385 );
nand ( n86387 , n86384 , n84614 , n406978 );
nand ( n408901 , n408894 , n86383 , n86386 , n86387 );
buf ( n408902 , n408901 );
and ( n86390 , n377757 , n396401 );
not ( n408904 , n377757 );
and ( n86392 , n408904 , n80732 );
or ( n408906 , n86390 , n86392 );
buf ( n408907 , n408906 );
not ( n86395 , n408907 );
buf ( n408909 , n45012 );
not ( n408910 , n408909 );
or ( n86398 , n86395 , n408910 );
buf ( n408912 , n407704 );
buf ( n408913 , n365149 );
nand ( n408914 , n408912 , n408913 );
buf ( n408915 , n408914 );
buf ( n408916 , n408915 );
nand ( n86404 , n86398 , n408916 );
buf ( n408918 , n86404 );
buf ( n408919 , n408918 );
xor ( n408920 , n408902 , n408919 );
xor ( n408921 , n408226 , n408254 );
xor ( n408922 , n408921 , n408311 );
buf ( n408923 , n408922 );
buf ( n408924 , n408923 );
and ( n86412 , n408920 , n408924 );
and ( n408926 , n408902 , n408919 );
or ( n408927 , n86412 , n408926 );
buf ( n408928 , n408927 );
buf ( n408929 , n408928 );
not ( n408930 , n397190 );
not ( n86418 , n408526 );
or ( n86419 , n408930 , n86418 );
buf ( n408933 , n377584 );
not ( n408934 , n408933 );
buf ( n408935 , n402185 );
not ( n86423 , n408935 );
or ( n408937 , n408934 , n86423 );
buf ( n86425 , n377592 );
buf ( n408939 , n31311 );
nand ( n408940 , n86425 , n408939 );
buf ( n408941 , n408940 );
buf ( n408942 , n408941 );
nand ( n86430 , n408937 , n408942 );
buf ( n408944 , n86430 );
buf ( n408945 , n408944 );
buf ( n408946 , n85179 );
nand ( n86434 , n408945 , n408946 );
buf ( n408948 , n86434 );
nand ( n408949 , n86419 , n408948 );
not ( n86437 , n45055 );
buf ( n408951 , n377122 );
not ( n86439 , n408951 );
buf ( n408953 , n400916 );
not ( n408954 , n408953 );
or ( n86442 , n86439 , n408954 );
buf ( n408956 , n342879 );
buf ( n408957 , n57463 );
nand ( n86445 , n408956 , n408957 );
buf ( n408959 , n86445 );
buf ( n408960 , n408959 );
nand ( n86448 , n86442 , n408960 );
buf ( n408962 , n86448 );
not ( n86450 , n408962 );
or ( n86451 , n86437 , n86450 );
buf ( n408965 , n86012 );
buf ( n408966 , n365242 );
nand ( n86454 , n408965 , n408966 );
buf ( n408968 , n86454 );
nand ( n408969 , n86451 , n408968 );
xor ( n86457 , n408949 , n408969 );
buf ( n408971 , n397190 );
not ( n408972 , n408971 );
buf ( n408973 , n408944 );
not ( n86461 , n408973 );
or ( n86462 , n408972 , n86461 );
buf ( n408976 , n398363 );
not ( n408977 , n408976 );
buf ( n408978 , n365384 );
not ( n86466 , n408978 );
or ( n408980 , n408977 , n86466 );
buf ( n408981 , n84042 );
buf ( n408982 , n377592 );
nand ( n408983 , n408981 , n408982 );
buf ( n408984 , n408983 );
buf ( n408985 , n408984 );
nand ( n408986 , n408980 , n408985 );
buf ( n408987 , n408986 );
buf ( n408988 , n408987 );
buf ( n408989 , n85179 );
nand ( n408990 , n408988 , n408989 );
buf ( n408991 , n408990 );
buf ( n408992 , n408991 );
nand ( n86480 , n86462 , n408992 );
buf ( n86481 , n86480 );
not ( n408995 , n86481 );
and ( n408996 , n377143 , n396401 );
not ( n86484 , n377143 );
buf ( n408998 , n402190 );
and ( n408999 , n86484 , n408998 );
or ( n86487 , n408996 , n408999 );
buf ( n409001 , n86487 );
not ( n409002 , n409001 );
buf ( n409003 , n402201 );
not ( n409004 , n409003 );
or ( n409005 , n409002 , n409004 );
buf ( n409006 , n408906 );
buf ( n409007 , n365149 );
nand ( n409008 , n409006 , n409007 );
buf ( n409009 , n409008 );
buf ( n409010 , n409009 );
nand ( n409011 , n409005 , n409010 );
buf ( n409012 , n409011 );
not ( n409013 , n409012 );
or ( n86501 , n408995 , n409013 );
buf ( n409015 , n86481 );
buf ( n409016 , n409012 );
or ( n86504 , n409015 , n409016 );
buf ( n409018 , n377349 );
not ( n409019 , n409018 );
buf ( n409020 , n409019 );
buf ( n409021 , n409020 );
not ( n409022 , n85756 );
buf ( n409023 , n409022 );
and ( n86511 , n409021 , n409023 );
not ( n86512 , n409021 );
buf ( n409026 , n44906 );
and ( n86514 , n86512 , n409026 );
nor ( n409028 , n86511 , n86514 );
buf ( n409029 , n409028 );
buf ( n409030 , n409029 );
not ( n409031 , n409030 );
buf ( n409032 , n368599 );
not ( n86520 , n409032 );
or ( n409034 , n409031 , n86520 );
buf ( n409035 , n408208 );
buf ( n409036 , n369444 );
nand ( n86524 , n409035 , n409036 );
buf ( n409038 , n86524 );
buf ( n409039 , n409038 );
nand ( n86527 , n409034 , n409039 );
buf ( n409041 , n86527 );
buf ( n409042 , n409041 );
not ( n409043 , n409042 );
buf ( n409044 , n377754 );
not ( n409045 , n409044 );
buf ( n409046 , n406246 );
not ( n86534 , n409046 );
or ( n409048 , n409045 , n86534 );
buf ( n409049 , n406950 );
buf ( n409050 , n377754 );
not ( n409051 , n409050 );
buf ( n409052 , n409051 );
buf ( n409053 , n409052 );
nand ( n409054 , n409049 , n409053 );
buf ( n409055 , n409054 );
buf ( n409056 , n409055 );
nand ( n86544 , n409048 , n409056 );
buf ( n86545 , n86544 );
buf ( n409059 , n86545 );
not ( n86547 , n409059 );
buf ( n409061 , n406260 );
not ( n409062 , n409061 );
or ( n86550 , n86547 , n409062 );
buf ( n409064 , n408293 );
buf ( n409065 , n44915 );
nand ( n86553 , n409064 , n409065 );
buf ( n409067 , n86553 );
buf ( n409068 , n409067 );
nand ( n86556 , n86550 , n409068 );
buf ( n86557 , n86556 );
buf ( n409071 , n86557 );
not ( n86559 , n409071 );
or ( n86560 , n409043 , n86559 );
buf ( n409074 , n86557 );
buf ( n409075 , n409041 );
or ( n86563 , n409074 , n409075 );
xor ( n409077 , n407768 , n408039 );
xor ( n409078 , n409077 , n408188 );
buf ( n409079 , n409078 );
buf ( n409080 , n409079 );
nand ( n409081 , n86563 , n409080 );
buf ( n409082 , n409081 );
buf ( n409083 , n409082 );
nand ( n409084 , n86560 , n409083 );
buf ( n409085 , n409084 );
buf ( n409086 , n409085 );
nand ( n409087 , n86504 , n409086 );
buf ( n409088 , n409087 );
nand ( n86576 , n86501 , n409088 );
and ( n409090 , n86457 , n86576 );
and ( n86578 , n408949 , n408969 );
or ( n409092 , n409090 , n86578 );
buf ( n409093 , n409092 );
xor ( n409094 , n408929 , n409093 );
buf ( n409095 , n379260 );
not ( n86583 , n409095 );
buf ( n409097 , n408557 );
not ( n86585 , n409097 );
or ( n86586 , n86583 , n86585 );
buf ( n409100 , n379274 );
not ( n86588 , n409100 );
buf ( n409102 , n381266 );
not ( n86590 , n409102 );
or ( n86591 , n86588 , n86590 );
buf ( n409105 , n351160 );
buf ( n409106 , n379271 );
nand ( n86594 , n409105 , n409106 );
buf ( n409108 , n86594 );
buf ( n409109 , n409108 );
nand ( n409110 , n86591 , n409109 );
buf ( n409111 , n409110 );
buf ( n409112 , n409111 );
buf ( n409113 , n379962 );
nand ( n86601 , n409112 , n409113 );
buf ( n409115 , n86601 );
buf ( n409116 , n409115 );
nand ( n86604 , n86586 , n409116 );
buf ( n86605 , n86604 );
buf ( n409119 , n86605 );
and ( n86607 , n409094 , n409119 );
and ( n409121 , n408929 , n409093 );
or ( n409122 , n86607 , n409121 );
buf ( n409123 , n409122 );
xor ( n409124 , n86380 , n409123 );
xor ( n409125 , n86004 , n408539 );
xor ( n86613 , n409125 , n408565 );
buf ( n409127 , n86613 );
and ( n409128 , n409124 , n409127 );
and ( n409129 , n86380 , n409123 );
or ( n86617 , n409128 , n409129 );
buf ( n409131 , n86617 );
and ( n86619 , n408861 , n409131 );
and ( n86620 , n408827 , n408860 );
or ( n409134 , n86619 , n86620 );
buf ( n409135 , n409134 );
buf ( n409136 , n409135 );
and ( n409137 , n408798 , n409136 );
and ( n409138 , n408793 , n408797 );
or ( n86626 , n409137 , n409138 );
buf ( n409140 , n86626 );
buf ( n409141 , n409140 );
and ( n86629 , n408688 , n409141 );
and ( n409143 , n407516 , n408687 );
or ( n86631 , n86629 , n409143 );
buf ( n409145 , n86631 );
buf ( n409146 , n409145 );
xor ( n409147 , n407512 , n409146 );
xor ( n409148 , n407611 , n408610 );
and ( n86636 , n409148 , n408684 );
and ( n409150 , n407611 , n408610 );
or ( n409151 , n86636 , n409150 );
buf ( n409152 , n409151 );
buf ( n409153 , n409152 );
xor ( n86641 , n408630 , n408663 );
and ( n409155 , n86641 , n408681 );
and ( n409156 , n408630 , n408663 );
or ( n86644 , n409155 , n409156 );
buf ( n409158 , n86644 );
buf ( n409159 , n409158 );
xor ( n409160 , n408404 , n408417 );
and ( n86648 , n409160 , n408436 );
and ( n409162 , n408404 , n408417 );
or ( n86650 , n86648 , n409162 );
buf ( n409164 , n86650 );
buf ( n409165 , n409164 );
xor ( n409166 , n406306 , n406340 );
xor ( n86654 , n409166 , n406369 );
buf ( n409168 , n86654 );
buf ( n409169 , n409168 );
xor ( n409170 , n409165 , n409169 );
buf ( n409171 , n56849 );
buf ( n409172 , n366380 );
not ( n409173 , n409172 );
buf ( n409174 , n378138 );
not ( n86662 , n409174 );
or ( n409176 , n409173 , n86662 );
buf ( n409177 , n378098 );
nand ( n409178 , n409176 , n409177 );
buf ( n409179 , n409178 );
buf ( n409180 , n409179 );
buf ( n409181 , n378135 );
buf ( n409182 , n342759 );
nand ( n409183 , n409181 , n409182 );
buf ( n409184 , n409183 );
buf ( n409185 , n409184 );
and ( n86673 , n409171 , n409180 , n409185 );
buf ( n409187 , n86673 );
buf ( n409188 , n409187 );
and ( n86676 , n409170 , n409188 );
and ( n86677 , n409165 , n409169 );
or ( n86678 , n86676 , n86677 );
buf ( n409192 , n86678 );
buf ( n409193 , n409192 );
buf ( n409194 , n379260 );
not ( n86682 , n409194 );
buf ( n409196 , n379274 );
not ( n86684 , n409196 );
buf ( n409198 , n386837 );
not ( n86686 , n409198 );
or ( n86687 , n86684 , n86686 );
buf ( n409201 , n32202 );
buf ( n409202 , n379271 );
nand ( n86690 , n409201 , n409202 );
buf ( n409204 , n86690 );
buf ( n409205 , n409204 );
nand ( n86693 , n86687 , n409205 );
buf ( n409207 , n86693 );
buf ( n409208 , n409207 );
not ( n86696 , n409208 );
or ( n409210 , n86682 , n86696 );
buf ( n409211 , n408371 );
buf ( n409212 , n379962 );
nand ( n409213 , n409211 , n409212 );
buf ( n409214 , n409213 );
buf ( n409215 , n409214 );
nand ( n409216 , n409210 , n409215 );
buf ( n409217 , n409216 );
buf ( n409218 , n409217 );
xor ( n409219 , n409193 , n409218 );
buf ( n409220 , n50782 );
buf ( n409221 , n408594 );
or ( n409222 , n409220 , n409221 );
buf ( n86710 , n377068 );
not ( n86711 , n86710 );
buf ( n86712 , n396289 );
not ( n86713 , n86712 );
or ( n86714 , n86711 , n86713 );
buf ( n409228 , n56849 );
buf ( n409229 , n377071 );
nand ( n409230 , n409228 , n409229 );
buf ( n409231 , n409230 );
buf ( n409232 , n409231 );
nand ( n86720 , n86714 , n409232 );
buf ( n409234 , n86720 );
buf ( n409235 , n409234 );
not ( n409236 , n409235 );
buf ( n409237 , n409236 );
buf ( n409238 , n409237 );
buf ( n409239 , n386027 );
or ( n409240 , n409238 , n409239 );
nand ( n86728 , n409222 , n409240 );
buf ( n86729 , n86728 );
buf ( n409243 , n86729 );
and ( n86731 , n409219 , n409243 );
and ( n409245 , n409193 , n409218 );
or ( n409246 , n86731 , n409245 );
buf ( n409247 , n409246 );
buf ( n409248 , n409247 );
buf ( n409249 , n379890 );
not ( n409250 , n409249 );
buf ( n409251 , n405711 );
not ( n409252 , n409251 );
or ( n409253 , n409250 , n409252 );
buf ( n409254 , n407583 );
buf ( n409255 , n379916 );
nand ( n409256 , n409254 , n409255 );
buf ( n409257 , n409256 );
buf ( n409258 , n409257 );
nand ( n86746 , n409253 , n409258 );
buf ( n409260 , n86746 );
buf ( n409261 , n409260 );
xor ( n409262 , n409248 , n409261 );
xor ( n86750 , n407529 , n407533 );
and ( n86751 , n86750 , n407561 );
and ( n409265 , n407529 , n407533 );
or ( n86753 , n86751 , n409265 );
buf ( n409267 , n86753 );
buf ( n409268 , n409267 );
buf ( n409269 , n409234 );
not ( n409270 , n409269 );
buf ( n409271 , n366399 );
not ( n409272 , n409271 );
or ( n409273 , n409270 , n409272 );
buf ( n409274 , n85122 );
not ( n86762 , n409274 );
buf ( n409276 , n366428 );
nand ( n409277 , n86762 , n409276 );
buf ( n409278 , n409277 );
buf ( n409279 , n409278 );
nand ( n409280 , n409273 , n409279 );
buf ( n409281 , n409280 );
buf ( n409282 , n409281 );
xor ( n409283 , n409268 , n409282 );
buf ( n409284 , n379263 );
not ( n409285 , n409284 );
buf ( n409286 , n85009 );
not ( n86774 , n409286 );
or ( n86775 , n409285 , n86774 );
buf ( n409289 , n409207 );
buf ( n409290 , n379299 );
nand ( n409291 , n409289 , n409290 );
buf ( n409292 , n409291 );
buf ( n409293 , n409292 );
nand ( n86781 , n86775 , n409293 );
buf ( n409295 , n86781 );
buf ( n409296 , n409295 );
xor ( n86784 , n409283 , n409296 );
buf ( n409298 , n86784 );
buf ( n86786 , n409298 );
and ( n86787 , n409262 , n86786 );
and ( n409301 , n409248 , n409261 );
or ( n409302 , n86787 , n409301 );
buf ( n409303 , n409302 );
buf ( n409304 , n409303 );
xor ( n86792 , n409159 , n409304 );
buf ( n409306 , n408655 );
not ( n86794 , n409306 );
buf ( n409308 , n363429 );
not ( n86796 , n409308 );
or ( n86797 , n86794 , n86796 );
buf ( n409311 , n46693 );
not ( n86799 , n409311 );
buf ( n409313 , n377071 );
not ( n86801 , n409313 );
and ( n409315 , n86799 , n86801 );
buf ( n409316 , n46693 );
buf ( n409317 , n377071 );
and ( n86805 , n409316 , n409317 );
nor ( n86806 , n409315 , n86805 );
buf ( n409320 , n86806 );
buf ( n409321 , n409320 );
not ( n409322 , n409321 );
buf ( n409323 , n58231 );
nand ( n86811 , n409322 , n409323 );
buf ( n409325 , n86811 );
buf ( n409326 , n409325 );
nand ( n86814 , n86797 , n409326 );
buf ( n409328 , n86814 );
buf ( n86816 , n409328 );
not ( n86817 , n405404 );
not ( n86818 , n86817 );
not ( n409332 , n405295 );
not ( n409333 , n405282 );
not ( n86821 , n409333 );
or ( n86822 , n409332 , n86821 );
not ( n409336 , n405295 );
nand ( n409337 , n409336 , n405282 );
nand ( n86825 , n86822 , n409337 );
not ( n409339 , n86825 );
or ( n409340 , n86818 , n409339 );
or ( n86828 , n86817 , n86825 );
nand ( n409342 , n409340 , n86828 );
buf ( n409343 , n409342 );
buf ( n409344 , n397190 );
not ( n86832 , n409344 );
buf ( n409346 , n404742 );
not ( n86834 , n409346 );
or ( n86835 , n86832 , n86834 );
buf ( n409349 , n85179 );
buf ( n409350 , n85025 );
nand ( n86838 , n409349 , n409350 );
buf ( n409352 , n86838 );
buf ( n409353 , n409352 );
nand ( n409354 , n86835 , n409353 );
buf ( n409355 , n409354 );
buf ( n409356 , n409355 );
xor ( n86844 , n409343 , n409356 );
xor ( n409358 , n406179 , n406204 );
and ( n409359 , n409358 , n406230 );
and ( n86847 , n406179 , n406204 );
or ( n409361 , n409359 , n86847 );
buf ( n409362 , n409361 );
buf ( n409363 , n409362 );
xor ( n409364 , n86844 , n409363 );
buf ( n409365 , n409364 );
buf ( n409366 , n409365 );
xor ( n409367 , n86816 , n409366 );
xor ( n409368 , n409268 , n409282 );
and ( n86856 , n409368 , n409296 );
and ( n409370 , n409268 , n409282 );
or ( n409371 , n86856 , n409370 );
buf ( n409372 , n409371 );
buf ( n409373 , n409372 );
xor ( n409374 , n409367 , n409373 );
buf ( n409375 , n409374 );
buf ( n409376 , n409375 );
xor ( n409377 , n86792 , n409376 );
buf ( n409378 , n409377 );
buf ( n409379 , n409378 );
xor ( n409380 , n409153 , n409379 );
xor ( n409381 , n407100 , n407105 );
xor ( n409382 , n409381 , n407135 );
buf ( n409383 , n409382 );
buf ( n409384 , n409383 );
buf ( n409385 , n58923 );
not ( n86873 , n409385 );
buf ( n409387 , n407234 );
not ( n86875 , n409387 );
or ( n409389 , n86873 , n86875 );
buf ( n409390 , n86328 );
buf ( n409391 , n58867 );
nand ( n86879 , n409390 , n409391 );
buf ( n409393 , n86879 );
buf ( n409394 , n409393 );
nand ( n409395 , n409389 , n409394 );
buf ( n409396 , n409395 );
buf ( n409397 , n409396 );
xor ( n86885 , n409384 , n409397 );
xor ( n409399 , n409193 , n409218 );
xor ( n86887 , n409399 , n409243 );
buf ( n409401 , n86887 );
buf ( n409402 , n409401 );
and ( n409403 , n86885 , n409402 );
and ( n86891 , n409384 , n409397 );
or ( n409405 , n409403 , n86891 );
buf ( n409406 , n409405 );
buf ( n409407 , n409406 );
xor ( n409408 , n409248 , n409261 );
xor ( n409409 , n409408 , n86786 );
buf ( n409410 , n409409 );
buf ( n409411 , n409410 );
xor ( n409412 , n409407 , n409411 );
buf ( n409413 , n379890 );
not ( n86901 , n409413 );
buf ( n409415 , n407598 );
not ( n409416 , n409415 );
or ( n86904 , n86901 , n409416 );
buf ( n409418 , n408874 );
buf ( n409419 , n379916 );
nand ( n86907 , n409418 , n409419 );
buf ( n409421 , n86907 );
buf ( n409422 , n409421 );
nand ( n86910 , n86904 , n409422 );
buf ( n409424 , n86910 );
buf ( n409425 , n409424 );
xor ( n86913 , n409165 , n409169 );
xor ( n86914 , n86913 , n409188 );
buf ( n409428 , n86914 );
buf ( n409429 , n409428 );
xor ( n86917 , n409425 , n409429 );
xor ( n409431 , n407632 , n407657 );
xor ( n409432 , n409431 , n407683 );
buf ( n409433 , n409432 );
buf ( n409434 , n409433 );
and ( n86922 , n86917 , n409434 );
and ( n409436 , n409425 , n409429 );
or ( n86924 , n86922 , n409436 );
buf ( n409438 , n86924 );
buf ( n409439 , n409438 );
xor ( n86927 , n407564 , n407568 );
xor ( n86928 , n86927 , n407606 );
buf ( n409442 , n86928 );
buf ( n409443 , n409442 );
xor ( n409444 , n409439 , n409443 );
buf ( n409445 , n380404 );
not ( n86933 , n409445 );
buf ( n409447 , n408804 );
not ( n409448 , n409447 );
or ( n86936 , n86933 , n409448 );
buf ( n409450 , n407210 );
buf ( n409451 , n380356 );
nand ( n86939 , n409450 , n409451 );
buf ( n86940 , n86939 );
buf ( n409454 , n86940 );
nand ( n86942 , n86936 , n409454 );
buf ( n409456 , n86942 );
buf ( n409457 , n409456 );
and ( n86945 , n409444 , n409457 );
and ( n86946 , n409439 , n409443 );
or ( n409460 , n86945 , n86946 );
buf ( n409461 , n409460 );
buf ( n409462 , n409461 );
and ( n86950 , n409412 , n409462 );
and ( n86951 , n409407 , n409411 );
or ( n409465 , n86950 , n86951 );
buf ( n409466 , n409465 );
buf ( n409467 , n409466 );
xor ( n409468 , n409380 , n409467 );
buf ( n409469 , n409468 );
buf ( n409470 , n409469 );
xor ( n409471 , n409147 , n409470 );
buf ( n409472 , n409471 );
buf ( n409473 , n409472 );
xor ( n409474 , n409407 , n409411 );
xor ( n86962 , n409474 , n409462 );
buf ( n86963 , n86962 );
buf ( n409477 , n86963 );
xor ( n86965 , n409384 , n409397 );
xor ( n409479 , n86965 , n409402 );
buf ( n409480 , n409479 );
buf ( n409481 , n409480 );
xor ( n86969 , n409425 , n409429 );
xor ( n86970 , n86969 , n409434 );
buf ( n409484 , n86970 );
buf ( n409485 , n409484 );
xor ( n86973 , n408439 , n408457 );
xor ( n86974 , n86973 , n408463 );
buf ( n409488 , n86974 );
buf ( n409489 , n409488 );
buf ( n409490 , n58923 );
not ( n86978 , n409490 );
buf ( n409492 , n408852 );
not ( n409493 , n409492 );
or ( n409494 , n86978 , n409493 );
buf ( n409495 , n379368 );
buf ( n409496 , n31260 );
and ( n86984 , n409495 , n409496 );
not ( n86985 , n409495 );
buf ( n409499 , n80834 );
and ( n409500 , n86985 , n409499 );
nor ( n86988 , n86984 , n409500 );
buf ( n409502 , n86988 );
buf ( n409503 , n409502 );
buf ( n409504 , n379353 );
nand ( n409505 , n409503 , n409504 );
buf ( n409506 , n409505 );
buf ( n409507 , n409506 );
nand ( n409508 , n409494 , n409507 );
buf ( n409509 , n409508 );
buf ( n409510 , n409509 );
xor ( n409511 , n409489 , n409510 );
buf ( n409512 , n378098 );
buf ( n409513 , n375901 );
and ( n409514 , n409512 , n409513 );
not ( n409515 , n409512 );
buf ( n409516 , n366659 );
and ( n409517 , n409515 , n409516 );
nor ( n87005 , n409514 , n409517 );
buf ( n409519 , n87005 );
buf ( n409520 , n409519 );
not ( n409521 , n409520 );
buf ( n409522 , n375896 );
not ( n409523 , n409522 );
or ( n409524 , n409521 , n409523 );
buf ( n409525 , n408700 );
buf ( n409526 , n375920 );
nand ( n409527 , n409525 , n409526 );
buf ( n409528 , n409527 );
buf ( n409529 , n409528 );
nand ( n409530 , n409524 , n409529 );
buf ( n409531 , n409530 );
buf ( n409532 , n409531 );
xor ( n409533 , n408741 , n408745 );
xor ( n87021 , n409533 , n408764 );
buf ( n409535 , n87021 );
buf ( n409536 , n409535 );
xor ( n409537 , n409532 , n409536 );
buf ( n409538 , n379890 );
not ( n87026 , n409538 );
buf ( n409540 , n408888 );
not ( n87028 , n409540 );
or ( n87029 , n87026 , n87028 );
buf ( n409543 , n379838 );
not ( n409544 , n409543 );
buf ( n409545 , n351228 );
not ( n87033 , n409545 );
or ( n409547 , n409544 , n87033 );
buf ( n409548 , n57233 );
buf ( n87036 , n398741 );
nand ( n87037 , n409548 , n87036 );
buf ( n87038 , n87037 );
buf ( n87039 , n87038 );
nand ( n87040 , n409547 , n87039 );
buf ( n87041 , n87040 );
buf ( n409555 , n87041 );
buf ( n409556 , n379916 );
nand ( n409557 , n409555 , n409556 );
buf ( n409558 , n409557 );
buf ( n409559 , n409558 );
nand ( n87047 , n87029 , n409559 );
buf ( n409561 , n87047 );
buf ( n409562 , n409561 );
and ( n409563 , n409537 , n409562 );
and ( n409564 , n409532 , n409536 );
or ( n87052 , n409563 , n409564 );
buf ( n409566 , n87052 );
buf ( n409567 , n409566 );
and ( n409568 , n409511 , n409567 );
and ( n87056 , n409489 , n409510 );
or ( n409570 , n409568 , n87056 );
buf ( n409571 , n409570 );
buf ( n409572 , n409571 );
xor ( n409573 , n409485 , n409572 );
xor ( n409574 , n408491 , n408508 );
xor ( n87062 , n409574 , n408534 );
buf ( n409576 , n87062 );
buf ( n409577 , n409576 );
buf ( n409578 , n377068 );
not ( n409579 , n409578 );
buf ( n87067 , n380923 );
not ( n87068 , n87067 );
or ( n87069 , n409579 , n87068 );
buf ( n87070 , n22619 );
buf ( n87071 , n377071 );
nand ( n87072 , n87070 , n87071 );
buf ( n87073 , n87072 );
buf ( n87074 , n87073 );
nand ( n87075 , n87069 , n87074 );
buf ( n87076 , n87075 );
buf ( n409590 , n87076 );
not ( n409591 , n409590 );
buf ( n409592 , n45553 );
not ( n409593 , n409592 );
or ( n409594 , n409591 , n409593 );
buf ( n409595 , n85991 );
buf ( n409596 , n56794 );
nand ( n87084 , n409595 , n409596 );
buf ( n409598 , n87084 );
buf ( n409599 , n409598 );
nand ( n87087 , n409594 , n409599 );
buf ( n409601 , n87087 );
buf ( n409602 , n409601 );
xor ( n409603 , n409577 , n409602 );
and ( n409604 , n378843 , n364978 );
not ( n87092 , n378843 );
and ( n409606 , n87092 , n386093 );
or ( n409607 , n409604 , n409606 );
buf ( n409608 , n409607 );
not ( n409609 , n409608 );
buf ( n409610 , n365024 );
not ( n87098 , n409610 );
or ( n409612 , n409609 , n87098 );
buf ( n409613 , n408728 );
buf ( n409614 , n365108 );
nand ( n87102 , n409613 , n409614 );
buf ( n409616 , n87102 );
buf ( n409617 , n409616 );
nand ( n409618 , n409612 , n409617 );
buf ( n409619 , n409618 );
buf ( n409620 , n409619 );
buf ( n409621 , n375920 );
buf ( n409622 , n378098 );
and ( n409623 , n409621 , n409622 );
buf ( n409624 , n409623 );
buf ( n409625 , n409624 );
xor ( n409626 , n409620 , n409625 );
xor ( n409627 , n408902 , n408919 );
xor ( n87115 , n409627 , n408924 );
buf ( n409629 , n87115 );
buf ( n409630 , n409629 );
and ( n87118 , n409626 , n409630 );
and ( n409632 , n409620 , n409625 );
or ( n409633 , n87118 , n409632 );
buf ( n409634 , n409633 );
buf ( n409635 , n409634 );
and ( n409636 , n409603 , n409635 );
and ( n87124 , n409577 , n409602 );
or ( n409638 , n409636 , n87124 );
buf ( n409639 , n409638 );
buf ( n409640 , n409639 );
xor ( n409641 , n408713 , n86256 );
xor ( n409642 , n409641 , n86261 );
buf ( n409643 , n409642 );
buf ( n409644 , n409643 );
xor ( n87132 , n409640 , n409644 );
buf ( n87133 , n379260 );
not ( n87134 , n87133 );
buf ( n87135 , n409111 );
not ( n87136 , n87135 );
or ( n87137 , n87134 , n87136 );
buf ( n409651 , n379274 );
not ( n409652 , n409651 );
buf ( n409653 , n364900 );
not ( n409654 , n409653 );
or ( n409655 , n409652 , n409654 );
buf ( n409656 , n352268 );
buf ( n409657 , n379271 );
nand ( n87145 , n409656 , n409657 );
buf ( n409659 , n87145 );
buf ( n409660 , n409659 );
nand ( n87148 , n409655 , n409660 );
buf ( n409662 , n87148 );
buf ( n409663 , n409662 );
buf ( n409664 , n379962 );
nand ( n87152 , n409663 , n409664 );
buf ( n409666 , n87152 );
buf ( n409667 , n409666 );
nand ( n87155 , n87137 , n409667 );
buf ( n409669 , n87155 );
buf ( n409670 , n409669 );
not ( n87158 , n409670 );
buf ( n409672 , n22619 );
buf ( n409673 , n364975 );
not ( n409674 , n409673 );
buf ( n409675 , n365663 );
nand ( n409676 , n409674 , n409675 );
buf ( n409677 , n409676 );
buf ( n409678 , n409677 );
buf ( n409679 , n378098 );
and ( n409680 , n409678 , n409679 );
buf ( n409681 , n364975 );
not ( n409682 , n409681 );
buf ( n409683 , n365663 );
nor ( n87171 , n409682 , n409683 );
buf ( n87172 , n87171 );
buf ( n409686 , n87172 );
nor ( n87174 , n409680 , n409686 );
buf ( n409688 , n87174 );
buf ( n409689 , n409688 );
nand ( n87177 , n409672 , n409689 );
buf ( n409691 , n87177 );
not ( n87179 , n409691 );
not ( n87180 , n87179 );
buf ( n87181 , n409012 );
buf ( n409695 , n86481 );
xor ( n409696 , n87181 , n409695 );
buf ( n409697 , n409085 );
xnor ( n87185 , n409696 , n409697 );
buf ( n409699 , n87185 );
buf ( n87187 , n409699 );
not ( n409701 , n87187 );
buf ( n409702 , n409701 );
not ( n87190 , n409702 );
or ( n87191 , n87180 , n87190 );
not ( n409705 , n409699 );
not ( n87193 , n409691 );
or ( n87194 , n409705 , n87193 );
buf ( n409708 , n397190 );
not ( n409709 , n409708 );
buf ( n409710 , n408987 );
not ( n409711 , n409710 );
or ( n87199 , n409709 , n409711 );
buf ( n409713 , n398363 );
not ( n409714 , n409713 );
buf ( n409715 , n48458 );
not ( n409716 , n409715 );
or ( n409717 , n409714 , n409716 );
buf ( n409718 , n368656 );
buf ( n87203 , n377592 );
nand ( n87204 , n409718 , n87203 );
buf ( n409721 , n87204 );
buf ( n409722 , n409721 );
nand ( n87207 , n409717 , n409722 );
buf ( n409724 , n87207 );
buf ( n409725 , n409724 );
buf ( n409726 , n85179 );
nand ( n87211 , n409725 , n409726 );
buf ( n409728 , n87211 );
buf ( n409729 , n409728 );
nand ( n87214 , n87199 , n409729 );
buf ( n409731 , n87214 );
buf ( n409732 , n409731 );
buf ( n409733 , n369809 );
not ( n87218 , n409733 );
buf ( n409735 , n393883 );
not ( n87220 , n409735 );
buf ( n409737 , n369372 );
not ( n87222 , n409737 );
or ( n87223 , n87220 , n87222 );
buf ( n409740 , n405370 );
buf ( n409741 , n369763 );
nand ( n87226 , n409740 , n409741 );
buf ( n409743 , n87226 );
buf ( n409744 , n409743 );
nand ( n87229 , n87223 , n409744 );
buf ( n409746 , n87229 );
buf ( n409747 , n409746 );
not ( n87232 , n409747 );
or ( n409749 , n87218 , n87232 );
buf ( n409750 , n393883 );
buf ( n409751 , n377379 );
and ( n409752 , n409750 , n409751 );
not ( n87237 , n409750 );
buf ( n409754 , n408201 );
and ( n87239 , n87237 , n409754 );
or ( n87240 , n409752 , n87239 );
buf ( n409757 , n87240 );
buf ( n409758 , n409757 );
not ( n409759 , n409758 );
buf ( n409760 , n369804 );
nand ( n409761 , n409759 , n409760 );
buf ( n409762 , n409761 );
buf ( n409763 , n409762 );
nand ( n87248 , n409749 , n409763 );
buf ( n87249 , n87248 );
buf ( n409766 , n87249 );
xor ( n87251 , n408171 , n408175 );
xor ( n409768 , n87251 , n408179 );
xor ( n409769 , n407959 , n407963 );
xor ( n87254 , n409769 , n408016 );
buf ( n409771 , n87254 );
buf ( n409772 , n409771 );
buf ( n409773 , n395810 );
buf ( n409774 , n394724 );
and ( n409775 , n409773 , n409774 );
buf ( n409776 , n395816 );
buf ( n409777 , n384421 );
and ( n409778 , n409776 , n409777 );
nor ( n87263 , n409775 , n409778 );
buf ( n409780 , n87263 );
buf ( n409781 , n409780 );
buf ( n409782 , n384414 );
or ( n409783 , n409781 , n409782 );
buf ( n409784 , n407841 );
buf ( n409785 , n395635 );
or ( n409786 , n409784 , n409785 );
nand ( n87271 , n409783 , n409786 );
buf ( n409788 , n87271 );
buf ( n409789 , n409788 );
xor ( n409790 , n409772 , n409789 );
xor ( n87275 , n407981 , n407982 );
xor ( n409792 , n87275 , n408011 );
buf ( n409793 , n409792 );
buf ( n409794 , n79312 );
buf ( n409795 , n382638 );
and ( n409796 , n409794 , n409795 );
buf ( n409797 , n79318 );
buf ( n409798 , n382647 );
and ( n87283 , n409797 , n409798 );
nor ( n87284 , n409796 , n87283 );
buf ( n409801 , n87284 );
buf ( n409802 , n409801 );
buf ( n409803 , n382849 );
or ( n87288 , n409802 , n409803 );
buf ( n409805 , n407950 );
buf ( n409806 , n384157 );
or ( n409807 , n409805 , n409806 );
nand ( n87292 , n87288 , n409807 );
buf ( n87293 , n87292 );
xor ( n87294 , n409793 , n87293 );
buf ( n409811 , n79114 );
buf ( n409812 , n384343 );
and ( n87297 , n409811 , n409812 );
buf ( n409814 , n400487 );
buf ( n409815 , n384089 );
and ( n87300 , n409814 , n409815 );
nor ( n409817 , n87297 , n87300 );
buf ( n409818 , n409817 );
buf ( n409819 , n409818 );
buf ( n409820 , n384354 );
or ( n409821 , n409819 , n409820 );
buf ( n409822 , n408142 );
buf ( n409823 , n384082 );
or ( n409824 , n409822 , n409823 );
nand ( n409825 , n409821 , n409824 );
buf ( n409826 , n409825 );
and ( n87311 , n87294 , n409826 );
and ( n409828 , n409793 , n87293 );
or ( n87313 , n87311 , n409828 );
buf ( n409830 , n87313 );
and ( n409831 , n409790 , n409830 );
and ( n409832 , n409772 , n409789 );
or ( n87317 , n409831 , n409832 );
buf ( n409834 , n87317 );
xor ( n87319 , n407816 , n407832 );
xor ( n409836 , n87319 , n407849 );
and ( n409837 , n409834 , n409836 );
buf ( n409838 , n75451 );
buf ( n409839 , n394724 );
and ( n409840 , n409838 , n409839 );
buf ( n409841 , n396596 );
buf ( n409842 , n384421 );
and ( n87327 , n409841 , n409842 );
nor ( n87328 , n409840 , n87327 );
buf ( n409845 , n87328 );
buf ( n409846 , n409845 );
buf ( n409847 , n384414 );
or ( n409848 , n409846 , n409847 );
buf ( n409849 , n409780 );
buf ( n409850 , n395635 );
or ( n87335 , n409849 , n409850 );
nand ( n87336 , n409848 , n87335 );
buf ( n409853 , n87336 );
xor ( n87338 , n85594 , n408008 );
buf ( n409855 , n87338 );
buf ( n409856 , n409855 );
buf ( n409857 , n80468 );
buf ( n409858 , n382638 );
and ( n409859 , n409857 , n409858 );
buf ( n409860 , n401921 );
buf ( n409861 , n62243 );
and ( n409862 , n409860 , n409861 );
nor ( n409863 , n409859 , n409862 );
buf ( n409864 , n409863 );
buf ( n409865 , n409864 );
buf ( n409866 , n382849 );
or ( n87351 , n409865 , n409866 );
buf ( n409868 , n409801 );
buf ( n409869 , n384157 );
or ( n87354 , n409868 , n409869 );
nand ( n409871 , n87351 , n87354 );
buf ( n409872 , n409871 );
buf ( n409873 , n409872 );
xor ( n409874 , n409856 , n409873 );
buf ( n409875 , n380734 );
buf ( n409876 , n406588 );
buf ( n409877 , n403772 );
and ( n87362 , n409876 , n409877 );
buf ( n409879 , n63664 );
buf ( n409880 , n403775 );
and ( n409881 , n409879 , n409880 );
nor ( n87366 , n87362 , n409881 );
buf ( n409883 , n87366 );
buf ( n409884 , n409883 );
or ( n87369 , n409875 , n409884 );
buf ( n409886 , n408116 );
buf ( n409887 , n380733 );
or ( n409888 , n409886 , n409887 );
nand ( n87373 , n87369 , n409888 );
buf ( n87374 , n87373 );
buf ( n409891 , n87374 );
buf ( n409892 , n376889 );
buf ( n409893 , n623 );
and ( n87378 , n409892 , n409893 );
buf ( n409895 , n376910 );
buf ( n409896 , n85590 );
and ( n87381 , n409895 , n409896 );
buf ( n409898 , n57800 );
nor ( n87383 , n87381 , n409898 );
buf ( n409900 , n87383 );
buf ( n409901 , n409900 );
buf ( n409902 , n376866 );
nor ( n409903 , n87378 , n409901 , n409902 );
buf ( n409904 , n409903 );
buf ( n409905 , n409904 );
xor ( n87390 , n409891 , n409905 );
buf ( n409907 , n57789 );
buf ( n409908 , n405813 );
and ( n87393 , n409907 , n409908 );
buf ( n87394 , n378470 );
buf ( n409911 , n405816 );
and ( n409912 , n87394 , n409911 );
nor ( n87397 , n87393 , n409912 );
buf ( n409914 , n87397 );
buf ( n409915 , n409914 );
not ( n87400 , n409915 );
buf ( n409917 , n87400 );
buf ( n409918 , n409917 );
not ( n87403 , n409918 );
buf ( n409920 , n378468 );
not ( n87405 , n409920 );
or ( n409922 , n87403 , n87405 );
buf ( n409923 , n378476 );
buf ( n409924 , n408000 );
or ( n409925 , n409923 , n409924 );
nand ( n409926 , n409922 , n409925 );
buf ( n409927 , n409926 );
buf ( n409928 , n409927 );
and ( n87413 , n87390 , n409928 );
and ( n87414 , n409891 , n409905 );
or ( n409931 , n87413 , n87414 );
buf ( n409932 , n409931 );
buf ( n409933 , n409932 );
and ( n409934 , n409874 , n409933 );
and ( n409935 , n409856 , n409873 );
or ( n87420 , n409934 , n409935 );
buf ( n409937 , n87420 );
xor ( n409938 , n409853 , n409937 );
buf ( n409939 , n400503 );
buf ( n409940 , n384343 );
and ( n409941 , n409939 , n409940 );
buf ( n409942 , n400509 );
buf ( n409943 , n384089 );
and ( n409944 , n409942 , n409943 );
nor ( n409945 , n409941 , n409944 );
buf ( n409946 , n409945 );
buf ( n409947 , n409946 );
buf ( n409948 , n384354 );
or ( n409949 , n409947 , n409948 );
buf ( n409950 , n409818 );
buf ( n409951 , n384082 );
or ( n87436 , n409950 , n409951 );
nand ( n409953 , n409949 , n87436 );
buf ( n409954 , n409953 );
buf ( n409955 , n409954 );
buf ( n409956 , n56623 );
buf ( n409957 , n623 );
or ( n409958 , n409956 , n409957 );
buf ( n409959 , n376921 );
buf ( n409960 , n376866 );
buf ( n409961 , n623 );
and ( n409962 , n409959 , n409960 , n409961 );
buf ( n409963 , n376931 );
nor ( n87448 , n409962 , n409963 );
buf ( n409965 , n87448 );
buf ( n409966 , n409965 );
nand ( n409967 , n409958 , n409966 );
buf ( n409968 , n409967 );
buf ( n409969 , n378341 );
buf ( n409970 , n57800 );
buf ( n409971 , n406746 );
and ( n87456 , n409970 , n409971 );
buf ( n409973 , n378284 );
buf ( n409974 , n406749 );
and ( n87459 , n409973 , n409974 );
nor ( n409976 , n87456 , n87459 );
buf ( n409977 , n409976 );
buf ( n409978 , n409977 );
or ( n409979 , n409969 , n409978 );
buf ( n409980 , n378262 );
buf ( n409981 , n408098 );
or ( n409982 , n409980 , n409981 );
nand ( n409983 , n409979 , n409982 );
buf ( n409984 , n409983 );
xor ( n87469 , n409968 , n409984 );
buf ( n409986 , n56517 );
buf ( n87471 , n85590 );
nor ( n87472 , n409986 , n87471 );
buf ( n87473 , n87472 );
buf ( n409990 , n87473 );
buf ( n409991 , n82201 );
buf ( n409992 , n403798 );
or ( n87477 , n409991 , n409992 );
buf ( n409994 , n406588 );
buf ( n409995 , n403795 );
or ( n87480 , n409994 , n409995 );
nand ( n87481 , n87477 , n87480 );
buf ( n409998 , n87481 );
buf ( n409999 , n409998 );
not ( n87484 , n409999 );
buf ( n410001 , n380735 );
not ( n410002 , n410001 );
or ( n87487 , n87484 , n410002 );
buf ( n410004 , n409883 );
buf ( n410005 , n380733 );
or ( n87490 , n410004 , n410005 );
nand ( n87491 , n87487 , n87490 );
buf ( n410008 , n87491 );
buf ( n410009 , n410008 );
and ( n87494 , n409990 , n410009 );
buf ( n410011 , n87494 );
and ( n87496 , n87469 , n410011 );
and ( n87497 , n409968 , n409984 );
or ( n87498 , n87496 , n87497 );
buf ( n410015 , n87498 );
xor ( n410016 , n409955 , n410015 );
xor ( n87501 , n408089 , n408106 );
xor ( n87502 , n87501 , n408124 );
buf ( n410019 , n87502 );
buf ( n410020 , n410019 );
and ( n410021 , n410016 , n410020 );
and ( n410022 , n409955 , n410015 );
or ( n87507 , n410021 , n410022 );
buf ( n410024 , n87507 );
and ( n87509 , n409938 , n410024 );
and ( n410026 , n409853 , n409937 );
or ( n87511 , n87509 , n410026 );
buf ( n410028 , n87511 );
buf ( n410029 , n396499 );
buf ( n410030 , n394840 );
and ( n410031 , n410029 , n410030 );
buf ( n410032 , n394816 );
buf ( n410033 , n395890 );
and ( n410034 , n410032 , n410033 );
nor ( n410035 , n410031 , n410034 );
buf ( n410036 , n410035 );
buf ( n410037 , n410036 );
buf ( n410038 , n394838 );
or ( n87523 , n410037 , n410038 );
buf ( n410040 , n408054 );
buf ( n410041 , n394835 );
or ( n410042 , n410040 , n410041 );
nand ( n87527 , n87523 , n410042 );
buf ( n87528 , n87527 );
buf ( n410045 , n87528 );
xor ( n87530 , n410028 , n410045 );
xor ( n410047 , n408134 , n408151 );
xor ( n410048 , n410047 , n408156 );
buf ( n410049 , n410048 );
buf ( n410050 , n410049 );
and ( n410051 , n87530 , n410050 );
and ( n87536 , n410028 , n410045 );
or ( n87537 , n410051 , n87536 );
buf ( n410054 , n87537 );
xor ( n87539 , n407816 , n407832 );
xor ( n410056 , n87539 , n407849 );
and ( n87541 , n410054 , n410056 );
and ( n87542 , n409834 , n410054 );
or ( n410059 , n409837 , n87541 , n87542 );
xor ( n410060 , n407816 , n407832 );
xor ( n87545 , n410060 , n407849 );
xor ( n410062 , n409834 , n410054 );
xor ( n410063 , n87545 , n410062 );
buf ( n410064 , n410063 );
xor ( n410065 , n408063 , n408161 );
xor ( n410066 , n410065 , n408167 );
buf ( n410067 , n410066 );
buf ( n410068 , n410067 );
xor ( n410069 , n410064 , n410068 );
xor ( n410070 , n409772 , n409789 );
xor ( n87555 , n410070 , n409830 );
buf ( n410072 , n87555 );
xor ( n410073 , n407904 , n407909 );
xor ( n87558 , n410073 , n407931 );
xor ( n87559 , n85661 , n408128 );
xor ( n87560 , n87558 , n87559 );
xor ( n87561 , n409793 , n87293 );
xor ( n87562 , n87561 , n409826 );
and ( n410079 , n87560 , n87562 );
xor ( n410080 , n409891 , n409905 );
xor ( n87565 , n410080 , n409928 );
buf ( n87566 , n87565 );
buf ( n87567 , n87566 );
buf ( n410084 , n81950 );
buf ( n410085 , n382638 );
and ( n87570 , n410084 , n410085 );
buf ( n410087 , n403589 );
buf ( n410088 , n382647 );
and ( n410089 , n410087 , n410088 );
nor ( n87574 , n87570 , n410089 );
buf ( n410091 , n87574 );
buf ( n410092 , n410091 );
buf ( n410093 , n382849 );
or ( n87578 , n410092 , n410093 );
buf ( n410095 , n409864 );
buf ( n410096 , n384157 );
or ( n87581 , n410095 , n410096 );
nand ( n410098 , n87578 , n87581 );
buf ( n410099 , n410098 );
buf ( n410100 , n410099 );
xor ( n410101 , n87567 , n410100 );
buf ( n410102 , n382849 );
buf ( n410103 , n81995 );
buf ( n410104 , n382835 );
and ( n410105 , n410103 , n410104 );
buf ( n410106 , n403645 );
buf ( n410107 , n382647 );
and ( n410108 , n410106 , n410107 );
nor ( n410109 , n410105 , n410108 );
buf ( n410110 , n410109 );
buf ( n410111 , n410110 );
or ( n410112 , n410102 , n410111 );
buf ( n410113 , n410091 );
buf ( n410114 , n384157 );
or ( n87599 , n410113 , n410114 );
nand ( n410116 , n410112 , n87599 );
buf ( n410117 , n410116 );
buf ( n410118 , n410117 );
buf ( n410119 , n380581 );
buf ( n410120 , n57789 );
buf ( n410121 , n406569 );
and ( n410122 , n410120 , n410121 );
buf ( n410123 , n378470 );
buf ( n410124 , n406572 );
and ( n410125 , n410123 , n410124 );
nor ( n87610 , n410122 , n410125 );
buf ( n87611 , n87610 );
buf ( n410128 , n87611 );
or ( n87613 , n410119 , n410128 );
buf ( n410130 , n409914 );
buf ( n410131 , n378476 );
or ( n87616 , n410130 , n410131 );
nand ( n87617 , n87613 , n87616 );
buf ( n410134 , n87617 );
buf ( n410135 , n410134 );
xor ( n87620 , n410118 , n410135 );
buf ( n410137 , n378424 );
buf ( n410138 , n409977 );
or ( n87623 , n410137 , n410138 );
buf ( n410140 , n378287 );
nand ( n410141 , n87623 , n410140 );
buf ( n410142 , n410141 );
buf ( n410143 , n410142 );
and ( n87628 , n87620 , n410143 );
and ( n87629 , n410118 , n410135 );
or ( n87630 , n87628 , n87629 );
buf ( n410147 , n87630 );
buf ( n410148 , n410147 );
and ( n87633 , n410101 , n410148 );
and ( n410150 , n87567 , n410100 );
or ( n87635 , n87633 , n410150 );
buf ( n410152 , n87635 );
buf ( n410153 , n396615 );
buf ( n410154 , n394724 );
and ( n410155 , n410153 , n410154 );
buf ( n410156 , n396621 );
buf ( n410157 , n384421 );
and ( n410158 , n410156 , n410157 );
nor ( n410159 , n410155 , n410158 );
buf ( n410160 , n410159 );
buf ( n410161 , n410160 );
buf ( n410162 , n384414 );
or ( n87647 , n410161 , n410162 );
buf ( n410164 , n409845 );
buf ( n410165 , n395635 );
or ( n410166 , n410164 , n410165 );
nand ( n87651 , n87647 , n410166 );
buf ( n87652 , n87651 );
xor ( n410169 , n410152 , n87652 );
xor ( n87654 , n409856 , n409873 );
xor ( n410171 , n87654 , n409933 );
buf ( n410172 , n410171 );
and ( n410173 , n410169 , n410172 );
and ( n410174 , n410152 , n87652 );
or ( n410175 , n410173 , n410174 );
xor ( n410176 , n409793 , n87293 );
xor ( n87658 , n410176 , n409826 );
and ( n410178 , n410175 , n87658 );
and ( n87660 , n87560 , n410175 );
or ( n87661 , n410079 , n410178 , n87660 );
xor ( n410181 , n410072 , n87661 );
buf ( n410182 , n74644 );
buf ( n410183 , n394840 );
and ( n410184 , n410182 , n410183 );
buf ( n87666 , n395683 );
buf ( n410186 , n395890 );
and ( n410187 , n87666 , n410186 );
nor ( n410188 , n410184 , n410187 );
buf ( n410189 , n410188 );
buf ( n410190 , n410189 );
buf ( n410191 , n394838 );
or ( n410192 , n410190 , n410191 );
buf ( n410193 , n410036 );
buf ( n410194 , n394835 );
or ( n410195 , n410193 , n410194 );
nand ( n410196 , n410192 , n410195 );
buf ( n410197 , n410196 );
xor ( n410198 , n409853 , n409937 );
xor ( n87680 , n410198 , n410024 );
and ( n410200 , n410197 , n87680 );
xor ( n410201 , n409955 , n410015 );
xor ( n410202 , n410201 , n410020 );
buf ( n410203 , n410202 );
buf ( n410204 , n410203 );
buf ( n410205 , n395810 );
buf ( n410206 , n394840 );
and ( n410207 , n410205 , n410206 );
buf ( n410208 , n395816 );
buf ( n410209 , n395890 );
and ( n410210 , n410208 , n410209 );
nor ( n410211 , n410207 , n410210 );
buf ( n410212 , n410211 );
buf ( n410213 , n410212 );
buf ( n410214 , n394838 );
or ( n87696 , n410213 , n410214 );
buf ( n410216 , n410189 );
buf ( n410217 , n394835 );
or ( n87699 , n410216 , n410217 );
nand ( n410219 , n87696 , n87699 );
buf ( n410220 , n410219 );
buf ( n410221 , n410220 );
xor ( n410222 , n410204 , n410221 );
buf ( n410223 , n79312 );
buf ( n410224 , n384343 );
and ( n410225 , n410223 , n410224 );
buf ( n410226 , n79318 );
buf ( n410227 , n384089 );
and ( n87709 , n410226 , n410227 );
nor ( n410229 , n410225 , n87709 );
buf ( n410230 , n410229 );
buf ( n410231 , n410230 );
buf ( n410232 , n384354 );
or ( n410233 , n410231 , n410232 );
buf ( n410234 , n409946 );
buf ( n410235 , n384082 );
or ( n410236 , n410234 , n410235 );
nand ( n87718 , n410233 , n410236 );
buf ( n410238 , n87718 );
xor ( n87720 , n409968 , n409984 );
xor ( n87721 , n87720 , n410011 );
and ( n410241 , n410238 , n87721 );
buf ( n410242 , n79114 );
buf ( n410243 , n394724 );
and ( n410244 , n410242 , n410243 );
buf ( n87726 , n400487 );
buf ( n410246 , n384421 );
and ( n410247 , n87726 , n410246 );
nor ( n410248 , n410244 , n410247 );
buf ( n410249 , n410248 );
buf ( n410250 , n410249 );
buf ( n410251 , n384414 );
or ( n410252 , n410250 , n410251 );
buf ( n410253 , n410160 );
buf ( n410254 , n395635 );
or ( n410255 , n410253 , n410254 );
nand ( n87737 , n410252 , n410255 );
buf ( n87738 , n87737 );
xor ( n410258 , n409968 , n409984 );
xor ( n87740 , n410258 , n410011 );
and ( n410260 , n87738 , n87740 );
and ( n87742 , n410238 , n87738 );
or ( n410262 , n410241 , n410260 , n87742 );
buf ( n410263 , n410262 );
and ( n410264 , n410222 , n410263 );
and ( n410265 , n410204 , n410221 );
or ( n87747 , n410264 , n410265 );
buf ( n410267 , n87747 );
xor ( n410268 , n409853 , n409937 );
xor ( n87750 , n410268 , n410024 );
and ( n410270 , n410267 , n87750 );
and ( n410271 , n410197 , n410267 );
or ( n87753 , n410200 , n410270 , n410271 );
and ( n87754 , n410181 , n87753 );
and ( n87755 , n410072 , n87661 );
or ( n87756 , n87754 , n87755 );
buf ( n410276 , n87756 );
and ( n410277 , n410069 , n410276 );
and ( n87759 , n410064 , n410068 );
or ( n87760 , n410277 , n87759 );
buf ( n410280 , n87760 );
xor ( n87762 , n410059 , n410280 );
xor ( n87763 , n409768 , n87762 );
buf ( n410283 , n87763 );
not ( n410284 , n369804 );
buf ( n410285 , n368584 );
not ( n410286 , n410285 );
buf ( n410287 , n410286 );
buf ( n410288 , n410287 );
not ( n87770 , n410288 );
buf ( n410290 , n377349 );
not ( n87772 , n410290 );
or ( n87773 , n87770 , n87772 );
buf ( n410293 , n377349 );
buf ( n410294 , n368581 );
buf ( n87776 , n410294 );
buf ( n410296 , n87776 );
buf ( n410297 , n410296 );
or ( n410298 , n410293 , n410297 );
buf ( n410299 , n410298 );
buf ( n410300 , n410299 );
nand ( n87782 , n87773 , n410300 );
buf ( n410302 , n87782 );
not ( n87784 , n410302 );
or ( n87785 , n410284 , n87784 );
buf ( n410305 , n369809 );
not ( n87787 , n410305 );
buf ( n410307 , n87787 );
or ( n87789 , n409757 , n410307 );
nand ( n87790 , n87785 , n87789 );
buf ( n410310 , n87790 );
xor ( n410311 , n410283 , n410310 );
xor ( n87793 , n410028 , n410045 );
xor ( n410313 , n87793 , n410050 );
buf ( n410314 , n410313 );
xor ( n87796 , n410072 , n87661 );
xor ( n87797 , n87796 , n87753 );
and ( n87798 , n410314 , n87797 );
buf ( n410318 , n75451 );
buf ( n410319 , n394840 );
and ( n87801 , n410318 , n410319 );
buf ( n410321 , n396596 );
buf ( n410322 , n395890 );
and ( n410323 , n410321 , n410322 );
nor ( n87805 , n87801 , n410323 );
buf ( n410325 , n87805 );
buf ( n410326 , n410325 );
buf ( n410327 , n394838 );
or ( n87809 , n410326 , n410327 );
buf ( n410329 , n410212 );
buf ( n410330 , n394835 );
or ( n87812 , n410329 , n410330 );
nand ( n410332 , n87809 , n87812 );
buf ( n410333 , n410332 );
buf ( n410334 , n410333 );
buf ( n410335 , n80468 );
buf ( n410336 , n384343 );
and ( n410337 , n410335 , n410336 );
buf ( n410338 , n401921 );
buf ( n410339 , n384089 );
and ( n87821 , n410338 , n410339 );
nor ( n87822 , n410337 , n87821 );
buf ( n410342 , n87822 );
buf ( n410343 , n410342 );
buf ( n410344 , n384354 );
or ( n87826 , n410343 , n410344 );
buf ( n410346 , n410230 );
buf ( n410347 , n384082 );
or ( n87829 , n410346 , n410347 );
nand ( n410349 , n87826 , n87829 );
buf ( n410350 , n410349 );
buf ( n410351 , n410350 );
xor ( n87833 , n409990 , n410009 );
buf ( n410353 , n87833 );
buf ( n410354 , n410353 );
xor ( n87836 , n410351 , n410354 );
buf ( n410356 , n382849 );
buf ( n410357 , n382638 );
buf ( n410358 , n403772 );
and ( n87840 , n410357 , n410358 );
buf ( n410360 , n403775 );
buf ( n410361 , n382647 );
and ( n87843 , n410360 , n410361 );
nor ( n87844 , n87840 , n87843 );
buf ( n410364 , n87844 );
buf ( n410365 , n410364 );
or ( n87847 , n410356 , n410365 );
buf ( n410367 , n410110 );
buf ( n410368 , n382634 );
or ( n410369 , n410367 , n410368 );
nand ( n87851 , n87847 , n410369 );
buf ( n410371 , n87851 );
buf ( n410372 , n410371 );
buf ( n410373 , n57768 );
buf ( n410374 , n623 );
and ( n87856 , n410373 , n410374 );
buf ( n410376 , n378270 );
buf ( n410377 , n85590 );
and ( n87859 , n410376 , n410377 );
buf ( n410379 , n57789 );
nor ( n410380 , n87859 , n410379 );
buf ( n410381 , n410380 );
buf ( n410382 , n410381 );
buf ( n410383 , n57800 );
nor ( n87865 , n87856 , n410382 , n410383 );
buf ( n410385 , n87865 );
buf ( n410386 , n410385 );
xor ( n410387 , n410372 , n410386 );
buf ( n410388 , n380581 );
buf ( n410389 , n57789 );
buf ( n410390 , n406746 );
and ( n87872 , n410389 , n410390 );
buf ( n410392 , n378470 );
buf ( n410393 , n406749 );
and ( n87875 , n410392 , n410393 );
nor ( n410395 , n87872 , n87875 );
buf ( n410396 , n410395 );
buf ( n410397 , n410396 );
or ( n410398 , n410388 , n410397 );
buf ( n87880 , n87611 );
buf ( n410400 , n378476 );
or ( n410401 , n87880 , n410400 );
nand ( n410402 , n410398 , n410401 );
buf ( n410403 , n410402 );
buf ( n410404 , n410403 );
and ( n410405 , n410387 , n410404 );
and ( n410406 , n410372 , n410386 );
or ( n87888 , n410405 , n410406 );
buf ( n410408 , n87888 );
buf ( n410409 , n410408 );
and ( n87891 , n87836 , n410409 );
and ( n410411 , n410351 , n410354 );
or ( n410412 , n87891 , n410411 );
buf ( n410413 , n410412 );
buf ( n410414 , n410413 );
xor ( n87896 , n410334 , n410414 );
xor ( n410416 , n87567 , n410100 );
xor ( n87898 , n410416 , n410148 );
buf ( n410418 , n87898 );
buf ( n410419 , n410418 );
and ( n410420 , n87896 , n410419 );
and ( n87902 , n410334 , n410414 );
or ( n410422 , n410420 , n87902 );
buf ( n410423 , n410422 );
xor ( n87905 , n410152 , n87652 );
xor ( n410425 , n87905 , n410172 );
and ( n410426 , n410423 , n410425 );
xor ( n87908 , n410204 , n410221 );
xor ( n410428 , n87908 , n410263 );
buf ( n410429 , n410428 );
xor ( n87911 , n410152 , n87652 );
xor ( n410431 , n87911 , n410172 );
and ( n410432 , n410429 , n410431 );
and ( n87914 , n410423 , n410429 );
or ( n410434 , n410426 , n410432 , n87914 );
buf ( n410435 , n410434 );
xor ( n87917 , n409793 , n87293 );
xor ( n410437 , n87917 , n409826 );
xor ( n410438 , n87560 , n410175 );
xor ( n87920 , n410437 , n410438 );
buf ( n410440 , n87920 );
xor ( n87922 , n410435 , n410440 );
xor ( n87923 , n409853 , n409937 );
xor ( n410443 , n87923 , n410024 );
xor ( n410444 , n410197 , n410267 );
xor ( n87926 , n410443 , n410444 );
buf ( n410446 , n87926 );
and ( n410447 , n87922 , n410446 );
and ( n87929 , n410435 , n410440 );
or ( n87930 , n410447 , n87929 );
buf ( n410450 , n87930 );
xor ( n410451 , n410072 , n87661 );
xor ( n87933 , n410451 , n87753 );
and ( n410453 , n410450 , n87933 );
and ( n87935 , n410314 , n410450 );
or ( n410455 , n87798 , n410453 , n87935 );
buf ( n410456 , n410455 );
xor ( n87938 , n410064 , n410068 );
xor ( n410458 , n87938 , n410276 );
buf ( n410459 , n410458 );
buf ( n410460 , n410459 );
xor ( n410461 , n410456 , n410460 );
buf ( n410462 , n406346 );
not ( n410463 , n410462 );
buf ( n410464 , n368561 );
not ( n410465 , n410464 );
or ( n87947 , n410463 , n410465 );
buf ( n410467 , n410296 );
buf ( n410468 , n377779 );
nand ( n410469 , n410467 , n410468 );
buf ( n410470 , n410469 );
buf ( n410471 , n410470 );
nand ( n410472 , n87947 , n410471 );
buf ( n410473 , n410472 );
buf ( n410474 , n410473 );
not ( n410475 , n410474 );
buf ( n410476 , n369801 );
not ( n87958 , n410476 );
or ( n410478 , n410475 , n87958 );
buf ( n410479 , n410302 );
buf ( n410480 , n369809 );
nand ( n410481 , n410479 , n410480 );
buf ( n410482 , n410481 );
buf ( n410483 , n410482 );
nand ( n410484 , n410478 , n410483 );
buf ( n410485 , n410484 );
buf ( n87967 , n410485 );
and ( n87968 , n410461 , n87967 );
and ( n410488 , n410456 , n410460 );
or ( n410489 , n87968 , n410488 );
buf ( n410490 , n410489 );
buf ( n410491 , n410490 );
and ( n87973 , n410311 , n410491 );
and ( n87974 , n410283 , n410310 );
or ( n410494 , n87973 , n87974 );
buf ( n410495 , n410494 );
buf ( n410496 , n410495 );
xor ( n410497 , n409766 , n410496 );
buf ( n410498 , n377143 );
not ( n87980 , n410498 );
buf ( n410500 , n406953 );
not ( n87982 , n410500 );
or ( n87983 , n87980 , n87982 );
buf ( n410503 , n406249 );
buf ( n410504 , n377153 );
nand ( n87986 , n410503 , n410504 );
buf ( n410506 , n87986 );
buf ( n410507 , n410506 );
nand ( n87989 , n87983 , n410507 );
buf ( n87990 , n87989 );
buf ( n410510 , n87990 );
not ( n87992 , n410510 );
buf ( n410512 , n406260 );
not ( n87994 , n410512 );
or ( n87995 , n87992 , n87994 );
buf ( n410515 , n86545 );
buf ( n410516 , n44915 );
nand ( n87998 , n410515 , n410516 );
buf ( n410518 , n87998 );
buf ( n410519 , n410518 );
nand ( n410520 , n87995 , n410519 );
buf ( n410521 , n410520 );
buf ( n410522 , n410521 );
and ( n88004 , n410497 , n410522 );
and ( n88005 , n409766 , n410496 );
or ( n88006 , n88004 , n88005 );
buf ( n410526 , n88006 );
buf ( n410527 , n410526 );
xor ( n88009 , n409732 , n410527 );
and ( n410529 , n396401 , n377122 );
not ( n410530 , n396401 );
and ( n88012 , n410530 , n57463 );
or ( n410532 , n410529 , n88012 );
buf ( n410533 , n410532 );
not ( n88015 , n410533 );
buf ( n410535 , n365181 );
not ( n88017 , n410535 );
or ( n88018 , n88015 , n88017 );
buf ( n410538 , n86487 );
buf ( n410539 , n365146 );
not ( n88021 , n410539 );
buf ( n410541 , n88021 );
buf ( n410542 , n410541 );
nand ( n88024 , n410538 , n410542 );
buf ( n410544 , n88024 );
buf ( n410545 , n410544 );
nand ( n88027 , n88018 , n410545 );
buf ( n410547 , n88027 );
buf ( n410548 , n410547 );
and ( n88030 , n88009 , n410548 );
and ( n410550 , n409732 , n410527 );
or ( n88032 , n88030 , n410550 );
buf ( n410552 , n88032 );
nand ( n410553 , n87194 , n410552 );
nand ( n88035 , n87191 , n410553 );
buf ( n410555 , n88035 );
not ( n88037 , n410555 );
or ( n88038 , n87158 , n88037 );
buf ( n410558 , n88035 );
buf ( n410559 , n409669 );
or ( n410560 , n410558 , n410559 );
xor ( n88042 , n408276 , n408280 );
xor ( n88043 , n88042 , n408306 );
buf ( n410563 , n88043 );
buf ( n410564 , n410563 );
xor ( n88046 , n408171 , n408175 );
xor ( n410566 , n88046 , n408179 );
and ( n88048 , n410059 , n410566 );
xor ( n410568 , n408171 , n408175 );
xor ( n88050 , n410568 , n408179 );
and ( n410570 , n410280 , n88050 );
and ( n410571 , n410059 , n410280 );
or ( n88053 , n88048 , n410570 , n410571 );
buf ( n410573 , n88053 );
xor ( n88055 , n85397 , n85437 );
xor ( n88056 , n88055 , n408035 );
xor ( n410576 , n408043 , n408182 );
xor ( n88058 , n88056 , n410576 );
buf ( n410578 , n88058 );
xor ( n410579 , n410573 , n410578 );
buf ( n410580 , n406346 );
not ( n410581 , n410580 );
buf ( n410582 , n44906 );
not ( n410583 , n410582 );
or ( n410584 , n410581 , n410583 );
buf ( n410585 , n409022 );
buf ( n410586 , n377779 );
nand ( n410587 , n410585 , n410586 );
buf ( n410588 , n410587 );
buf ( n410589 , n410588 );
nand ( n410590 , n410584 , n410589 );
buf ( n410591 , n410590 );
buf ( n410592 , n410591 );
not ( n410593 , n410592 );
buf ( n410594 , n368599 );
not ( n410595 , n410594 );
or ( n410596 , n410593 , n410595 );
buf ( n410597 , n409029 );
buf ( n410598 , n369444 );
nand ( n410599 , n410597 , n410598 );
buf ( n410600 , n410599 );
buf ( n410601 , n410600 );
nand ( n410602 , n410596 , n410601 );
buf ( n410603 , n410602 );
buf ( n410604 , n410603 );
and ( n88086 , n410579 , n410604 );
and ( n410606 , n410573 , n410578 );
or ( n88088 , n88086 , n410606 );
buf ( n410608 , n88088 );
buf ( n410609 , n410608 );
not ( n88091 , n410609 );
not ( n410611 , n369809 );
not ( n88093 , n408268 );
or ( n88094 , n410611 , n88093 );
nand ( n410614 , n409746 , n369804 );
nand ( n410615 , n88094 , n410614 );
buf ( n410616 , n410615 );
not ( n410617 , n410616 );
buf ( n410618 , n410617 );
buf ( n410619 , n410618 );
nand ( n410620 , n88091 , n410619 );
buf ( n410621 , n410620 );
buf ( n410622 , n410621 );
not ( n88104 , n410622 );
buf ( n410624 , n86557 );
not ( n410625 , n410624 );
xnor ( n88107 , n409041 , n409079 );
buf ( n410627 , n88107 );
not ( n410628 , n410627 );
and ( n88110 , n410625 , n410628 );
buf ( n410630 , n86557 );
buf ( n410631 , n88107 );
and ( n88113 , n410630 , n410631 );
nor ( n88114 , n88110 , n88113 );
buf ( n410634 , n88114 );
buf ( n410635 , n410634 );
not ( n88117 , n410635 );
buf ( n410637 , n88117 );
buf ( n410638 , n410637 );
not ( n88120 , n410638 );
or ( n410640 , n88104 , n88120 );
buf ( n410641 , n410608 );
buf ( n410642 , n410615 );
nand ( n410643 , n410641 , n410642 );
buf ( n410644 , n410643 );
buf ( n410645 , n410644 );
nand ( n88127 , n410640 , n410645 );
buf ( n410647 , n88127 );
buf ( n410648 , n410647 );
xor ( n410649 , n410564 , n410648 );
buf ( n410650 , n58984 );
not ( n410651 , n410650 );
buf ( n410652 , n400916 );
not ( n88134 , n410652 );
or ( n410654 , n410651 , n88134 );
buf ( n410655 , n65351 );
buf ( n410656 , n408722 );
nand ( n88138 , n410655 , n410656 );
buf ( n410658 , n88138 );
buf ( n410659 , n410658 );
nand ( n88141 , n410654 , n410659 );
buf ( n410661 , n88141 );
buf ( n410662 , n410661 );
not ( n410663 , n410662 );
buf ( n410664 , n45055 );
not ( n410665 , n410664 );
or ( n88147 , n410663 , n410665 );
buf ( n410667 , n408962 );
buf ( n410668 , n365242 );
nand ( n410669 , n410667 , n410668 );
buf ( n410670 , n410669 );
buf ( n410671 , n410670 );
nand ( n410672 , n88147 , n410671 );
buf ( n410673 , n410672 );
buf ( n410674 , n410673 );
and ( n410675 , n410649 , n410674 );
and ( n410676 , n410564 , n410648 );
or ( n88158 , n410675 , n410676 );
buf ( n410678 , n88158 );
buf ( n410679 , n410678 );
nand ( n88161 , n410560 , n410679 );
buf ( n88162 , n88161 );
buf ( n88163 , n88162 );
nand ( n88164 , n88038 , n88163 );
buf ( n88165 , n88164 );
buf ( n88166 , n88165 );
xor ( n88167 , n408929 , n409093 );
xor ( n410687 , n88167 , n409119 );
buf ( n410688 , n410687 );
buf ( n410689 , n410688 );
xor ( n410690 , n88166 , n410689 );
xor ( n88172 , n408949 , n408969 );
xor ( n410692 , n88172 , n86576 );
buf ( n410693 , n410692 );
buf ( n410694 , n377094 );
not ( n88176 , n410694 );
buf ( n410696 , n380923 );
not ( n410697 , n410696 );
or ( n88179 , n88176 , n410697 );
buf ( n410699 , n22619 );
buf ( n410700 , n56687 );
nand ( n410701 , n410699 , n410700 );
buf ( n410702 , n410701 );
buf ( n410703 , n410702 );
nand ( n410704 , n88179 , n410703 );
buf ( n410705 , n410704 );
buf ( n410706 , n410705 );
not ( n88188 , n410706 );
buf ( n410708 , n384501 );
not ( n410709 , n410708 );
or ( n88191 , n88188 , n410709 );
buf ( n410711 , n87076 );
buf ( n410712 , n56794 );
nand ( n88194 , n410711 , n410712 );
buf ( n410714 , n88194 );
buf ( n410715 , n410714 );
nand ( n88197 , n88191 , n410715 );
buf ( n88198 , n88197 );
buf ( n410718 , n88198 );
xor ( n88200 , n410693 , n410718 );
buf ( n410720 , n379890 );
not ( n88202 , n410720 );
buf ( n410722 , n87041 );
not ( n410723 , n410722 );
or ( n410724 , n88202 , n410723 );
buf ( n410725 , n379838 );
not ( n410726 , n410725 );
buf ( n410727 , n45336 );
not ( n88209 , n410727 );
or ( n88210 , n410726 , n88209 );
buf ( n410730 , n378543 );
not ( n88212 , n410730 );
buf ( n410732 , n398741 );
nand ( n88214 , n88212 , n410732 );
buf ( n410734 , n88214 );
buf ( n410735 , n410734 );
nand ( n88217 , n88210 , n410735 );
buf ( n410737 , n88217 );
buf ( n88219 , n410737 );
buf ( n88220 , n379916 );
nand ( n88221 , n88219 , n88220 );
buf ( n88222 , n88221 );
buf ( n410742 , n88222 );
nand ( n88224 , n410724 , n410742 );
buf ( n410744 , n88224 );
buf ( n410745 , n410744 );
and ( n410746 , n88200 , n410745 );
and ( n88228 , n410693 , n410718 );
or ( n88229 , n410746 , n88228 );
buf ( n410749 , n88229 );
buf ( n410750 , n410749 );
and ( n88232 , n410690 , n410750 );
and ( n88233 , n88166 , n410689 );
or ( n88234 , n88232 , n88233 );
buf ( n410754 , n88234 );
buf ( n410755 , n410754 );
and ( n410756 , n87132 , n410755 );
and ( n88238 , n409640 , n409644 );
or ( n410758 , n410756 , n88238 );
buf ( n410759 , n410758 );
buf ( n410760 , n410759 );
and ( n88242 , n409573 , n410760 );
and ( n410762 , n409485 , n409572 );
or ( n410763 , n88242 , n410762 );
buf ( n410764 , n410763 );
buf ( n410765 , n410764 );
xor ( n410766 , n409481 , n410765 );
xor ( n410767 , n409439 , n409443 );
xor ( n410768 , n410767 , n409457 );
buf ( n410769 , n410768 );
buf ( n410770 , n410769 );
and ( n88247 , n410766 , n410770 );
and ( n88248 , n409481 , n410765 );
or ( n410773 , n88247 , n88248 );
buf ( n410774 , n410773 );
buf ( n410775 , n410774 );
xor ( n410776 , n409477 , n410775 );
xor ( n410777 , n407516 , n408687 );
xor ( n88254 , n410777 , n409141 );
buf ( n410779 , n88254 );
buf ( n410780 , n410779 );
and ( n88257 , n410776 , n410780 );
and ( n410782 , n409477 , n410775 );
or ( n410783 , n88257 , n410782 );
buf ( n410784 , n410783 );
buf ( n410785 , n410784 );
nand ( n88262 , n409473 , n410785 );
buf ( n410787 , n88262 );
xor ( n88264 , n409477 , n410775 );
xor ( n88265 , n88264 , n410780 );
buf ( n410790 , n88265 );
buf ( n410791 , n410790 );
xor ( n88268 , n408793 , n408797 );
xor ( n88269 , n88268 , n409136 );
buf ( n410794 , n88269 );
buf ( n410795 , n410794 );
xor ( n88272 , n409481 , n410765 );
xor ( n88273 , n88272 , n410770 );
buf ( n410798 , n88273 );
buf ( n410799 , n410798 );
xor ( n88276 , n410795 , n410799 );
xor ( n88277 , n408779 , n408783 );
xor ( n88278 , n88277 , n408788 );
buf ( n410803 , n88278 );
buf ( n410804 , n410803 );
xor ( n88281 , n408827 , n408860 );
xor ( n88282 , n88281 , n409131 );
buf ( n410807 , n88282 );
buf ( n410808 , n410807 );
xor ( n88285 , n410804 , n410808 );
xor ( n88286 , n409485 , n409572 );
xor ( n88287 , n88286 , n410760 );
buf ( n410812 , n88287 );
buf ( n410813 , n410812 );
and ( n410814 , n88285 , n410813 );
and ( n88291 , n410804 , n410808 );
or ( n410816 , n410814 , n88291 );
buf ( n410817 , n410816 );
buf ( n410818 , n410817 );
and ( n88295 , n88276 , n410818 );
and ( n88296 , n410795 , n410799 );
or ( n88297 , n88295 , n88296 );
buf ( n410822 , n88297 );
buf ( n410823 , n410822 );
nand ( n88300 , n410791 , n410823 );
buf ( n410825 , n88300 );
nand ( n88302 , n410787 , n410825 );
not ( n410827 , n88302 );
not ( n88304 , n410827 );
xor ( n88305 , n410795 , n410799 );
xor ( n88306 , n88305 , n410818 );
buf ( n410831 , n88306 );
buf ( n410832 , n410831 );
not ( n88309 , n410832 );
buf ( n410834 , n88309 );
buf ( n410835 , n410834 );
xor ( n88312 , n86380 , n409123 );
xor ( n410837 , n88312 , n409127 );
buf ( n410838 , n410837 );
buf ( n410839 , n380404 );
not ( n410840 , n410839 );
buf ( n410841 , n380368 );
not ( n88318 , n410841 );
buf ( n410843 , n45125 );
not ( n410844 , n410843 );
or ( n88321 , n88318 , n410844 );
buf ( n410846 , n45113 );
buf ( n410847 , n380364 );
nand ( n410848 , n410846 , n410847 );
buf ( n410849 , n410848 );
buf ( n410850 , n410849 );
nand ( n410851 , n88321 , n410850 );
buf ( n410852 , n410851 );
buf ( n410853 , n410852 );
not ( n410854 , n410853 );
or ( n88331 , n410840 , n410854 );
buf ( n410856 , n408819 );
buf ( n410857 , n380356 );
nand ( n88334 , n410856 , n410857 );
buf ( n410859 , n88334 );
buf ( n410860 , n410859 );
nand ( n410861 , n88331 , n410860 );
buf ( n410862 , n410861 );
buf ( n410863 , n410862 );
or ( n410864 , n410838 , n410863 );
buf ( n410865 , n410864 );
buf ( n410866 , n410865 );
xor ( n88343 , n409577 , n409602 );
xor ( n410868 , n88343 , n409635 );
buf ( n410869 , n410868 );
buf ( n410870 , n410869 );
buf ( n410871 , n58923 );
not ( n88348 , n410871 );
buf ( n410873 , n409502 );
not ( n410874 , n410873 );
or ( n88351 , n88348 , n410874 );
and ( n410876 , n365440 , n407228 );
not ( n88353 , n365440 );
and ( n88354 , n88353 , n379368 );
or ( n410879 , n410876 , n88354 );
buf ( n410880 , n410879 );
buf ( n410881 , n58867 );
nand ( n410882 , n410880 , n410881 );
buf ( n410883 , n410882 );
buf ( n410884 , n410883 );
nand ( n410885 , n88351 , n410884 );
buf ( n410886 , n410885 );
buf ( n410887 , n410886 );
xor ( n88364 , n410870 , n410887 );
buf ( n410889 , n379260 );
not ( n88366 , n410889 );
buf ( n410891 , n409662 );
not ( n88368 , n410891 );
or ( n410893 , n88366 , n88368 );
buf ( n410894 , n379274 );
not ( n410895 , n410894 );
buf ( n410896 , n60751 );
not ( n88373 , n410896 );
or ( n410898 , n410895 , n88373 );
buf ( n410899 , n45802 );
buf ( n410900 , n379271 );
nand ( n410901 , n410899 , n410900 );
buf ( n410902 , n410901 );
buf ( n410903 , n410902 );
nand ( n88380 , n410898 , n410903 );
buf ( n410905 , n88380 );
buf ( n410906 , n410905 );
buf ( n410907 , n379962 );
nand ( n410908 , n410906 , n410907 );
buf ( n410909 , n410908 );
buf ( n410910 , n410909 );
nand ( n410911 , n410893 , n410910 );
buf ( n410912 , n410911 );
buf ( n410913 , n410912 );
buf ( n410914 , n377068 );
buf ( n88391 , n386093 );
and ( n88392 , n410914 , n88391 );
not ( n410917 , n410914 );
buf ( n410918 , n364978 );
and ( n88395 , n410917 , n410918 );
nor ( n410920 , n88392 , n88395 );
buf ( n410921 , n410920 );
buf ( n410922 , n410921 );
not ( n410923 , n410922 );
buf ( n410924 , n365024 );
not ( n88401 , n410924 );
or ( n410926 , n410923 , n88401 );
buf ( n410927 , n409607 );
buf ( n410928 , n365108 );
nand ( n410929 , n410927 , n410928 );
buf ( n410930 , n410929 );
buf ( n410931 , n410930 );
nand ( n410932 , n410926 , n410931 );
buf ( n410933 , n410932 );
buf ( n410934 , n410933 );
xor ( n410935 , n410913 , n410934 );
buf ( n410936 , n379260 );
not ( n410937 , n410936 );
buf ( n410938 , n410905 );
not ( n88415 , n410938 );
or ( n410940 , n410937 , n88415 );
buf ( n410941 , n379274 );
not ( n88418 , n410941 );
buf ( n410943 , n402185 );
not ( n410944 , n410943 );
or ( n410945 , n88418 , n410944 );
buf ( n410946 , n351345 );
buf ( n410947 , n379271 );
nand ( n410948 , n410946 , n410947 );
buf ( n410949 , n410948 );
buf ( n410950 , n410949 );
nand ( n410951 , n410945 , n410950 );
buf ( n410952 , n410951 );
buf ( n410953 , n410952 );
buf ( n410954 , n379962 );
nand ( n410955 , n410953 , n410954 );
buf ( n410956 , n410955 );
buf ( n410957 , n410956 );
nand ( n88434 , n410940 , n410957 );
buf ( n410959 , n88434 );
buf ( n88436 , n410959 );
buf ( n410961 , n45491 );
not ( n88438 , n410961 );
buf ( n410963 , n379515 );
nor ( n410964 , n88438 , n410963 );
buf ( n410965 , n410964 );
buf ( n410966 , n410965 );
xor ( n410967 , n88436 , n410966 );
buf ( n410968 , n378843 );
not ( n410969 , n410968 );
buf ( n410970 , n394065 );
not ( n88447 , n410970 );
or ( n410972 , n410969 , n88447 );
buf ( n410973 , n65349 );
buf ( n410974 , n378843 );
not ( n88451 , n410974 );
buf ( n410976 , n88451 );
buf ( n410977 , n410976 );
nand ( n410978 , n410973 , n410977 );
buf ( n410979 , n410978 );
buf ( n410980 , n410979 );
nand ( n410981 , n410972 , n410980 );
buf ( n410982 , n410981 );
buf ( n410983 , n410982 );
not ( n88460 , n410983 );
buf ( n410985 , n45055 );
not ( n88462 , n410985 );
or ( n88463 , n88460 , n88462 );
buf ( n410988 , n410661 );
buf ( n410989 , n365242 );
nand ( n88466 , n410988 , n410989 );
buf ( n410991 , n88466 );
buf ( n410992 , n410991 );
nand ( n88469 , n88463 , n410992 );
buf ( n410994 , n88469 );
buf ( n410995 , n410994 );
and ( n410996 , n410967 , n410995 );
and ( n88473 , n88436 , n410966 );
or ( n88474 , n410996 , n88473 );
buf ( n410999 , n88474 );
buf ( n411000 , n410999 );
and ( n411001 , n410935 , n411000 );
and ( n88478 , n410913 , n410934 );
or ( n88479 , n411001 , n88478 );
buf ( n411004 , n88479 );
buf ( n411005 , n411004 );
xor ( n411006 , n409620 , n409625 );
xor ( n88483 , n411006 , n409630 );
buf ( n411008 , n88483 );
buf ( n411009 , n411008 );
xor ( n88486 , n411005 , n411009 );
xor ( n411011 , n410573 , n410578 );
xor ( n411012 , n411011 , n410604 );
buf ( n411013 , n411012 );
buf ( n411014 , n411013 );
buf ( n411015 , n397190 );
not ( n411016 , n411015 );
buf ( n411017 , n409724 );
not ( n88494 , n411017 );
or ( n88495 , n411016 , n88494 );
buf ( n411020 , n85179 );
buf ( n411021 , n398363 );
not ( n411022 , n411021 );
buf ( n411023 , n48791 );
not ( n88500 , n411023 );
or ( n411025 , n411022 , n88500 );
buf ( n411026 , n351044 );
buf ( n411027 , n377592 );
nand ( n411028 , n411026 , n411027 );
buf ( n411029 , n411028 );
buf ( n411030 , n411029 );
nand ( n411031 , n411025 , n411030 );
buf ( n411032 , n411031 );
buf ( n411033 , n411032 );
nand ( n411034 , n411020 , n411033 );
buf ( n411035 , n411034 );
buf ( n411036 , n411035 );
nand ( n88513 , n88495 , n411036 );
buf ( n411038 , n88513 );
buf ( n411039 , n411038 );
xor ( n88516 , n411014 , n411039 );
buf ( n411041 , n377754 );
not ( n411042 , n411041 );
buf ( n411043 , n85756 );
not ( n411044 , n411043 );
or ( n88521 , n411042 , n411044 );
buf ( n411046 , n409022 );
buf ( n411047 , n409052 );
nand ( n88524 , n411046 , n411047 );
buf ( n411049 , n88524 );
buf ( n411050 , n411049 );
nand ( n88527 , n88521 , n411050 );
buf ( n411052 , n88527 );
buf ( n411053 , n411052 );
not ( n88530 , n411053 );
buf ( n411055 , n368599 );
not ( n411056 , n411055 );
or ( n88533 , n88530 , n411056 );
buf ( n411058 , n410591 );
buf ( n411059 , n368621 );
nand ( n411060 , n411058 , n411059 );
buf ( n411061 , n411060 );
buf ( n411062 , n411061 );
nand ( n411063 , n88533 , n411062 );
buf ( n411064 , n411063 );
buf ( n411065 , n411064 );
buf ( n411066 , n76050 );
not ( n88543 , n411066 );
buf ( n411068 , n411032 );
not ( n88545 , n411068 );
or ( n411070 , n88543 , n88545 );
buf ( n411071 , n398363 );
not ( n88548 , n411071 );
buf ( n411073 , n406930 );
not ( n88550 , n411073 );
or ( n88551 , n88548 , n88550 );
buf ( n411076 , n406933 );
buf ( n411077 , n377592 );
nand ( n88554 , n411076 , n411077 );
buf ( n411079 , n88554 );
buf ( n411080 , n411079 );
nand ( n88557 , n88551 , n411080 );
buf ( n411082 , n88557 );
buf ( n411083 , n411082 );
buf ( n411084 , n85179 );
nand ( n88561 , n411083 , n411084 );
buf ( n411086 , n88561 );
buf ( n411087 , n411086 );
nand ( n88564 , n411070 , n411087 );
buf ( n411089 , n88564 );
buf ( n411090 , n411089 );
xor ( n88567 , n411065 , n411090 );
buf ( n88568 , n57463 );
not ( n88569 , n88568 );
buf ( n88570 , n405357 );
not ( n88571 , n88570 );
or ( n88572 , n88569 , n88571 );
buf ( n411097 , n406950 );
not ( n411098 , n411097 );
buf ( n411099 , n377122 );
nand ( n411100 , n411098 , n411099 );
buf ( n411101 , n411100 );
buf ( n411102 , n411101 );
nand ( n88579 , n88572 , n411102 );
buf ( n88580 , n88579 );
buf ( n411105 , n88580 );
not ( n88582 , n411105 );
buf ( n411107 , n404115 );
not ( n88584 , n411107 );
or ( n88585 , n88582 , n88584 );
buf ( n411110 , n87990 );
buf ( n411111 , n44915 );
nand ( n88588 , n411110 , n411111 );
buf ( n411113 , n88588 );
buf ( n411114 , n411113 );
nand ( n88591 , n88585 , n411114 );
buf ( n411116 , n88591 );
buf ( n411117 , n411116 );
and ( n411118 , n88567 , n411117 );
and ( n88595 , n411065 , n411090 );
or ( n411120 , n411118 , n88595 );
buf ( n411121 , n411120 );
buf ( n411122 , n411121 );
and ( n411123 , n88516 , n411122 );
and ( n411124 , n411014 , n411039 );
or ( n88601 , n411123 , n411124 );
buf ( n411126 , n88601 );
buf ( n411127 , n411126 );
and ( n88604 , n410608 , n410615 );
not ( n411129 , n410608 );
and ( n411130 , n411129 , n410618 );
or ( n411131 , n88604 , n411130 );
and ( n88608 , n411131 , n410637 );
not ( n411133 , n411131 );
and ( n88610 , n411133 , n410634 );
or ( n88611 , n88608 , n88610 );
buf ( n411136 , n88611 );
xor ( n88613 , n411127 , n411136 );
xor ( n88614 , n409732 , n410527 );
xor ( n88615 , n88614 , n410548 );
buf ( n411140 , n88615 );
buf ( n411141 , n411140 );
and ( n88618 , n88613 , n411141 );
and ( n88619 , n411127 , n411136 );
or ( n88620 , n88618 , n88619 );
buf ( n411145 , n88620 );
buf ( n411146 , n411145 );
xor ( n88623 , n410564 , n410648 );
xor ( n88624 , n88623 , n410674 );
buf ( n411149 , n88624 );
buf ( n411150 , n411149 );
xor ( n88627 , n411146 , n411150 );
buf ( n411152 , n379890 );
not ( n88629 , n411152 );
buf ( n411154 , n410737 );
not ( n88631 , n411154 );
or ( n411156 , n88629 , n88631 );
buf ( n411157 , n379838 );
not ( n411158 , n411157 );
buf ( n411159 , n381266 );
not ( n411160 , n411159 );
or ( n88637 , n411158 , n411160 );
buf ( n411162 , n351160 );
buf ( n411163 , n398741 );
nand ( n88640 , n411162 , n411163 );
buf ( n411165 , n88640 );
buf ( n411166 , n411165 );
nand ( n88643 , n88637 , n411166 );
buf ( n411168 , n88643 );
buf ( n411169 , n411168 );
buf ( n411170 , n379912 );
buf ( n411171 , n411170 );
nand ( n88648 , n411169 , n411171 );
buf ( n411173 , n88648 );
buf ( n411174 , n411173 );
nand ( n411175 , n411156 , n411174 );
buf ( n411176 , n411175 );
buf ( n411177 , n411176 );
and ( n88654 , n88627 , n411177 );
and ( n411179 , n411146 , n411150 );
or ( n88656 , n88654 , n411179 );
buf ( n411181 , n88656 );
buf ( n411182 , n411181 );
and ( n88659 , n88486 , n411182 );
and ( n411184 , n411005 , n411009 );
or ( n88661 , n88659 , n411184 );
buf ( n411186 , n88661 );
buf ( n411187 , n411186 );
and ( n411188 , n88364 , n411187 );
and ( n88665 , n410870 , n410887 );
or ( n411190 , n411188 , n88665 );
buf ( n411191 , n411190 );
buf ( n411192 , n411191 );
and ( n411193 , n410866 , n411192 );
buf ( n88670 , n410862 );
buf ( n88671 , n410837 );
and ( n88672 , n88670 , n88671 );
buf ( n88673 , n88672 );
buf ( n88674 , n88673 );
nor ( n88675 , n411193 , n88674 );
buf ( n88676 , n88675 );
buf ( n411201 , n88676 );
not ( n88678 , n411201 );
buf ( n411203 , n88678 );
buf ( n411204 , n411203 );
not ( n88681 , n411204 );
xor ( n88682 , n410804 , n410808 );
xor ( n88683 , n88682 , n410813 );
buf ( n411208 , n88683 );
buf ( n411209 , n411208 );
not ( n411210 , n411209 );
or ( n411211 , n88681 , n411210 );
buf ( n411212 , n411208 );
buf ( n411213 , n411203 );
or ( n411214 , n411212 , n411213 );
xor ( n88691 , n409489 , n409510 );
xor ( n411216 , n88691 , n409567 );
buf ( n411217 , n411216 );
buf ( n411218 , n411217 );
xor ( n88695 , n409640 , n409644 );
xor ( n88696 , n88695 , n410755 );
buf ( n411221 , n88696 );
buf ( n411222 , n411221 );
xor ( n88699 , n411218 , n411222 );
xor ( n88700 , n409532 , n409536 );
xor ( n411225 , n88700 , n409562 );
buf ( n411226 , n411225 );
buf ( n411227 , n411226 );
xor ( n411228 , n88166 , n410689 );
xor ( n411229 , n411228 , n410750 );
buf ( n411230 , n411229 );
buf ( n411231 , n411230 );
xor ( n411232 , n411227 , n411231 );
buf ( n411233 , n380356 );
not ( n88706 , n411233 );
buf ( n411235 , n410852 );
not ( n411236 , n411235 );
or ( n88709 , n88706 , n411236 );
buf ( n411238 , n380368 );
not ( n411239 , n411238 );
buf ( n411240 , n386359 );
not ( n88713 , n411240 );
or ( n88714 , n411239 , n88713 );
buf ( n88715 , n352212 );
buf ( n411244 , n380364 );
nand ( n88717 , n88715 , n411244 );
buf ( n411246 , n88717 );
buf ( n411247 , n411246 );
nand ( n88720 , n88714 , n411247 );
buf ( n411249 , n88720 );
buf ( n411250 , n411249 );
buf ( n411251 , n380404 );
nand ( n411252 , n411250 , n411251 );
buf ( n411253 , n411252 );
buf ( n411254 , n411253 );
nand ( n88727 , n88709 , n411254 );
buf ( n88728 , n88727 );
buf ( n411257 , n88728 );
and ( n88730 , n411232 , n411257 );
and ( n411259 , n411227 , n411231 );
or ( n88732 , n88730 , n411259 );
buf ( n411261 , n88732 );
buf ( n411262 , n411261 );
and ( n88735 , n88699 , n411262 );
and ( n411264 , n411218 , n411222 );
or ( n88737 , n88735 , n411264 );
buf ( n411266 , n88737 );
buf ( n411267 , n411266 );
nand ( n88740 , n411214 , n411267 );
buf ( n411269 , n88740 );
buf ( n411270 , n411269 );
nand ( n88743 , n411211 , n411270 );
buf ( n411272 , n88743 );
buf ( n411273 , n411272 );
not ( n411274 , n411273 );
buf ( n411275 , n411274 );
buf ( n411276 , n411275 );
nand ( n411277 , n410835 , n411276 );
buf ( n411278 , n411277 );
buf ( n411279 , n411278 );
not ( n411280 , n411279 );
buf ( n411281 , n410831 );
buf ( n411282 , n411272 );
nand ( n411283 , n411281 , n411282 );
buf ( n411284 , n411283 );
buf ( n411285 , n411284 );
buf ( n411286 , n58923 );
not ( n88759 , n411286 );
buf ( n411288 , n410879 );
not ( n411289 , n411288 );
or ( n411290 , n88759 , n411289 );
buf ( n411291 , n379368 );
not ( n88764 , n411291 );
buf ( n411293 , n382496 );
not ( n411294 , n411293 );
or ( n88767 , n88764 , n411294 );
buf ( n411296 , n378736 );
buf ( n411297 , n407228 );
nand ( n411298 , n411296 , n411297 );
buf ( n411299 , n411298 );
buf ( n411300 , n411299 );
nand ( n88773 , n88767 , n411300 );
buf ( n411302 , n88773 );
buf ( n411303 , n411302 );
buf ( n411304 , n379353 );
nand ( n411305 , n411303 , n411304 );
buf ( n411306 , n411305 );
buf ( n411307 , n411306 );
nand ( n88780 , n411290 , n411307 );
buf ( n411309 , n88780 );
buf ( n411310 , n411309 );
buf ( n411311 , n378098 );
not ( n411312 , n411311 );
buf ( n411313 , n380923 );
not ( n411314 , n411313 );
or ( n411315 , n411312 , n411314 );
buf ( n411316 , n22619 );
buf ( n411317 , n379515 );
nand ( n88790 , n411316 , n411317 );
buf ( n411319 , n88790 );
buf ( n411320 , n411319 );
nand ( n411321 , n411315 , n411320 );
buf ( n411322 , n411321 );
buf ( n411323 , n411322 );
not ( n411324 , n411323 );
buf ( n411325 , n365725 );
not ( n88798 , n411325 );
or ( n88799 , n411324 , n88798 );
buf ( n411328 , n410705 );
buf ( n411329 , n56794 );
nand ( n88802 , n411328 , n411329 );
buf ( n411331 , n88802 );
buf ( n411332 , n411331 );
nand ( n411333 , n88799 , n411332 );
buf ( n411334 , n411333 );
buf ( n411335 , n411334 );
and ( n411336 , n58984 , n402191 );
not ( n88809 , n58984 );
and ( n88810 , n88809 , n80732 );
or ( n88811 , n411336 , n88810 );
buf ( n411340 , n88811 );
not ( n411341 , n411340 );
buf ( n411342 , n402201 );
not ( n411343 , n411342 );
or ( n88816 , n411341 , n411343 );
buf ( n411345 , n410532 );
buf ( n411346 , n365149 );
nand ( n411347 , n411345 , n411346 );
buf ( n411348 , n411347 );
buf ( n411349 , n411348 );
nand ( n88822 , n88816 , n411349 );
buf ( n411351 , n88822 );
buf ( n411352 , n411351 );
xor ( n88825 , n409766 , n410496 );
xor ( n411354 , n88825 , n410522 );
buf ( n411355 , n411354 );
buf ( n411356 , n411355 );
xor ( n411357 , n411352 , n411356 );
buf ( n411358 , n379260 );
not ( n88831 , n411358 );
buf ( n411360 , n410952 );
not ( n411361 , n411360 );
or ( n88834 , n88831 , n411361 );
and ( n88835 , n379274 , n365384 );
not ( n411364 , n379274 );
buf ( n411365 , n365384 );
not ( n88838 , n411365 );
buf ( n88839 , n88838 );
and ( n411368 , n411364 , n88839 );
or ( n88841 , n88835 , n411368 );
buf ( n411370 , n88841 );
buf ( n411371 , n379962 );
nand ( n411372 , n411370 , n411371 );
buf ( n411373 , n411372 );
buf ( n411374 , n411373 );
nand ( n88847 , n88834 , n411374 );
buf ( n411376 , n88847 );
buf ( n411377 , n411376 );
and ( n88850 , n411357 , n411377 );
and ( n411379 , n411352 , n411356 );
or ( n411380 , n88850 , n411379 );
buf ( n411381 , n411380 );
buf ( n411382 , n411381 );
buf ( n411383 , n386091 );
not ( n88856 , n411383 );
buf ( n411385 , n377094 );
not ( n411386 , n411385 );
buf ( n411387 , n396004 );
not ( n88860 , n411387 );
or ( n411389 , n411386 , n88860 );
buf ( n411390 , n76415 );
buf ( n411391 , n56687 );
nand ( n411392 , n411390 , n411391 );
buf ( n411393 , n411392 );
buf ( n411394 , n411393 );
nand ( n411395 , n411389 , n411394 );
buf ( n411396 , n411395 );
buf ( n411397 , n411396 );
not ( n411398 , n411397 );
or ( n411399 , n88856 , n411398 );
buf ( n411400 , n410921 );
buf ( n411401 , n365108 );
nand ( n411402 , n411400 , n411401 );
buf ( n411403 , n411402 );
buf ( n88876 , n411403 );
nand ( n88877 , n411399 , n88876 );
buf ( n411406 , n88877 );
buf ( n411407 , n411406 );
xor ( n88880 , n411382 , n411407 );
xor ( n411409 , n411014 , n411039 );
xor ( n88882 , n411409 , n411122 );
buf ( n411411 , n88882 );
buf ( n411412 , n411411 );
xor ( n411413 , n410283 , n410310 );
xor ( n411414 , n411413 , n410491 );
buf ( n411415 , n411414 );
buf ( n411416 , n411415 );
xor ( n88889 , n410456 , n410460 );
xor ( n411418 , n88889 , n87967 );
buf ( n411419 , n411418 );
buf ( n411420 , n411419 );
buf ( n411421 , n76050 );
not ( n411422 , n411421 );
buf ( n411423 , n411082 );
not ( n411424 , n411423 );
or ( n411425 , n411422 , n411424 );
buf ( n411426 , n398363 );
not ( n411427 , n411426 );
buf ( n88900 , n408201 );
not ( n88901 , n88900 );
or ( n88902 , n411427 , n88901 );
not ( n411431 , n377583 );
buf ( n88904 , n411431 );
buf ( n411433 , n88904 );
buf ( n411434 , n352381 );
nand ( n411435 , n411433 , n411434 );
buf ( n411436 , n411435 );
buf ( n411437 , n411436 );
nand ( n411438 , n88902 , n411437 );
buf ( n411439 , n411438 );
buf ( n411440 , n411439 );
buf ( n411441 , n85179 );
nand ( n88914 , n411440 , n411441 );
buf ( n411443 , n88914 );
buf ( n411444 , n411443 );
nand ( n411445 , n411425 , n411444 );
buf ( n411446 , n411445 );
buf ( n411447 , n411446 );
xor ( n411448 , n411420 , n411447 );
buf ( n411449 , n377143 );
not ( n88922 , n411449 );
buf ( n411451 , n85756 );
not ( n411452 , n411451 );
or ( n88925 , n88922 , n411452 );
buf ( n411454 , n409022 );
buf ( n411455 , n377153 );
nand ( n88928 , n411454 , n411455 );
buf ( n411457 , n88928 );
buf ( n411458 , n411457 );
nand ( n411459 , n88925 , n411458 );
buf ( n411460 , n411459 );
buf ( n411461 , n411460 );
not ( n411462 , n411461 );
buf ( n411463 , n368599 );
not ( n411464 , n411463 );
or ( n411465 , n411462 , n411464 );
buf ( n411466 , n411052 );
buf ( n411467 , n368621 );
nand ( n88940 , n411466 , n411467 );
buf ( n411469 , n88940 );
buf ( n411470 , n411469 );
nand ( n88943 , n411465 , n411470 );
buf ( n411472 , n88943 );
buf ( n411473 , n411472 );
and ( n88946 , n411448 , n411473 );
and ( n88947 , n411420 , n411447 );
or ( n88948 , n88946 , n88947 );
buf ( n411477 , n88948 );
buf ( n411478 , n411477 );
xor ( n88951 , n411416 , n411478 );
buf ( n411480 , n379260 );
not ( n88953 , n411480 );
buf ( n411482 , n88841 );
not ( n88955 , n411482 );
or ( n88956 , n88953 , n88955 );
buf ( n411485 , n379274 );
not ( n88958 , n411485 );
buf ( n411487 , n48458 );
not ( n88960 , n411487 );
or ( n411489 , n88958 , n88960 );
buf ( n411490 , n368656 );
buf ( n411491 , n379271 );
nand ( n411492 , n411490 , n411491 );
buf ( n411493 , n411492 );
buf ( n411494 , n411493 );
nand ( n411495 , n411489 , n411494 );
buf ( n411496 , n411495 );
buf ( n411497 , n411496 );
buf ( n411498 , n379962 );
nand ( n88971 , n411497 , n411498 );
buf ( n411500 , n88971 );
buf ( n411501 , n411500 );
nand ( n88974 , n88956 , n411501 );
buf ( n411503 , n88974 );
buf ( n411504 , n411503 );
and ( n88977 , n88951 , n411504 );
and ( n411506 , n411416 , n411478 );
or ( n411507 , n88977 , n411506 );
buf ( n411508 , n411507 );
buf ( n411509 , n411508 );
xor ( n411510 , n411412 , n411509 );
buf ( n411511 , n76415 );
buf ( n411512 , n22899 );
not ( n411513 , n411512 );
buf ( n411514 , n386040 );
not ( n88987 , n411514 );
or ( n411516 , n411513 , n88987 );
buf ( n88989 , n378098 );
nand ( n88990 , n411516 , n88989 );
buf ( n88991 , n88990 );
buf ( n88992 , n88991 );
buf ( n411521 , n85938 );
buf ( n411522 , n342848 );
nand ( n88995 , n411521 , n411522 );
buf ( n411524 , n88995 );
buf ( n411525 , n411524 );
and ( n411526 , n411511 , n88992 , n411525 );
buf ( n411527 , n411526 );
buf ( n411528 , n411527 );
and ( n89001 , n411510 , n411528 );
and ( n89002 , n411412 , n411509 );
or ( n411531 , n89001 , n89002 );
buf ( n411532 , n411531 );
buf ( n411533 , n411532 );
and ( n89006 , n88880 , n411533 );
and ( n89007 , n411382 , n411407 );
or ( n89008 , n89006 , n89007 );
buf ( n411537 , n89008 );
buf ( n411538 , n411537 );
xor ( n89011 , n411335 , n411538 );
buf ( n411540 , n410552 );
buf ( n411541 , n409702 );
xor ( n411542 , n411540 , n411541 );
buf ( n411543 , n409691 );
xnor ( n411544 , n411542 , n411543 );
buf ( n411545 , n411544 );
buf ( n411546 , n411545 );
and ( n89019 , n89011 , n411546 );
and ( n411548 , n411335 , n411538 );
or ( n89021 , n89019 , n411548 );
buf ( n411550 , n89021 );
buf ( n411551 , n411550 );
xor ( n89024 , n411310 , n411551 );
xor ( n411553 , n410678 , n409669 );
xor ( n411554 , n411553 , n88035 );
buf ( n411555 , n411554 );
and ( n411556 , n89024 , n411555 );
and ( n411557 , n411310 , n411551 );
or ( n89030 , n411556 , n411557 );
buf ( n411559 , n89030 );
buf ( n411560 , n411559 );
xor ( n89033 , n410693 , n410718 );
xor ( n411562 , n89033 , n410745 );
buf ( n411563 , n411562 );
buf ( n411564 , n411563 );
buf ( n411565 , n380356 );
not ( n89038 , n411565 );
buf ( n411567 , n411249 );
not ( n411568 , n411567 );
or ( n89041 , n89038 , n411568 );
buf ( n411570 , n380368 );
not ( n411571 , n411570 );
buf ( n411572 , n365474 );
not ( n411573 , n411572 );
or ( n89046 , n411571 , n411573 );
buf ( n411575 , n31260 );
buf ( n411576 , n380364 );
nand ( n89049 , n411575 , n411576 );
buf ( n411578 , n89049 );
buf ( n411579 , n411578 );
nand ( n411580 , n89046 , n411579 );
buf ( n411581 , n411580 );
buf ( n411582 , n411581 );
buf ( n411583 , n380404 );
nand ( n411584 , n411582 , n411583 );
buf ( n411585 , n411584 );
buf ( n411586 , n411585 );
nand ( n411587 , n89041 , n411586 );
buf ( n411588 , n411587 );
buf ( n411589 , n411588 );
xor ( n89062 , n411564 , n411589 );
xor ( n89063 , n410913 , n410934 );
xor ( n89064 , n89063 , n411000 );
buf ( n411593 , n89064 );
buf ( n411594 , n411593 );
buf ( n411595 , n58923 );
not ( n411596 , n411595 );
buf ( n411597 , n411302 );
not ( n411598 , n411597 );
or ( n411599 , n411596 , n411598 );
buf ( n411600 , n407228 );
not ( n411601 , n411600 );
buf ( n411602 , n57233 );
not ( n89074 , n411602 );
or ( n411604 , n411601 , n89074 );
buf ( n411605 , n83069 );
buf ( n411606 , n407228 );
or ( n411607 , n411605 , n411606 );
buf ( n411608 , n411607 );
buf ( n411609 , n411608 );
nand ( n411610 , n411604 , n411609 );
buf ( n411611 , n411610 );
buf ( n411612 , n411611 );
buf ( n411613 , n379353 );
nand ( n89085 , n411612 , n411613 );
buf ( n411615 , n89085 );
buf ( n411616 , n411615 );
nand ( n89088 , n411599 , n411616 );
buf ( n411618 , n89088 );
buf ( n411619 , n411618 );
xor ( n89091 , n411594 , n411619 );
buf ( n411621 , n411168 );
buf ( n411622 , n379890 );
and ( n89094 , n411621 , n411622 );
buf ( n411624 , n379838 );
not ( n411625 , n411624 );
buf ( n411626 , n32234 );
not ( n411627 , n411626 );
or ( n411628 , n411625 , n411627 );
buf ( n411629 , n352268 );
buf ( n411630 , n398741 );
nand ( n411631 , n411629 , n411630 );
buf ( n411632 , n411631 );
buf ( n411633 , n411632 );
nand ( n411634 , n411628 , n411633 );
buf ( n411635 , n411634 );
buf ( n411636 , n411635 );
not ( n411637 , n411636 );
buf ( n411638 , n59424 );
nor ( n89110 , n411637 , n411638 );
buf ( n411640 , n89110 );
buf ( n411641 , n411640 );
nor ( n411642 , n89094 , n411641 );
buf ( n411643 , n411642 );
buf ( n411644 , n411643 );
not ( n411645 , n411644 );
buf ( n411646 , n379368 );
not ( n89118 , n411646 );
buf ( n411648 , n378543 );
not ( n411649 , n411648 );
or ( n89121 , n89118 , n411649 );
buf ( n411651 , n351195 );
buf ( n411652 , n407228 );
nand ( n411653 , n411651 , n411652 );
buf ( n411654 , n411653 );
buf ( n411655 , n411654 );
nand ( n411656 , n89121 , n411655 );
buf ( n411657 , n411656 );
buf ( n411658 , n411657 );
not ( n89130 , n411658 );
buf ( n411660 , n89130 );
buf ( n411661 , n411660 );
not ( n89133 , n411661 );
buf ( n411663 , n379350 );
not ( n89135 , n411663 );
and ( n89136 , n89133 , n89135 );
buf ( n411666 , n411611 );
buf ( n411667 , n58923 );
and ( n89139 , n411666 , n411667 );
nor ( n89140 , n89136 , n89139 );
buf ( n411670 , n89140 );
buf ( n411671 , n411670 );
not ( n89143 , n411671 );
or ( n89144 , n411645 , n89143 );
xor ( n89145 , n411127 , n411136 );
xor ( n89146 , n89145 , n411141 );
buf ( n411676 , n89146 );
buf ( n411677 , n411676 );
nand ( n89149 , n89144 , n411677 );
buf ( n411679 , n89149 );
buf ( n411680 , n411679 );
buf ( n411681 , n411643 );
not ( n89153 , n411681 );
buf ( n411683 , n411670 );
not ( n89155 , n411683 );
buf ( n411685 , n89155 );
buf ( n411686 , n411685 );
nand ( n89158 , n89153 , n411686 );
buf ( n411688 , n89158 );
buf ( n411689 , n411688 );
nand ( n411690 , n411680 , n411689 );
buf ( n411691 , n411690 );
buf ( n411692 , n411691 );
and ( n89164 , n89091 , n411692 );
and ( n89165 , n411594 , n411619 );
or ( n89166 , n89164 , n89165 );
buf ( n411696 , n89166 );
buf ( n411697 , n411696 );
and ( n89169 , n89062 , n411697 );
and ( n411699 , n411564 , n411589 );
or ( n89171 , n89169 , n411699 );
buf ( n411701 , n89171 );
buf ( n411702 , n411701 );
xor ( n411703 , n411560 , n411702 );
xor ( n89175 , n410870 , n410887 );
xor ( n411705 , n89175 , n411187 );
buf ( n411706 , n411705 );
buf ( n411707 , n411706 );
and ( n89179 , n411703 , n411707 );
and ( n89180 , n411560 , n411702 );
or ( n411710 , n89179 , n89180 );
buf ( n411711 , n411710 );
buf ( n411712 , n411711 );
buf ( n411713 , n410837 );
buf ( n411714 , n410862 );
xor ( n89186 , n411713 , n411714 );
buf ( n411716 , n411191 );
xor ( n411717 , n89186 , n411716 );
buf ( n411718 , n411717 );
buf ( n411719 , n411718 );
xor ( n89191 , n411712 , n411719 );
xor ( n89192 , n411218 , n411222 );
xor ( n411722 , n89192 , n411262 );
buf ( n411723 , n411722 );
buf ( n411724 , n411723 );
xor ( n89196 , n89191 , n411724 );
buf ( n411726 , n89196 );
buf ( n411727 , n411726 );
xor ( n89199 , n411227 , n411231 );
xor ( n411729 , n89199 , n411257 );
buf ( n411730 , n411729 );
buf ( n411731 , n411730 );
xor ( n411732 , n411005 , n411009 );
xor ( n411733 , n411732 , n411182 );
buf ( n411734 , n411733 );
buf ( n411735 , n411734 );
buf ( n411736 , n377068 );
not ( n89208 , n411736 );
buf ( n411738 , n394065 );
not ( n411739 , n411738 );
or ( n89211 , n89208 , n411739 );
buf ( n411741 , n377071 );
buf ( n411742 , n65349 );
nand ( n89214 , n411741 , n411742 );
buf ( n411744 , n89214 );
buf ( n411745 , n411744 );
nand ( n89217 , n89211 , n411745 );
buf ( n89218 , n89217 );
buf ( n411748 , n89218 );
not ( n89220 , n411748 );
buf ( n411750 , n400929 );
not ( n411751 , n411750 );
or ( n411752 , n89220 , n411751 );
buf ( n411753 , n410982 );
buf ( n411754 , n365242 );
nand ( n411755 , n411753 , n411754 );
buf ( n411756 , n411755 );
buf ( n411757 , n411756 );
nand ( n89229 , n411752 , n411757 );
buf ( n411759 , n89229 );
buf ( n411760 , n411759 );
buf ( n411761 , n378843 );
not ( n89233 , n411761 );
buf ( n411763 , n45050 );
not ( n411764 , n411763 );
or ( n89236 , n89233 , n411764 );
buf ( n411766 , n410976 );
buf ( n411767 , n402190 );
nand ( n89239 , n411766 , n411767 );
buf ( n411769 , n89239 );
buf ( n411770 , n411769 );
nand ( n89242 , n89236 , n411770 );
buf ( n89243 , n89242 );
buf ( n411773 , n89243 );
not ( n89245 , n411773 );
not ( n411775 , n45010 );
buf ( n411776 , n411775 );
not ( n89248 , n411776 );
or ( n411778 , n89245 , n89248 );
buf ( n411779 , n88811 );
buf ( n411780 , n410541 );
nand ( n89252 , n411779 , n411780 );
buf ( n411782 , n89252 );
buf ( n411783 , n411782 );
nand ( n411784 , n411778 , n411783 );
buf ( n411785 , n411784 );
buf ( n411786 , n411785 );
xor ( n411787 , n410072 , n87661 );
xor ( n89259 , n411787 , n87753 );
xor ( n411789 , n410314 , n410450 );
xor ( n411790 , n89259 , n411789 );
buf ( n411791 , n411790 );
buf ( n411792 , n377754 );
not ( n411793 , n411792 );
buf ( n411794 , n368584 );
not ( n89266 , n411794 );
or ( n89267 , n411793 , n89266 );
buf ( n411797 , n368561 );
not ( n89269 , n411797 );
buf ( n411799 , n409052 );
nand ( n411800 , n89269 , n411799 );
buf ( n411801 , n411800 );
buf ( n411802 , n411801 );
nand ( n89274 , n89267 , n411802 );
buf ( n411804 , n89274 );
buf ( n411805 , n411804 );
not ( n411806 , n411805 );
buf ( n411807 , n369801 );
not ( n411808 , n411807 );
or ( n411809 , n411806 , n411808 );
buf ( n411810 , n410473 );
buf ( n411811 , n369809 );
nand ( n411812 , n411810 , n411811 );
buf ( n411813 , n411812 );
buf ( n411814 , n411813 );
nand ( n89286 , n411809 , n411814 );
buf ( n411816 , n89286 );
buf ( n89288 , n411816 );
xor ( n89289 , n411791 , n89288 );
buf ( n411819 , n76050 );
not ( n411820 , n411819 );
buf ( n411821 , n411439 );
not ( n411822 , n411821 );
or ( n89294 , n411820 , n411822 );
buf ( n411824 , n398363 );
not ( n411825 , n411824 );
buf ( n411826 , n377349 );
not ( n89298 , n411826 );
or ( n89299 , n411825 , n89298 );
buf ( n411829 , n409020 );
buf ( n411830 , n88904 );
nand ( n89302 , n411829 , n411830 );
buf ( n411832 , n89302 );
buf ( n411833 , n411832 );
nand ( n89305 , n89299 , n411833 );
buf ( n411835 , n89305 );
buf ( n411836 , n411835 );
buf ( n411837 , n85179 );
nand ( n89309 , n411836 , n411837 );
buf ( n411839 , n89309 );
buf ( n411840 , n411839 );
nand ( n89312 , n89294 , n411840 );
buf ( n411842 , n89312 );
buf ( n411843 , n411842 );
and ( n89315 , n89289 , n411843 );
and ( n411845 , n411791 , n89288 );
or ( n89317 , n89315 , n411845 );
buf ( n411847 , n89317 );
buf ( n411848 , n411847 );
buf ( n411849 , n379260 );
not ( n411850 , n411849 );
buf ( n411851 , n411496 );
not ( n89323 , n411851 );
or ( n411853 , n411850 , n89323 );
not ( n411854 , n379274 );
not ( n89326 , n48791 );
or ( n411856 , n411854 , n89326 );
buf ( n411857 , n351044 );
buf ( n411858 , n379271 );
nand ( n411859 , n411857 , n411858 );
buf ( n411860 , n411859 );
nand ( n411861 , n411856 , n411860 );
nand ( n89333 , n411861 , n379962 );
buf ( n411863 , n89333 );
nand ( n411864 , n411853 , n411863 );
buf ( n411865 , n411864 );
buf ( n411866 , n411865 );
xor ( n89338 , n411848 , n411866 );
and ( n89339 , n58984 , n369183 );
not ( n411869 , n58984 );
and ( n89341 , n411869 , n406249 );
or ( n411871 , n89339 , n89341 );
buf ( n411872 , n411871 );
not ( n89344 , n411872 );
buf ( n411874 , n404115 );
not ( n411875 , n411874 );
or ( n89347 , n89344 , n411875 );
buf ( n411877 , n88580 );
buf ( n411878 , n44915 );
nand ( n89350 , n411877 , n411878 );
buf ( n89351 , n89350 );
buf ( n411881 , n89351 );
nand ( n89353 , n89347 , n411881 );
buf ( n411883 , n89353 );
buf ( n411884 , n411883 );
and ( n89356 , n89338 , n411884 );
and ( n411886 , n411848 , n411866 );
or ( n411887 , n89356 , n411886 );
buf ( n411888 , n411887 );
buf ( n411889 , n411888 );
xor ( n89361 , n411786 , n411889 );
xor ( n89362 , n411065 , n411090 );
xor ( n411892 , n89362 , n411117 );
buf ( n411893 , n411892 );
buf ( n411894 , n411893 );
and ( n411895 , n89361 , n411894 );
and ( n411896 , n411786 , n411889 );
or ( n89368 , n411895 , n411896 );
buf ( n411898 , n89368 );
buf ( n89370 , n411898 );
xor ( n89371 , n411760 , n89370 );
xor ( n411901 , n411352 , n411356 );
xor ( n411902 , n411901 , n411377 );
buf ( n411903 , n411902 );
buf ( n411904 , n411903 );
and ( n411905 , n89371 , n411904 );
and ( n89377 , n411760 , n89370 );
or ( n411907 , n411905 , n89377 );
buf ( n411908 , n411907 );
buf ( n411909 , n411908 );
xor ( n89381 , n88436 , n410966 );
xor ( n411911 , n89381 , n410995 );
buf ( n411912 , n411911 );
buf ( n411913 , n411912 );
xor ( n411914 , n411909 , n411913 );
buf ( n411915 , n379890 );
not ( n89387 , n411915 );
buf ( n411917 , n411635 );
not ( n411918 , n411917 );
or ( n89390 , n89387 , n411918 );
buf ( n411920 , n379838 );
not ( n411921 , n411920 );
buf ( n411922 , n74977 );
not ( n89394 , n411922 );
or ( n411924 , n411921 , n89394 );
buf ( n411925 , n398741 );
buf ( n411926 , n45802 );
nand ( n89398 , n411925 , n411926 );
buf ( n411928 , n89398 );
buf ( n411929 , n411928 );
nand ( n89401 , n411924 , n411929 );
buf ( n89402 , n89401 );
buf ( n411932 , n89402 );
buf ( n411933 , n411170 );
nand ( n411934 , n411932 , n411933 );
buf ( n411935 , n411934 );
buf ( n411936 , n411935 );
nand ( n411937 , n89390 , n411936 );
buf ( n411938 , n411937 );
buf ( n411939 , n411938 );
not ( n89411 , n411939 );
buf ( n411941 , n379515 );
buf ( n411942 , n396004 );
and ( n89414 , n411941 , n411942 );
not ( n411944 , n411941 );
buf ( n411945 , n386093 );
and ( n89417 , n411944 , n411945 );
nor ( n411947 , n89414 , n89417 );
buf ( n411948 , n411947 );
buf ( n411949 , n411948 );
not ( n411950 , n411949 );
buf ( n411951 , n365021 );
not ( n411952 , n411951 );
or ( n89424 , n411950 , n411952 );
buf ( n411954 , n411396 );
buf ( n411955 , n365108 );
nand ( n89427 , n411954 , n411955 );
buf ( n411957 , n89427 );
buf ( n411958 , n411957 );
nand ( n89430 , n89424 , n411958 );
buf ( n411960 , n89430 );
buf ( n411961 , n411960 );
not ( n89433 , n411961 );
or ( n411963 , n89411 , n89433 );
buf ( n411964 , n411938 );
buf ( n411965 , n411960 );
or ( n411966 , n411964 , n411965 );
buf ( n411967 , n365010 );
buf ( n411968 , n378098 );
nand ( n89440 , n411967 , n411968 );
buf ( n411970 , n89440 );
buf ( n411971 , n411970 );
not ( n411972 , n411971 );
xor ( n89444 , n411416 , n411478 );
xor ( n411974 , n89444 , n411504 );
buf ( n411975 , n411974 );
buf ( n411976 , n411975 );
not ( n89448 , n411976 );
buf ( n411978 , n89448 );
buf ( n411979 , n411978 );
not ( n89451 , n411979 );
or ( n89452 , n411972 , n89451 );
xor ( n89453 , n410152 , n87652 );
xor ( n89454 , n89453 , n410172 );
xor ( n89455 , n410423 , n410429 );
xor ( n89456 , n89454 , n89455 );
buf ( n411986 , n89456 );
xor ( n89458 , n409968 , n409984 );
xor ( n89459 , n89458 , n410011 );
xor ( n89460 , n410238 , n87738 );
xor ( n89461 , n89459 , n89460 );
buf ( n411991 , n89461 );
xor ( n89463 , n410118 , n410135 );
xor ( n89464 , n89463 , n410143 );
buf ( n411994 , n89464 );
buf ( n411995 , n411994 );
buf ( n411996 , n400503 );
buf ( n411997 , n394724 );
and ( n89469 , n411996 , n411997 );
buf ( n411999 , n400509 );
buf ( n412000 , n384421 );
and ( n89472 , n411999 , n412000 );
nor ( n89473 , n89469 , n89472 );
buf ( n412003 , n89473 );
buf ( n412004 , n412003 );
buf ( n412005 , n384414 );
or ( n412006 , n412004 , n412005 );
buf ( n412007 , n410249 );
buf ( n412008 , n395635 );
or ( n89480 , n412007 , n412008 );
nand ( n412010 , n412006 , n89480 );
buf ( n412011 , n412010 );
buf ( n412012 , n412011 );
xor ( n412013 , n411995 , n412012 );
buf ( n412014 , n378262 );
buf ( n412015 , n85590 );
nor ( n412016 , n412014 , n412015 );
buf ( n412017 , n412016 );
buf ( n412018 , n412017 );
buf ( n412019 , n382638 );
buf ( n412020 , n403795 );
and ( n89492 , n412019 , n412020 );
buf ( n412022 , n382647 );
buf ( n412023 , n403798 );
and ( n89495 , n412022 , n412023 );
nor ( n89496 , n89492 , n89495 );
buf ( n412026 , n89496 );
buf ( n89498 , n412026 );
not ( n412028 , n89498 );
buf ( n412029 , n412028 );
buf ( n412030 , n412029 );
not ( n89502 , n412030 );
buf ( n412032 , n382655 );
not ( n89504 , n412032 );
or ( n412034 , n89502 , n89504 );
buf ( n412035 , n410364 );
buf ( n412036 , n382634 );
or ( n89505 , n412035 , n412036 );
nand ( n89506 , n412034 , n89505 );
buf ( n412039 , n89506 );
buf ( n412040 , n412039 );
and ( n89509 , n412018 , n412040 );
buf ( n412042 , n89509 );
buf ( n412043 , n380734 );
buf ( n412044 , n406588 );
buf ( n412045 , n405813 );
and ( n89514 , n412044 , n412045 );
buf ( n412047 , n63664 );
buf ( n412048 , n405816 );
and ( n89517 , n412047 , n412048 );
nor ( n412050 , n89514 , n89517 );
buf ( n412051 , n412050 );
buf ( n412052 , n412051 );
or ( n412053 , n412043 , n412052 );
buf ( n412054 , n409998 );
not ( n89523 , n412054 );
buf ( n89524 , n89523 );
buf ( n412057 , n89524 );
buf ( n412058 , n380733 );
or ( n412059 , n412057 , n412058 );
nand ( n412060 , n412053 , n412059 );
buf ( n412061 , n412060 );
xor ( n89530 , n412042 , n412061 );
buf ( n412063 , n378287 );
buf ( n412064 , n623 );
or ( n89533 , n412063 , n412064 );
buf ( n412066 , n378280 );
buf ( n412067 , n57800 );
buf ( n412068 , n623 );
and ( n412069 , n412066 , n412067 , n412068 );
buf ( n412070 , n378295 );
not ( n412071 , n412070 );
buf ( n412072 , n412071 );
buf ( n412073 , n412072 );
nor ( n89542 , n412069 , n412073 );
buf ( n412075 , n89542 );
buf ( n412076 , n412075 );
nand ( n89545 , n89533 , n412076 );
buf ( n412078 , n89545 );
and ( n89547 , n89530 , n412078 );
and ( n412080 , n412042 , n412061 );
or ( n412081 , n89547 , n412080 );
buf ( n412082 , n412081 );
and ( n412083 , n412013 , n412082 );
and ( n89552 , n411995 , n412012 );
or ( n412085 , n412083 , n89552 );
buf ( n412086 , n412085 );
buf ( n412087 , n412086 );
xor ( n412088 , n411991 , n412087 );
buf ( n412089 , n384354 );
buf ( n412090 , n81995 );
buf ( n412091 , n382627 );
and ( n89560 , n412090 , n412091 );
buf ( n412093 , n403645 );
buf ( n412094 , n62026 );
and ( n412095 , n412093 , n412094 );
nor ( n89564 , n89560 , n412095 );
buf ( n412097 , n89564 );
buf ( n412098 , n412097 );
or ( n412099 , n412089 , n412098 );
buf ( n412100 , n81950 );
buf ( n412101 , n382627 );
and ( n412102 , n412100 , n412101 );
buf ( n412103 , n403589 );
buf ( n412104 , n62026 );
and ( n412105 , n412103 , n412104 );
nor ( n412106 , n412102 , n412105 );
buf ( n412107 , n412106 );
buf ( n412108 , n412107 );
buf ( n412109 , n384082 );
or ( n89578 , n412108 , n412109 );
nand ( n412111 , n412099 , n89578 );
buf ( n412112 , n412111 );
buf ( n412113 , n412112 );
buf ( n412114 , n380734 );
buf ( n412115 , n406588 );
buf ( n412116 , n406569 );
and ( n89585 , n412115 , n412116 );
buf ( n412118 , n82201 );
buf ( n412119 , n406572 );
and ( n89588 , n412118 , n412119 );
nor ( n89589 , n89585 , n89588 );
buf ( n412122 , n89589 );
buf ( n412123 , n412122 );
or ( n412124 , n412114 , n412123 );
buf ( n412125 , n412051 );
buf ( n412126 , n380733 );
or ( n412127 , n412125 , n412126 );
nand ( n412128 , n412124 , n412127 );
buf ( n412129 , n412128 );
buf ( n412130 , n412129 );
xor ( n412131 , n412113 , n412130 );
buf ( n412132 , n410396 );
buf ( n412133 , n394774 );
or ( n412134 , n412132 , n412133 );
buf ( n89603 , n378473 );
nand ( n89604 , n412134 , n89603 );
buf ( n89605 , n89604 );
buf ( n412138 , n89605 );
and ( n89607 , n412131 , n412138 );
and ( n412140 , n412113 , n412130 );
or ( n412141 , n89607 , n412140 );
buf ( n412142 , n412141 );
buf ( n89611 , n412107 );
buf ( n89612 , n384354 );
or ( n89613 , n89611 , n89612 );
buf ( n412146 , n410342 );
buf ( n412147 , n384082 );
or ( n412148 , n412146 , n412147 );
nand ( n89617 , n89613 , n412148 );
buf ( n89618 , n89617 );
xor ( n412151 , n412142 , n89618 );
xor ( n89620 , n410372 , n410386 );
xor ( n412153 , n89620 , n410404 );
buf ( n412154 , n412153 );
and ( n89623 , n412151 , n412154 );
and ( n89624 , n412142 , n89618 );
or ( n412157 , n89623 , n89624 );
buf ( n412158 , n412157 );
buf ( n412159 , n396615 );
buf ( n412160 , n394840 );
and ( n412161 , n412159 , n412160 );
buf ( n412162 , n396621 );
buf ( n412163 , n395890 );
and ( n412164 , n412162 , n412163 );
nor ( n89633 , n412161 , n412164 );
buf ( n89634 , n89633 );
buf ( n412167 , n89634 );
buf ( n412168 , n394838 );
or ( n89637 , n412167 , n412168 );
buf ( n412170 , n410325 );
buf ( n412171 , n394835 );
or ( n412172 , n412170 , n412171 );
nand ( n412173 , n89637 , n412172 );
buf ( n412174 , n412173 );
buf ( n412175 , n412174 );
xor ( n89644 , n412158 , n412175 );
xor ( n89645 , n410351 , n410354 );
xor ( n89646 , n89645 , n410409 );
buf ( n412179 , n89646 );
buf ( n412180 , n412179 );
and ( n412181 , n89644 , n412180 );
and ( n89650 , n412158 , n412175 );
or ( n89651 , n412181 , n89650 );
buf ( n412184 , n89651 );
buf ( n412185 , n412184 );
and ( n412186 , n412088 , n412185 );
and ( n89655 , n411991 , n412087 );
or ( n89656 , n412186 , n89655 );
buf ( n412189 , n89656 );
buf ( n412190 , n412189 );
xor ( n89659 , n411986 , n412190 );
xor ( n89660 , n411995 , n412012 );
xor ( n89661 , n89660 , n412082 );
buf ( n412194 , n89661 );
buf ( n412195 , n384414 );
buf ( n412196 , n79312 );
buf ( n412197 , n394724 );
and ( n89666 , n412196 , n412197 );
buf ( n412199 , n79318 );
buf ( n412200 , n384421 );
and ( n89669 , n412199 , n412200 );
nor ( n412202 , n89666 , n89669 );
buf ( n412203 , n412202 );
buf ( n412204 , n412203 );
or ( n412205 , n412195 , n412204 );
buf ( n89674 , n412003 );
buf ( n412207 , n395635 );
or ( n412208 , n89674 , n412207 );
nand ( n412209 , n412205 , n412208 );
buf ( n412210 , n412209 );
xor ( n89679 , n412042 , n412061 );
xor ( n412212 , n89679 , n412078 );
and ( n412213 , n412210 , n412212 );
buf ( n412214 , n394840 );
buf ( n412215 , n79114 );
and ( n412216 , n412214 , n412215 );
not ( n89685 , n412214 );
buf ( n412218 , n400487 );
and ( n412219 , n89685 , n412218 );
nor ( n89688 , n412216 , n412219 );
buf ( n412221 , n89688 );
buf ( n412222 , n412221 );
buf ( n412223 , n394838 );
or ( n412224 , n412222 , n412223 );
buf ( n412225 , n89634 );
buf ( n412226 , n394835 );
or ( n89695 , n412225 , n412226 );
nand ( n89696 , n412224 , n89695 );
buf ( n412229 , n89696 );
xor ( n412230 , n412042 , n412061 );
xor ( n89699 , n412230 , n412078 );
and ( n412232 , n412229 , n89699 );
and ( n412233 , n412210 , n412229 );
or ( n89702 , n412213 , n412232 , n412233 );
xor ( n412235 , n412194 , n89702 );
xor ( n412236 , n412158 , n412175 );
xor ( n412237 , n412236 , n412180 );
buf ( n412238 , n412237 );
and ( n412239 , n412235 , n412238 );
and ( n412240 , n412194 , n89702 );
or ( n89709 , n412239 , n412240 );
buf ( n412242 , n89709 );
xor ( n412243 , n410334 , n410414 );
xor ( n412244 , n412243 , n410419 );
buf ( n412245 , n412244 );
buf ( n412246 , n412245 );
xor ( n89715 , n412242 , n412246 );
xor ( n89716 , n411991 , n412087 );
xor ( n412249 , n89716 , n412185 );
buf ( n412250 , n412249 );
buf ( n412251 , n412250 );
and ( n89720 , n89715 , n412251 );
and ( n89721 , n412242 , n412246 );
or ( n412254 , n89720 , n89721 );
buf ( n412255 , n412254 );
buf ( n412256 , n412255 );
and ( n412257 , n89659 , n412256 );
and ( n412258 , n411986 , n412190 );
or ( n89727 , n412257 , n412258 );
buf ( n412260 , n89727 );
buf ( n89729 , n412260 );
xor ( n412262 , n410435 , n410440 );
xor ( n89731 , n412262 , n410446 );
buf ( n412264 , n89731 );
buf ( n412265 , n412264 );
xor ( n89734 , n89729 , n412265 );
buf ( n412267 , n76050 );
not ( n412268 , n412267 );
buf ( n412269 , n411835 );
not ( n89738 , n412269 );
or ( n89739 , n412268 , n89738 );
buf ( n412272 , n377583 );
not ( n89741 , n412272 );
buf ( n412274 , n377776 );
not ( n412275 , n412274 );
or ( n89744 , n89741 , n412275 );
buf ( n412277 , n377776 );
not ( n89746 , n412277 );
buf ( n412279 , n89746 );
buf ( n412280 , n412279 );
buf ( n412281 , n88904 );
nand ( n89750 , n412280 , n412281 );
buf ( n412283 , n89750 );
buf ( n412284 , n412283 );
nand ( n89753 , n89744 , n412284 );
buf ( n412286 , n89753 );
buf ( n412287 , n412286 );
buf ( n412288 , n85179 );
nand ( n89757 , n412287 , n412288 );
buf ( n412290 , n89757 );
buf ( n412291 , n412290 );
nand ( n412292 , n89739 , n412291 );
buf ( n412293 , n412292 );
buf ( n412294 , n412293 );
and ( n412295 , n89734 , n412294 );
and ( n89764 , n89729 , n412265 );
or ( n89765 , n412295 , n89764 );
buf ( n412298 , n89765 );
buf ( n412299 , n412298 );
not ( n89768 , n412299 );
buf ( n412301 , n377122 );
not ( n412302 , n412301 );
buf ( n412303 , n44906 );
not ( n89772 , n412303 );
or ( n412305 , n412302 , n89772 );
buf ( n412306 , n409022 );
buf ( n412307 , n57463 );
nand ( n412308 , n412306 , n412307 );
buf ( n412309 , n412308 );
buf ( n412310 , n412309 );
nand ( n412311 , n412305 , n412310 );
buf ( n412312 , n412311 );
buf ( n412313 , n412312 );
not ( n89782 , n412313 );
buf ( n412315 , n368599 );
not ( n89784 , n412315 );
or ( n89785 , n89782 , n89784 );
buf ( n412318 , n411460 );
buf ( n412319 , n368593 );
not ( n412320 , n412319 );
buf ( n412321 , n412320 );
buf ( n412322 , n412321 );
nand ( n89791 , n412318 , n412322 );
buf ( n412324 , n89791 );
buf ( n412325 , n412324 );
nand ( n412326 , n89785 , n412325 );
buf ( n412327 , n412326 );
buf ( n412328 , n412327 );
not ( n89797 , n412328 );
or ( n89798 , n89768 , n89797 );
buf ( n412331 , n412327 );
buf ( n412332 , n412298 );
or ( n89801 , n412331 , n412332 );
xor ( n89802 , n411791 , n89288 );
xor ( n89803 , n89802 , n411843 );
buf ( n412336 , n89803 );
buf ( n412337 , n412336 );
nand ( n89806 , n89801 , n412337 );
buf ( n412339 , n89806 );
buf ( n412340 , n412339 );
nand ( n412341 , n89798 , n412340 );
buf ( n412342 , n412341 );
buf ( n412343 , n412342 );
xor ( n89812 , n411420 , n411447 );
xor ( n89813 , n89812 , n411473 );
buf ( n412346 , n89813 );
buf ( n412347 , n412346 );
xor ( n89816 , n412343 , n412347 );
buf ( n412349 , n342475 );
buf ( n412350 , n402190 );
nor ( n412351 , n412349 , n412350 );
buf ( n412352 , n412351 );
buf ( n412353 , n412352 );
buf ( n412354 , n379515 );
or ( n89823 , n412353 , n412354 );
buf ( n412356 , n342475 );
buf ( n89825 , n402190 );
nand ( n89826 , n412356 , n89825 );
buf ( n412359 , n89826 );
buf ( n412360 , n412359 );
nand ( n89829 , n89823 , n412360 );
buf ( n412362 , n89829 );
buf ( n412363 , n412362 );
buf ( n412364 , n394065 );
nor ( n89833 , n412363 , n412364 );
buf ( n412366 , n89833 );
buf ( n412367 , n412366 );
and ( n89836 , n89816 , n412367 );
and ( n89837 , n412343 , n412347 );
or ( n412370 , n89836 , n89837 );
buf ( n412371 , n412370 );
buf ( n412372 , n412371 );
nand ( n89841 , n89452 , n412372 );
buf ( n412374 , n89841 );
buf ( n412375 , n412374 );
buf ( n412376 , n411970 );
not ( n89845 , n412376 );
buf ( n412378 , n411975 );
nand ( n89847 , n89845 , n412378 );
buf ( n412380 , n89847 );
buf ( n412381 , n412380 );
nand ( n89850 , n412375 , n412381 );
buf ( n412383 , n89850 );
buf ( n412384 , n412383 );
nand ( n89853 , n411966 , n412384 );
buf ( n412386 , n89853 );
buf ( n412387 , n412386 );
nand ( n89856 , n411963 , n412387 );
buf ( n412389 , n89856 );
buf ( n412390 , n412389 );
and ( n89859 , n411914 , n412390 );
and ( n89860 , n411909 , n411913 );
or ( n89861 , n89859 , n89860 );
buf ( n412394 , n89861 );
buf ( n412395 , n412394 );
xor ( n89864 , n411146 , n411150 );
xor ( n89865 , n89864 , n411177 );
buf ( n412398 , n89865 );
buf ( n412399 , n412398 );
xor ( n412400 , n412395 , n412399 );
xor ( n412401 , n411335 , n411538 );
xor ( n89870 , n412401 , n411546 );
buf ( n412403 , n89870 );
buf ( n412404 , n412403 );
and ( n89873 , n412400 , n412404 );
and ( n89874 , n412395 , n412399 );
or ( n89875 , n89873 , n89874 );
buf ( n412408 , n89875 );
buf ( n412409 , n412408 );
xor ( n412410 , n411735 , n412409 );
xor ( n89879 , n411310 , n411551 );
xor ( n412412 , n89879 , n411555 );
buf ( n412413 , n412412 );
buf ( n412414 , n412413 );
and ( n89883 , n412410 , n412414 );
and ( n412416 , n411735 , n412409 );
or ( n89885 , n89883 , n412416 );
buf ( n412418 , n89885 );
buf ( n412419 , n412418 );
xor ( n89888 , n411731 , n412419 );
xor ( n89889 , n411560 , n411702 );
xor ( n89890 , n89889 , n411707 );
buf ( n412423 , n89890 );
buf ( n412424 , n412423 );
and ( n412425 , n89888 , n412424 );
and ( n89894 , n411731 , n412419 );
or ( n412427 , n412425 , n89894 );
buf ( n412428 , n412427 );
buf ( n412429 , n412428 );
nand ( n412430 , n411727 , n412429 );
buf ( n412431 , n412430 );
buf ( n412432 , n412431 );
not ( n89901 , n412432 );
xor ( n412434 , n411712 , n411719 );
and ( n412435 , n412434 , n411724 );
and ( n89904 , n411712 , n411719 );
or ( n412437 , n412435 , n89904 );
buf ( n412438 , n412437 );
not ( n89907 , n412438 );
not ( n412440 , n411266 );
and ( n89909 , n88676 , n412440 );
not ( n412442 , n88676 );
and ( n89911 , n412442 , n411266 );
nor ( n412444 , n89909 , n89911 );
and ( n89913 , n412444 , n411208 );
not ( n412446 , n412444 );
not ( n89915 , n411208 );
and ( n89916 , n412446 , n89915 );
nor ( n412449 , n89913 , n89916 );
not ( n412450 , n412449 );
nand ( n89919 , n89907 , n412450 );
buf ( n412452 , n89919 );
nand ( n412453 , n89901 , n412452 );
buf ( n412454 , n412453 );
buf ( n412455 , n412454 );
nand ( n412456 , n412438 , n412449 );
buf ( n412457 , n412456 );
nand ( n89926 , n411285 , n412455 , n412457 );
buf ( n412459 , n89926 );
buf ( n412460 , n412459 );
not ( n89929 , n412460 );
or ( n412462 , n411280 , n89929 );
xor ( n412463 , n411564 , n411589 );
xor ( n89932 , n412463 , n411697 );
buf ( n412465 , n89932 );
buf ( n412466 , n412465 );
buf ( n412467 , n380356 );
not ( n89936 , n412467 );
buf ( n412469 , n411581 );
not ( n89938 , n412469 );
or ( n89939 , n89936 , n89938 );
buf ( n412472 , n380368 );
not ( n412473 , n412472 );
buf ( n412474 , n386837 );
not ( n412475 , n412474 );
or ( n412476 , n412473 , n412475 );
buf ( n412477 , n32202 );
buf ( n412478 , n380368 );
not ( n412479 , n412478 );
buf ( n412480 , n412479 );
buf ( n89943 , n412480 );
nand ( n89944 , n412477 , n89943 );
buf ( n412483 , n89944 );
buf ( n412484 , n412483 );
nand ( n89947 , n412476 , n412484 );
buf ( n412486 , n89947 );
buf ( n412487 , n412486 );
buf ( n412488 , n380404 );
nand ( n89951 , n412487 , n412488 );
buf ( n412490 , n89951 );
buf ( n412491 , n412490 );
nand ( n412492 , n89939 , n412491 );
buf ( n412493 , n412492 );
buf ( n412494 , n412493 );
xor ( n412495 , n411382 , n411407 );
xor ( n89958 , n412495 , n411533 );
buf ( n412497 , n89958 );
buf ( n412498 , n412497 );
buf ( n412499 , n380356 );
not ( n89962 , n412499 );
buf ( n412501 , n412486 );
not ( n412502 , n412501 );
or ( n89965 , n89962 , n412502 );
buf ( n412504 , n380368 );
not ( n412505 , n412504 );
buf ( n412506 , n382496 );
not ( n89969 , n412506 );
or ( n412508 , n412505 , n89969 );
buf ( n412509 , n378736 );
buf ( n412510 , n412480 );
nand ( n412511 , n412509 , n412510 );
buf ( n412512 , n412511 );
buf ( n412513 , n412512 );
nand ( n412514 , n412508 , n412513 );
buf ( n412515 , n412514 );
buf ( n412516 , n412515 );
buf ( n412517 , n380404 );
nand ( n89980 , n412516 , n412517 );
buf ( n89981 , n89980 );
buf ( n412520 , n89981 );
nand ( n89983 , n89965 , n412520 );
buf ( n412522 , n89983 );
buf ( n412523 , n412522 );
xor ( n412524 , n412498 , n412523 );
xor ( n89987 , n411412 , n411509 );
xor ( n89988 , n89987 , n411528 );
buf ( n412527 , n89988 );
xor ( n89990 , n377094 , n65349 );
buf ( n412529 , n89990 );
not ( n412530 , n412529 );
buf ( n412531 , n400929 );
not ( n89994 , n412531 );
or ( n89995 , n412530 , n89994 );
buf ( n412534 , n89218 );
buf ( n412535 , n365242 );
nand ( n89998 , n412534 , n412535 );
buf ( n412537 , n89998 );
buf ( n412538 , n412537 );
nand ( n90001 , n89995 , n412538 );
buf ( n412540 , n90001 );
buf ( n412541 , n412540 );
not ( n90004 , n412541 );
buf ( n412543 , n90004 );
buf ( n412544 , n412543 );
not ( n412545 , n412544 );
buf ( n412546 , n379890 );
not ( n90009 , n412546 );
buf ( n412548 , n89402 );
not ( n412549 , n412548 );
or ( n90012 , n90009 , n412549 );
buf ( n412551 , n379838 );
not ( n412552 , n412551 );
buf ( n412553 , n402185 );
not ( n412554 , n412553 );
or ( n412555 , n412552 , n412554 );
buf ( n412556 , n398741 );
buf ( n412557 , n31311 );
nand ( n412558 , n412556 , n412557 );
buf ( n412559 , n412558 );
buf ( n412560 , n412559 );
nand ( n90023 , n412555 , n412560 );
buf ( n412562 , n90023 );
buf ( n412563 , n412562 );
buf ( n412564 , n411170 );
nand ( n412565 , n412563 , n412564 );
buf ( n412566 , n412565 );
buf ( n412567 , n412566 );
nand ( n412568 , n90012 , n412567 );
buf ( n412569 , n412568 );
buf ( n412570 , n412569 );
not ( n412571 , n412570 );
buf ( n412572 , n412571 );
buf ( n412573 , n412572 );
not ( n412574 , n412573 );
or ( n412575 , n412545 , n412574 );
not ( n90038 , n58770 );
not ( n412577 , n90038 );
not ( n412578 , n411861 );
or ( n412579 , n412577 , n412578 );
buf ( n412580 , n377571 );
not ( n412581 , n412580 );
buf ( n412582 , n369372 );
not ( n412583 , n412582 );
or ( n90046 , n412581 , n412583 );
buf ( n412585 , n379268 );
buf ( n412586 , n352353 );
nand ( n412587 , n412585 , n412586 );
buf ( n412588 , n412587 );
buf ( n412589 , n412588 );
nand ( n412590 , n90046 , n412589 );
buf ( n412591 , n412590 );
nand ( n412592 , n412591 , n379962 );
nand ( n412593 , n412579 , n412592 );
buf ( n412594 , n377140 );
not ( n90057 , n412594 );
buf ( n412596 , n368561 );
not ( n90059 , n412596 );
or ( n90060 , n90057 , n90059 );
buf ( n412599 , n410287 );
buf ( n412600 , n377140 );
not ( n90063 , n412600 );
buf ( n412602 , n90063 );
buf ( n412603 , n412602 );
nand ( n412604 , n412599 , n412603 );
buf ( n412605 , n412604 );
buf ( n412606 , n412605 );
nand ( n90069 , n90060 , n412606 );
buf ( n412608 , n90069 );
buf ( n412609 , n412608 );
not ( n90072 , n412609 );
buf ( n412611 , n369801 );
not ( n412612 , n412611 );
or ( n90075 , n90072 , n412612 );
buf ( n412614 , n411804 );
buf ( n412615 , n369809 );
nand ( n412616 , n412614 , n412615 );
buf ( n412617 , n412616 );
buf ( n412618 , n412617 );
nand ( n90081 , n90075 , n412618 );
buf ( n412620 , n90081 );
xor ( n90083 , n411986 , n412190 );
xor ( n412622 , n90083 , n412256 );
buf ( n412623 , n412622 );
not ( n412624 , n76050 );
not ( n412625 , n412286 );
or ( n90088 , n412624 , n412625 );
buf ( n412627 , n407553 );
buf ( n412628 , n351013 );
not ( n90091 , n412628 );
buf ( n90092 , n90091 );
buf ( n412631 , n90092 );
not ( n90094 , n412631 );
buf ( n412633 , n49582 );
not ( n412634 , n412633 );
or ( n90097 , n90094 , n412634 );
buf ( n412636 , n377612 );
buf ( n412637 , n377754 );
nand ( n412638 , n412636 , n412637 );
buf ( n412639 , n412638 );
buf ( n412640 , n412639 );
nand ( n412641 , n90097 , n412640 );
buf ( n412642 , n412641 );
buf ( n412643 , n412642 );
nand ( n90106 , n412627 , n412643 );
buf ( n412645 , n90106 );
nand ( n90108 , n90088 , n412645 );
xor ( n90109 , n412623 , n90108 );
buf ( n412648 , n80468 );
buf ( n412649 , n384421 );
not ( n90112 , n412649 );
buf ( n90113 , n90112 );
buf ( n412652 , n90113 );
and ( n90115 , n412648 , n412652 );
buf ( n412654 , n401921 );
buf ( n412655 , n384421 );
and ( n90118 , n412654 , n412655 );
nor ( n90119 , n90115 , n90118 );
buf ( n412658 , n90119 );
buf ( n412659 , n412658 );
buf ( n412660 , n384414 );
or ( n412661 , n412659 , n412660 );
buf ( n90124 , n412203 );
buf ( n412663 , n395635 );
or ( n412664 , n90124 , n412663 );
nand ( n412665 , n412661 , n412664 );
buf ( n412666 , n412665 );
buf ( n412667 , n412666 );
xor ( n412668 , n412018 , n412040 );
buf ( n412669 , n412668 );
buf ( n412670 , n412669 );
xor ( n412671 , n412667 , n412670 );
buf ( n412672 , n382849 );
buf ( n412673 , n382638 );
buf ( n412674 , n405813 );
and ( n90137 , n412673 , n412674 );
buf ( n412676 , n382647 );
buf ( n412677 , n405816 );
and ( n90140 , n412676 , n412677 );
nor ( n412679 , n90137 , n90140 );
buf ( n412680 , n412679 );
buf ( n412681 , n412680 );
or ( n412682 , n412672 , n412681 );
buf ( n412683 , n412026 );
buf ( n412684 , n382634 );
or ( n90147 , n412683 , n412684 );
nand ( n412686 , n412682 , n90147 );
buf ( n412687 , n412686 );
buf ( n412688 , n57969 );
buf ( n412689 , n623 );
and ( n412690 , n412688 , n412689 );
buf ( n412691 , n378458 );
buf ( n412692 , n85590 );
and ( n90155 , n412691 , n412692 );
buf ( n412694 , n406588 );
nor ( n90157 , n90155 , n412694 );
buf ( n412696 , n90157 );
buf ( n412697 , n412696 );
buf ( n412698 , n57789 );
nor ( n90161 , n412690 , n412697 , n412698 );
buf ( n412700 , n90161 );
xor ( n90163 , n412687 , n412700 );
buf ( n412702 , n406588 );
buf ( n412703 , n406746 );
and ( n412704 , n412702 , n412703 );
buf ( n412705 , n82201 );
buf ( n412706 , n406749 );
and ( n412707 , n412705 , n412706 );
nor ( n90170 , n412704 , n412707 );
buf ( n412709 , n90170 );
buf ( n412710 , n412709 );
not ( n90173 , n412710 );
buf ( n412712 , n90173 );
buf ( n412713 , n412712 );
not ( n90176 , n412713 );
buf ( n412715 , n380735 );
not ( n412716 , n412715 );
or ( n90179 , n90176 , n412716 );
buf ( n412718 , n412122 );
buf ( n412719 , n380733 );
or ( n412720 , n412718 , n412719 );
nand ( n412721 , n90179 , n412720 );
buf ( n412722 , n412721 );
and ( n412723 , n90163 , n412722 );
and ( n412724 , n412687 , n412700 );
or ( n90187 , n412723 , n412724 );
buf ( n412726 , n90187 );
and ( n412727 , n412671 , n412726 );
and ( n90190 , n412667 , n412670 );
or ( n412729 , n412727 , n90190 );
buf ( n412730 , n412729 );
xor ( n412731 , n412142 , n89618 );
xor ( n90194 , n412731 , n412154 );
and ( n90195 , n412730 , n90194 );
buf ( n412734 , n378473 );
buf ( n412735 , n623 );
or ( n412736 , n412734 , n412735 );
buf ( n412737 , n378468 );
buf ( n412738 , n57789 );
buf ( n412739 , n623 );
and ( n412740 , n412737 , n412738 , n412739 );
buf ( n412741 , n378480 );
nor ( n412742 , n412740 , n412741 );
buf ( n412743 , n412742 );
buf ( n412744 , n412743 );
nand ( n412745 , n412736 , n412744 );
buf ( n412746 , n412745 );
buf ( n412747 , n384354 );
buf ( n412748 , n382627 );
buf ( n412749 , n403772 );
and ( n412750 , n412748 , n412749 );
buf ( n412751 , n403775 );
buf ( n412752 , n384089 );
and ( n412753 , n412751 , n412752 );
nor ( n90216 , n412750 , n412753 );
buf ( n412755 , n90216 );
buf ( n412756 , n412755 );
or ( n90219 , n412747 , n412756 );
buf ( n412758 , n412097 );
buf ( n412759 , n384082 );
or ( n412760 , n412758 , n412759 );
nand ( n90223 , n90219 , n412760 );
buf ( n412762 , n90223 );
xor ( n412763 , n412746 , n412762 );
buf ( n412764 , n378476 );
buf ( n412765 , n85590 );
nor ( n412766 , n412764 , n412765 );
buf ( n412767 , n412766 );
buf ( n412768 , n412767 );
buf ( n412769 , n382849 );
buf ( n412770 , n382638 );
buf ( n412771 , n406569 );
and ( n90234 , n412770 , n412771 );
buf ( n412773 , n382647 );
buf ( n412774 , n406572 );
and ( n90237 , n412773 , n412774 );
nor ( n412776 , n90234 , n90237 );
buf ( n412777 , n412776 );
buf ( n412778 , n412777 );
or ( n412779 , n412769 , n412778 );
buf ( n412780 , n412680 );
buf ( n412781 , n382634 );
or ( n412782 , n412780 , n412781 );
nand ( n412783 , n412779 , n412782 );
buf ( n412784 , n412783 );
buf ( n412785 , n412784 );
and ( n90245 , n412768 , n412785 );
buf ( n412787 , n90245 );
and ( n412788 , n412763 , n412787 );
and ( n412789 , n412746 , n412762 );
or ( n90249 , n412788 , n412789 );
buf ( n412791 , n90249 );
buf ( n412792 , n400503 );
buf ( n412793 , n394840 );
and ( n90253 , n412792 , n412793 );
buf ( n412795 , n400509 );
buf ( n412796 , n384408 );
and ( n90256 , n412795 , n412796 );
nor ( n412798 , n90253 , n90256 );
buf ( n412799 , n412798 );
buf ( n412800 , n412799 );
buf ( n412801 , n394838 );
or ( n90261 , n412800 , n412801 );
buf ( n412803 , n412221 );
buf ( n412804 , n394835 );
or ( n412805 , n412803 , n412804 );
nand ( n90265 , n90261 , n412805 );
buf ( n412807 , n90265 );
buf ( n412808 , n412807 );
xor ( n90268 , n412791 , n412808 );
xor ( n412810 , n412113 , n412130 );
xor ( n90270 , n412810 , n412138 );
buf ( n412812 , n90270 );
buf ( n412813 , n412812 );
and ( n412814 , n90268 , n412813 );
and ( n412815 , n412791 , n412808 );
or ( n90275 , n412814 , n412815 );
buf ( n412817 , n90275 );
xor ( n412818 , n412142 , n89618 );
xor ( n90278 , n412818 , n412154 );
and ( n412820 , n412817 , n90278 );
and ( n412821 , n412730 , n412817 );
or ( n90281 , n90195 , n412820 , n412821 );
xor ( n412823 , n412194 , n89702 );
xor ( n412824 , n412823 , n412238 );
and ( n90284 , n90281 , n412824 );
xor ( n90285 , n412667 , n412670 );
xor ( n412827 , n90285 , n412726 );
buf ( n412828 , n412827 );
buf ( n412829 , n81950 );
buf ( n412830 , n90113 );
and ( n412831 , n412829 , n412830 );
buf ( n412832 , n403589 );
buf ( n412833 , n384421 );
and ( n412834 , n412832 , n412833 );
nor ( n90294 , n412831 , n412834 );
buf ( n412836 , n90294 );
buf ( n412837 , n412836 );
buf ( n412838 , n384414 );
or ( n412839 , n412837 , n412838 );
buf ( n412840 , n412658 );
buf ( n412841 , n395635 );
or ( n412842 , n412840 , n412841 );
nand ( n412843 , n412839 , n412842 );
buf ( n412844 , n412843 );
xor ( n412845 , n412687 , n412700 );
xor ( n412846 , n412845 , n412722 );
and ( n90306 , n412844 , n412846 );
buf ( n412848 , n81995 );
buf ( n412849 , n90113 );
and ( n90309 , n412848 , n412849 );
buf ( n412851 , n403645 );
buf ( n412852 , n384421 );
and ( n412853 , n412851 , n412852 );
nor ( n90313 , n90309 , n412853 );
buf ( n412855 , n90313 );
buf ( n412856 , n412855 );
buf ( n412857 , n384414 );
or ( n90317 , n412856 , n412857 );
buf ( n412859 , n412836 );
buf ( n412860 , n395635 );
or ( n90320 , n412859 , n412860 );
nand ( n90321 , n90317 , n90320 );
buf ( n90322 , n90321 );
buf ( n412864 , n90322 );
buf ( n412865 , n384354 );
buf ( n412866 , n382627 );
buf ( n412867 , n403795 );
and ( n90327 , n412866 , n412867 );
buf ( n412869 , n62026 );
buf ( n412870 , n403798 );
and ( n90330 , n412869 , n412870 );
nor ( n90331 , n90327 , n90330 );
buf ( n412873 , n90331 );
buf ( n412874 , n412873 );
or ( n412875 , n412865 , n412874 );
buf ( n412876 , n412755 );
buf ( n412877 , n384082 );
or ( n412878 , n412876 , n412877 );
nand ( n90338 , n412875 , n412878 );
buf ( n412880 , n90338 );
buf ( n412881 , n412880 );
xor ( n412882 , n412864 , n412881 );
buf ( n412883 , n412709 );
buf ( n412884 , n380733 );
or ( n412885 , n412883 , n412884 );
buf ( n412886 , n60226 );
nand ( n90346 , n412885 , n412886 );
buf ( n412888 , n90346 );
buf ( n412889 , n412888 );
and ( n90349 , n412882 , n412889 );
and ( n412891 , n412864 , n412881 );
or ( n412892 , n90349 , n412891 );
buf ( n412893 , n412892 );
xor ( n90353 , n412687 , n412700 );
xor ( n412895 , n90353 , n412722 );
and ( n412896 , n412893 , n412895 );
and ( n90356 , n412844 , n412893 );
or ( n90357 , n90306 , n412896 , n90356 );
xor ( n412899 , n412828 , n90357 );
xor ( n412900 , n412791 , n412808 );
xor ( n90360 , n412900 , n412813 );
buf ( n412902 , n90360 );
and ( n90362 , n412899 , n412902 );
and ( n90363 , n412828 , n90357 );
or ( n412905 , n90362 , n90363 );
buf ( n412906 , n412905 );
xor ( n412907 , n412042 , n412061 );
xor ( n90367 , n412907 , n412078 );
xor ( n90368 , n412210 , n412229 );
xor ( n412910 , n90367 , n90368 );
buf ( n90370 , n412910 );
xor ( n90371 , n412906 , n90370 );
xor ( n412913 , n412142 , n89618 );
xor ( n412914 , n412913 , n412154 );
xor ( n90374 , n412730 , n412817 );
xor ( n412916 , n412914 , n90374 );
buf ( n412917 , n412916 );
and ( n412918 , n90371 , n412917 );
and ( n90378 , n412906 , n90370 );
or ( n412920 , n412918 , n90378 );
buf ( n412921 , n412920 );
xor ( n90381 , n412194 , n89702 );
xor ( n412923 , n90381 , n412238 );
and ( n412924 , n412921 , n412923 );
and ( n412925 , n90281 , n412921 );
or ( n90385 , n90284 , n412924 , n412925 );
buf ( n412927 , n90385 );
xor ( n412928 , n412242 , n412246 );
xor ( n412929 , n412928 , n412251 );
buf ( n412930 , n412929 );
buf ( n412931 , n412930 );
xor ( n412932 , n412927 , n412931 );
buf ( n90392 , n377140 );
not ( n90393 , n90392 );
buf ( n90394 , n411431 );
not ( n90395 , n90394 );
or ( n90396 , n90393 , n90395 );
buf ( n412938 , n377612 );
not ( n412939 , n412938 );
buf ( n412940 , n412939 );
buf ( n412941 , n412940 );
buf ( n412942 , n412602 );
nand ( n412943 , n412941 , n412942 );
buf ( n412944 , n412943 );
buf ( n412945 , n412944 );
nand ( n412946 , n90396 , n412945 );
buf ( n412947 , n412946 );
buf ( n412948 , n412947 );
not ( n90408 , n412948 );
buf ( n412950 , n407553 );
not ( n90410 , n412950 );
or ( n412952 , n90408 , n90410 );
buf ( n412953 , n57147 );
not ( n90413 , n412953 );
buf ( n412955 , n412642 );
nand ( n412956 , n90413 , n412955 );
buf ( n412957 , n412956 );
buf ( n412958 , n412957 );
nand ( n90418 , n412952 , n412958 );
buf ( n412960 , n90418 );
buf ( n412961 , n412960 );
and ( n412962 , n412932 , n412961 );
and ( n90422 , n412927 , n412931 );
or ( n90423 , n412962 , n90422 );
buf ( n412965 , n90423 );
and ( n412966 , n90109 , n412965 );
and ( n90426 , n412623 , n90108 );
or ( n412968 , n412966 , n90426 );
xor ( n412969 , n412620 , n412968 );
xor ( n90429 , n89729 , n412265 );
xor ( n412971 , n90429 , n412294 );
buf ( n412972 , n412971 );
and ( n90432 , n412969 , n412972 );
and ( n90433 , n412620 , n412968 );
or ( n90434 , n90432 , n90433 );
xor ( n90435 , n412593 , n90434 );
and ( n90436 , n378843 , n406953 );
not ( n90437 , n378843 );
and ( n90438 , n90437 , n406249 );
or ( n90439 , n90436 , n90438 );
buf ( n412981 , n90439 );
not ( n90441 , n412981 );
buf ( n412983 , n404115 );
not ( n90443 , n412983 );
or ( n90444 , n90441 , n90443 );
buf ( n412986 , n411871 );
buf ( n412987 , n44915 );
nand ( n412988 , n412986 , n412987 );
buf ( n412989 , n412988 );
buf ( n412990 , n412989 );
nand ( n90450 , n90444 , n412990 );
buf ( n412992 , n90450 );
and ( n90452 , n90435 , n412992 );
and ( n90453 , n412593 , n90434 );
or ( n90454 , n90452 , n90453 );
buf ( n412996 , n90454 );
buf ( n412997 , n379890 );
not ( n412998 , n412997 );
buf ( n412999 , n412562 );
not ( n413000 , n412999 );
or ( n90460 , n412998 , n413000 );
buf ( n413002 , n379838 );
not ( n90462 , n413002 );
buf ( n413004 , n365384 );
not ( n413005 , n413004 );
or ( n413006 , n90462 , n413005 );
buf ( n413007 , n84042 );
buf ( n413008 , n398741 );
nand ( n413009 , n413007 , n413008 );
buf ( n413010 , n413009 );
buf ( n413011 , n413010 );
nand ( n413012 , n413006 , n413011 );
buf ( n413013 , n413012 );
buf ( n413014 , n413013 );
buf ( n413015 , n411170 );
nand ( n413016 , n413014 , n413015 );
buf ( n413017 , n413016 );
buf ( n413018 , n413017 );
nand ( n413019 , n90460 , n413018 );
buf ( n413020 , n413019 );
buf ( n413021 , n413020 );
xor ( n413022 , n412996 , n413021 );
xor ( n413023 , n411848 , n411866 );
xor ( n90483 , n413023 , n411884 );
buf ( n413025 , n90483 );
buf ( n413026 , n413025 );
and ( n90486 , n413022 , n413026 );
and ( n413028 , n412996 , n413021 );
or ( n90488 , n90486 , n413028 );
buf ( n413030 , n90488 );
buf ( n413031 , n413030 );
nand ( n90491 , n412575 , n413031 );
buf ( n413033 , n90491 );
buf ( n413034 , n413033 );
buf ( n413035 , n412572 );
not ( n413036 , n413035 );
buf ( n413037 , n412540 );
nand ( n90497 , n413036 , n413037 );
buf ( n90498 , n90497 );
buf ( n413040 , n90498 );
nand ( n413041 , n413034 , n413040 );
buf ( n413042 , n413041 );
xor ( n413043 , n412527 , n413042 );
xor ( n413044 , n411760 , n89370 );
xor ( n90504 , n413044 , n411904 );
buf ( n413046 , n90504 );
and ( n413047 , n413043 , n413046 );
and ( n90507 , n412527 , n413042 );
or ( n413049 , n413047 , n90507 );
buf ( n413050 , n413049 );
and ( n90510 , n412524 , n413050 );
and ( n413052 , n412498 , n412523 );
or ( n413053 , n90510 , n413052 );
buf ( n413054 , n413053 );
buf ( n413055 , n413054 );
xor ( n90515 , n412494 , n413055 );
xor ( n90516 , n411594 , n411619 );
xor ( n90517 , n90516 , n411692 );
buf ( n413059 , n90517 );
buf ( n413060 , n413059 );
and ( n413061 , n90515 , n413060 );
and ( n413062 , n412494 , n413055 );
or ( n90522 , n413061 , n413062 );
buf ( n413064 , n90522 );
buf ( n413065 , n413064 );
xor ( n90525 , n412466 , n413065 );
xor ( n90526 , n411735 , n412409 );
xor ( n90527 , n90526 , n412414 );
buf ( n413069 , n90527 );
buf ( n413070 , n413069 );
and ( n413071 , n90525 , n413070 );
and ( n90531 , n412466 , n413065 );
or ( n90532 , n413071 , n90531 );
buf ( n413074 , n90532 );
buf ( n413075 , n413074 );
xor ( n90535 , n411731 , n412419 );
xor ( n413077 , n90535 , n412424 );
buf ( n413078 , n413077 );
buf ( n413079 , n413078 );
xor ( n90539 , n413075 , n413079 );
xor ( n413081 , n411909 , n411913 );
xor ( n90541 , n413081 , n412390 );
buf ( n413083 , n90541 );
buf ( n413084 , n413083 );
not ( n90544 , n413084 );
xor ( n90545 , n411676 , n411643 );
buf ( n413087 , n90545 );
not ( n90547 , n413087 );
buf ( n413089 , n411685 );
not ( n90549 , n413089 );
and ( n90550 , n90547 , n90549 );
buf ( n413092 , n411685 );
buf ( n413093 , n90545 );
and ( n90553 , n413092 , n413093 );
nor ( n90554 , n90550 , n90553 );
buf ( n413096 , n90554 );
buf ( n413097 , n413096 );
nand ( n90557 , n90544 , n413097 );
buf ( n413099 , n90557 );
not ( n90559 , n413099 );
buf ( n413101 , n58923 );
not ( n90561 , n413101 );
buf ( n413103 , n411657 );
not ( n90563 , n413103 );
or ( n90564 , n90561 , n90563 );
buf ( n413106 , n379368 );
not ( n90566 , n413106 );
buf ( n413108 , n381266 );
not ( n413109 , n413108 );
or ( n90569 , n90566 , n413109 );
buf ( n413111 , n351160 );
buf ( n413112 , n407228 );
nand ( n413113 , n413111 , n413112 );
buf ( n413114 , n413113 );
buf ( n413115 , n413114 );
nand ( n413116 , n90569 , n413115 );
buf ( n413117 , n413116 );
buf ( n413118 , n413117 );
buf ( n413119 , n379353 );
nand ( n413120 , n413118 , n413119 );
buf ( n413121 , n413120 );
buf ( n413122 , n413121 );
nand ( n413123 , n90564 , n413122 );
buf ( n413124 , n413123 );
buf ( n413125 , n413124 );
not ( n90585 , n413125 );
xor ( n413127 , n411960 , n411938 );
xor ( n413128 , n413127 , n412383 );
buf ( n413129 , n413128 );
not ( n413130 , n413129 );
or ( n413131 , n90585 , n413130 );
buf ( n413132 , n413128 );
buf ( n413133 , n413124 );
or ( n90593 , n413132 , n413133 );
xor ( n413135 , n411786 , n411889 );
xor ( n413136 , n413135 , n411894 );
buf ( n413137 , n413136 );
buf ( n413138 , n413137 );
not ( n413139 , n413138 );
buf ( n413140 , n411970 );
buf ( n413141 , n412371 );
xor ( n90601 , n413140 , n413141 );
buf ( n413143 , n411975 );
xor ( n90603 , n90601 , n413143 );
buf ( n413145 , n90603 );
buf ( n413146 , n413145 );
not ( n90606 , n413146 );
buf ( n413148 , n90606 );
buf ( n413149 , n413148 );
not ( n90609 , n413149 );
or ( n413151 , n413139 , n90609 );
buf ( n413152 , n413137 );
not ( n90612 , n413152 );
buf ( n413154 , n90612 );
not ( n413155 , n413154 );
not ( n90615 , n413145 );
or ( n413157 , n413155 , n90615 );
buf ( n413158 , n377068 );
not ( n90618 , n413158 );
buf ( n413160 , n22956 );
not ( n413161 , n413160 );
or ( n413162 , n90618 , n413161 );
buf ( n413163 , n402190 );
buf ( n413164 , n377071 );
nand ( n90624 , n413163 , n413164 );
buf ( n413166 , n90624 );
buf ( n413167 , n413166 );
nand ( n90627 , n413162 , n413167 );
buf ( n413169 , n90627 );
buf ( n90629 , n413169 );
not ( n90630 , n90629 );
buf ( n90631 , n411775 );
not ( n90632 , n90631 );
or ( n90633 , n90630 , n90632 );
buf ( n90634 , n89243 );
buf ( n90635 , n407713 );
nand ( n90636 , n90634 , n90635 );
buf ( n90637 , n90636 );
buf ( n90638 , n90637 );
nand ( n90639 , n90633 , n90638 );
buf ( n90640 , n90639 );
not ( n413182 , n90640 );
buf ( n413183 , n406249 );
buf ( n413184 , n342934 );
nand ( n413185 , n413183 , n413184 );
buf ( n413186 , n413185 );
buf ( n413187 , n413186 );
buf ( n413188 , n342934 );
buf ( n413189 , n342965 );
or ( n90649 , n413188 , n413189 );
buf ( n413191 , n378098 );
nand ( n90651 , n90649 , n413191 );
buf ( n413193 , n90651 );
buf ( n413194 , n413193 );
buf ( n413195 , n22954 );
nand ( n90655 , n413187 , n413194 , n413195 );
buf ( n413197 , n90655 );
buf ( n413198 , n413197 );
not ( n90658 , n413198 );
not ( n90659 , n90439 );
not ( n90660 , n44915 );
or ( n90661 , n90659 , n90660 );
and ( n90662 , n377068 , n369183 );
not ( n90663 , n377068 );
and ( n90664 , n90663 , n405357 );
or ( n90665 , n90662 , n90664 );
nand ( n90666 , n90665 , n404115 );
nand ( n90667 , n90661 , n90666 );
buf ( n413209 , n90667 );
not ( n90669 , n413209 );
buf ( n413211 , n90669 );
buf ( n413212 , n413211 );
not ( n90672 , n413212 );
or ( n90673 , n90658 , n90672 );
xor ( n90674 , n412620 , n412968 );
xor ( n90675 , n90674 , n412972 );
buf ( n413217 , n90675 );
nand ( n90677 , n90673 , n413217 );
buf ( n90678 , n90677 );
buf ( n413220 , n90678 );
buf ( n413221 , n90667 );
buf ( n413222 , n413197 );
not ( n90682 , n413222 );
buf ( n413224 , n90682 );
buf ( n413225 , n413224 );
nand ( n90685 , n413221 , n413225 );
buf ( n413227 , n90685 );
buf ( n413228 , n413227 );
nand ( n90688 , n413220 , n413228 );
buf ( n413230 , n90688 );
buf ( n413231 , n413230 );
not ( n90691 , n413231 );
buf ( n413233 , n379890 );
not ( n90693 , n413233 );
buf ( n413235 , n413013 );
not ( n413236 , n413235 );
or ( n90696 , n90693 , n413236 );
buf ( n413238 , n379838 );
not ( n413239 , n413238 );
buf ( n413240 , n408236 );
not ( n90700 , n413240 );
or ( n90701 , n413239 , n90700 );
buf ( n413243 , n368656 );
buf ( n413244 , n398741 );
nand ( n90704 , n413243 , n413244 );
buf ( n413246 , n90704 );
buf ( n413247 , n413246 );
nand ( n90707 , n90701 , n413247 );
buf ( n413249 , n90707 );
buf ( n413250 , n413249 );
buf ( n413251 , n411170 );
nand ( n413252 , n413250 , n413251 );
buf ( n413253 , n413252 );
buf ( n413254 , n413253 );
nand ( n413255 , n90696 , n413254 );
buf ( n413256 , n413255 );
buf ( n413257 , n413256 );
not ( n90717 , n413257 );
buf ( n413259 , n90717 );
buf ( n413260 , n413259 );
buf ( n413261 , n412298 );
buf ( n413262 , n412327 );
xor ( n413263 , n413261 , n413262 );
buf ( n413264 , n412336 );
xnor ( n413265 , n413263 , n413264 );
buf ( n413266 , n413265 );
buf ( n413267 , n413266 );
nand ( n413268 , n413260 , n413267 );
buf ( n413269 , n413268 );
buf ( n413270 , n413269 );
not ( n90730 , n413270 );
or ( n90731 , n90691 , n90730 );
buf ( n413273 , n413256 );
buf ( n413274 , n413266 );
not ( n90734 , n413274 );
buf ( n413276 , n90734 );
buf ( n413277 , n413276 );
nand ( n413278 , n413273 , n413277 );
buf ( n413279 , n413278 );
buf ( n413280 , n413279 );
nand ( n90740 , n90731 , n413280 );
buf ( n413282 , n90740 );
not ( n90742 , n413282 );
or ( n90743 , n413182 , n90742 );
not ( n90744 , n90640 );
not ( n90745 , n90744 );
not ( n90746 , n413282 );
not ( n413288 , n90746 );
or ( n90748 , n90745 , n413288 );
xor ( n413290 , n412343 , n412347 );
xor ( n413291 , n413290 , n412367 );
buf ( n413292 , n413291 );
nand ( n90752 , n90748 , n413292 );
nand ( n413294 , n90743 , n90752 );
nand ( n90754 , n413157 , n413294 );
buf ( n413296 , n90754 );
nand ( n413297 , n413151 , n413296 );
buf ( n413298 , n413297 );
buf ( n413299 , n413298 );
nand ( n413300 , n90593 , n413299 );
buf ( n413301 , n413300 );
buf ( n413302 , n413301 );
nand ( n413303 , n413131 , n413302 );
buf ( n413304 , n413303 );
not ( n413305 , n413304 );
or ( n413306 , n90559 , n413305 );
buf ( n413307 , n413096 );
not ( n413308 , n413307 );
buf ( n413309 , n413083 );
nand ( n90769 , n413308 , n413309 );
buf ( n413311 , n90769 );
nand ( n90771 , n413306 , n413311 );
buf ( n413313 , n90771 );
xor ( n90773 , n412395 , n412399 );
xor ( n90774 , n90773 , n412404 );
buf ( n413316 , n90774 );
buf ( n413317 , n413316 );
xor ( n90777 , n413313 , n413317 );
xor ( n90778 , n412494 , n413055 );
xor ( n90779 , n90778 , n413060 );
buf ( n413321 , n90779 );
buf ( n413322 , n413321 );
and ( n413323 , n90777 , n413322 );
and ( n90783 , n413313 , n413317 );
or ( n413325 , n413323 , n90783 );
buf ( n413326 , n413325 );
buf ( n413327 , n413326 );
xor ( n90787 , n412466 , n413065 );
xor ( n90788 , n90787 , n413070 );
buf ( n413330 , n90788 );
buf ( n413331 , n413330 );
xor ( n90791 , n413327 , n413331 );
xor ( n413333 , n412498 , n412523 );
xor ( n413334 , n413333 , n413050 );
buf ( n413335 , n413334 );
buf ( n413336 , n413335 );
not ( n90796 , n413336 );
xor ( n413338 , n413083 , n413096 );
xor ( n413339 , n413338 , n413304 );
buf ( n413340 , n413339 );
not ( n413341 , n413340 );
buf ( n413342 , n413341 );
buf ( n413343 , n413342 );
not ( n90803 , n413343 );
or ( n413345 , n90796 , n90803 );
buf ( n413346 , n413335 );
not ( n90806 , n413346 );
buf ( n90807 , n90806 );
not ( n90808 , n90807 );
not ( n90809 , n413339 );
or ( n90810 , n90808 , n90809 );
buf ( n413352 , n380356 );
not ( n90812 , n413352 );
buf ( n413354 , n412515 );
not ( n413355 , n413354 );
or ( n90815 , n90812 , n413355 );
buf ( n413357 , n380368 );
not ( n90817 , n413357 );
buf ( n413359 , n31194 );
not ( n413360 , n413359 );
or ( n413361 , n90817 , n413360 );
buf ( n413362 , n57233 );
buf ( n413363 , n412480 );
nand ( n413364 , n413362 , n413363 );
buf ( n413365 , n413364 );
buf ( n413366 , n413365 );
nand ( n90826 , n413361 , n413366 );
buf ( n413368 , n90826 );
buf ( n413369 , n413368 );
buf ( n413370 , n380404 );
nand ( n90830 , n413369 , n413370 );
buf ( n413372 , n90830 );
buf ( n413373 , n413372 );
nand ( n90833 , n90815 , n413373 );
buf ( n413375 , n90833 );
xor ( n90835 , n412527 , n413042 );
xor ( n90836 , n90835 , n413046 );
xor ( n413378 , n413375 , n90836 );
buf ( n413379 , n58923 );
not ( n90839 , n413379 );
buf ( n413381 , n413117 );
not ( n90841 , n413381 );
or ( n90842 , n90839 , n90841 );
and ( n413384 , n32234 , n379368 );
not ( n413385 , n32234 );
and ( n90845 , n413385 , n407228 );
or ( n413387 , n413384 , n90845 );
buf ( n413388 , n413387 );
buf ( n413389 , n379353 );
nand ( n413390 , n413388 , n413389 );
buf ( n413391 , n413390 );
buf ( n413392 , n413391 );
nand ( n413393 , n90842 , n413392 );
buf ( n413394 , n413393 );
buf ( n413395 , n413394 );
buf ( n413396 , n380356 );
not ( n90856 , n413396 );
buf ( n413398 , n413368 );
not ( n413399 , n413398 );
or ( n413400 , n90856 , n413399 );
buf ( n413401 , n412480 );
not ( n90861 , n413401 );
buf ( n413403 , n351195 );
not ( n413404 , n413403 );
or ( n90864 , n90861 , n413404 );
buf ( n413406 , n351195 );
buf ( n413407 , n412480 );
or ( n90867 , n413406 , n413407 );
nand ( n413409 , n90864 , n90867 );
buf ( n413410 , n413409 );
buf ( n413411 , n413410 );
buf ( n413412 , n380404 );
nand ( n413413 , n413411 , n413412 );
buf ( n413414 , n413413 );
buf ( n413415 , n413414 );
nand ( n90875 , n413400 , n413415 );
buf ( n413417 , n90875 );
buf ( n413418 , n413417 );
or ( n413419 , n413395 , n413418 );
buf ( n413420 , n378098 );
not ( n413421 , n413420 );
buf ( n413422 , n394065 );
not ( n90882 , n413422 );
or ( n413424 , n413421 , n90882 );
buf ( n413425 , n65349 );
buf ( n413426 , n379515 );
nand ( n90886 , n413425 , n413426 );
buf ( n413428 , n90886 );
buf ( n413429 , n413428 );
nand ( n413430 , n413424 , n413429 );
buf ( n413431 , n413430 );
buf ( n413432 , n413431 );
not ( n413433 , n413432 );
buf ( n413434 , n400929 );
not ( n413435 , n413434 );
or ( n90895 , n413433 , n413435 );
buf ( n413437 , n89990 );
buf ( n413438 , n365242 );
nand ( n90898 , n413437 , n413438 );
buf ( n413440 , n90898 );
buf ( n90900 , n413440 );
nand ( n90901 , n90895 , n90900 );
buf ( n90902 , n90901 );
buf ( n413444 , n90902 );
not ( n90904 , n413444 );
xor ( n413446 , n412996 , n413021 );
xor ( n90906 , n413446 , n413026 );
buf ( n413448 , n90906 );
buf ( n413449 , n413448 );
not ( n413450 , n413449 );
or ( n413451 , n90904 , n413450 );
buf ( n413452 , n413448 );
buf ( n413453 , n90902 );
or ( n413454 , n413452 , n413453 );
not ( n413455 , n379260 );
not ( n90915 , n412591 );
or ( n413457 , n413455 , n90915 );
buf ( n413458 , n377571 );
not ( n90918 , n413458 );
buf ( n413460 , n408201 );
not ( n90920 , n413460 );
or ( n90921 , n90918 , n90920 );
buf ( n413463 , n352381 );
buf ( n413464 , n379271 );
nand ( n90924 , n413463 , n413464 );
buf ( n413466 , n90924 );
buf ( n413467 , n413466 );
nand ( n90927 , n90921 , n413467 );
buf ( n413469 , n90927 );
buf ( n90929 , n413469 );
buf ( n413471 , n379962 );
nand ( n90931 , n90929 , n413471 );
buf ( n413473 , n90931 );
nand ( n90933 , n413457 , n413473 );
buf ( n413475 , n90933 );
not ( n90935 , n413475 );
buf ( n413477 , n58984 );
not ( n413478 , n413477 );
buf ( n413479 , n23037 );
not ( n90939 , n413479 );
buf ( n90940 , n90939 );
buf ( n413482 , n90940 );
not ( n90942 , n413482 );
or ( n413484 , n413478 , n90942 );
buf ( n413485 , n409022 );
buf ( n413486 , n408722 );
nand ( n90946 , n413485 , n413486 );
buf ( n413488 , n90946 );
buf ( n413489 , n413488 );
nand ( n90949 , n413484 , n413489 );
buf ( n90950 , n90949 );
not ( n413492 , n90950 );
buf ( n413493 , n48356 );
buf ( n413494 , n368593 );
and ( n413495 , n413493 , n413494 );
buf ( n413496 , n413495 );
not ( n90956 , n413496 );
or ( n413498 , n413492 , n90956 );
nand ( n90958 , n412312 , n369444 );
nand ( n413500 , n413498 , n90958 );
buf ( n413501 , n413500 );
not ( n90961 , n413501 );
or ( n413503 , n90935 , n90961 );
or ( n413504 , n413500 , n90933 );
buf ( n413505 , n379260 );
not ( n413506 , n413505 );
buf ( n413507 , n413469 );
not ( n90967 , n413507 );
or ( n413509 , n413506 , n90967 );
buf ( n413510 , n377571 );
not ( n90970 , n413510 );
buf ( n413512 , n377349 );
not ( n413513 , n413512 );
or ( n413514 , n90970 , n413513 );
buf ( n413515 , n409020 );
buf ( n413516 , n379268 );
nand ( n413517 , n413515 , n413516 );
buf ( n413518 , n413517 );
buf ( n413519 , n413518 );
nand ( n413520 , n413514 , n413519 );
buf ( n413521 , n413520 );
buf ( n413522 , n413521 );
buf ( n413523 , n379962 );
nand ( n413524 , n413522 , n413523 );
buf ( n413525 , n413524 );
buf ( n413526 , n413525 );
nand ( n413527 , n413509 , n413526 );
buf ( n413528 , n413527 );
not ( n413529 , n413528 );
buf ( n413530 , n377122 );
not ( n413531 , n413530 );
buf ( n413532 , n368561 );
not ( n413533 , n413532 );
or ( n90985 , n413531 , n413533 );
buf ( n413535 , n410287 );
buf ( n413536 , n57463 );
nand ( n413537 , n413535 , n413536 );
buf ( n413538 , n413537 );
buf ( n413539 , n413538 );
nand ( n413540 , n90985 , n413539 );
buf ( n413541 , n413540 );
buf ( n413542 , n413541 );
not ( n413543 , n413542 );
buf ( n413544 , n369801 );
not ( n413545 , n413544 );
or ( n413546 , n413543 , n413545 );
buf ( n413547 , n412608 );
buf ( n413548 , n369809 );
nand ( n413549 , n413547 , n413548 );
buf ( n413550 , n413549 );
buf ( n413551 , n413550 );
nand ( n91003 , n413546 , n413551 );
buf ( n413553 , n91003 );
not ( n91005 , n413553 );
or ( n91006 , n413529 , n91005 );
not ( n413556 , n413528 );
not ( n413557 , n413556 );
not ( n91009 , n413553 );
not ( n413559 , n91009 );
or ( n413560 , n413557 , n413559 );
xor ( n91012 , n412623 , n90108 );
xor ( n413562 , n91012 , n412965 );
nand ( n91014 , n413560 , n413562 );
nand ( n91015 , n91006 , n91014 );
nand ( n91016 , n413504 , n91015 );
buf ( n413566 , n91016 );
nand ( n91018 , n413503 , n413566 );
buf ( n413568 , n91018 );
buf ( n413569 , n413568 );
buf ( n413570 , n45052 );
buf ( n413571 , n378098 );
and ( n91023 , n413570 , n413571 );
buf ( n413573 , n91023 );
buf ( n413574 , n413573 );
xor ( n91026 , n413569 , n413574 );
xor ( n91027 , n412593 , n90434 );
xor ( n413577 , n91027 , n412992 );
buf ( n413578 , n413577 );
and ( n91030 , n91026 , n413578 );
and ( n91031 , n413569 , n413574 );
or ( n413581 , n91030 , n91031 );
buf ( n413582 , n413581 );
buf ( n413583 , n413582 );
nand ( n413584 , n413454 , n413583 );
buf ( n413585 , n413584 );
buf ( n413586 , n413585 );
nand ( n413587 , n413451 , n413586 );
buf ( n413588 , n413587 );
buf ( n413589 , n413588 );
nand ( n91041 , n413419 , n413589 );
buf ( n413591 , n91041 );
buf ( n413592 , n413591 );
buf ( n413593 , n413394 );
buf ( n413594 , n413417 );
nand ( n91046 , n413593 , n413594 );
buf ( n413596 , n91046 );
buf ( n413597 , n413596 );
nand ( n91049 , n413592 , n413597 );
buf ( n413599 , n91049 );
and ( n91051 , n413378 , n413599 );
and ( n413601 , n413375 , n90836 );
or ( n413602 , n91051 , n413601 );
nand ( n91054 , n90810 , n413602 );
buf ( n413604 , n91054 );
nand ( n413605 , n413345 , n413604 );
buf ( n413606 , n413605 );
buf ( n413607 , n413606 );
xor ( n91059 , n413313 , n413317 );
xor ( n413609 , n91059 , n413322 );
buf ( n413610 , n413609 );
buf ( n413611 , n413610 );
xor ( n413612 , n413607 , n413611 );
buf ( n413613 , n413124 );
buf ( n413614 , n413298 );
xor ( n91066 , n413613 , n413614 );
buf ( n413616 , n413128 );
xnor ( n91068 , n91066 , n413616 );
buf ( n413618 , n91068 );
buf ( n413619 , n413618 );
not ( n91071 , n413619 );
xor ( n413621 , n413375 , n90836 );
xor ( n91073 , n413621 , n413599 );
buf ( n413623 , n91073 );
not ( n91075 , n413623 );
buf ( n413625 , n91075 );
buf ( n413626 , n413625 );
not ( n91078 , n413626 );
or ( n91079 , n91071 , n91078 );
xor ( n91080 , n413137 , n413294 );
xnor ( n91081 , n91080 , n413148 );
buf ( n413631 , n91081 );
buf ( n413632 , n412569 );
buf ( n413633 , n412543 );
xor ( n413634 , n413632 , n413633 );
buf ( n413635 , n413030 );
xor ( n413636 , n413634 , n413635 );
buf ( n413637 , n413636 );
buf ( n413638 , n413637 );
or ( n413639 , n413631 , n413638 );
buf ( n413640 , n413639 );
buf ( n413641 , n413640 );
buf ( n413642 , n413637 );
not ( n91094 , n413642 );
buf ( n413644 , n91081 );
not ( n413645 , n413644 );
or ( n413646 , n91094 , n413645 );
buf ( n413647 , n58923 );
not ( n91099 , n413647 );
buf ( n413649 , n413387 );
not ( n413650 , n413649 );
or ( n91102 , n91099 , n413650 );
and ( n413652 , n31093 , n379365 );
not ( n413653 , n31093 );
and ( n91105 , n413653 , n379368 );
or ( n413655 , n413652 , n91105 );
buf ( n413656 , n413655 );
buf ( n413657 , n379353 );
nand ( n413658 , n413656 , n413657 );
buf ( n413659 , n413658 );
buf ( n413660 , n413659 );
nand ( n413661 , n91102 , n413660 );
buf ( n413662 , n413661 );
buf ( n413663 , n413662 );
not ( n413664 , n413663 );
not ( n91116 , n45010 );
buf ( n413666 , n91116 );
not ( n413667 , n413666 );
and ( n413668 , n377094 , n22956 );
not ( n91120 , n377094 );
and ( n91121 , n91120 , n402190 );
or ( n91122 , n413668 , n91121 );
buf ( n413672 , n91122 );
not ( n91124 , n413672 );
or ( n91125 , n413667 , n91124 );
buf ( n413675 , n365146 );
not ( n91127 , n413675 );
buf ( n413677 , n413169 );
nand ( n91129 , n91127 , n413677 );
buf ( n91130 , n91129 );
buf ( n413680 , n91130 );
nand ( n413681 , n91125 , n413680 );
buf ( n413682 , n413681 );
buf ( n413683 , n413682 );
buf ( n413684 , n379890 );
not ( n91136 , n413684 );
buf ( n413686 , n413249 );
not ( n91138 , n413686 );
or ( n413688 , n91136 , n91138 );
and ( n413689 , n351043 , n398741 );
not ( n413690 , n351043 );
and ( n91142 , n413690 , n379838 );
or ( n413692 , n413689 , n91142 );
buf ( n413693 , n413692 );
buf ( n413694 , n411170 );
nand ( n413695 , n413693 , n413694 );
buf ( n413696 , n413695 );
buf ( n413697 , n413696 );
nand ( n413698 , n413688 , n413697 );
buf ( n413699 , n413698 );
buf ( n91151 , n413699 );
not ( n91152 , n91151 );
and ( n413702 , n413500 , n90933 );
not ( n91154 , n413500 );
not ( n413704 , n90933 );
and ( n91156 , n91154 , n413704 );
nor ( n91157 , n413702 , n91156 );
xnor ( n91158 , n91015 , n91157 );
buf ( n413708 , n91158 );
not ( n91160 , n413708 );
buf ( n91161 , n91160 );
buf ( n91162 , n91161 );
not ( n91163 , n91162 );
or ( n91164 , n91152 , n91163 );
buf ( n91165 , n413699 );
not ( n413715 , n91165 );
buf ( n413716 , n413715 );
buf ( n413717 , n413716 );
not ( n413718 , n413717 );
buf ( n413719 , n91158 );
not ( n413720 , n413719 );
or ( n413721 , n413718 , n413720 );
buf ( n91173 , n378843 );
not ( n91174 , n91173 );
buf ( n413724 , n90940 );
not ( n91176 , n413724 );
or ( n413726 , n91174 , n91176 );
buf ( n413727 , n378843 );
not ( n91179 , n413727 );
buf ( n413729 , n409022 );
nand ( n413730 , n91179 , n413729 );
buf ( n413731 , n413730 );
buf ( n413732 , n413731 );
nand ( n413733 , n413726 , n413732 );
buf ( n413734 , n413733 );
buf ( n413735 , n413734 );
not ( n413736 , n413735 );
buf ( n413737 , n368599 );
not ( n91189 , n413737 );
or ( n413739 , n413736 , n91189 );
nand ( n413740 , n90950 , n369444 );
buf ( n413741 , n413740 );
nand ( n413742 , n413739 , n413741 );
buf ( n413743 , n413742 );
xor ( n91195 , n412927 , n412931 );
xor ( n413745 , n91195 , n412961 );
buf ( n413746 , n413745 );
buf ( n413747 , n413746 );
buf ( n413748 , n379260 );
not ( n413749 , n413748 );
buf ( n413750 , n413521 );
not ( n413751 , n413750 );
or ( n91203 , n413749 , n413751 );
buf ( n413753 , n377571 );
not ( n91205 , n413753 );
buf ( n413755 , n377776 );
not ( n413756 , n413755 );
or ( n413757 , n91205 , n413756 );
buf ( n413758 , n351027 );
buf ( n413759 , n379268 );
nand ( n413760 , n413758 , n413759 );
buf ( n413761 , n413760 );
buf ( n413762 , n413761 );
nand ( n413763 , n413757 , n413762 );
buf ( n413764 , n413763 );
buf ( n413765 , n413764 );
buf ( n413766 , n65117 );
nand ( n413767 , n413765 , n413766 );
buf ( n413768 , n413767 );
buf ( n413769 , n413768 );
nand ( n413770 , n91203 , n413769 );
buf ( n413771 , n413770 );
buf ( n413772 , n413771 );
xor ( n413773 , n413747 , n413772 );
buf ( n413774 , n58984 );
not ( n91226 , n413774 );
buf ( n413776 , n368584 );
not ( n413777 , n413776 );
or ( n91229 , n91226 , n413777 );
buf ( n413779 , n410287 );
buf ( n413780 , n408722 );
nand ( n91232 , n413779 , n413780 );
buf ( n413782 , n91232 );
buf ( n413783 , n413782 );
nand ( n91235 , n91229 , n413783 );
buf ( n413785 , n91235 );
buf ( n413786 , n413785 );
not ( n413787 , n413786 );
buf ( n91239 , n369801 );
not ( n91240 , n91239 );
or ( n91241 , n413787 , n91240 );
buf ( n413791 , n410307 );
not ( n413792 , n413791 );
buf ( n413793 , n413541 );
nand ( n413794 , n413792 , n413793 );
buf ( n413795 , n413794 );
buf ( n413796 , n413795 );
nand ( n413797 , n91241 , n413796 );
buf ( n413798 , n413797 );
buf ( n413799 , n413798 );
and ( n91251 , n413773 , n413799 );
and ( n91252 , n413747 , n413772 );
or ( n91253 , n91251 , n91252 );
buf ( n413803 , n91253 );
or ( n91255 , n413743 , n413803 );
xor ( n91256 , n91009 , n413562 );
xor ( n413806 , n91256 , n413556 );
nand ( n91258 , n91255 , n413806 );
nand ( n413808 , n413803 , n413743 );
nand ( n413809 , n91258 , n413808 );
buf ( n413810 , n413809 );
nand ( n91262 , n413721 , n413810 );
buf ( n91263 , n91262 );
buf ( n413813 , n91263 );
nand ( n91265 , n91164 , n413813 );
buf ( n413815 , n91265 );
buf ( n413816 , n413815 );
xor ( n413817 , n413683 , n413816 );
buf ( n413818 , n58923 );
not ( n91270 , n413818 );
buf ( n413820 , n413655 );
not ( n91272 , n413820 );
or ( n91273 , n91270 , n91272 );
buf ( n413823 , n379368 );
not ( n91275 , n413823 );
buf ( n413825 , n402185 );
not ( n91277 , n413825 );
or ( n413827 , n91275 , n91277 );
buf ( n413828 , n351345 );
buf ( n413829 , n379365 );
nand ( n413830 , n413828 , n413829 );
buf ( n413831 , n413830 );
buf ( n413832 , n413831 );
nand ( n413833 , n413827 , n413832 );
buf ( n413834 , n413833 );
buf ( n413835 , n413834 );
buf ( n413836 , n379353 );
nand ( n413837 , n413835 , n413836 );
buf ( n413838 , n413837 );
buf ( n413839 , n413838 );
nand ( n91291 , n91273 , n413839 );
buf ( n413841 , n91291 );
buf ( n413842 , n413841 );
and ( n413843 , n413817 , n413842 );
and ( n91295 , n413683 , n413816 );
or ( n91296 , n413843 , n91295 );
buf ( n413846 , n91296 );
buf ( n413847 , n413846 );
not ( n91299 , n413847 );
or ( n91300 , n413664 , n91299 );
buf ( n413850 , n413662 );
not ( n91302 , n413850 );
buf ( n413852 , n91302 );
not ( n91304 , n413852 );
buf ( n413854 , n413846 );
not ( n91306 , n413854 );
buf ( n413856 , n91306 );
not ( n91308 , n413856 );
or ( n91309 , n91304 , n91308 );
xor ( n91310 , n90640 , n413282 );
xor ( n413860 , n91310 , n413292 );
nand ( n91312 , n91309 , n413860 );
buf ( n413862 , n91312 );
nand ( n91314 , n91300 , n413862 );
buf ( n413864 , n91314 );
buf ( n413865 , n413864 );
nand ( n91317 , n413646 , n413865 );
buf ( n413867 , n91317 );
buf ( n413868 , n413867 );
nand ( n91320 , n413641 , n413868 );
buf ( n413870 , n91320 );
buf ( n91322 , n413870 );
buf ( n413872 , n91322 );
nand ( n413873 , n91079 , n413872 );
buf ( n413874 , n413873 );
buf ( n413875 , n413874 );
buf ( n413876 , n413618 );
not ( n91328 , n413876 );
buf ( n413878 , n91073 );
nand ( n91330 , n91328 , n413878 );
buf ( n413880 , n91330 );
buf ( n413881 , n413880 );
nand ( n413882 , n413875 , n413881 );
buf ( n413883 , n413882 );
buf ( n413884 , n413883 );
not ( n413885 , n413884 );
not ( n91337 , n413602 );
not ( n91338 , n90807 );
or ( n413888 , n91337 , n91338 );
not ( n91340 , n413335 );
or ( n413890 , n413602 , n91340 );
nand ( n91342 , n413888 , n413890 );
and ( n91343 , n91342 , n413339 );
not ( n413893 , n91342 );
and ( n91345 , n413893 , n413342 );
nor ( n413895 , n91343 , n91345 );
buf ( n413896 , n413895 );
nand ( n413897 , n413885 , n413896 );
buf ( n413898 , n413897 );
buf ( n413899 , n413898 );
not ( n413900 , n413899 );
buf ( n91352 , n413637 );
buf ( n91353 , n413864 );
xor ( n91354 , n91352 , n91353 );
buf ( n413904 , n91081 );
xnor ( n413905 , n91354 , n413904 );
buf ( n413906 , n413905 );
buf ( n413907 , n413906 );
buf ( n413908 , n413582 );
not ( n91360 , n413908 );
buf ( n413910 , n91360 );
and ( n91362 , n90902 , n413910 );
not ( n413912 , n90902 );
and ( n91364 , n413912 , n413582 );
nor ( n91365 , n91362 , n91364 );
xor ( n413915 , n91365 , n413448 );
buf ( n413916 , n413915 );
not ( n413917 , n413916 );
buf ( n413918 , n413917 );
buf ( n413919 , n413918 );
not ( n413920 , n413919 );
buf ( n413921 , n413410 );
buf ( n413922 , n380356 );
and ( n413923 , n413921 , n413922 );
buf ( n413924 , n380368 );
buf ( n413925 , n351160 );
xor ( n413926 , n413924 , n413925 );
buf ( n413927 , n413926 );
buf ( n413928 , n413927 );
not ( n91380 , n413928 );
buf ( n413930 , n385064 );
nor ( n413931 , n91380 , n413930 );
buf ( n413932 , n413931 );
buf ( n413933 , n413932 );
nor ( n413934 , n413923 , n413933 );
buf ( n413935 , n413934 );
buf ( n413936 , n413935 );
not ( n413937 , n413936 );
buf ( n413938 , n413937 );
buf ( n413939 , n413938 );
not ( n413940 , n413939 );
or ( n91392 , n413920 , n413940 );
buf ( n413942 , n413915 );
not ( n413943 , n413942 );
buf ( n413944 , n413935 );
not ( n413945 , n413944 );
or ( n91397 , n413943 , n413945 );
buf ( n413947 , n379890 );
not ( n413948 , n413947 );
buf ( n413949 , n413692 );
not ( n91401 , n413949 );
or ( n413951 , n413948 , n91401 );
buf ( n413952 , n379838 );
not ( n91404 , n413952 );
buf ( n413954 , n369372 );
not ( n413955 , n413954 );
or ( n413956 , n91404 , n413955 );
buf ( n413957 , n398741 );
buf ( n413958 , n352353 );
nand ( n413959 , n413957 , n413958 );
buf ( n413960 , n413959 );
buf ( n413961 , n413960 );
nand ( n413962 , n413956 , n413961 );
buf ( n413963 , n413962 );
buf ( n413964 , n413963 );
buf ( n413965 , n411170 );
nand ( n91417 , n413964 , n413965 );
buf ( n413967 , n91417 );
buf ( n413968 , n413967 );
nand ( n91420 , n413951 , n413968 );
buf ( n413970 , n91420 );
buf ( n413971 , n413970 );
not ( n91423 , n413971 );
buf ( n91424 , n44970 );
buf ( n91425 , n378098 );
nand ( n91426 , n91424 , n91425 );
buf ( n91427 , n91426 );
buf ( n413977 , n91427 );
not ( n91429 , n413977 );
buf ( n91430 , n91429 );
buf ( n413980 , n91430 );
not ( n413981 , n413980 );
or ( n91433 , n91423 , n413981 );
buf ( n413983 , n413970 );
not ( n413984 , n413983 );
buf ( n413985 , n413984 );
buf ( n413986 , n413985 );
not ( n413987 , n413986 );
buf ( n413988 , n91427 );
not ( n413989 , n413988 );
or ( n91441 , n413987 , n413989 );
not ( n413991 , n377094 );
not ( n91443 , n365136 );
or ( n91444 , n413991 , n91443 );
buf ( n413994 , n405357 );
buf ( n413995 , n377094 );
not ( n91447 , n413995 );
buf ( n413997 , n91447 );
buf ( n413998 , n413997 );
nand ( n91450 , n413994 , n413998 );
buf ( n414000 , n91450 );
nand ( n414001 , n91444 , n414000 );
buf ( n414002 , n414001 );
not ( n91454 , n414002 );
buf ( n414004 , n84022 );
not ( n91456 , n414004 );
or ( n414006 , n91454 , n91456 );
buf ( n414007 , n90665 );
buf ( n414008 , n44915 );
nand ( n414009 , n414007 , n414008 );
buf ( n414010 , n414009 );
buf ( n414011 , n414010 );
nand ( n91463 , n414006 , n414011 );
buf ( n414013 , n91463 );
buf ( n414014 , n414013 );
nand ( n414015 , n91441 , n414014 );
buf ( n414016 , n414015 );
buf ( n414017 , n414016 );
nand ( n91469 , n91433 , n414017 );
buf ( n414019 , n91469 );
buf ( n414020 , n414019 );
buf ( n414021 , n402201 );
not ( n91473 , n414021 );
buf ( n414023 , n378098 );
not ( n414024 , n414023 );
buf ( n414025 , n45050 );
not ( n414026 , n414025 );
or ( n414027 , n414024 , n414026 );
buf ( n414028 , n408998 );
buf ( n414029 , n379515 );
nand ( n414030 , n414028 , n414029 );
buf ( n414031 , n414030 );
buf ( n414032 , n414031 );
nand ( n414033 , n414027 , n414032 );
buf ( n414034 , n414033 );
buf ( n414035 , n414034 );
not ( n414036 , n414035 );
or ( n414037 , n91473 , n414036 );
buf ( n414038 , n407713 );
buf ( n414039 , n91122 );
nand ( n91491 , n414038 , n414039 );
buf ( n91492 , n91491 );
buf ( n414042 , n91492 );
nand ( n91494 , n414037 , n414042 );
buf ( n414044 , n91494 );
buf ( n414045 , n414044 );
xor ( n91497 , n414020 , n414045 );
buf ( n414047 , n58923 );
not ( n414048 , n414047 );
buf ( n414049 , n413834 );
not ( n91501 , n414049 );
or ( n91502 , n414048 , n91501 );
and ( n91503 , n379368 , n365384 );
not ( n91504 , n379368 );
and ( n414054 , n91504 , n351062 );
or ( n91506 , n91503 , n414054 );
buf ( n414056 , n91506 );
buf ( n414057 , n379350 );
not ( n414058 , n414057 );
buf ( n414059 , n414058 );
buf ( n414060 , n414059 );
nand ( n91512 , n414056 , n414060 );
buf ( n414062 , n91512 );
buf ( n414063 , n414062 );
nand ( n91515 , n91502 , n414063 );
buf ( n414065 , n91515 );
buf ( n414066 , n414065 );
and ( n91518 , n91497 , n414066 );
and ( n91519 , n414020 , n414045 );
or ( n91520 , n91518 , n91519 );
buf ( n414070 , n91520 );
buf ( n414071 , n414070 );
not ( n91523 , n414071 );
buf ( n414073 , n91523 );
buf ( n414074 , n414073 );
not ( n414075 , n414074 );
xor ( n91527 , n413569 , n413574 );
xor ( n91528 , n91527 , n413578 );
buf ( n414078 , n91528 );
buf ( n414079 , n414078 );
not ( n414080 , n414079 );
buf ( n414081 , n414080 );
buf ( n414082 , n414081 );
not ( n414083 , n414082 );
or ( n414084 , n414075 , n414083 );
buf ( n414085 , n413259 );
not ( n414086 , n414085 );
buf ( n414087 , n413276 );
not ( n91539 , n414087 );
or ( n414089 , n414086 , n91539 );
buf ( n91541 , n413256 );
buf ( n91542 , n413266 );
nand ( n91543 , n91541 , n91542 );
buf ( n91544 , n91543 );
buf ( n91545 , n91544 );
nand ( n91546 , n414089 , n91545 );
buf ( n91547 , n91546 );
buf ( n414097 , n91547 );
buf ( n414098 , n413230 );
not ( n91550 , n414098 );
buf ( n414100 , n91550 );
buf ( n414101 , n414100 );
and ( n91553 , n414097 , n414101 );
not ( n414103 , n414097 );
buf ( n414104 , n413230 );
and ( n414105 , n414103 , n414104 );
nor ( n91557 , n91553 , n414105 );
buf ( n414107 , n91557 );
buf ( n414108 , n414107 );
not ( n414109 , n414108 );
buf ( n414110 , n414109 );
buf ( n414111 , n414110 );
nand ( n414112 , n414084 , n414111 );
buf ( n414113 , n414112 );
buf ( n414114 , n414113 );
buf ( n414115 , n414070 );
buf ( n414116 , n414078 );
nand ( n91566 , n414115 , n414116 );
buf ( n414118 , n91566 );
buf ( n414119 , n414118 );
nand ( n414120 , n414114 , n414119 );
buf ( n414121 , n414120 );
buf ( n414122 , n414121 );
nand ( n414123 , n91397 , n414122 );
buf ( n414124 , n414123 );
buf ( n414125 , n414124 );
nand ( n91575 , n91392 , n414125 );
buf ( n414127 , n91575 );
buf ( n91577 , n414127 );
not ( n414129 , n91577 );
buf ( n414130 , n414129 );
buf ( n414131 , n414130 );
buf ( n414132 , n413394 );
buf ( n414133 , n413588 );
xor ( n414134 , n414132 , n414133 );
buf ( n414135 , n413417 );
xnor ( n414136 , n414134 , n414135 );
buf ( n414137 , n414136 );
buf ( n414138 , n414137 );
and ( n414139 , n414131 , n414138 );
buf ( n414140 , n414139 );
buf ( n414141 , n414140 );
or ( n91591 , n413907 , n414141 );
buf ( n414143 , n414137 );
buf ( n414144 , n414130 );
or ( n414145 , n414143 , n414144 );
buf ( n414146 , n414145 );
buf ( n414147 , n414146 );
nand ( n91597 , n91591 , n414147 );
buf ( n414149 , n91597 );
not ( n414150 , n414149 );
not ( n414151 , n413618 );
not ( n91601 , n414151 );
not ( n414153 , n413870 );
or ( n414154 , n91601 , n414153 );
not ( n91604 , n413870 );
nand ( n414156 , n91604 , n413618 );
nand ( n414157 , n414154 , n414156 );
and ( n91607 , n414157 , n91073 );
not ( n91608 , n414157 );
not ( n414160 , n91073 );
and ( n91610 , n91608 , n414160 );
nor ( n414162 , n91607 , n91610 );
nand ( n91612 , n414150 , n414162 );
not ( n414164 , n91612 );
buf ( n414165 , n414121 );
not ( n91615 , n414165 );
buf ( n414167 , n413935 );
not ( n91617 , n414167 );
and ( n91618 , n91615 , n91617 );
buf ( n414170 , n413935 );
buf ( n414171 , n414121 );
and ( n91621 , n414170 , n414171 );
nor ( n91622 , n91618 , n91621 );
buf ( n414174 , n91622 );
buf ( n414175 , n414174 );
buf ( n414176 , n413918 );
and ( n414177 , n414175 , n414176 );
not ( n91627 , n414175 );
buf ( n414179 , n413915 );
and ( n91629 , n91627 , n414179 );
nor ( n91630 , n414177 , n91629 );
buf ( n414182 , n91630 );
not ( n91632 , n413662 );
not ( n91633 , n413856 );
or ( n91634 , n91632 , n91633 );
buf ( n414186 , n413846 );
buf ( n414187 , n413852 );
nand ( n91637 , n414186 , n414187 );
buf ( n91638 , n91637 );
nand ( n91639 , n91634 , n91638 );
or ( n91640 , n91639 , n413860 );
nand ( n414192 , n91639 , n413860 );
nand ( n91642 , n91640 , n414192 );
xor ( n414194 , n413683 , n413816 );
xor ( n91644 , n414194 , n413842 );
buf ( n414196 , n91644 );
buf ( n414197 , n414196 );
buf ( n414198 , n380356 );
not ( n91648 , n414198 );
buf ( n414200 , n413927 );
not ( n414201 , n414200 );
or ( n91651 , n91648 , n414201 );
and ( n414203 , n380368 , n32234 );
not ( n91653 , n380368 );
and ( n91654 , n91653 , n352268 );
or ( n91655 , n414203 , n91654 );
buf ( n414207 , n91655 );
buf ( n414208 , n380401 );
nand ( n91658 , n414207 , n414208 );
buf ( n414210 , n91658 );
buf ( n414211 , n414210 );
nand ( n91661 , n91651 , n414211 );
buf ( n414213 , n91661 );
buf ( n414214 , n414213 );
or ( n91664 , n414197 , n414214 );
xor ( n91665 , n91427 , n413970 );
xor ( n91666 , n91665 , n414013 );
not ( n414218 , n91666 );
buf ( n414219 , n351043 );
buf ( n414220 , n379365 );
xor ( n414221 , n414219 , n414220 );
buf ( n414222 , n414221 );
not ( n414223 , n414222 );
not ( n91673 , n379350 );
and ( n414225 , n414223 , n91673 );
buf ( n414226 , n379368 );
not ( n91676 , n414226 );
buf ( n414228 , n408236 );
not ( n414229 , n414228 );
or ( n414230 , n91676 , n414229 );
buf ( n414231 , n352314 );
buf ( n91681 , n379365 );
nand ( n91682 , n414231 , n91681 );
buf ( n91683 , n91682 );
buf ( n414235 , n91683 );
nand ( n91685 , n414230 , n414235 );
buf ( n91686 , n91685 );
and ( n414238 , n91686 , n58923 );
nor ( n91688 , n414225 , n414238 );
buf ( n414240 , n91688 );
not ( n91690 , n414240 );
not ( n91691 , n378098 );
not ( n91692 , n406246 );
or ( n91693 , n91691 , n91692 );
buf ( n414245 , n405357 );
buf ( n414246 , n379515 );
nand ( n91696 , n414245 , n414246 );
buf ( n414248 , n91696 );
nand ( n91698 , n91693 , n414248 );
not ( n91699 , n91698 );
not ( n91700 , n84022 );
or ( n91701 , n91699 , n91700 );
not ( n414253 , n365076 );
nand ( n414254 , n414253 , n414001 );
nand ( n414255 , n91701 , n414254 );
not ( n414256 , n414255 );
buf ( n414257 , n414256 );
not ( n91707 , n414257 );
or ( n414259 , n91690 , n91707 );
buf ( n414260 , n413764 );
buf ( n414261 , n379260 );
and ( n414262 , n414260 , n414261 );
buf ( n414263 , n377571 );
not ( n91713 , n414263 );
buf ( n414265 , n90092 );
not ( n414266 , n414265 );
or ( n91716 , n91713 , n414266 );
buf ( n414268 , n351013 );
buf ( n414269 , n379268 );
nand ( n91719 , n414268 , n414269 );
buf ( n414271 , n91719 );
buf ( n414272 , n414271 );
nand ( n91722 , n91716 , n414272 );
buf ( n414274 , n91722 );
buf ( n414275 , n414274 );
not ( n91725 , n414275 );
buf ( n414277 , n379296 );
nor ( n91727 , n91725 , n414277 );
buf ( n414279 , n91727 );
buf ( n414280 , n414279 );
nor ( n414281 , n414262 , n414280 );
buf ( n414282 , n414281 );
buf ( n414283 , n414282 );
not ( n414284 , n377122 );
not ( n414285 , n411431 );
or ( n414286 , n414284 , n414285 );
buf ( n414287 , n57463 );
buf ( n414288 , n49582 );
nand ( n91738 , n414287 , n414288 );
buf ( n414290 , n91738 );
nand ( n91740 , n414286 , n414290 );
buf ( n414292 , n91740 );
not ( n414293 , n414292 );
buf ( n414294 , n407553 );
not ( n414295 , n414294 );
or ( n414296 , n414293 , n414295 );
buf ( n414297 , n412947 );
buf ( n414298 , n377579 );
nand ( n414299 , n414297 , n414298 );
buf ( n414300 , n414299 );
buf ( n414301 , n414300 );
nand ( n91751 , n414296 , n414301 );
buf ( n414303 , n91751 );
buf ( n414304 , n414303 );
xor ( n414305 , n412194 , n89702 );
xor ( n91755 , n414305 , n412238 );
xor ( n414307 , n90281 , n412921 );
xor ( n414308 , n91755 , n414307 );
buf ( n414309 , n414308 );
not ( n414310 , n414309 );
buf ( n414311 , n414310 );
buf ( n414312 , n414311 );
and ( n91762 , n414304 , n414312 );
not ( n414314 , n414304 );
buf ( n414315 , n414308 );
and ( n91765 , n414314 , n414315 );
nor ( n414317 , n91762 , n91765 );
buf ( n414318 , n414317 );
buf ( n414319 , n414318 );
xor ( n91769 , n414283 , n414319 );
buf ( n414321 , n91769 );
not ( n91771 , n414321 );
buf ( n414323 , n365075 );
buf ( n414324 , n378098 );
nand ( n91774 , n414323 , n414324 );
buf ( n414326 , n91774 );
buf ( n414327 , n414326 );
not ( n91777 , n414327 );
buf ( n414329 , n91777 );
not ( n91779 , n414329 );
or ( n414331 , n91771 , n91779 );
buf ( n414332 , n414321 );
not ( n91782 , n414332 );
buf ( n414334 , n91782 );
buf ( n414335 , n414334 );
not ( n91785 , n414335 );
buf ( n414337 , n414326 );
not ( n414338 , n414337 );
or ( n91788 , n91785 , n414338 );
buf ( n414340 , n379260 );
not ( n414341 , n414340 );
buf ( n414342 , n414274 );
not ( n91792 , n414342 );
or ( n414344 , n414341 , n91792 );
xor ( n91794 , n350988 , n377571 );
buf ( n414346 , n91794 );
buf ( n414347 , n379293 );
nand ( n91797 , n414346 , n414347 );
buf ( n414349 , n91797 );
buf ( n91799 , n414349 );
nand ( n91800 , n414344 , n91799 );
buf ( n91801 , n91800 );
buf ( n91802 , n91801 );
xor ( n91803 , n412828 , n90357 );
xor ( n414355 , n91803 , n412902 );
buf ( n414356 , n79312 );
buf ( n414357 , n394840 );
and ( n91807 , n414356 , n414357 );
buf ( n414359 , n79318 );
buf ( n414360 , n384408 );
and ( n91810 , n414359 , n414360 );
nor ( n414362 , n91807 , n91810 );
buf ( n414363 , n414362 );
buf ( n414364 , n414363 );
buf ( n414365 , n394838 );
or ( n91815 , n414364 , n414365 );
buf ( n414367 , n412799 );
buf ( n414368 , n394835 );
or ( n91818 , n414367 , n414368 );
nand ( n91819 , n91815 , n91818 );
buf ( n414371 , n91819 );
xor ( n91821 , n412746 , n412762 );
xor ( n414373 , n91821 , n412787 );
and ( n91823 , n414371 , n414373 );
xor ( n91824 , n412768 , n412785 );
buf ( n414376 , n91824 );
buf ( n414377 , n414376 );
buf ( n414378 , n384354 );
buf ( n414379 , n382627 );
buf ( n414380 , n405813 );
and ( n414381 , n414379 , n414380 );
buf ( n414382 , n62026 );
buf ( n414383 , n405816 );
and ( n414384 , n414382 , n414383 );
nor ( n414385 , n414381 , n414384 );
buf ( n414386 , n414385 );
buf ( n414387 , n414386 );
or ( n414388 , n414378 , n414387 );
buf ( n414389 , n412873 );
buf ( n414390 , n384082 );
or ( n414391 , n414389 , n414390 );
nand ( n91841 , n414388 , n414391 );
buf ( n414393 , n91841 );
buf ( n414394 , n380696 );
buf ( n414395 , n623 );
and ( n91845 , n414394 , n414395 );
buf ( n414397 , n380697 );
buf ( n414398 , n85590 );
and ( n91848 , n414397 , n414398 );
buf ( n414400 , n382638 );
nor ( n414401 , n91848 , n414400 );
buf ( n414402 , n414401 );
buf ( n414403 , n414402 );
buf ( n414404 , n406588 );
nor ( n91854 , n91845 , n414403 , n414404 );
buf ( n414406 , n91854 );
xor ( n91856 , n414393 , n414406 );
buf ( n414408 , n382849 );
buf ( n414409 , n382638 );
buf ( n414410 , n406746 );
and ( n91860 , n414409 , n414410 );
buf ( n414412 , n382647 );
buf ( n414413 , n406749 );
and ( n91863 , n414412 , n414413 );
nor ( n414415 , n91860 , n91863 );
buf ( n414416 , n414415 );
buf ( n414417 , n414416 );
or ( n91867 , n414408 , n414417 );
buf ( n414419 , n412777 );
buf ( n414420 , n382634 );
or ( n91870 , n414419 , n414420 );
nand ( n414422 , n91867 , n91870 );
buf ( n414423 , n414422 );
and ( n91873 , n91856 , n414423 );
and ( n414425 , n414393 , n414406 );
or ( n414426 , n91873 , n414425 );
buf ( n414427 , n414426 );
xor ( n414428 , n414377 , n414427 );
buf ( n414429 , n380730 );
buf ( n414430 , n623 );
and ( n91880 , n414429 , n414430 );
buf ( n414432 , n91880 );
buf ( n414433 , n414432 );
buf ( n414434 , n90113 );
buf ( n414435 , n403795 );
and ( n91885 , n414434 , n414435 );
buf ( n414437 , n403798 );
buf ( n414438 , n384421 );
and ( n91888 , n414437 , n414438 );
nor ( n414440 , n91885 , n91888 );
buf ( n414441 , n414440 );
buf ( n414442 , n414441 );
buf ( n414443 , n384414 );
or ( n414444 , n414442 , n414443 );
buf ( n414445 , n403772 );
buf ( n414446 , n90113 );
and ( n91891 , n414445 , n414446 );
buf ( n414448 , n403775 );
buf ( n414449 , n384421 );
and ( n91894 , n414448 , n414449 );
nor ( n414451 , n91891 , n91894 );
buf ( n414452 , n414451 );
buf ( n414453 , n414452 );
buf ( n414454 , n395635 );
or ( n91899 , n414453 , n414454 );
nand ( n414456 , n414444 , n91899 );
buf ( n414457 , n414456 );
buf ( n414458 , n414457 );
and ( n414459 , n414433 , n414458 );
buf ( n414460 , n414459 );
buf ( n414461 , n414460 );
buf ( n414462 , n414452 );
buf ( n414463 , n384414 );
or ( n414464 , n414462 , n414463 );
buf ( n414465 , n412855 );
buf ( n414466 , n395635 );
or ( n91911 , n414465 , n414466 );
nand ( n414468 , n414464 , n91911 );
buf ( n414469 , n414468 );
buf ( n414470 , n414469 );
xor ( n414471 , n414461 , n414470 );
buf ( n414472 , n60226 );
buf ( n414473 , n623 );
or ( n91918 , n414472 , n414473 );
buf ( n414475 , n380735 );
buf ( n414476 , n406588 );
buf ( n414477 , n623 );
and ( n414478 , n414475 , n414476 , n414477 );
buf ( n91923 , n380744 );
not ( n91924 , n91923 );
buf ( n91925 , n91924 );
buf ( n414482 , n91925 );
nor ( n91927 , n414478 , n414482 );
buf ( n91928 , n91927 );
buf ( n414485 , n91928 );
nand ( n91930 , n91918 , n414485 );
buf ( n91931 , n91930 );
buf ( n414488 , n91931 );
and ( n91933 , n414471 , n414488 );
and ( n91934 , n414461 , n414470 );
or ( n91935 , n91933 , n91934 );
buf ( n414492 , n91935 );
buf ( n414493 , n414492 );
and ( n91938 , n414428 , n414493 );
and ( n91939 , n414377 , n414427 );
or ( n91940 , n91938 , n91939 );
buf ( n414497 , n91940 );
xor ( n91942 , n412746 , n412762 );
xor ( n91943 , n91942 , n412787 );
and ( n414500 , n414497 , n91943 );
and ( n414501 , n414371 , n414497 );
or ( n91946 , n91823 , n414500 , n414501 );
xor ( n414503 , n412864 , n412881 );
xor ( n91948 , n414503 , n412889 );
buf ( n414505 , n91948 );
buf ( n414506 , n80468 );
buf ( n414507 , n394840 );
and ( n414508 , n414506 , n414507 );
buf ( n414509 , n401921 );
buf ( n414510 , n384408 );
and ( n414511 , n414509 , n414510 );
nor ( n414512 , n414508 , n414511 );
buf ( n414513 , n414512 );
buf ( n414514 , n414513 );
buf ( n414515 , n394838 );
or ( n91960 , n414514 , n414515 );
buf ( n414517 , n414363 );
buf ( n414518 , n394835 );
or ( n414519 , n414517 , n414518 );
nand ( n91964 , n91960 , n414519 );
buf ( n91965 , n91964 );
xor ( n414522 , n414505 , n91965 );
buf ( n414523 , n81950 );
buf ( n414524 , n394840 );
and ( n414525 , n414523 , n414524 );
buf ( n414526 , n403589 );
buf ( n414527 , n384408 );
and ( n414528 , n414526 , n414527 );
nor ( n91973 , n414525 , n414528 );
buf ( n414530 , n91973 );
buf ( n91975 , n414530 );
buf ( n91976 , n394838 );
or ( n91977 , n91975 , n91976 );
buf ( n91978 , n414513 );
buf ( n414535 , n394835 );
or ( n414536 , n91978 , n414535 );
nand ( n414537 , n91977 , n414536 );
buf ( n414538 , n414537 );
xor ( n414539 , n414393 , n414406 );
xor ( n414540 , n414539 , n414423 );
and ( n91985 , n414538 , n414540 );
xor ( n414542 , n414433 , n414458 );
buf ( n414543 , n414542 );
buf ( n414544 , n414543 );
buf ( n414545 , n384354 );
buf ( n414546 , n382627 );
buf ( n414547 , n406569 );
and ( n91992 , n414546 , n414547 );
buf ( n414549 , n384089 );
buf ( n414550 , n406572 );
and ( n414551 , n414549 , n414550 );
nor ( n414552 , n91992 , n414551 );
buf ( n414553 , n414552 );
buf ( n414554 , n414553 );
or ( n414555 , n414545 , n414554 );
buf ( n414556 , n414386 );
buf ( n414557 , n384082 );
or ( n414558 , n414556 , n414557 );
nand ( n92003 , n414555 , n414558 );
buf ( n414560 , n92003 );
buf ( n414561 , n414560 );
xor ( n92006 , n414544 , n414561 );
buf ( n414563 , n382634 );
buf ( n414564 , n414416 );
or ( n92009 , n414563 , n414564 );
buf ( n414566 , n382659 );
nand ( n414567 , n92009 , n414566 );
buf ( n414568 , n414567 );
buf ( n414569 , n414568 );
and ( n414570 , n92006 , n414569 );
and ( n92015 , n414544 , n414561 );
or ( n92016 , n414570 , n92015 );
buf ( n414573 , n92016 );
xor ( n92018 , n414393 , n414406 );
xor ( n414575 , n92018 , n414423 );
and ( n92020 , n414573 , n414575 );
and ( n414577 , n414538 , n414573 );
or ( n414578 , n91985 , n92020 , n414577 );
and ( n92023 , n414522 , n414578 );
and ( n414580 , n414505 , n91965 );
or ( n414581 , n92023 , n414580 );
buf ( n414582 , n414581 );
xor ( n414583 , n412687 , n412700 );
xor ( n92028 , n414583 , n412722 );
xor ( n414585 , n412844 , n412893 );
xor ( n92030 , n92028 , n414585 );
buf ( n414587 , n92030 );
xor ( n92032 , n414582 , n414587 );
xor ( n92033 , n412746 , n412762 );
xor ( n414590 , n92033 , n412787 );
xor ( n414591 , n414371 , n414497 );
xor ( n92036 , n414590 , n414591 );
buf ( n414593 , n92036 );
and ( n414594 , n92032 , n414593 );
and ( n92039 , n414582 , n414587 );
or ( n414596 , n414594 , n92039 );
buf ( n414597 , n414596 );
xor ( n92042 , n91946 , n414597 );
xor ( n92043 , n414355 , n92042 );
buf ( n92044 , n92043 );
buf ( n414601 , n379260 );
not ( n92046 , n414601 );
buf ( n414603 , n91794 );
not ( n414604 , n414603 );
or ( n92049 , n92046 , n414604 );
buf ( n414606 , n379293 );
buf ( n414607 , n377119 );
not ( n92052 , n414607 );
buf ( n414609 , n23104 );
not ( n414610 , n414609 );
buf ( n414611 , n414610 );
buf ( n414612 , n414611 );
not ( n414613 , n414612 );
or ( n92058 , n92052 , n414613 );
buf ( n414615 , n377571 );
buf ( n414616 , n30931 );
not ( n92061 , n414616 );
buf ( n414618 , n92061 );
buf ( n414619 , n414618 );
nand ( n414620 , n414615 , n414619 );
buf ( n414621 , n414620 );
buf ( n414622 , n414621 );
nand ( n92067 , n92058 , n414622 );
buf ( n414624 , n92067 );
buf ( n414625 , n414624 );
nand ( n414626 , n414606 , n414625 );
buf ( n414627 , n414626 );
buf ( n414628 , n414627 );
nand ( n414629 , n92049 , n414628 );
buf ( n414630 , n414629 );
buf ( n414631 , n414630 );
xor ( n92076 , n92044 , n414631 );
xor ( n414633 , n414377 , n414427 );
xor ( n92078 , n414633 , n414493 );
buf ( n414635 , n92078 );
xor ( n414636 , n414505 , n91965 );
xor ( n92081 , n414636 , n414578 );
and ( n414638 , n414635 , n92081 );
buf ( n414639 , n382610 );
buf ( n414640 , n623 );
and ( n92085 , n414639 , n414640 );
buf ( n414642 , n382642 );
buf ( n414643 , n85590 );
and ( n414644 , n414642 , n414643 );
buf ( n414645 , n382627 );
nor ( n414646 , n414644 , n414645 );
buf ( n414647 , n414646 );
buf ( n414648 , n414647 );
buf ( n414649 , n382835 );
nor ( n92094 , n92085 , n414648 , n414649 );
buf ( n92095 , n92094 );
buf ( n414652 , n384414 );
buf ( n414653 , n90113 );
buf ( n414654 , n405813 );
and ( n414655 , n414653 , n414654 );
buf ( n414656 , n384421 );
buf ( n414657 , n405816 );
and ( n414658 , n414656 , n414657 );
nor ( n92103 , n414655 , n414658 );
buf ( n414660 , n92103 );
buf ( n414661 , n414660 );
or ( n92106 , n414652 , n414661 );
buf ( n414663 , n414441 );
buf ( n414664 , n395635 );
or ( n92109 , n414663 , n414664 );
nand ( n414666 , n92106 , n92109 );
buf ( n414667 , n414666 );
xor ( n92112 , n92095 , n414667 );
buf ( n414669 , n384414 );
buf ( n414670 , n90113 );
buf ( n414671 , n406569 );
and ( n414672 , n414670 , n414671 );
buf ( n414673 , n384421 );
buf ( n414674 , n406572 );
and ( n92119 , n414673 , n414674 );
nor ( n92120 , n414672 , n92119 );
buf ( n414677 , n92120 );
buf ( n414678 , n414677 );
or ( n414679 , n414669 , n414678 );
buf ( n414680 , n414660 );
buf ( n414681 , n395635 );
or ( n92126 , n414680 , n414681 );
nand ( n414683 , n414679 , n92126 );
buf ( n414684 , n414683 );
buf ( n414685 , n414684 );
buf ( n414686 , n382634 );
buf ( n414687 , n85590 );
nor ( n92132 , n414686 , n414687 );
buf ( n92133 , n92132 );
buf ( n414690 , n92133 );
and ( n414691 , n414685 , n414690 );
buf ( n414692 , n414691 );
and ( n414693 , n92112 , n414692 );
and ( n92138 , n92095 , n414667 );
or ( n414695 , n414693 , n92138 );
buf ( n414696 , n414695 );
buf ( n414697 , n81995 );
buf ( n414698 , n394840 );
and ( n92143 , n414697 , n414698 );
buf ( n414700 , n403645 );
buf ( n414701 , n384408 );
and ( n92146 , n414700 , n414701 );
nor ( n92147 , n92143 , n92146 );
buf ( n414704 , n92147 );
buf ( n414705 , n414704 );
buf ( n414706 , n394838 );
or ( n92151 , n414705 , n414706 );
buf ( n414708 , n414530 );
buf ( n414709 , n394835 );
or ( n92154 , n414708 , n414709 );
nand ( n414711 , n92151 , n92154 );
buf ( n414712 , n414711 );
buf ( n414713 , n414712 );
xor ( n414714 , n414696 , n414713 );
xor ( n92159 , n414544 , n414561 );
xor ( n92160 , n92159 , n414569 );
buf ( n414717 , n92160 );
buf ( n414718 , n414717 );
and ( n414719 , n414714 , n414718 );
and ( n92164 , n414696 , n414713 );
or ( n92165 , n414719 , n92164 );
buf ( n414722 , n92165 );
buf ( n414723 , n414722 );
xor ( n414724 , n414461 , n414470 );
xor ( n92169 , n414724 , n414488 );
buf ( n414726 , n92169 );
buf ( n414727 , n414726 );
xor ( n92172 , n414723 , n414727 );
xor ( n414729 , n414393 , n414406 );
xor ( n92174 , n414729 , n414423 );
xor ( n414731 , n414538 , n414573 );
xor ( n92176 , n92174 , n414731 );
buf ( n414733 , n92176 );
and ( n92178 , n92172 , n414733 );
and ( n92179 , n414723 , n414727 );
or ( n92180 , n92178 , n92179 );
buf ( n414737 , n92180 );
xor ( n414738 , n414505 , n91965 );
xor ( n414739 , n414738 , n414578 );
and ( n414740 , n414737 , n414739 );
and ( n92185 , n414635 , n414737 );
or ( n414742 , n414638 , n414740 , n92185 );
buf ( n414743 , n414742 );
xor ( n414744 , n414582 , n414587 );
xor ( n414745 , n414744 , n414593 );
buf ( n414746 , n414745 );
buf ( n414747 , n414746 );
xor ( n414748 , n414743 , n414747 );
buf ( n414749 , n379472 );
not ( n414750 , n414749 );
buf ( n414751 , n414611 );
not ( n414752 , n414751 );
or ( n92197 , n414750 , n414752 );
buf ( n414754 , n379472 );
not ( n92199 , n414754 );
buf ( n92200 , n92199 );
buf ( n414757 , n92200 );
buf ( n414758 , n377571 );
nand ( n414759 , n414757 , n414758 );
buf ( n414760 , n414759 );
buf ( n414761 , n414760 );
nand ( n414762 , n92197 , n414761 );
buf ( n414763 , n414762 );
buf ( n414764 , n414763 );
not ( n92209 , n414764 );
buf ( n414766 , n379293 );
not ( n414767 , n414766 );
or ( n92212 , n92209 , n414767 );
buf ( n414769 , n414624 );
buf ( n414770 , n379260 );
nand ( n92215 , n414769 , n414770 );
buf ( n414772 , n92215 );
buf ( n414773 , n414772 );
nand ( n414774 , n92212 , n414773 );
buf ( n414775 , n414774 );
buf ( n414776 , n414775 );
and ( n414777 , n414748 , n414776 );
and ( n414778 , n414743 , n414747 );
or ( n414779 , n414777 , n414778 );
buf ( n414780 , n414779 );
buf ( n414781 , n414780 );
and ( n92226 , n92076 , n414781 );
and ( n92227 , n92044 , n414631 );
or ( n414784 , n92226 , n92227 );
buf ( n414785 , n414784 );
buf ( n414786 , n414785 );
xor ( n414787 , n91802 , n414786 );
xor ( n414788 , n412906 , n90370 );
xor ( n92233 , n414788 , n412917 );
buf ( n414790 , n92233 );
buf ( n414791 , n414790 );
xor ( n92236 , n412828 , n90357 );
xor ( n414793 , n92236 , n412902 );
and ( n92238 , n91946 , n414793 );
xor ( n414795 , n412828 , n90357 );
xor ( n92240 , n414795 , n412902 );
and ( n92241 , n414597 , n92240 );
and ( n414798 , n91946 , n414597 );
or ( n414799 , n92238 , n92241 , n414798 );
buf ( n414800 , n414799 );
xnor ( n414801 , n414791 , n414800 );
buf ( n414802 , n414801 );
buf ( n414803 , n407553 );
not ( n414804 , n414803 );
buf ( n414805 , n379472 );
not ( n92250 , n414805 );
buf ( n414807 , n411431 );
not ( n414808 , n414807 );
or ( n92253 , n92250 , n414808 );
buf ( n414810 , n412940 );
buf ( n414811 , n92200 );
nand ( n414812 , n414810 , n414811 );
buf ( n414813 , n414812 );
buf ( n414814 , n414813 );
nand ( n92259 , n92253 , n414814 );
buf ( n414816 , n92259 );
buf ( n414817 , n414816 );
not ( n414818 , n414817 );
or ( n92263 , n414804 , n414818 );
nand ( n414820 , n377579 , n91740 );
buf ( n414821 , n414820 );
nand ( n414822 , n92263 , n414821 );
buf ( n414823 , n414822 );
not ( n92268 , n414823 );
xor ( n414825 , n414802 , n92268 );
buf ( n414826 , n414825 );
and ( n92271 , n414787 , n414826 );
and ( n92272 , n91802 , n414786 );
or ( n92273 , n92271 , n92272 );
buf ( n414830 , n92273 );
buf ( n414831 , n414830 );
nand ( n414832 , n91788 , n414831 );
buf ( n414833 , n414832 );
nand ( n92278 , n414331 , n414833 );
buf ( n414835 , n92278 );
nand ( n92280 , n414259 , n414835 );
buf ( n414837 , n92280 );
buf ( n92282 , n414837 );
buf ( n414839 , n91688 );
not ( n92284 , n414839 );
buf ( n414841 , n414256 );
not ( n414842 , n414841 );
buf ( n414843 , n414842 );
buf ( n414844 , n414843 );
nand ( n414845 , n92284 , n414844 );
buf ( n414846 , n414845 );
buf ( n414847 , n414846 );
and ( n92292 , n92282 , n414847 );
buf ( n414849 , n92292 );
not ( n92294 , n414849 );
and ( n92295 , n414218 , n92294 );
buf ( n92296 , n414849 );
buf ( n92297 , n91666 );
nand ( n92298 , n92296 , n92297 );
buf ( n92299 , n92298 );
xor ( n414856 , n413743 , n413803 );
xor ( n92301 , n414856 , n413806 );
and ( n414858 , n92299 , n92301 );
nor ( n414859 , n92295 , n414858 );
buf ( n414860 , n414859 );
not ( n92305 , n414860 );
buf ( n414862 , n92305 );
not ( n92307 , n414862 );
buf ( n414864 , n414303 );
not ( n414865 , n414864 );
buf ( n414866 , n414282 );
not ( n92311 , n414866 );
buf ( n92312 , n92311 );
buf ( n414869 , n92312 );
not ( n92314 , n414869 );
or ( n414871 , n414865 , n92314 );
buf ( n414872 , n414303 );
not ( n92317 , n414872 );
buf ( n414874 , n92317 );
buf ( n414875 , n414874 );
not ( n414876 , n414875 );
buf ( n414877 , n414282 );
not ( n92322 , n414877 );
or ( n414879 , n414876 , n92322 );
buf ( n414880 , n414308 );
nand ( n414881 , n414879 , n414880 );
buf ( n414882 , n414881 );
buf ( n414883 , n414882 );
nand ( n414884 , n414871 , n414883 );
buf ( n414885 , n414884 );
buf ( n414886 , n414885 );
buf ( n414887 , n342965 );
buf ( n414888 , n90940 );
not ( n414889 , n414888 );
buf ( n414890 , n365062 );
not ( n92335 , n414890 );
or ( n414892 , n414889 , n92335 );
buf ( n414893 , n378098 );
nand ( n92338 , n414892 , n414893 );
buf ( n414895 , n92338 );
buf ( n414896 , n414895 );
buf ( n414897 , n23037 );
buf ( n414898 , n342445 );
nand ( n414899 , n414897 , n414898 );
buf ( n414900 , n414899 );
buf ( n414901 , n414900 );
and ( n414902 , n414887 , n414896 , n414901 );
buf ( n414903 , n414902 );
buf ( n414904 , n414903 );
xor ( n414905 , n414886 , n414904 );
xor ( n414906 , n413747 , n413772 );
xor ( n92351 , n414906 , n413799 );
buf ( n414908 , n92351 );
buf ( n414909 , n414908 );
and ( n414910 , n414905 , n414909 );
and ( n92355 , n414886 , n414904 );
or ( n414912 , n414910 , n92355 );
buf ( n414913 , n414912 );
buf ( n414914 , n414913 );
and ( n92359 , n413963 , n379890 );
and ( n414916 , n377379 , n398741 );
not ( n414917 , n377379 );
and ( n92362 , n414917 , n379838 );
or ( n92363 , n414916 , n92362 );
and ( n414920 , n92363 , n411170 );
nor ( n414921 , n92359 , n414920 );
buf ( n414922 , n414921 );
not ( n414923 , n414922 );
buf ( n414924 , n414923 );
buf ( n414925 , n414924 );
not ( n92370 , n414925 );
buf ( n414927 , n377068 );
not ( n92372 , n414927 );
buf ( n414929 , n85756 );
not ( n92374 , n414929 );
or ( n92375 , n92372 , n92374 );
buf ( n414932 , n377068 );
not ( n414933 , n414932 );
buf ( n414934 , n23037 );
nand ( n92379 , n414933 , n414934 );
buf ( n414936 , n92379 );
buf ( n414937 , n414936 );
nand ( n92382 , n92375 , n414937 );
buf ( n414939 , n92382 );
buf ( n414940 , n414939 );
not ( n92385 , n414940 );
buf ( n414942 , n413496 );
not ( n414943 , n414942 );
or ( n92388 , n92385 , n414943 );
buf ( n414945 , n368593 );
not ( n92390 , n414945 );
buf ( n414947 , n413734 );
nand ( n92392 , n92390 , n414947 );
buf ( n92393 , n92392 );
buf ( n414950 , n92393 );
nand ( n92395 , n92388 , n414950 );
buf ( n414952 , n92395 );
buf ( n414953 , n414952 );
not ( n414954 , n414953 );
or ( n92399 , n92370 , n414954 );
or ( n414956 , n414924 , n414952 );
buf ( n414957 , n92363 );
buf ( n414958 , n379890 );
and ( n414959 , n414957 , n414958 );
not ( n414960 , n352404 );
buf ( n414961 , n379253 );
not ( n414962 , n414961 );
buf ( n414963 , n414962 );
not ( n92408 , n414963 );
or ( n414965 , n414960 , n92408 );
nand ( n92410 , n377349 , n379253 );
nand ( n92411 , n414965 , n92410 );
buf ( n414968 , n92411 );
buf ( n414969 , n411170 );
and ( n414970 , n414968 , n414969 );
buf ( n414971 , n414970 );
buf ( n414972 , n414971 );
nor ( n92417 , n414959 , n414972 );
buf ( n92418 , n92417 );
buf ( n414975 , n92418 );
not ( n92420 , n414975 );
buf ( n414977 , n378843 );
not ( n414978 , n414977 );
buf ( n414979 , n368561 );
not ( n414980 , n414979 );
or ( n414981 , n414978 , n414980 );
buf ( n414982 , n410296 );
buf ( n414983 , n410976 );
nand ( n414984 , n414982 , n414983 );
buf ( n414985 , n414984 );
buf ( n414986 , n414985 );
nand ( n92431 , n414981 , n414986 );
buf ( n414988 , n92431 );
buf ( n414989 , n414988 );
not ( n92434 , n414989 );
buf ( n414991 , n369801 );
not ( n92436 , n414991 );
or ( n414993 , n92434 , n92436 );
buf ( n414994 , n413785 );
buf ( n414995 , n369809 );
nand ( n414996 , n414994 , n414995 );
buf ( n414997 , n414996 );
buf ( n414998 , n414997 );
nand ( n92443 , n414993 , n414998 );
buf ( n415000 , n92443 );
buf ( n92445 , n415000 );
nand ( n92446 , n92420 , n92445 );
buf ( n92447 , n92446 );
buf ( n415004 , n415000 );
not ( n92449 , n415004 );
buf ( n92450 , n92449 );
not ( n415007 , n92450 );
not ( n92452 , n92418 );
or ( n415009 , n415007 , n92452 );
not ( n415010 , n414799 );
not ( n92455 , n414823 );
or ( n415012 , n415010 , n92455 );
or ( n92457 , n414823 , n414799 );
nand ( n92458 , n92457 , n414790 );
nand ( n415015 , n415012 , n92458 );
nand ( n92460 , n415009 , n415015 );
nand ( n415017 , n92447 , n92460 );
nand ( n415018 , n414956 , n415017 );
buf ( n415019 , n415018 );
nand ( n415020 , n92399 , n415019 );
buf ( n415021 , n415020 );
buf ( n415022 , n415021 );
xor ( n415023 , n414914 , n415022 );
buf ( n415024 , n58923 );
not ( n92469 , n415024 );
buf ( n415026 , n91506 );
not ( n415027 , n415026 );
or ( n415028 , n92469 , n415027 );
buf ( n415029 , n91686 );
buf ( n415030 , n414059 );
nand ( n92475 , n415029 , n415030 );
buf ( n415032 , n92475 );
buf ( n415033 , n415032 );
nand ( n92478 , n415028 , n415033 );
buf ( n92479 , n92478 );
buf ( n415036 , n92479 );
and ( n415037 , n415023 , n415036 );
and ( n415038 , n414914 , n415022 );
or ( n92483 , n415037 , n415038 );
buf ( n415040 , n92483 );
not ( n92485 , n415040 );
or ( n415042 , n92307 , n92485 );
buf ( n415043 , n415040 );
not ( n92488 , n415043 );
buf ( n415045 , n92488 );
not ( n92490 , n415045 );
not ( n92491 , n414859 );
or ( n92492 , n92490 , n92491 );
buf ( n415049 , n90675 );
buf ( n415050 , n413224 );
xor ( n92495 , n415049 , n415050 );
buf ( n415052 , n90667 );
xnor ( n92497 , n92495 , n415052 );
buf ( n415054 , n92497 );
buf ( n415055 , n415054 );
not ( n415056 , n415055 );
buf ( n415057 , n415056 );
nand ( n92502 , n92492 , n415057 );
nand ( n92503 , n415042 , n92502 );
buf ( n415060 , n92503 );
nand ( n92505 , n91664 , n415060 );
buf ( n415062 , n92505 );
buf ( n415063 , n414213 );
buf ( n415064 , n414196 );
nand ( n415065 , n415063 , n415064 );
buf ( n415066 , n415065 );
and ( n415067 , n415062 , n415066 );
and ( n92512 , n91642 , n415067 );
or ( n415069 , n414182 , n92512 );
or ( n415070 , n91642 , n415067 );
nand ( n92515 , n415069 , n415070 );
buf ( n415072 , n92515 );
not ( n415073 , n415072 );
xor ( n92518 , n414131 , n414138 );
buf ( n415075 , n92518 );
xor ( n92520 , n415075 , n413906 );
buf ( n415077 , n92520 );
nand ( n92522 , n415073 , n415077 );
buf ( n415079 , n92522 );
not ( n415080 , n415079 );
xor ( n92525 , n415015 , n92450 );
xnor ( n92526 , n92525 , n92418 );
not ( n415083 , n92526 );
buf ( n415084 , n23034 );
buf ( n415085 , n22484 );
buf ( n415086 , n410296 );
or ( n415087 , n415085 , n415086 );
buf ( n415088 , n378098 );
nand ( n92533 , n415087 , n415088 );
buf ( n415090 , n92533 );
buf ( n415091 , n415090 );
buf ( n415092 , n22484 );
buf ( n415093 , n410287 );
nand ( n415094 , n415092 , n415093 );
buf ( n415095 , n415094 );
buf ( n415096 , n415095 );
nand ( n415097 , n415084 , n415091 , n415096 );
buf ( n415098 , n415097 );
not ( n92543 , n415098 );
and ( n92544 , n92411 , n379890 );
and ( n415101 , n351027 , n414963 );
not ( n415102 , n351027 );
and ( n92547 , n415102 , n379253 );
or ( n415104 , n415101 , n92547 );
buf ( n415105 , n415104 );
buf ( n415106 , n379912 );
and ( n92551 , n415105 , n415106 );
buf ( n415108 , n92551 );
nor ( n415109 , n92544 , n415108 );
not ( n92554 , n415109 );
and ( n415111 , n92543 , n92554 );
buf ( n415112 , n415098 );
buf ( n415113 , n415109 );
nand ( n92558 , n415112 , n415113 );
buf ( n415115 , n92558 );
buf ( n415116 , n377068 );
not ( n92561 , n415116 );
buf ( n415118 , n368584 );
not ( n415119 , n415118 );
or ( n92564 , n92561 , n415119 );
not ( n415121 , n377065 );
nand ( n415122 , n343193 , n415121 );
buf ( n415123 , n415122 );
nand ( n92568 , n92564 , n415123 );
buf ( n415125 , n92568 );
buf ( n415126 , n415125 );
not ( n92571 , n415126 );
buf ( n415128 , n369801 );
not ( n415129 , n415128 );
or ( n92574 , n92571 , n415129 );
buf ( n415131 , n414988 );
buf ( n415132 , n369809 );
nand ( n92577 , n415131 , n415132 );
buf ( n415134 , n92577 );
buf ( n415135 , n415134 );
nand ( n92580 , n92574 , n415135 );
buf ( n92581 , n92580 );
and ( n415138 , n415115 , n92581 );
nor ( n92583 , n415111 , n415138 );
not ( n415140 , n92583 );
nand ( n92585 , n415083 , n415140 );
not ( n415142 , n92585 );
buf ( n415143 , n377094 );
not ( n92588 , n415143 );
buf ( n415145 , n85756 );
not ( n415146 , n415145 );
or ( n92591 , n92588 , n415146 );
buf ( n415148 , n409022 );
buf ( n415149 , n413997 );
nand ( n415150 , n415148 , n415149 );
buf ( n415151 , n415150 );
buf ( n415152 , n415151 );
nand ( n92597 , n92591 , n415152 );
buf ( n415154 , n92597 );
buf ( n415155 , n415154 );
not ( n415156 , n415155 );
buf ( n415157 , n415156 );
buf ( n415158 , n415157 );
not ( n415159 , n415158 );
buf ( n415160 , n368596 );
not ( n92605 , n415160 );
and ( n415162 , n415159 , n92605 );
buf ( n415163 , n414939 );
not ( n92608 , n415163 );
buf ( n415165 , n368593 );
nor ( n415166 , n92608 , n415165 );
buf ( n415167 , n415166 );
buf ( n415168 , n415167 );
nor ( n92613 , n415162 , n415168 );
buf ( n415170 , n92613 );
buf ( n415171 , n415170 );
not ( n415172 , n415171 );
or ( n92617 , n415142 , n415172 );
nand ( n92618 , n92526 , n92583 );
nand ( n92619 , n92617 , n92618 );
not ( n92620 , n92619 );
not ( n415177 , n415017 );
not ( n415178 , n415177 );
not ( n92623 , n414924 );
not ( n92624 , n414952 );
not ( n92625 , n92624 );
or ( n92626 , n92623 , n92625 );
nand ( n92627 , n414952 , n414921 );
nand ( n415184 , n92626 , n92627 );
not ( n415185 , n415184 );
and ( n92630 , n415178 , n415185 );
and ( n415187 , n415177 , n415184 );
nor ( n415188 , n92630 , n415187 );
not ( n415189 , n415188 );
nand ( n415190 , n92620 , n415189 );
buf ( n415191 , n415190 );
not ( n415192 , n415188 );
not ( n415193 , n92619 );
or ( n92638 , n415192 , n415193 );
xor ( n415195 , n414886 , n414904 );
xor ( n415196 , n415195 , n414909 );
buf ( n415197 , n415196 );
nand ( n415198 , n92638 , n415197 );
buf ( n415199 , n415198 );
nand ( n415200 , n415191 , n415199 );
buf ( n415201 , n415200 );
buf ( n415202 , n415201 );
not ( n415203 , n415202 );
xor ( n415204 , n414914 , n415022 );
xor ( n92649 , n415204 , n415036 );
buf ( n415206 , n92649 );
buf ( n415207 , n415206 );
not ( n92652 , n415207 );
buf ( n415209 , n92652 );
buf ( n415210 , n415209 );
not ( n92655 , n415210 );
or ( n92656 , n415203 , n92655 );
buf ( n415213 , n415201 );
not ( n92658 , n415213 );
buf ( n415215 , n415206 );
nand ( n92660 , n92658 , n415215 );
buf ( n415217 , n92660 );
buf ( n415218 , n415217 );
nand ( n415219 , n92656 , n415218 );
buf ( n415220 , n415219 );
buf ( n415221 , n415220 );
buf ( n415222 , n380356 );
not ( n92667 , n415222 );
and ( n415224 , n74977 , n380368 );
not ( n92669 , n74977 );
buf ( n415226 , n380368 );
not ( n415227 , n415226 );
buf ( n415228 , n415227 );
and ( n415229 , n92669 , n415228 );
or ( n415230 , n415224 , n415229 );
buf ( n415231 , n415230 );
not ( n92676 , n415231 );
or ( n415233 , n92667 , n92676 );
and ( n92678 , n31311 , n415228 );
not ( n415235 , n31311 );
and ( n415236 , n415235 , n380368 );
or ( n92681 , n92678 , n415236 );
buf ( n415238 , n92681 );
buf ( n415239 , n380401 );
nand ( n92684 , n415238 , n415239 );
buf ( n415241 , n92684 );
buf ( n415242 , n415241 );
nand ( n92687 , n415233 , n415242 );
buf ( n415244 , n92687 );
buf ( n415245 , n415244 );
not ( n415246 , n415245 );
buf ( n415247 , n415246 );
buf ( n415248 , n415247 );
and ( n415249 , n415221 , n415248 );
not ( n92694 , n415221 );
buf ( n415251 , n415244 );
and ( n415252 , n92694 , n415251 );
nor ( n92697 , n415249 , n415252 );
buf ( n92698 , n92697 );
buf ( n415255 , n92698 );
not ( n92700 , n415255 );
buf ( n92701 , n92700 );
buf ( n415258 , n92701 );
buf ( n415259 , n92301 );
buf ( n415260 , n91666 );
xor ( n415261 , n415259 , n415260 );
buf ( n415262 , n414849 );
xor ( n415263 , n415261 , n415262 );
buf ( n415264 , n415263 );
buf ( n92709 , n415264 );
buf ( n415266 , n380356 );
not ( n92711 , n415266 );
buf ( n415268 , n92681 );
not ( n415269 , n415268 );
or ( n415270 , n92711 , n415269 );
and ( n92715 , n415228 , n351062 );
not ( n92716 , n415228 );
and ( n415273 , n92716 , n365384 );
or ( n92718 , n92715 , n415273 );
buf ( n415275 , n92718 );
buf ( n415276 , n380401 );
nand ( n92721 , n415275 , n415276 );
buf ( n415278 , n92721 );
buf ( n415279 , n415278 );
nand ( n92724 , n415270 , n415279 );
buf ( n415281 , n92724 );
buf ( n415282 , n415281 );
not ( n92727 , n415282 );
xor ( n415284 , n92278 , n91688 );
buf ( n415285 , n414843 );
not ( n415286 , n415285 );
buf ( n415287 , n415286 );
xor ( n92732 , n415284 , n415287 );
buf ( n415289 , n92732 );
not ( n92734 , n415289 );
or ( n92735 , n92727 , n92734 );
buf ( n415292 , n415281 );
buf ( n415293 , n92732 );
or ( n92738 , n415292 , n415293 );
buf ( n415295 , n414326 );
not ( n415296 , n415295 );
buf ( n415297 , n414334 );
not ( n92742 , n415297 );
buf ( n415299 , n414830 );
not ( n92744 , n415299 );
or ( n92745 , n92742 , n92744 );
buf ( n415302 , n414830 );
buf ( n415303 , n414334 );
or ( n415304 , n415302 , n415303 );
nand ( n92749 , n92745 , n415304 );
buf ( n92750 , n92749 );
buf ( n415307 , n92750 );
not ( n92752 , n415307 );
and ( n92753 , n415296 , n92752 );
buf ( n415310 , n414326 );
buf ( n415311 , n92750 );
and ( n92756 , n415310 , n415311 );
nor ( n415313 , n92753 , n92756 );
buf ( n415314 , n415313 );
buf ( n415315 , n415314 );
not ( n92760 , n415315 );
buf ( n415317 , n414222 );
not ( n415318 , n415317 );
buf ( n415319 , n415318 );
buf ( n415320 , n415319 );
buf ( n415321 , n58923 );
and ( n92766 , n415320 , n415321 );
and ( n92767 , n352353 , n379365 );
not ( n415324 , n352353 );
and ( n92769 , n415324 , n379368 );
or ( n92770 , n92767 , n92769 );
buf ( n415327 , n92770 );
buf ( n415328 , n414059 );
and ( n415329 , n415327 , n415328 );
buf ( n415330 , n415329 );
buf ( n415331 , n415330 );
nor ( n415332 , n92766 , n415331 );
buf ( n415333 , n415332 );
buf ( n415334 , n415333 );
not ( n92779 , n415334 );
or ( n92780 , n92760 , n92779 );
xor ( n415337 , n91802 , n414786 );
xor ( n92782 , n415337 , n414826 );
buf ( n415339 , n92782 );
buf ( n415340 , n415339 );
not ( n92785 , n415340 );
buf ( n415342 , n92785 );
buf ( n415343 , n415342 );
not ( n92788 , n415343 );
buf ( n415345 , n379890 );
not ( n92790 , n415345 );
buf ( n415347 , n415104 );
not ( n92792 , n415347 );
or ( n92793 , n92790 , n92792 );
buf ( n415350 , n414963 );
buf ( n415351 , n90092 );
and ( n92796 , n415350 , n415351 );
not ( n92797 , n415350 );
buf ( n415354 , n377754 );
and ( n92799 , n92797 , n415354 );
nor ( n92800 , n92796 , n92799 );
buf ( n415357 , n92800 );
buf ( n415358 , n415357 );
buf ( n415359 , n379912 );
nand ( n415360 , n415358 , n415359 );
buf ( n415361 , n415360 );
buf ( n415362 , n415361 );
nand ( n92807 , n92793 , n415362 );
buf ( n415364 , n92807 );
buf ( n415365 , n415364 );
not ( n92810 , n415365 );
buf ( n415367 , n368590 );
buf ( n415368 , n378098 );
nand ( n415369 , n415367 , n415368 );
buf ( n415370 , n415369 );
buf ( n415371 , n415370 );
not ( n92816 , n415371 );
buf ( n415373 , n92816 );
buf ( n415374 , n415373 );
not ( n92819 , n415374 );
or ( n415376 , n92810 , n92819 );
buf ( n415377 , n415364 );
not ( n92822 , n415377 );
buf ( n415379 , n92822 );
buf ( n415380 , n415379 );
not ( n92825 , n415380 );
buf ( n415382 , n415370 );
not ( n92827 , n415382 );
or ( n92828 , n92825 , n92827 );
buf ( n415385 , n377094 );
not ( n92830 , n415385 );
buf ( n415387 , n368561 );
not ( n92832 , n415387 );
or ( n92833 , n92830 , n92832 );
buf ( n92834 , n410296 );
buf ( n415391 , n413997 );
nand ( n415392 , n92834 , n415391 );
buf ( n415393 , n415392 );
buf ( n415394 , n415393 );
nand ( n415395 , n92833 , n415394 );
buf ( n415396 , n415395 );
buf ( n415397 , n415396 );
not ( n92842 , n415397 );
buf ( n415399 , n369801 );
not ( n92844 , n415399 );
or ( n92845 , n92842 , n92844 );
buf ( n415402 , n49588 );
not ( n92847 , n415402 );
buf ( n415404 , n415125 );
nand ( n92849 , n92847 , n415404 );
buf ( n415406 , n92849 );
buf ( n415407 , n415406 );
nand ( n92852 , n92845 , n415407 );
buf ( n415409 , n92852 );
buf ( n415410 , n415409 );
nand ( n415411 , n92828 , n415410 );
buf ( n415412 , n415411 );
buf ( n415413 , n415412 );
nand ( n92858 , n415376 , n415413 );
buf ( n415415 , n92858 );
buf ( n415416 , n415415 );
not ( n92861 , n415416 );
buf ( n415418 , n92861 );
buf ( n415419 , n415418 );
not ( n415420 , n415419 );
or ( n415421 , n92788 , n415420 );
xor ( n92866 , n414743 , n414747 );
xor ( n415423 , n92866 , n414776 );
buf ( n415424 , n415423 );
buf ( n415425 , n415424 );
xor ( n415426 , n414505 , n91965 );
xor ( n92871 , n415426 , n414578 );
xor ( n92872 , n414635 , n414737 );
xor ( n415429 , n92871 , n92872 );
buf ( n415430 , n415429 );
buf ( n415431 , n382627 );
buf ( n415432 , n406746 );
and ( n415433 , n415431 , n415432 );
buf ( n415434 , n384089 );
buf ( n415435 , n406749 );
and ( n92880 , n415434 , n415435 );
nor ( n92881 , n415433 , n92880 );
buf ( n415438 , n92881 );
buf ( n415439 , n415438 );
buf ( n415440 , n384082 );
or ( n92885 , n415439 , n415440 );
buf ( n415442 , n384092 );
nand ( n92887 , n92885 , n415442 );
buf ( n415444 , n92887 );
buf ( n415445 , n403795 );
buf ( n415446 , n394840 );
and ( n92891 , n415445 , n415446 );
buf ( n415448 , n403798 );
buf ( n415449 , n384408 );
and ( n92894 , n415448 , n415449 );
nor ( n92895 , n92891 , n92894 );
buf ( n415452 , n92895 );
buf ( n415453 , n415452 );
buf ( n415454 , n394838 );
or ( n415455 , n415453 , n415454 );
buf ( n415456 , n403772 );
buf ( n415457 , n394840 );
and ( n92902 , n415456 , n415457 );
buf ( n415459 , n403775 );
buf ( n415460 , n384408 );
and ( n92905 , n415459 , n415460 );
nor ( n92906 , n92902 , n92905 );
buf ( n415463 , n92906 );
buf ( n415464 , n415463 );
buf ( n415465 , n394835 );
or ( n92910 , n415464 , n415465 );
nand ( n92911 , n415455 , n92910 );
buf ( n415468 , n92911 );
xor ( n92913 , n415444 , n415468 );
xor ( n92914 , n414685 , n414690 );
buf ( n415471 , n92914 );
and ( n92916 , n92913 , n415471 );
and ( n415473 , n415444 , n415468 );
or ( n415474 , n92916 , n415473 );
xor ( n92919 , n92095 , n414667 );
xor ( n415476 , n92919 , n414692 );
and ( n92921 , n415474 , n415476 );
buf ( n415478 , n415463 );
buf ( n415479 , n394838 );
or ( n415480 , n415478 , n415479 );
buf ( n415481 , n414704 );
buf ( n415482 , n394835 );
or ( n92927 , n415481 , n415482 );
nand ( n92928 , n415480 , n92927 );
buf ( n415485 , n92928 );
buf ( n415486 , n415485 );
buf ( n415487 , n384354 );
buf ( n415488 , n415438 );
or ( n92933 , n415487 , n415488 );
buf ( n415490 , n414553 );
buf ( n415491 , n384082 );
or ( n92936 , n415490 , n415491 );
nand ( n92937 , n92933 , n92936 );
buf ( n415494 , n92937 );
buf ( n415495 , n415494 );
xor ( n415496 , n415486 , n415495 );
buf ( n415497 , n382659 );
buf ( n415498 , n623 );
or ( n92943 , n415497 , n415498 );
buf ( n415500 , n382655 );
buf ( n415501 , n382835 );
buf ( n415502 , n623 );
and ( n92947 , n415500 , n415501 , n415502 );
buf ( n92948 , n382667 );
not ( n92949 , n92948 );
buf ( n415506 , n92949 );
buf ( n415507 , n415506 );
nor ( n415508 , n92947 , n415507 );
buf ( n415509 , n415508 );
buf ( n415510 , n415509 );
nand ( n415511 , n92943 , n415510 );
buf ( n415512 , n415511 );
buf ( n415513 , n415512 );
xor ( n415514 , n415496 , n415513 );
buf ( n415515 , n415514 );
xor ( n415516 , n92095 , n414667 );
xor ( n415517 , n415516 , n414692 );
and ( n92962 , n415515 , n415517 );
and ( n415519 , n415474 , n415515 );
or ( n415520 , n92921 , n92962 , n415519 );
buf ( n415521 , n415520 );
xor ( n415522 , n415486 , n415495 );
and ( n92967 , n415522 , n415513 );
and ( n92968 , n415486 , n415495 );
or ( n92969 , n92967 , n92968 );
buf ( n415526 , n92969 );
buf ( n415527 , n415526 );
xor ( n92972 , n415521 , n415527 );
xor ( n415529 , n414696 , n414713 );
xor ( n92974 , n415529 , n414718 );
buf ( n415531 , n92974 );
buf ( n415532 , n415531 );
and ( n92977 , n92972 , n415532 );
and ( n415534 , n415521 , n415527 );
or ( n92979 , n92977 , n415534 );
buf ( n415536 , n92979 );
buf ( n415537 , n415536 );
xor ( n92982 , n414723 , n414727 );
xor ( n92983 , n92982 , n414733 );
buf ( n415540 , n92983 );
buf ( n415541 , n415540 );
xor ( n415542 , n415537 , n415541 );
buf ( n415543 , n379890 );
not ( n415544 , n415543 );
buf ( n415545 , n379253 );
not ( n92990 , n415545 );
buf ( n415547 , n414618 );
not ( n92992 , n415547 );
or ( n92993 , n92990 , n92992 );
buf ( n92994 , n377119 );
buf ( n92995 , n379250 );
nand ( n92996 , n92994 , n92995 );
buf ( n92997 , n92996 );
buf ( n415554 , n92997 );
nand ( n92999 , n92993 , n415554 );
buf ( n415556 , n92999 );
buf ( n415557 , n415556 );
not ( n415558 , n415557 );
or ( n93003 , n415544 , n415558 );
buf ( n415560 , n379253 );
buf ( n415561 , n379472 );
and ( n93006 , n415560 , n415561 );
not ( n93007 , n415560 );
buf ( n415564 , n92200 );
and ( n93009 , n93007 , n415564 );
nor ( n415566 , n93006 , n93009 );
buf ( n415567 , n415566 );
buf ( n415568 , n415567 );
buf ( n415569 , n379912 );
nand ( n415570 , n415568 , n415569 );
buf ( n415571 , n415570 );
buf ( n415572 , n415571 );
nand ( n93017 , n93003 , n415572 );
buf ( n415574 , n93017 );
buf ( n415575 , n415574 );
and ( n93020 , n415542 , n415575 );
and ( n93021 , n415537 , n415541 );
or ( n93022 , n93020 , n93021 );
buf ( n415579 , n93022 );
buf ( n415580 , n415579 );
xor ( n93025 , n415430 , n415580 );
buf ( n415582 , n379293 );
not ( n415583 , n415582 );
buf ( n415584 , n378840 );
not ( n415585 , n415584 );
buf ( n415586 , n57145 );
not ( n93031 , n415586 );
or ( n415588 , n415585 , n93031 );
buf ( n415589 , n377571 );
buf ( n415590 , n378840 );
not ( n93035 , n415590 );
buf ( n415592 , n93035 );
buf ( n415593 , n415592 );
nand ( n415594 , n415589 , n415593 );
buf ( n415595 , n415594 );
buf ( n415596 , n415595 );
nand ( n93041 , n415588 , n415596 );
buf ( n415598 , n93041 );
buf ( n415599 , n415598 );
not ( n93044 , n415599 );
or ( n93045 , n415583 , n93044 );
buf ( n415602 , n414763 );
buf ( n415603 , n379260 );
nand ( n93048 , n415602 , n415603 );
buf ( n415605 , n93048 );
buf ( n415606 , n415605 );
nand ( n93051 , n93045 , n415606 );
buf ( n415608 , n93051 );
buf ( n415609 , n415608 );
and ( n93054 , n93025 , n415609 );
and ( n93055 , n415430 , n415580 );
or ( n415612 , n93054 , n93055 );
buf ( n415613 , n415612 );
buf ( n415614 , n415613 );
xor ( n93059 , n415425 , n415614 );
buf ( n415616 , n407553 );
not ( n415617 , n415616 );
buf ( n415618 , n377065 );
not ( n415619 , n415618 );
buf ( n415620 , n49582 );
not ( n415621 , n415620 );
buf ( n415622 , n415621 );
buf ( n415623 , n415622 );
not ( n415624 , n415623 );
or ( n93069 , n415619 , n415624 );
buf ( n415626 , n377583 );
buf ( n415627 , n415121 );
nand ( n93072 , n415626 , n415627 );
buf ( n415629 , n93072 );
buf ( n415630 , n415629 );
nand ( n93075 , n93069 , n415630 );
buf ( n93076 , n93075 );
buf ( n415633 , n93076 );
not ( n93078 , n415633 );
or ( n415635 , n415617 , n93078 );
buf ( n415636 , n57147 );
not ( n93081 , n415636 );
buf ( n415638 , n378843 );
not ( n415639 , n415638 );
buf ( n415640 , n415622 );
not ( n93085 , n415640 );
or ( n415642 , n415639 , n93085 );
buf ( n415643 , n49582 );
buf ( n415644 , n410976 );
nand ( n415645 , n415643 , n415644 );
buf ( n415646 , n415645 );
buf ( n415647 , n415646 );
nand ( n415648 , n415642 , n415647 );
buf ( n415649 , n415648 );
buf ( n415650 , n415649 );
nand ( n415651 , n93081 , n415650 );
buf ( n415652 , n415651 );
buf ( n415653 , n415652 );
nand ( n93098 , n415635 , n415653 );
buf ( n93099 , n93098 );
buf ( n415656 , n93099 );
and ( n93101 , n93059 , n415656 );
and ( n415658 , n415425 , n415614 );
or ( n415659 , n93101 , n415658 );
buf ( n415660 , n415659 );
buf ( n415661 , n415660 );
xor ( n415662 , n92044 , n414631 );
xor ( n93107 , n415662 , n414781 );
buf ( n415664 , n93107 );
buf ( n415665 , n415664 );
buf ( n415666 , n415649 );
not ( n415667 , n415666 );
buf ( n415668 , n407553 );
not ( n93113 , n415668 );
or ( n415670 , n415667 , n93113 );
buf ( n415671 , n414816 );
buf ( n415672 , n377579 );
nand ( n93117 , n415671 , n415672 );
buf ( n415674 , n93117 );
buf ( n415675 , n415674 );
nand ( n415676 , n415670 , n415675 );
buf ( n415677 , n415676 );
buf ( n415678 , n415677 );
or ( n415679 , n415665 , n415678 );
buf ( n415680 , n415679 );
buf ( n415681 , n415680 );
and ( n415682 , n415661 , n415681 );
buf ( n415683 , n415677 );
buf ( n415684 , n415664 );
and ( n93129 , n415683 , n415684 );
buf ( n415686 , n93129 );
buf ( n415687 , n415686 );
nor ( n415688 , n415682 , n415687 );
buf ( n415689 , n415688 );
buf ( n415690 , n415689 );
not ( n93135 , n415690 );
buf ( n415692 , n93135 );
buf ( n415693 , n415692 );
nand ( n93138 , n415421 , n415693 );
buf ( n93139 , n93138 );
buf ( n415696 , n93139 );
buf ( n415697 , n415415 );
buf ( n415698 , n415339 );
nand ( n93143 , n415697 , n415698 );
buf ( n415700 , n93143 );
buf ( n415701 , n415700 );
nand ( n415702 , n415696 , n415701 );
buf ( n415703 , n415702 );
buf ( n415704 , n415703 );
nand ( n415705 , n92780 , n415704 );
buf ( n415706 , n415705 );
buf ( n415707 , n415706 );
buf ( n415708 , n415314 );
not ( n415709 , n415708 );
buf ( n415710 , n415709 );
buf ( n415711 , n415710 );
buf ( n415712 , n415333 );
not ( n415713 , n415712 );
buf ( n415714 , n415713 );
buf ( n415715 , n415714 );
nand ( n93160 , n415711 , n415715 );
buf ( n415717 , n93160 );
buf ( n415718 , n415717 );
nand ( n93163 , n415707 , n415718 );
buf ( n415720 , n93163 );
buf ( n415721 , n415720 );
nand ( n93166 , n92738 , n415721 );
buf ( n415723 , n93166 );
buf ( n415724 , n415723 );
nand ( n93169 , n92735 , n415724 );
buf ( n415726 , n93169 );
buf ( n415727 , n415726 );
or ( n93172 , n92709 , n415727 );
buf ( n93173 , n93172 );
buf ( n415730 , n93173 );
and ( n93175 , n415258 , n415730 );
buf ( n415732 , n415726 );
buf ( n415733 , n415264 );
and ( n415734 , n415732 , n415733 );
buf ( n415735 , n415734 );
buf ( n415736 , n415735 );
nor ( n93181 , n93175 , n415736 );
buf ( n93182 , n93181 );
buf ( n415739 , n93182 );
not ( n415740 , n415739 );
not ( n93185 , n415244 );
not ( n93186 , n415201 );
or ( n93187 , n93185 , n93186 );
buf ( n415744 , n415244 );
buf ( n415745 , n415201 );
nor ( n93190 , n415744 , n415745 );
buf ( n415747 , n93190 );
or ( n93192 , n415747 , n415209 );
nand ( n93193 , n93187 , n93192 );
buf ( n415750 , n93193 );
not ( n93195 , n415750 );
buf ( n415752 , n415045 );
not ( n415753 , n415752 );
buf ( n415754 , n415057 );
not ( n415755 , n415754 );
or ( n415756 , n415753 , n415755 );
buf ( n415757 , n415040 );
buf ( n415758 , n415054 );
nand ( n415759 , n415757 , n415758 );
buf ( n415760 , n415759 );
buf ( n415761 , n415760 );
nand ( n93206 , n415756 , n415761 );
buf ( n415763 , n93206 );
buf ( n415764 , n415763 );
buf ( n415765 , n414859 );
and ( n415766 , n415764 , n415765 );
not ( n93211 , n415764 );
buf ( n415768 , n414862 );
and ( n415769 , n93211 , n415768 );
nor ( n415770 , n415766 , n415769 );
buf ( n415771 , n415770 );
buf ( n415772 , n415771 );
not ( n415773 , n415772 );
or ( n93218 , n93195 , n415773 );
buf ( n415775 , n415771 );
buf ( n415776 , n93193 );
or ( n93221 , n415775 , n415776 );
nand ( n93222 , n93218 , n93221 );
buf ( n415779 , n93222 );
buf ( n415780 , n415779 );
buf ( n415781 , n413699 );
buf ( n415782 , n91161 );
xor ( n93227 , n415781 , n415782 );
buf ( n415784 , n413809 );
xor ( n415785 , n93227 , n415784 );
buf ( n415786 , n415785 );
buf ( n415787 , n415786 );
xor ( n93232 , n414020 , n414045 );
xor ( n93233 , n93232 , n414066 );
buf ( n415790 , n93233 );
buf ( n415791 , n415790 );
xor ( n93236 , n415787 , n415791 );
buf ( n415793 , n380356 );
not ( n415794 , n415793 );
buf ( n415795 , n91655 );
not ( n415796 , n415795 );
or ( n415797 , n415794 , n415796 );
buf ( n415798 , n415230 );
buf ( n415799 , n380401 );
nand ( n93244 , n415798 , n415799 );
buf ( n415801 , n93244 );
buf ( n415802 , n415801 );
nand ( n415803 , n415797 , n415802 );
buf ( n415804 , n415803 );
buf ( n415805 , n415804 );
xor ( n93250 , n93236 , n415805 );
buf ( n415807 , n93250 );
buf ( n415808 , n415807 );
not ( n93253 , n415808 );
buf ( n415810 , n93253 );
buf ( n415811 , n415810 );
and ( n415812 , n415780 , n415811 );
not ( n415813 , n415780 );
buf ( n415814 , n415807 );
and ( n415815 , n415813 , n415814 );
nor ( n415816 , n415812 , n415815 );
buf ( n415817 , n415816 );
buf ( n415818 , n415817 );
not ( n93263 , n415818 );
or ( n93264 , n415740 , n93263 );
xor ( n415821 , n415732 , n415733 );
buf ( n415822 , n415821 );
xor ( n415823 , n415822 , n92698 );
buf ( n415824 , n415823 );
xor ( n415825 , n92619 , n415197 );
and ( n415826 , n415825 , n415189 );
not ( n93271 , n415825 );
and ( n415828 , n93271 , n415188 );
nor ( n415829 , n415826 , n415828 );
buf ( n415830 , n415829 );
buf ( n415831 , n378098 );
not ( n415832 , n415831 );
buf ( n415833 , n85756 );
not ( n415834 , n415833 );
or ( n415835 , n415832 , n415834 );
buf ( n415836 , n409022 );
buf ( n415837 , n379515 );
nand ( n93282 , n415836 , n415837 );
buf ( n415839 , n93282 );
buf ( n415840 , n415839 );
nand ( n415841 , n415835 , n415840 );
buf ( n415842 , n415841 );
buf ( n415843 , n415842 );
not ( n415844 , n415843 );
buf ( n415845 , n368599 );
not ( n93290 , n415845 );
or ( n415847 , n415844 , n93290 );
buf ( n93292 , n415154 );
buf ( n93293 , n412321 );
nand ( n93294 , n93292 , n93293 );
buf ( n415851 , n93294 );
buf ( n415852 , n415851 );
nand ( n93297 , n415847 , n415852 );
buf ( n415854 , n93297 );
buf ( n415855 , n415854 );
buf ( n415856 , n58923 );
not ( n93301 , n415856 );
buf ( n415858 , n92770 );
not ( n93303 , n415858 );
or ( n415860 , n93301 , n93303 );
and ( n93305 , n408201 , n379368 );
not ( n93306 , n408201 );
and ( n93307 , n93306 , n379365 );
or ( n93308 , n93305 , n93307 );
buf ( n415865 , n93308 );
buf ( n415866 , n414059 );
nand ( n93311 , n415865 , n415866 );
buf ( n415868 , n93311 );
buf ( n415869 , n415868 );
nand ( n93314 , n415860 , n415869 );
buf ( n93315 , n93314 );
buf ( n415872 , n93315 );
or ( n415873 , n415855 , n415872 );
buf ( n415874 , n415873 );
buf ( n415875 , n415874 );
buf ( n415876 , n415109 );
buf ( n415877 , n415098 );
xor ( n93322 , n415876 , n415877 );
buf ( n415879 , n92581 );
xor ( n93324 , n93322 , n415879 );
buf ( n415881 , n93324 );
buf ( n415882 , n415881 );
and ( n93327 , n415875 , n415882 );
buf ( n415884 , n415854 );
buf ( n415885 , n93315 );
and ( n93330 , n415884 , n415885 );
buf ( n415887 , n93330 );
buf ( n415888 , n415887 );
nor ( n93333 , n93327 , n415888 );
buf ( n415890 , n93333 );
and ( n93335 , n92526 , n415140 );
not ( n93336 , n92526 );
and ( n93337 , n93336 , n92583 );
nor ( n93338 , n93335 , n93337 );
not ( n93339 , n415171 );
and ( n93340 , n93338 , n93339 );
not ( n93341 , n93338 );
and ( n93342 , n93341 , n415171 );
nor ( n93343 , n93340 , n93342 );
xor ( n415900 , n415890 , n93343 );
buf ( n415901 , n92718 );
buf ( n415902 , n380356 );
and ( n415903 , n415901 , n415902 );
buf ( n415904 , n380368 );
not ( n93349 , n415904 );
buf ( n415906 , n408236 );
not ( n93351 , n415906 );
or ( n415908 , n93349 , n93351 );
buf ( n415909 , n368656 );
buf ( n415910 , n415228 );
nand ( n93355 , n415909 , n415910 );
buf ( n415912 , n93355 );
buf ( n415913 , n415912 );
nand ( n93358 , n415908 , n415913 );
buf ( n93359 , n93358 );
buf ( n415916 , n93359 );
not ( n415917 , n415916 );
buf ( n93362 , n380401 );
not ( n93363 , n93362 );
buf ( n93364 , n93363 );
buf ( n93365 , n93364 );
nor ( n415922 , n415917 , n93365 );
buf ( n415923 , n415922 );
buf ( n415924 , n415923 );
nor ( n415925 , n415903 , n415924 );
buf ( n415926 , n415925 );
and ( n93371 , n415900 , n415926 );
and ( n93372 , n415890 , n93343 );
or ( n415929 , n93371 , n93372 );
buf ( n415930 , n415929 );
xor ( n415931 , n415830 , n415930 );
buf ( n415932 , n415720 );
buf ( n415933 , n415281 );
xor ( n93378 , n415932 , n415933 );
buf ( n415935 , n92732 );
xnor ( n93380 , n93378 , n415935 );
buf ( n93381 , n93380 );
buf ( n415938 , n93381 );
and ( n415939 , n415931 , n415938 );
and ( n415940 , n415830 , n415930 );
or ( n93385 , n415939 , n415940 );
buf ( n415942 , n93385 );
buf ( n93387 , n415942 );
nand ( n415944 , n415824 , n93387 );
buf ( n415945 , n415944 );
not ( n93390 , n415945 );
and ( n93391 , n415703 , n415333 );
not ( n93392 , n415703 );
and ( n415949 , n93392 , n415714 );
or ( n415950 , n93391 , n415949 );
and ( n415951 , n415950 , n415314 );
not ( n93396 , n415950 );
and ( n415953 , n93396 , n415710 );
nor ( n415954 , n415951 , n415953 );
buf ( n93399 , n415954 );
buf ( n415956 , n415339 );
not ( n415957 , n415956 );
buf ( n415958 , n415689 );
not ( n415959 , n415958 );
or ( n93404 , n415957 , n415959 );
buf ( n415961 , n415689 );
buf ( n415962 , n415339 );
or ( n93407 , n415961 , n415962 );
nand ( n415964 , n93404 , n93407 );
buf ( n415965 , n415964 );
buf ( n415966 , n415965 );
not ( n93411 , n415966 );
buf ( n415968 , n415418 );
not ( n415969 , n415968 );
and ( n415970 , n93411 , n415969 );
buf ( n415971 , n415418 );
buf ( n415972 , n415965 );
and ( n415973 , n415971 , n415972 );
nor ( n415974 , n415970 , n415973 );
buf ( n415975 , n415974 );
buf ( n415976 , n415975 );
buf ( n415977 , n379890 );
not ( n93422 , n415977 );
buf ( n415979 , n415357 );
not ( n93424 , n415979 );
or ( n415981 , n93422 , n93424 );
buf ( n415982 , n412602 );
not ( n93427 , n415982 );
buf ( n415984 , n379253 );
not ( n415985 , n415984 );
or ( n93430 , n93427 , n415985 );
buf ( n415987 , n350988 );
buf ( n93432 , n415987 );
buf ( n415989 , n93432 );
buf ( n415990 , n415989 );
buf ( n415991 , n414963 );
nand ( n415992 , n415990 , n415991 );
buf ( n415993 , n415992 );
buf ( n415994 , n415993 );
nand ( n415995 , n93430 , n415994 );
buf ( n415996 , n415995 );
buf ( n415997 , n415996 );
buf ( n415998 , n411170 );
nand ( n415999 , n415997 , n415998 );
buf ( n416000 , n415999 );
buf ( n416001 , n416000 );
nand ( n416002 , n415981 , n416001 );
buf ( n416003 , n416002 );
buf ( n416004 , n410296 );
not ( n416005 , n49582 );
nand ( n93450 , n416005 , n369789 );
and ( n93451 , n93450 , n378098 );
and ( n93452 , n377583 , n343053 );
nor ( n416009 , n93451 , n93452 );
buf ( n416010 , n416009 );
and ( n416011 , n416004 , n416010 );
buf ( n416012 , n416011 );
xor ( n93457 , n416003 , n416012 );
buf ( n416014 , n379890 );
not ( n416015 , n416014 );
buf ( n416016 , n415996 );
not ( n93461 , n416016 );
or ( n93462 , n416015 , n93461 );
buf ( n416019 , n415556 );
buf ( n416020 , n411170 );
nand ( n93465 , n416019 , n416020 );
buf ( n416022 , n93465 );
buf ( n416023 , n416022 );
nand ( n416024 , n93462 , n416023 );
buf ( n416025 , n416024 );
not ( n416026 , n416025 );
or ( n416027 , n49588 , n379515 );
nand ( n416028 , n416026 , n416027 );
not ( n93473 , n416028 );
buf ( n416030 , n377065 );
not ( n416031 , n416030 );
buf ( n416032 , n57145 );
not ( n416033 , n416032 );
or ( n93478 , n416031 , n416033 );
buf ( n416035 , n414611 );
not ( n93480 , n416035 );
buf ( n416037 , n93480 );
buf ( n416038 , n416037 );
buf ( n416039 , n415121 );
nand ( n416040 , n416038 , n416039 );
buf ( n416041 , n416040 );
buf ( n416042 , n416041 );
nand ( n416043 , n93478 , n416042 );
buf ( n416044 , n416043 );
buf ( n416045 , n416044 );
not ( n416046 , n416045 );
buf ( n416047 , n379293 );
not ( n93492 , n416047 );
or ( n93493 , n416046 , n93492 );
buf ( n416050 , n379260 );
buf ( n416051 , n415598 );
nand ( n416052 , n416050 , n416051 );
buf ( n416053 , n416052 );
buf ( n416054 , n416053 );
nand ( n416055 , n93493 , n416054 );
buf ( n416056 , n416055 );
buf ( n93501 , n416056 );
xor ( n93502 , n415537 , n415541 );
xor ( n416059 , n93502 , n415575 );
buf ( n416060 , n416059 );
buf ( n416061 , n416060 );
xor ( n93506 , n93501 , n416061 );
buf ( n416063 , n412940 );
buf ( n416064 , n57158 );
buf ( n416065 , n377571 );
or ( n416066 , n416064 , n416065 );
buf ( n416067 , n378098 );
nand ( n416068 , n416066 , n416067 );
buf ( n416069 , n416068 );
buf ( n416070 , n416069 );
buf ( n416071 , n57158 );
buf ( n416072 , n377571 );
nand ( n93517 , n416071 , n416072 );
buf ( n416074 , n93517 );
buf ( n416075 , n416074 );
and ( n93520 , n416063 , n416070 , n416075 );
buf ( n93521 , n93520 );
buf ( n416078 , n93521 );
and ( n416079 , n93506 , n416078 );
and ( n93524 , n93501 , n416061 );
or ( n416081 , n416079 , n93524 );
buf ( n416082 , n416081 );
not ( n416083 , n416082 );
or ( n93528 , n93473 , n416083 );
not ( n416085 , n416027 );
nand ( n416086 , n416085 , n416025 );
nand ( n416087 , n93528 , n416086 );
and ( n93532 , n93457 , n416087 );
and ( n93533 , n416003 , n416012 );
or ( n93534 , n93532 , n93533 );
xor ( n93535 , n415683 , n415684 );
buf ( n416092 , n93535 );
buf ( n416093 , n416092 );
buf ( n416094 , n415660 );
xor ( n416095 , n416093 , n416094 );
buf ( n416096 , n416095 );
xor ( n93541 , n93534 , n416096 );
buf ( n416098 , n58923 );
not ( n416099 , n416098 );
buf ( n416100 , n93308 );
not ( n416101 , n416100 );
or ( n416102 , n416099 , n416101 );
buf ( n416103 , n379368 );
not ( n93548 , n416103 );
buf ( n416105 , n377349 );
not ( n93550 , n416105 );
or ( n416107 , n93548 , n93550 );
buf ( n93552 , n409020 );
buf ( n93553 , n379365 );
nand ( n93554 , n93552 , n93553 );
buf ( n93555 , n93554 );
buf ( n416112 , n93555 );
nand ( n416113 , n416107 , n416112 );
buf ( n416114 , n416113 );
buf ( n416115 , n416114 );
buf ( n93560 , n414059 );
nand ( n416117 , n416115 , n93560 );
buf ( n416118 , n416117 );
buf ( n416119 , n416118 );
nand ( n93564 , n416102 , n416119 );
buf ( n416121 , n93564 );
and ( n416122 , n93541 , n416121 );
and ( n93567 , n93534 , n416096 );
or ( n416124 , n416122 , n93567 );
buf ( n416125 , n416124 );
not ( n93570 , n416125 );
buf ( n93571 , n93570 );
buf ( n416128 , n93571 );
xor ( n93573 , n415976 , n416128 );
buf ( n416130 , n93359 );
buf ( n416131 , n380356 );
and ( n93576 , n416130 , n416131 );
buf ( n416133 , n351043 );
buf ( n416134 , n380368 );
xor ( n416135 , n416133 , n416134 );
buf ( n416136 , n416135 );
buf ( n416137 , n416136 );
not ( n416138 , n416137 );
buf ( n93583 , n93364 );
nor ( n93584 , n416138 , n93583 );
buf ( n416141 , n93584 );
buf ( n416142 , n416141 );
nor ( n93587 , n93576 , n416142 );
buf ( n416144 , n93587 );
buf ( n416145 , n416144 );
and ( n416146 , n93573 , n416145 );
and ( n93591 , n415976 , n416128 );
or ( n416148 , n416146 , n93591 );
buf ( n416149 , n416148 );
buf ( n416150 , n416149 );
xor ( n93595 , n93399 , n416150 );
xor ( n416152 , n415890 , n93343 );
xor ( n93597 , n416152 , n415926 );
buf ( n416154 , n93597 );
and ( n93599 , n93595 , n416154 );
and ( n416156 , n93399 , n416150 );
or ( n93601 , n93599 , n416156 );
buf ( n416158 , n93601 );
buf ( n416159 , n416158 );
not ( n93604 , n416159 );
xor ( n416161 , n415830 , n415930 );
xor ( n416162 , n416161 , n415938 );
buf ( n416163 , n416162 );
buf ( n416164 , n416163 );
not ( n416165 , n416164 );
or ( n416166 , n93604 , n416165 );
buf ( n93611 , n415364 );
buf ( n416168 , n415409 );
xor ( n416169 , n93611 , n416168 );
buf ( n416170 , n415370 );
xnor ( n93615 , n416169 , n416170 );
buf ( n416172 , n93615 );
buf ( n416173 , n416172 );
buf ( n416174 , n380356 );
not ( n93619 , n416174 );
buf ( n416176 , n416136 );
not ( n93621 , n416176 );
or ( n416178 , n93619 , n93621 );
buf ( n416179 , n380368 );
not ( n93624 , n416179 );
buf ( n416181 , n406930 );
not ( n93626 , n416181 );
or ( n416183 , n93624 , n93626 );
buf ( n416184 , n49172 );
buf ( n416185 , n380364 );
nand ( n416186 , n416184 , n416185 );
buf ( n416187 , n416186 );
buf ( n416188 , n416187 );
nand ( n416189 , n416183 , n416188 );
buf ( n416190 , n416189 );
buf ( n416191 , n416190 );
buf ( n416192 , n380401 );
nand ( n416193 , n416191 , n416192 );
buf ( n416194 , n416193 );
buf ( n416195 , n416194 );
nand ( n416196 , n416178 , n416195 );
buf ( n416197 , n416196 );
buf ( n416198 , n416197 );
or ( n416199 , n416173 , n416198 );
xor ( n93644 , n415425 , n415614 );
xor ( n416201 , n93644 , n415656 );
buf ( n416202 , n416201 );
buf ( n416203 , n416202 );
buf ( n416204 , n378098 );
not ( n416205 , n416204 );
buf ( n416206 , n368561 );
not ( n93651 , n416206 );
or ( n93652 , n416205 , n93651 );
buf ( n416209 , n410296 );
buf ( n416210 , n379515 );
nand ( n416211 , n416209 , n416210 );
buf ( n416212 , n416211 );
buf ( n416213 , n416212 );
nand ( n93658 , n93652 , n416213 );
buf ( n93659 , n93658 );
buf ( n416216 , n93659 );
not ( n416217 , n416216 );
buf ( n416218 , n369801 );
not ( n416219 , n416218 );
or ( n416220 , n416217 , n416219 );
buf ( n93665 , n415396 );
buf ( n416222 , n369809 );
nand ( n416223 , n93665 , n416222 );
buf ( n416224 , n416223 );
buf ( n416225 , n416224 );
nand ( n93670 , n416220 , n416225 );
buf ( n93671 , n93670 );
buf ( n416228 , n93671 );
xor ( n416229 , n416203 , n416228 );
buf ( n416230 , n58923 );
not ( n416231 , n416230 );
buf ( n416232 , n416114 );
not ( n93677 , n416232 );
or ( n93678 , n416231 , n93677 );
buf ( n416235 , n379368 );
not ( n93680 , n416235 );
buf ( n416237 , n377776 );
not ( n416238 , n416237 );
or ( n93683 , n93680 , n416238 );
buf ( n416240 , n351027 );
buf ( n416241 , n379365 );
nand ( n93686 , n416240 , n416241 );
buf ( n416243 , n93686 );
buf ( n416244 , n416243 );
nand ( n416245 , n93683 , n416244 );
buf ( n416246 , n416245 );
buf ( n416247 , n416246 );
buf ( n416248 , n414059 );
nand ( n93693 , n416247 , n416248 );
buf ( n416250 , n93693 );
buf ( n416251 , n416250 );
nand ( n416252 , n93678 , n416251 );
buf ( n416253 , n416252 );
buf ( n416254 , n416253 );
and ( n93699 , n416229 , n416254 );
and ( n93700 , n416203 , n416228 );
or ( n416257 , n93699 , n93700 );
buf ( n416258 , n416257 );
buf ( n416259 , n416258 );
nand ( n416260 , n416199 , n416259 );
buf ( n416261 , n416260 );
buf ( n416262 , n416261 );
buf ( n93707 , n416197 );
buf ( n416264 , n416172 );
nand ( n416265 , n93707 , n416264 );
buf ( n416266 , n416265 );
buf ( n416267 , n416266 );
nand ( n416268 , n416262 , n416267 );
buf ( n416269 , n416268 );
buf ( n416270 , n416269 );
not ( n93715 , n416270 );
buf ( n416272 , n93315 );
buf ( n416273 , n415881 );
xor ( n93718 , n416272 , n416273 );
buf ( n416275 , n415854 );
xor ( n93720 , n93718 , n416275 );
buf ( n416277 , n93720 );
buf ( n416278 , n416277 );
not ( n416279 , n416278 );
or ( n93724 , n93715 , n416279 );
buf ( n416281 , n416269 );
not ( n416282 , n416281 );
buf ( n416283 , n416282 );
buf ( n416284 , n416283 );
not ( n416285 , n416284 );
buf ( n93730 , n416277 );
not ( n93731 , n93730 );
buf ( n93732 , n93731 );
buf ( n416289 , n93732 );
not ( n93734 , n416289 );
or ( n416291 , n416285 , n93734 );
xor ( n93736 , n415976 , n416128 );
xor ( n416293 , n93736 , n416145 );
buf ( n416294 , n416293 );
buf ( n416295 , n416294 );
not ( n416296 , n416295 );
buf ( n416297 , n416296 );
buf ( n416298 , n416297 );
nand ( n416299 , n416291 , n416298 );
buf ( n416300 , n416299 );
buf ( n416301 , n416300 );
nand ( n416302 , n93724 , n416301 );
buf ( n416303 , n416302 );
buf ( n416304 , n416303 );
not ( n416305 , n416304 );
xor ( n93750 , n93399 , n416150 );
xor ( n416307 , n93750 , n416154 );
buf ( n416308 , n416307 );
buf ( n416309 , n416308 );
nand ( n416310 , n416305 , n416309 );
buf ( n416311 , n416310 );
not ( n416312 , n416311 );
buf ( n416313 , n416258 );
buf ( n416314 , n416172 );
xor ( n93759 , n416313 , n416314 );
buf ( n416316 , n416197 );
xnor ( n416317 , n93759 , n416316 );
buf ( n416318 , n416317 );
buf ( n416319 , n416318 );
not ( n416320 , n416319 );
xor ( n93765 , n415430 , n415580 );
xor ( n93766 , n93765 , n415609 );
buf ( n416323 , n93766 );
buf ( n416324 , n416323 );
buf ( n416325 , n407553 );
not ( n93770 , n416325 );
buf ( n416327 , n377094 );
not ( n416328 , n416327 );
buf ( n416329 , n415622 );
not ( n93774 , n416329 );
or ( n93775 , n416328 , n93774 );
buf ( n416332 , n377583 );
buf ( n416333 , n413997 );
nand ( n416334 , n416332 , n416333 );
buf ( n416335 , n416334 );
buf ( n416336 , n416335 );
nand ( n93781 , n93775 , n416336 );
buf ( n93782 , n93781 );
buf ( n416339 , n93782 );
not ( n93784 , n416339 );
or ( n416341 , n93770 , n93784 );
buf ( n93786 , n93076 );
buf ( n93787 , n76050 );
nand ( n93788 , n93786 , n93787 );
buf ( n416345 , n93788 );
buf ( n416346 , n416345 );
nand ( n93791 , n416341 , n416346 );
buf ( n416348 , n93791 );
buf ( n416349 , n416348 );
xor ( n93794 , n416324 , n416349 );
buf ( n416351 , n58923 );
not ( n416352 , n416351 );
buf ( n416353 , n416246 );
not ( n416354 , n416353 );
or ( n93799 , n416352 , n416354 );
buf ( n416356 , n379368 );
not ( n416357 , n416356 );
buf ( n416358 , n409052 );
not ( n93803 , n416358 );
or ( n416360 , n416357 , n93803 );
buf ( n416361 , n377754 );
buf ( n416362 , n379365 );
nand ( n93807 , n416361 , n416362 );
buf ( n416364 , n93807 );
buf ( n416365 , n416364 );
nand ( n93810 , n416360 , n416365 );
buf ( n416367 , n93810 );
buf ( n416368 , n416367 );
buf ( n416369 , n414059 );
nand ( n416370 , n416368 , n416369 );
buf ( n416371 , n416370 );
buf ( n416372 , n416371 );
nand ( n93817 , n93799 , n416372 );
buf ( n416374 , n93817 );
buf ( n416375 , n416374 );
and ( n416376 , n93794 , n416375 );
and ( n93821 , n416324 , n416349 );
or ( n93822 , n416376 , n93821 );
buf ( n416379 , n93822 );
buf ( n93824 , n416379 );
xor ( n416381 , n416003 , n416012 );
xor ( n93826 , n416381 , n416087 );
buf ( n416383 , n93826 );
xor ( n416384 , n93824 , n416383 );
xor ( n93829 , n416203 , n416228 );
xor ( n93830 , n93829 , n416254 );
buf ( n416387 , n93830 );
buf ( n416388 , n416387 );
and ( n93833 , n416384 , n416388 );
and ( n93834 , n93824 , n416383 );
or ( n93835 , n93833 , n93834 );
buf ( n416392 , n93835 );
not ( n93837 , n416392 );
xor ( n93838 , n93534 , n416096 );
xor ( n93839 , n93838 , n416121 );
buf ( n416396 , n93839 );
not ( n93841 , n416396 );
buf ( n416398 , n93841 );
not ( n93843 , n416398 );
or ( n93844 , n93837 , n93843 );
not ( n93845 , n416392 );
nand ( n416402 , n93845 , n93839 );
nand ( n93847 , n93844 , n416402 );
buf ( n416404 , n93847 );
not ( n416405 , n416404 );
and ( n93850 , n416320 , n416405 );
buf ( n416407 , n416318 );
buf ( n416408 , n93847 );
and ( n93853 , n416407 , n416408 );
nor ( n416410 , n93850 , n93853 );
buf ( n416411 , n416410 );
buf ( n416412 , n416411 );
xor ( n416413 , n415521 , n415527 );
xor ( n93858 , n416413 , n415532 );
buf ( n416415 , n93858 );
buf ( n416416 , n416415 );
buf ( n416417 , n415567 );
not ( n93862 , n416417 );
buf ( n416419 , n379890 );
not ( n93864 , n416419 );
or ( n416421 , n93862 , n93864 );
buf ( n93866 , n379912 );
and ( n93867 , n379250 , n378840 );
not ( n416424 , n379250 );
and ( n93869 , n416424 , n415592 );
or ( n416426 , n93867 , n93869 );
buf ( n416427 , n416426 );
nand ( n416428 , n93866 , n416427 );
buf ( n416429 , n416428 );
buf ( n416430 , n416429 );
nand ( n416431 , n416421 , n416430 );
buf ( n416432 , n416431 );
buf ( n416433 , n416432 );
xor ( n93878 , n416416 , n416433 );
buf ( n416435 , n405813 );
buf ( n416436 , n394840 );
and ( n416437 , n416435 , n416436 );
buf ( n416438 , n405816 );
buf ( n416439 , n384408 );
and ( n93884 , n416438 , n416439 );
nor ( n93885 , n416437 , n93884 );
buf ( n416442 , n93885 );
buf ( n416443 , n416442 );
buf ( n416444 , n394838 );
or ( n93889 , n416443 , n416444 );
buf ( n416446 , n415452 );
buf ( n416447 , n394835 );
or ( n93892 , n416446 , n416447 );
nand ( n416449 , n93889 , n93892 );
buf ( n416450 , n416449 );
buf ( n416451 , n63425 );
buf ( n416452 , n623 );
and ( n416453 , n416451 , n416452 );
buf ( n416454 , n382627 );
buf ( n416455 , n63425 );
not ( n416456 , n416455 );
buf ( n416457 , n416456 );
buf ( n416458 , n416457 );
buf ( n416459 , n85590 );
and ( n93904 , n416458 , n416459 );
buf ( n416461 , n90113 );
nor ( n93906 , n93904 , n416461 );
buf ( n416463 , n93906 );
buf ( n416464 , n416463 );
nor ( n93909 , n416453 , n416454 , n416464 );
buf ( n416466 , n93909 );
xor ( n416467 , n416450 , n416466 );
buf ( n416468 , n384414 );
buf ( n416469 , n90113 );
buf ( n416470 , n406746 );
and ( n416471 , n416469 , n416470 );
buf ( n416472 , n384421 );
buf ( n416473 , n406749 );
and ( n93918 , n416472 , n416473 );
nor ( n93919 , n416471 , n93918 );
buf ( n416476 , n93919 );
buf ( n416477 , n416476 );
or ( n416478 , n416468 , n416477 );
buf ( n416479 , n414677 );
buf ( n416480 , n395635 );
or ( n93925 , n416479 , n416480 );
nand ( n93926 , n416478 , n93925 );
buf ( n416483 , n93926 );
and ( n416484 , n416467 , n416483 );
and ( n93929 , n416450 , n416466 );
or ( n93930 , n416484 , n93929 );
xor ( n416487 , n415444 , n415468 );
xor ( n416488 , n416487 , n415471 );
and ( n93933 , n93930 , n416488 );
buf ( n416490 , n394840 );
buf ( n416491 , n406569 );
and ( n416492 , n416490 , n416491 );
buf ( n416493 , n384408 );
buf ( n416494 , n406572 );
and ( n93939 , n416493 , n416494 );
nor ( n93940 , n416492 , n93939 );
buf ( n416497 , n93940 );
buf ( n416498 , n416497 );
buf ( n416499 , n394838 );
or ( n93944 , n416498 , n416499 );
buf ( n416501 , n416442 );
buf ( n416502 , n394835 );
or ( n416503 , n416501 , n416502 );
nand ( n93948 , n93944 , n416503 );
buf ( n416505 , n93948 );
buf ( n416506 , n416505 );
buf ( n416507 , n384082 );
buf ( n416508 , n85590 );
nor ( n416509 , n416507 , n416508 );
buf ( n416510 , n416509 );
buf ( n416511 , n416510 );
and ( n416512 , n416506 , n416511 );
buf ( n416513 , n416512 );
xor ( n416514 , n416450 , n416466 );
xor ( n93959 , n416514 , n416483 );
and ( n416516 , n416513 , n93959 );
buf ( n416517 , n384092 );
buf ( n416518 , n623 );
or ( n416519 , n416517 , n416518 );
buf ( n416520 , n384085 );
buf ( n416521 , n384343 );
buf ( n416522 , n623 );
and ( n93967 , n416520 , n416521 , n416522 );
buf ( n416524 , n384097 );
not ( n416525 , n416524 );
buf ( n416526 , n416525 );
buf ( n416527 , n416526 );
nor ( n93972 , n93967 , n416527 );
buf ( n416529 , n93972 );
buf ( n416530 , n416529 );
nand ( n416531 , n416519 , n416530 );
buf ( n416532 , n416531 );
xor ( n93977 , n416450 , n416466 );
xor ( n416534 , n93977 , n416483 );
and ( n416535 , n416532 , n416534 );
and ( n416536 , n416513 , n416532 );
or ( n93981 , n416516 , n416535 , n416536 );
xor ( n93982 , n415444 , n415468 );
xor ( n93983 , n93982 , n415471 );
and ( n93984 , n93981 , n93983 );
and ( n93985 , n93930 , n93981 );
or ( n416542 , n93933 , n93984 , n93985 );
buf ( n93987 , n416542 );
xor ( n416544 , n92095 , n414667 );
xor ( n93989 , n416544 , n414692 );
xor ( n416546 , n415474 , n415515 );
xor ( n416547 , n93989 , n416546 );
buf ( n416548 , n416547 );
xor ( n93993 , n93987 , n416548 );
buf ( n416550 , n379912 );
not ( n416551 , n416550 );
buf ( n416552 , n377065 );
not ( n93997 , n416552 );
buf ( n416554 , n379250 );
not ( n93999 , n416554 );
or ( n94000 , n93997 , n93999 );
buf ( n416557 , n379253 );
buf ( n416558 , n415121 );
nand ( n416559 , n416557 , n416558 );
buf ( n416560 , n416559 );
buf ( n416561 , n416560 );
nand ( n416562 , n94000 , n416561 );
buf ( n416563 , n416562 );
buf ( n416564 , n416563 );
not ( n416565 , n416564 );
or ( n416566 , n416551 , n416565 );
buf ( n416567 , n416426 );
buf ( n416568 , n379890 );
nand ( n416569 , n416567 , n416568 );
buf ( n416570 , n416569 );
buf ( n416571 , n416570 );
nand ( n416572 , n416566 , n416571 );
buf ( n416573 , n416572 );
buf ( n416574 , n416573 );
and ( n416575 , n93993 , n416574 );
and ( n94020 , n93987 , n416548 );
or ( n416577 , n416575 , n94020 );
buf ( n416578 , n416577 );
buf ( n416579 , n416578 );
and ( n94024 , n93878 , n416579 );
and ( n94025 , n416416 , n416433 );
or ( n94026 , n94024 , n94025 );
buf ( n416583 , n94026 );
buf ( n416584 , n416583 );
buf ( n416585 , n378098 );
buf ( n416586 , n49582 );
and ( n416587 , n416585 , n416586 );
not ( n94032 , n416585 );
buf ( n416589 , n411431 );
and ( n416590 , n94032 , n416589 );
nor ( n416591 , n416587 , n416590 );
buf ( n416592 , n416591 );
buf ( n416593 , n416592 );
not ( n94038 , n416593 );
buf ( n416595 , n407553 );
not ( n416596 , n416595 );
or ( n416597 , n94038 , n416596 );
buf ( n416598 , n57147 );
not ( n94043 , n416598 );
buf ( n416600 , n93782 );
nand ( n416601 , n94043 , n416600 );
buf ( n416602 , n416601 );
buf ( n416603 , n416602 );
nand ( n416604 , n416597 , n416603 );
buf ( n416605 , n416604 );
buf ( n416606 , n416605 );
xor ( n94051 , n416584 , n416606 );
buf ( n416608 , n58923 );
not ( n94053 , n416608 );
buf ( n416610 , n379368 );
buf ( n416611 , n350988 );
xor ( n94056 , n416610 , n416611 );
buf ( n416613 , n94056 );
buf ( n416614 , n416613 );
not ( n94059 , n416614 );
or ( n94060 , n94053 , n94059 );
xor ( n94061 , n379368 , n377119 );
buf ( n416618 , n94061 );
buf ( n416619 , n414059 );
nand ( n94064 , n416618 , n416619 );
buf ( n416621 , n94064 );
buf ( n416622 , n416621 );
nand ( n94067 , n94060 , n416622 );
buf ( n416624 , n94067 );
buf ( n416625 , n416624 );
not ( n416626 , n416625 );
buf ( n416627 , n377094 );
not ( n94072 , n416627 );
buf ( n416629 , n57145 );
not ( n94074 , n416629 );
or ( n416631 , n94072 , n94074 );
buf ( n94076 , n416037 );
buf ( n94077 , n413997 );
nand ( n94078 , n94076 , n94077 );
buf ( n94079 , n94078 );
buf ( n416636 , n94079 );
nand ( n94081 , n416631 , n416636 );
buf ( n94082 , n94081 );
buf ( n416639 , n94082 );
not ( n416640 , n416639 );
buf ( n416641 , n379293 );
not ( n94086 , n416641 );
or ( n94087 , n416640 , n94086 );
buf ( n416644 , n416044 );
buf ( n416645 , n379260 );
nand ( n416646 , n416644 , n416645 );
buf ( n416647 , n416646 );
buf ( n416648 , n416647 );
nand ( n416649 , n94087 , n416648 );
buf ( n416650 , n416649 );
buf ( n416651 , n416650 );
not ( n416652 , n416651 );
or ( n94097 , n416626 , n416652 );
buf ( n416654 , n416624 );
buf ( n416655 , n416650 );
or ( n94100 , n416654 , n416655 );
xor ( n94101 , n93987 , n416548 );
xor ( n416658 , n94101 , n416574 );
buf ( n416659 , n416658 );
buf ( n416660 , n416659 );
buf ( n416661 , n58923 );
not ( n94106 , n416661 );
buf ( n416663 , n94061 );
not ( n416664 , n416663 );
or ( n416665 , n94106 , n416664 );
and ( n94110 , n379472 , n379365 );
not ( n416667 , n379472 );
and ( n416668 , n416667 , n379368 );
or ( n94113 , n94110 , n416668 );
buf ( n416670 , n94113 );
buf ( n416671 , n414059 );
nand ( n94116 , n416670 , n416671 );
buf ( n416673 , n94116 );
buf ( n416674 , n416673 );
nand ( n416675 , n416665 , n416674 );
buf ( n416676 , n416675 );
buf ( n416677 , n416676 );
xor ( n416678 , n416660 , n416677 );
buf ( n416679 , n377571 );
not ( n416680 , n379287 );
nand ( n94125 , n416680 , n379250 );
buf ( n416682 , n94125 );
buf ( n416683 , n378098 );
and ( n94128 , n416682 , n416683 );
buf ( n416685 , n379287 );
buf ( n416686 , n379253 );
and ( n416687 , n416685 , n416686 );
nor ( n94132 , n94128 , n416687 );
buf ( n94133 , n94132 );
buf ( n416690 , n94133 );
and ( n416691 , n416679 , n416690 );
buf ( n416692 , n416691 );
buf ( n416693 , n416692 );
and ( n416694 , n416678 , n416693 );
and ( n416695 , n416660 , n416677 );
or ( n94140 , n416694 , n416695 );
buf ( n416697 , n94140 );
buf ( n416698 , n416697 );
nand ( n416699 , n94100 , n416698 );
buf ( n416700 , n416699 );
buf ( n416701 , n416700 );
nand ( n94146 , n94097 , n416701 );
buf ( n416703 , n94146 );
buf ( n416704 , n416703 );
and ( n416705 , n94051 , n416704 );
and ( n94150 , n416584 , n416606 );
or ( n416707 , n416705 , n94150 );
buf ( n416708 , n416707 );
buf ( n416709 , n416708 );
xor ( n94154 , n416025 , n416027 );
xnor ( n94155 , n94154 , n416082 );
buf ( n416712 , n94155 );
xor ( n416713 , n416709 , n416712 );
xor ( n94158 , n416324 , n416349 );
xor ( n416715 , n94158 , n416375 );
buf ( n416716 , n416715 );
buf ( n416717 , n416716 );
and ( n94162 , n416713 , n416717 );
and ( n416719 , n416709 , n416712 );
or ( n416720 , n94162 , n416719 );
buf ( n416721 , n416720 );
buf ( n416722 , n416721 );
not ( n416723 , n416722 );
buf ( n416724 , n416723 );
buf ( n416725 , n416724 );
not ( n416726 , n416725 );
buf ( n416727 , n416190 );
buf ( n416728 , n380356 );
and ( n416729 , n416727 , n416728 );
buf ( n416730 , n380368 );
not ( n416731 , n416730 );
buf ( n416732 , n408201 );
not ( n416733 , n416732 );
or ( n416734 , n416731 , n416733 );
buf ( n416735 , n380364 );
buf ( n416736 , n352381 );
nand ( n416737 , n416735 , n416736 );
buf ( n416738 , n416737 );
buf ( n416739 , n416738 );
nand ( n416740 , n416734 , n416739 );
buf ( n416741 , n416740 );
buf ( n416742 , n416741 );
buf ( n416743 , n380401 );
and ( n94188 , n416742 , n416743 );
buf ( n416745 , n94188 );
buf ( n416746 , n416745 );
nor ( n94191 , n416729 , n416746 );
buf ( n94192 , n94191 );
buf ( n416749 , n94192 );
not ( n94194 , n416749 );
or ( n416751 , n416726 , n94194 );
xor ( n416752 , n93824 , n416383 );
xor ( n94197 , n416752 , n416388 );
buf ( n416754 , n94197 );
buf ( n416755 , n416754 );
nand ( n94200 , n416751 , n416755 );
buf ( n94201 , n94200 );
buf ( n416758 , n94201 );
buf ( n416759 , n94192 );
not ( n94204 , n416759 );
buf ( n416761 , n416721 );
nand ( n94206 , n94204 , n416761 );
buf ( n416763 , n94206 );
buf ( n416764 , n416763 );
and ( n94209 , n416758 , n416764 );
buf ( n94210 , n94209 );
buf ( n416767 , n94210 );
nand ( n416768 , n416412 , n416767 );
buf ( n416769 , n416768 );
not ( n416770 , n416769 );
buf ( n94215 , n416650 );
buf ( n416772 , n416624 );
xor ( n94217 , n94215 , n416772 );
buf ( n416774 , n416697 );
xnor ( n416775 , n94217 , n416774 );
buf ( n416776 , n416775 );
buf ( n416777 , n416776 );
not ( n416778 , n416777 );
buf ( n416779 , n416778 );
buf ( n416780 , n416779 );
not ( n416781 , n416780 );
xor ( n94226 , n416416 , n416433 );
xor ( n416783 , n94226 , n416579 );
buf ( n416784 , n416783 );
buf ( n416785 , n416784 );
buf ( n416786 , n377579 );
buf ( n416787 , n378098 );
and ( n94232 , n416786 , n416787 );
buf ( n94233 , n94232 );
buf ( n416790 , n94233 );
xor ( n416791 , n416785 , n416790 );
xor ( n94236 , n415444 , n415468 );
xor ( n416793 , n94236 , n415471 );
xor ( n416794 , n93930 , n93981 );
xor ( n416795 , n416793 , n416794 );
buf ( n416796 , n416795 );
xor ( n416797 , n416506 , n416511 );
buf ( n416798 , n416797 );
buf ( n416799 , n416798 );
buf ( n416800 , n416476 );
buf ( n416801 , n395635 );
or ( n94246 , n416800 , n416801 );
buf ( n416803 , n384424 );
nand ( n416804 , n94246 , n416803 );
buf ( n416805 , n416804 );
buf ( n416806 , n416805 );
xor ( n94251 , n416799 , n416806 );
buf ( n416808 , n384398 );
buf ( n416809 , n623 );
and ( n94254 , n416808 , n416809 );
buf ( n416811 , n90113 );
buf ( n416812 , n384398 );
not ( n94257 , n416812 );
buf ( n94258 , n94257 );
buf ( n416815 , n94258 );
buf ( n416816 , n85590 );
and ( n94261 , n416815 , n416816 );
buf ( n416818 , n394840 );
nor ( n416819 , n94261 , n416818 );
buf ( n416820 , n416819 );
buf ( n416821 , n416820 );
nor ( n416822 , n94254 , n416811 , n416821 );
buf ( n416823 , n416822 );
buf ( n416824 , n416823 );
buf ( n416825 , n394840 );
buf ( n416826 , n406746 );
and ( n94271 , n416825 , n416826 );
buf ( n416828 , n384408 );
buf ( n416829 , n406749 );
and ( n416830 , n416828 , n416829 );
nor ( n416831 , n94271 , n416830 );
buf ( n416832 , n416831 );
buf ( n416833 , n416832 );
buf ( n416834 , n394838 );
or ( n416835 , n416833 , n416834 );
buf ( n416836 , n416497 );
buf ( n416837 , n394835 );
or ( n416838 , n416836 , n416837 );
nand ( n416839 , n416835 , n416838 );
buf ( n416840 , n416839 );
buf ( n416841 , n416840 );
xor ( n94286 , n416824 , n416841 );
buf ( n416843 , n384424 );
buf ( n416844 , n623 );
or ( n416845 , n416843 , n416844 );
buf ( n416846 , n384417 );
buf ( n416847 , n90113 );
buf ( n416848 , n623 );
and ( n416849 , n416846 , n416847 , n416848 );
buf ( n94294 , n384429 );
not ( n416851 , n94294 );
buf ( n416852 , n416851 );
buf ( n416853 , n416852 );
nor ( n416854 , n416849 , n416853 );
buf ( n416855 , n416854 );
buf ( n416856 , n416855 );
nand ( n416857 , n416845 , n416856 );
buf ( n416858 , n416857 );
buf ( n416859 , n416858 );
and ( n416860 , n94286 , n416859 );
and ( n94305 , n416824 , n416841 );
or ( n416862 , n416860 , n94305 );
buf ( n416863 , n416862 );
buf ( n416864 , n416863 );
and ( n416865 , n94251 , n416864 );
and ( n416866 , n416799 , n416806 );
or ( n94311 , n416865 , n416866 );
buf ( n416868 , n94311 );
buf ( n416869 , n416868 );
xor ( n94314 , n416450 , n416466 );
xor ( n416871 , n94314 , n416483 );
xor ( n416872 , n416513 , n416532 );
xor ( n416873 , n416871 , n416872 );
buf ( n416874 , n416873 );
xor ( n416875 , n416869 , n416874 );
buf ( n416876 , n342352 );
not ( n416877 , n416876 );
buf ( n416878 , n379876 );
buf ( n416879 , n379856 );
nor ( n416880 , n416878 , n416879 );
buf ( n416881 , n416880 );
buf ( n416882 , n416881 );
buf ( n416883 , n379515 );
or ( n94328 , n416882 , n416883 );
buf ( n416885 , n379876 );
buf ( n416886 , n379856 );
nand ( n94331 , n416885 , n416886 );
buf ( n416888 , n94331 );
buf ( n416889 , n416888 );
nand ( n94334 , n94328 , n416889 );
buf ( n416891 , n94334 );
buf ( n416892 , n416891 );
nor ( n416893 , n416877 , n416892 );
buf ( n416894 , n416893 );
buf ( n416895 , n416894 );
and ( n416896 , n416875 , n416895 );
and ( n416897 , n416869 , n416874 );
or ( n94342 , n416896 , n416897 );
buf ( n416899 , n94342 );
buf ( n416900 , n416899 );
xor ( n94345 , n416796 , n416900 );
buf ( n416902 , n377094 );
not ( n416903 , n416902 );
buf ( n416904 , n379250 );
not ( n94349 , n416904 );
or ( n416906 , n416903 , n94349 );
buf ( n416907 , n377094 );
not ( n416908 , n416907 );
buf ( n416909 , n342352 );
nand ( n416910 , n416908 , n416909 );
buf ( n416911 , n416910 );
buf ( n416912 , n416911 );
nand ( n94357 , n416906 , n416912 );
buf ( n94358 , n94357 );
buf ( n416915 , n94358 );
not ( n416916 , n416915 );
buf ( n416917 , n379912 );
not ( n416918 , n416917 );
or ( n94363 , n416916 , n416918 );
buf ( n416920 , n416563 );
buf ( n416921 , n379890 );
nand ( n94366 , n416920 , n416921 );
buf ( n416923 , n94366 );
buf ( n416924 , n416923 );
nand ( n94369 , n94363 , n416924 );
buf ( n416926 , n94369 );
buf ( n416927 , n416926 );
and ( n416928 , n94345 , n416927 );
and ( n416929 , n416796 , n416900 );
or ( n416930 , n416928 , n416929 );
buf ( n416931 , n416930 );
buf ( n416932 , n416931 );
nand ( n94377 , n90038 , n378098 );
not ( n94378 , n94377 );
buf ( n416935 , n94378 );
not ( n416936 , n416935 );
and ( n416937 , n94113 , n58923 );
buf ( n416938 , n379856 );
not ( n416939 , n416938 );
buf ( n416940 , n415592 );
not ( n416941 , n416940 );
or ( n94386 , n416939 , n416941 );
buf ( n416943 , n378840 );
buf ( n94388 , n379318 );
nand ( n416945 , n416943 , n94388 );
buf ( n416946 , n416945 );
buf ( n416947 , n416946 );
nand ( n416948 , n94386 , n416947 );
buf ( n416949 , n416948 );
buf ( n416950 , n416949 );
not ( n94395 , n416950 );
buf ( n416952 , n379350 );
nor ( n94397 , n94395 , n416952 );
buf ( n94398 , n94397 );
nor ( n416955 , n416937 , n94398 );
not ( n94400 , n416955 );
buf ( n94401 , n94400 );
not ( n94402 , n94401 );
or ( n94403 , n416936 , n94402 );
buf ( n416960 , n416955 );
not ( n94405 , n416960 );
buf ( n416962 , n94377 );
not ( n416963 , n416962 );
or ( n94408 , n94405 , n416963 );
buf ( n416965 , n58923 );
not ( n416966 , n416965 );
buf ( n416967 , n416949 );
not ( n416968 , n416967 );
or ( n416969 , n416966 , n416968 );
buf ( n416970 , n379350 );
not ( n94415 , n416970 );
buf ( n416972 , n94415 );
buf ( n416973 , n416972 );
buf ( n416974 , n377065 );
buf ( n416975 , n379856 );
and ( n94420 , n416974 , n416975 );
not ( n94421 , n416974 );
buf ( n416978 , n379859 );
and ( n94423 , n94421 , n416978 );
nor ( n416980 , n94420 , n94423 );
buf ( n416981 , n416980 );
buf ( n94426 , n416981 );
nand ( n94427 , n416973 , n94426 );
buf ( n94428 , n94427 );
buf ( n416985 , n94428 );
nand ( n416986 , n416969 , n416985 );
buf ( n416987 , n416986 );
not ( n416988 , n416987 );
buf ( n416989 , n378098 );
not ( n416990 , n416989 );
buf ( n416991 , n379250 );
not ( n94436 , n416991 );
or ( n94437 , n416990 , n94436 );
buf ( n416994 , n342352 );
buf ( n416995 , n379515 );
nand ( n416996 , n416994 , n416995 );
buf ( n416997 , n416996 );
buf ( n416998 , n416997 );
nand ( n416999 , n94437 , n416998 );
buf ( n417000 , n416999 );
not ( n94445 , n417000 );
not ( n417002 , n379912 );
or ( n417003 , n94445 , n417002 );
buf ( n417004 , n94358 );
buf ( n417005 , n379887 );
nand ( n417006 , n417004 , n417005 );
buf ( n417007 , n417006 );
nand ( n417008 , n417003 , n417007 );
not ( n94453 , n417008 );
or ( n417010 , n416988 , n94453 );
buf ( n417011 , n417008 );
buf ( n417012 , n416987 );
nor ( n94457 , n417011 , n417012 );
buf ( n417014 , n94457 );
buf ( n417015 , n58920 );
not ( n94460 , n417015 );
buf ( n417017 , n416981 );
not ( n94462 , n417017 );
or ( n94463 , n94460 , n94462 );
buf ( n417020 , n416972 );
and ( n417021 , n377091 , n379318 );
not ( n417022 , n377091 );
and ( n94467 , n417022 , n379856 );
or ( n417024 , n417021 , n94467 );
buf ( n417025 , n417024 );
nand ( n417026 , n417020 , n417025 );
buf ( n417027 , n417026 );
buf ( n417028 , n417027 );
nand ( n417029 , n94463 , n417028 );
buf ( n417030 , n417029 );
buf ( n417031 , n417030 );
not ( n94476 , n417031 );
buf ( n417033 , n94476 );
buf ( n417034 , n417033 );
buf ( n417035 , n379322 );
not ( n417036 , n417035 );
buf ( n417037 , n379339 );
not ( n417038 , n417037 );
or ( n417039 , n417036 , n417038 );
buf ( n417040 , n379322 );
buf ( n417041 , n379339 );
or ( n417042 , n417040 , n417041 );
buf ( n417043 , n378098 );
nand ( n94488 , n417042 , n417043 );
buf ( n94489 , n94488 );
buf ( n417046 , n94489 );
nand ( n94491 , n417039 , n417046 );
buf ( n417048 , n94491 );
not ( n417049 , n417048 );
nand ( n417050 , n379856 , n417049 );
not ( n94495 , n417050 );
buf ( n417052 , n384411 );
buf ( n417053 , n623 );
nand ( n94498 , n417052 , n417053 );
buf ( n94499 , n94498 );
buf ( n417056 , n94499 );
not ( n417057 , n417056 );
buf ( n417058 , n416832 );
buf ( n417059 , n394835 );
or ( n417060 , n417058 , n417059 );
buf ( n417061 , n394838 );
nand ( n94506 , n417060 , n417061 );
buf ( n94507 , n94506 );
buf ( n417064 , n94507 );
nand ( n94509 , n417057 , n417064 );
buf ( n417066 , n94509 );
not ( n94511 , n417066 );
and ( n94512 , n94495 , n94511 );
buf ( n94513 , n417066 );
buf ( n417070 , n417050 );
nand ( n417071 , n94513 , n417070 );
buf ( n417072 , n417071 );
xor ( n417073 , n416824 , n416841 );
xor ( n94518 , n417073 , n416859 );
buf ( n417075 , n94518 );
and ( n417076 , n417072 , n417075 );
nor ( n417077 , n94512 , n417076 );
buf ( n417078 , n417077 );
nand ( n94523 , n417034 , n417078 );
buf ( n94524 , n94523 );
xor ( n417081 , n416799 , n416806 );
xor ( n417082 , n417081 , n416864 );
buf ( n417083 , n417082 );
and ( n417084 , n94524 , n417083 );
buf ( n417085 , n417077 );
not ( n417086 , n417085 );
buf ( n417087 , n417086 );
and ( n417088 , n417030 , n417087 );
nor ( n94533 , n417084 , n417088 );
or ( n94534 , n417014 , n94533 );
nand ( n94535 , n417010 , n94534 );
buf ( n417092 , n94535 );
nand ( n94537 , n94408 , n417092 );
buf ( n94538 , n94537 );
buf ( n417095 , n94538 );
nand ( n417096 , n94403 , n417095 );
buf ( n417097 , n417096 );
buf ( n417098 , n417097 );
xor ( n417099 , n416932 , n417098 );
buf ( n417100 , n378098 );
not ( n417101 , n417100 );
buf ( n417102 , n57145 );
not ( n417103 , n417102 );
or ( n94548 , n417101 , n417103 );
buf ( n417105 , n377571 );
buf ( n417106 , n379515 );
nand ( n94551 , n417105 , n417106 );
buf ( n417108 , n94551 );
buf ( n417109 , n417108 );
nand ( n94554 , n94548 , n417109 );
buf ( n94555 , n94554 );
buf ( n417112 , n94555 );
not ( n94557 , n417112 );
buf ( n417114 , n379293 );
not ( n417115 , n417114 );
or ( n417116 , n94557 , n417115 );
buf ( n417117 , n94082 );
buf ( n417118 , n379260 );
nand ( n417119 , n417117 , n417118 );
buf ( n417120 , n417119 );
buf ( n94565 , n417120 );
nand ( n417122 , n417116 , n94565 );
buf ( n417123 , n417122 );
buf ( n417124 , n417123 );
and ( n94569 , n417099 , n417124 );
and ( n94570 , n416932 , n417098 );
or ( n94571 , n94569 , n94570 );
buf ( n417128 , n94571 );
buf ( n417129 , n417128 );
xor ( n417130 , n416791 , n417129 );
buf ( n417131 , n417130 );
buf ( n417132 , n417131 );
not ( n417133 , n417132 );
or ( n417134 , n416781 , n417133 );
xor ( n94579 , n416660 , n416677 );
xor ( n417136 , n94579 , n416693 );
buf ( n417137 , n417136 );
buf ( n417138 , n417137 );
xor ( n417139 , n416932 , n417098 );
xor ( n417140 , n417139 , n417124 );
buf ( n417141 , n417140 );
buf ( n417142 , n417141 );
xor ( n94587 , n417138 , n417142 );
buf ( n417144 , n380356 );
not ( n94589 , n417144 );
buf ( n417146 , n380368 );
not ( n417147 , n417146 );
buf ( n417148 , n90092 );
not ( n417149 , n417148 );
or ( n94594 , n417147 , n417149 );
buf ( n417151 , n380364 );
buf ( n417152 , n351013 );
nand ( n94597 , n417151 , n417152 );
buf ( n94598 , n94597 );
buf ( n417155 , n94598 );
nand ( n417156 , n94594 , n417155 );
buf ( n417157 , n417156 );
buf ( n417158 , n417157 );
not ( n417159 , n417158 );
or ( n417160 , n94589 , n417159 );
buf ( n417161 , n380364 );
buf ( n417162 , n415989 );
not ( n94607 , n417162 );
buf ( n417164 , n94607 );
buf ( n417165 , n417164 );
and ( n94610 , n417161 , n417165 );
not ( n94611 , n417161 );
buf ( n417168 , n377140 );
and ( n94613 , n94611 , n417168 );
or ( n94614 , n94610 , n94613 );
buf ( n417171 , n94614 );
buf ( n417172 , n417171 );
not ( n94616 , n417172 );
buf ( n417174 , n380398 );
nand ( n417175 , n94616 , n417174 );
buf ( n417176 , n417175 );
buf ( n417177 , n417176 );
nand ( n417178 , n417160 , n417177 );
buf ( n417179 , n417178 );
buf ( n417180 , n417179 );
and ( n417181 , n94587 , n417180 );
and ( n94623 , n417138 , n417142 );
or ( n417183 , n417181 , n94623 );
buf ( n417184 , n417183 );
buf ( n417185 , n417184 );
buf ( n417186 , n417131 );
not ( n417187 , n417186 );
buf ( n417188 , n416776 );
nand ( n417189 , n417187 , n417188 );
buf ( n417190 , n417189 );
buf ( n417191 , n417190 );
nand ( n417192 , n417185 , n417191 );
buf ( n417193 , n417192 );
buf ( n417194 , n417193 );
nand ( n417195 , n417134 , n417194 );
buf ( n417196 , n417195 );
buf ( n417197 , n417196 );
xor ( n94635 , n416796 , n416900 );
xor ( n417199 , n94635 , n416927 );
buf ( n417200 , n417199 );
buf ( n417201 , n417200 );
xor ( n417202 , n416869 , n416874 );
xor ( n94640 , n417202 , n416895 );
buf ( n417204 , n94640 );
buf ( n417205 , n417204 );
buf ( n417206 , n379515 );
buf ( n417207 , n379318 );
and ( n94645 , n417206 , n417207 );
not ( n94646 , n417206 );
buf ( n417210 , n379856 );
and ( n417211 , n94646 , n417210 );
nor ( n417212 , n94645 , n417211 );
buf ( n417213 , n417212 );
buf ( n417214 , n417213 );
not ( n417215 , n417214 );
buf ( n417216 , n416972 );
not ( n417217 , n417216 );
or ( n417218 , n417215 , n417217 );
buf ( n417219 , n417024 );
buf ( n94656 , n58920 );
nand ( n94657 , n417219 , n94656 );
buf ( n94658 , n94657 );
buf ( n417223 , n94658 );
nand ( n417224 , n417218 , n417223 );
buf ( n417225 , n417224 );
buf ( n417226 , n379339 );
buf ( n417227 , C1 );
buf ( n417228 , n417227 );
nand ( n417229 , n417226 , n417228 );
buf ( n417230 , n417229 );
buf ( n417231 , n417230 );
buf ( n417232 , n394835 );
buf ( n417233 , n85590 );
nor ( n417234 , n417232 , n417233 );
buf ( n417235 , n417234 );
buf ( n417236 , n417235 );
not ( n417237 , n417236 );
buf ( n417238 , n384408 );
nand ( n94668 , n417237 , n417238 );
buf ( n417240 , n94668 );
buf ( n417241 , n417240 );
nand ( n417242 , n417231 , n417241 );
buf ( n417243 , n417242 );
buf ( n417244 , n417243 );
buf ( n417245 , n394838 );
buf ( n417246 , n623 );
or ( n417247 , n417245 , n417246 );
buf ( n417248 , n394845 );
nand ( n417249 , n417247 , n417248 );
buf ( n417250 , n417249 );
buf ( n417251 , n417250 );
and ( n94678 , n417244 , n417251 );
buf ( n417253 , n417230 );
buf ( n417254 , n417240 );
nor ( n94681 , n417253 , n417254 );
buf ( n417256 , n94681 );
buf ( n94683 , n417256 );
nor ( n417258 , n94678 , n94683 );
buf ( n417259 , n417258 );
buf ( n417260 , n94507 );
not ( n417261 , n417260 );
buf ( n417262 , n94499 );
not ( n417263 , n417262 );
or ( n417264 , n417261 , n417263 );
buf ( n417265 , n94499 );
buf ( n417266 , n94507 );
or ( n417267 , n417265 , n417266 );
nand ( n94690 , n417264 , n417267 );
buf ( n417269 , n94690 );
not ( n417270 , n417269 );
nand ( n417271 , n417259 , n417270 );
not ( n417272 , n417271 );
buf ( n417273 , n379347 );
buf ( n417274 , n379515 );
nor ( n417275 , n417273 , n417274 );
buf ( n417276 , n417275 );
not ( n94695 , n417276 );
or ( n417278 , n417272 , n94695 );
buf ( n417279 , n417259 );
not ( n417280 , n417279 );
buf ( n417281 , n417280 );
nand ( n417282 , n417269 , n417281 );
nand ( n417283 , n417278 , n417282 );
or ( n417284 , n417225 , n417283 );
buf ( n417285 , n417284 );
xor ( n417286 , n417075 , n417066 );
and ( n417287 , n417050 , n417286 );
not ( n417288 , n417050 );
not ( n417289 , n417286 );
and ( n417290 , n417288 , n417289 );
nor ( n417291 , n417287 , n417290 );
buf ( n417292 , n417291 );
and ( n417293 , n417285 , n417292 );
and ( n417294 , n417225 , n417283 );
buf ( n417295 , n417294 );
nor ( n417296 , n417293 , n417295 );
buf ( n417297 , n417296 );
buf ( n417298 , n417297 );
buf ( n417299 , n379890 );
buf ( n417300 , n378098 );
nand ( n417301 , n417299 , n417300 );
buf ( n417302 , n417301 );
buf ( n417303 , n417302 );
nand ( n417304 , n417298 , n417303 );
buf ( n417305 , n417304 );
not ( n417306 , n417305 );
and ( n417307 , n417083 , n417077 );
not ( n417308 , n417083 );
and ( n417309 , n417308 , n417087 );
or ( n417310 , n417307 , n417309 );
buf ( n417311 , n417310 );
buf ( n417312 , n417030 );
and ( n417313 , n417311 , n417312 );
not ( n417314 , n417311 );
buf ( n417315 , n417033 );
and ( n417316 , n417314 , n417315 );
nor ( n417317 , n417313 , n417316 );
buf ( n417318 , n417317 );
not ( n417319 , n417318 );
or ( n417320 , n417306 , n417319 );
not ( n417321 , n417302 );
buf ( n417322 , n417297 );
not ( n417323 , n417322 );
buf ( n417324 , n417323 );
nand ( n417325 , n417321 , n417324 );
nand ( n417326 , n417320 , n417325 );
buf ( n417327 , n417326 );
xor ( n417328 , n417205 , n417327 );
buf ( n417329 , n380356 );
not ( n417330 , n417329 );
buf ( n417331 , n380368 );
not ( n417332 , n417331 );
buf ( n417333 , n414618 );
not ( n417334 , n417333 );
or ( n417335 , n417332 , n417334 );
buf ( n417336 , n30931 );
buf ( n417337 , n380364 );
nand ( n417338 , n417336 , n417337 );
buf ( n417339 , n417338 );
buf ( n417340 , n417339 );
nand ( n417341 , n417335 , n417340 );
buf ( n417342 , n417341 );
buf ( n417343 , n417342 );
not ( n417344 , n417343 );
or ( n417345 , n417330 , n417344 );
buf ( n417346 , n380368 );
not ( n417347 , n417346 );
buf ( n417348 , n92200 );
not ( n417349 , n417348 );
or ( n417350 , n417347 , n417349 );
buf ( n417351 , n379472 );
buf ( n417352 , n380364 );
nand ( n417353 , n417351 , n417352 );
buf ( n417354 , n417353 );
buf ( n417355 , n417354 );
nand ( n417356 , n417350 , n417355 );
buf ( n417357 , n417356 );
buf ( n417358 , n417357 );
buf ( n417359 , n380398 );
nand ( n417360 , n417358 , n417359 );
buf ( n417361 , n417360 );
buf ( n417362 , n417361 );
nand ( n417363 , n417345 , n417362 );
buf ( n417364 , n417363 );
buf ( n417365 , n417364 );
and ( n417366 , n417328 , n417365 );
and ( n417367 , n417205 , n417327 );
or ( n417368 , n417366 , n417367 );
buf ( n417369 , n417368 );
buf ( n417370 , n417369 );
xor ( n417371 , n417201 , n417370 );
buf ( n417372 , n94535 );
not ( n417373 , n94378 );
not ( n417374 , n94400 );
or ( n417375 , n417373 , n417374 );
or ( n417376 , n94378 , n94400 );
nand ( n417377 , n417375 , n417376 );
buf ( n417378 , n417377 );
xnor ( n417379 , n417372 , n417378 );
buf ( n417380 , n417379 );
buf ( n417381 , n417380 );
and ( n417382 , n417371 , n417381 );
and ( n417383 , n417201 , n417370 );
or ( n417384 , n417382 , n417383 );
buf ( n417385 , n417384 );
buf ( n417386 , n417385 );
xor ( n417387 , n417138 , n417142 );
xor ( n417388 , n417387 , n417180 );
buf ( n417389 , n417388 );
buf ( n94698 , n417389 );
xor ( n94699 , n417386 , n94698 );
not ( n417392 , n417342 );
not ( n417393 , n380398 );
or ( n417394 , n417392 , n417393 );
or ( n417395 , n417171 , n384940 );
nand ( n417396 , n417394 , n417395 );
buf ( n417397 , n417396 );
buf ( n417398 , n417302 );
buf ( n417399 , n417324 );
xor ( n94706 , n417398 , n417399 );
buf ( n417401 , n417318 );
xor ( n94708 , n94706 , n417401 );
buf ( n94709 , n94708 );
buf ( n94710 , n94709 );
buf ( n417405 , n417357 );
buf ( n417406 , n380356 );
and ( n94713 , n417405 , n417406 );
not ( n417408 , n380398 );
buf ( n417409 , n380364 );
buf ( n417410 , n378840 );
and ( n417411 , n417409 , n417410 );
not ( n417412 , n417409 );
buf ( n417413 , n415592 );
and ( n94720 , n417412 , n417413 );
nor ( n417415 , n417411 , n94720 );
buf ( n417416 , n417415 );
nor ( n417417 , n417408 , n417416 );
buf ( n417418 , n417417 );
nor ( n94725 , n94713 , n417418 );
buf ( n94726 , n94725 );
buf ( n417421 , n94726 );
or ( n417422 , n94710 , n417421 );
buf ( n417423 , n417422 );
buf ( n417424 , n417423 );
buf ( n417425 , n94709 );
buf ( n417426 , n94726 );
nand ( n417427 , n417425 , n417426 );
buf ( n417428 , n417427 );
buf ( n417429 , n417428 );
buf ( n417430 , n417225 );
not ( n417431 , n417291 );
and ( n417432 , n417283 , n417431 );
not ( n417433 , n417283 );
and ( n417434 , n417433 , n417291 );
nor ( n417435 , n417432 , n417434 );
buf ( n417436 , n417435 );
xnor ( n417437 , n417430 , n417436 );
buf ( n417438 , n417437 );
buf ( n417439 , n417438 );
buf ( n417440 , n380398 );
not ( n417441 , n417440 );
buf ( n417442 , n380361 );
buf ( n417443 , n377091 );
xor ( n417444 , n417442 , n417443 );
buf ( n417445 , n417444 );
buf ( n417446 , n417445 );
not ( n417447 , n417446 );
buf ( n417448 , n417447 );
buf ( n417449 , n417448 );
not ( n417450 , n417449 );
or ( n417451 , n417441 , n417450 );
buf ( n417452 , n380361 );
buf ( n417453 , n377065 );
and ( n417454 , n417452 , n417453 );
not ( n417455 , n417452 );
buf ( n417456 , n415121 );
and ( n417457 , n417455 , n417456 );
nor ( n417458 , n417454 , n417457 );
buf ( n417459 , n417458 );
buf ( n417460 , n417459 );
buf ( n417461 , n384940 );
or ( n417462 , n417460 , n417461 );
nand ( n417463 , n417451 , n417462 );
buf ( n417464 , n417463 );
buf ( n417465 , n417464 );
buf ( n417466 , C0 );
buf ( n417467 , n417466 );
buf ( n417468 , n417240 );
not ( n417469 , n417468 );
buf ( n417470 , n417250 );
not ( n417471 , n417470 );
or ( n417472 , n417469 , n417471 );
buf ( n417473 , n417250 );
buf ( n417474 , n417240 );
or ( n417475 , n417473 , n417474 );
nand ( n417476 , n417472 , n417475 );
buf ( n417477 , n417476 );
buf ( n417478 , n417477 );
not ( n417479 , n417478 );
buf ( n417480 , n417230 );
not ( n417481 , n417480 );
or ( n417482 , n417479 , n417481 );
buf ( n417483 , n417477 );
buf ( n417484 , n417230 );
or ( n417485 , n417483 , n417484 );
nand ( n417486 , n417482 , n417485 );
buf ( n417487 , n417486 );
buf ( n417488 , n417487 );
xor ( n417489 , n417467 , n417488 );
buf ( n417490 , n380398 );
not ( n417491 , n417490 );
buf ( n417492 , n379515 );
not ( n417493 , n417492 );
or ( n417494 , n417491 , n417493 );
buf ( n417495 , n417445 );
buf ( n417496 , n384940 );
or ( n417497 , n417495 , n417496 );
nand ( n417498 , n417494 , n417497 );
buf ( n417499 , n417498 );
buf ( n417500 , n417499 );
and ( n94732 , n417489 , n417500 );
or ( n417502 , n94732 , C0 );
buf ( n417503 , n417502 );
buf ( n417504 , n417503 );
xor ( n417505 , n417465 , n417504 );
not ( n94737 , n417282 );
nand ( n94738 , n94737 , n417276 );
not ( n417508 , n417271 );
nand ( n417509 , n417508 , n417276 );
not ( n417510 , n417276 );
nor ( n417511 , n417259 , n417269 );
nand ( n417512 , n417510 , n417511 );
nor ( n417513 , n417281 , n417270 );
nand ( n417514 , n417510 , n417513 );
nand ( n417515 , n94738 , n417509 , n417512 , n417514 );
buf ( n417516 , n417515 );
and ( n417517 , n417505 , n417516 );
and ( n417518 , n417465 , n417504 );
or ( n417519 , n417517 , n417518 );
buf ( n417520 , n417519 );
buf ( n94740 , n417520 );
xor ( n94741 , n417439 , n94740 );
buf ( n417523 , n417416 );
buf ( n417524 , n384940 );
or ( n417525 , n417523 , n417524 );
buf ( n417526 , n417459 );
not ( n417527 , n417526 );
buf ( n417528 , n380398 );
nand ( n417529 , n417527 , n417528 );
buf ( n417530 , n417529 );
buf ( n94750 , n417530 );
nand ( n94751 , n417525 , n94750 );
buf ( n417533 , n94751 );
buf ( n417534 , n417533 );
and ( n94754 , n94741 , n417534 );
and ( n417536 , n417439 , n94740 );
or ( n417537 , n94754 , n417536 );
buf ( n417538 , n417537 );
buf ( n417539 , n417538 );
nand ( n417540 , n417429 , n417539 );
buf ( n417541 , n417540 );
buf ( n417542 , n417541 );
nand ( n94762 , n417424 , n417542 );
buf ( n94763 , n94762 );
buf ( n417545 , n94763 );
not ( n417546 , n417545 );
buf ( n417547 , n417546 );
buf ( n417548 , n417547 );
xor ( n94768 , n417205 , n417327 );
xor ( n94769 , n94768 , n417365 );
buf ( n417551 , n94769 );
buf ( n417552 , n417551 );
buf ( n417553 , n417008 );
buf ( n417554 , n416987 );
xor ( n417555 , n417553 , n417554 );
buf ( n417556 , n417555 );
buf ( n417557 , n417556 );
buf ( n417558 , n94533 );
xnor ( n94774 , n417557 , n417558 );
buf ( n417560 , n94774 );
buf ( n417561 , n417560 );
nor ( n94777 , n417552 , n417561 );
buf ( n417563 , n94777 );
buf ( n417564 , n417563 );
or ( n94780 , n417548 , n417564 );
buf ( n417566 , n417551 );
buf ( n417567 , n417560 );
nand ( n94783 , n417566 , n417567 );
buf ( n417569 , n94783 );
buf ( n417570 , n417569 );
nand ( n94786 , n94780 , n417570 );
buf ( n417572 , n94786 );
buf ( n417573 , n417572 );
xor ( n94789 , n417397 , n417573 );
xor ( n94790 , n417201 , n417370 );
xor ( n94791 , n94790 , n417381 );
buf ( n417577 , n94791 );
buf ( n417578 , n417577 );
and ( n94794 , n94789 , n417578 );
and ( n94795 , n417397 , n417573 );
or ( n94796 , n94794 , n94795 );
buf ( n417582 , n94796 );
buf ( n417583 , n417582 );
and ( n94799 , n94699 , n417583 );
and ( n94800 , n417386 , n94698 );
or ( n94801 , n94799 , n94800 );
buf ( n417587 , n94801 );
not ( n94803 , n417587 );
buf ( n417589 , n416776 );
not ( n94805 , n417589 );
buf ( n417591 , n417131 );
not ( n94807 , n417591 );
or ( n94808 , n94805 , n94807 );
buf ( n417594 , n416776 );
buf ( n417595 , n417131 );
or ( n94811 , n417594 , n417595 );
nand ( n94812 , n94808 , n94811 );
buf ( n417598 , n94812 );
not ( n94814 , n417598 );
nand ( n94815 , n94814 , n417184 );
not ( n94816 , n417184 );
nand ( n94817 , n94816 , n417598 );
buf ( n417603 , n380368 );
not ( n94819 , n417603 );
buf ( n417605 , n377776 );
not ( n94821 , n417605 );
or ( n94822 , n94819 , n94821 );
buf ( n417608 , n412279 );
buf ( n417609 , n380364 );
nand ( n94825 , n417608 , n417609 );
buf ( n417611 , n94825 );
buf ( n417612 , n417611 );
nand ( n94828 , n94822 , n417612 );
buf ( n417614 , n94828 );
buf ( n417615 , n417614 );
buf ( n417616 , n380356 );
and ( n94831 , n417615 , n417616 );
buf ( n417618 , n417157 );
not ( n417619 , n417618 );
buf ( n417620 , n93364 );
nor ( n94833 , n417619 , n417620 );
buf ( n417622 , n94833 );
buf ( n417623 , n417622 );
nor ( n417624 , n94831 , n417623 );
buf ( n417625 , n417624 );
nand ( n417626 , n94815 , n94817 , n417625 );
not ( n94835 , n417626 );
or ( n94836 , n94803 , n94835 );
not ( n94837 , n417625 );
not ( n94838 , n417184 );
nand ( n94839 , n94838 , n94814 );
nand ( n94840 , n417184 , n417598 );
nand ( n94841 , n94837 , n94839 , n94840 );
nand ( n94842 , n94836 , n94841 );
buf ( n417635 , n94842 );
xor ( n94844 , n417197 , n417635 );
xor ( n94845 , n416584 , n416606 );
xor ( n94846 , n94845 , n416704 );
buf ( n417639 , n94846 );
buf ( n417640 , n417639 );
buf ( n417641 , n380356 );
not ( n417642 , n417641 );
buf ( n417643 , n380368 );
not ( n94850 , n417643 );
buf ( n417645 , n377349 );
not ( n417646 , n417645 );
or ( n94852 , n94850 , n417646 );
buf ( n417648 , n409020 );
buf ( n417649 , n380364 );
nand ( n94855 , n417648 , n417649 );
buf ( n417651 , n94855 );
buf ( n417652 , n417651 );
nand ( n94858 , n94852 , n417652 );
buf ( n417654 , n94858 );
buf ( n417655 , n417654 );
not ( n94861 , n417655 );
or ( n94862 , n417642 , n94861 );
buf ( n417658 , n417614 );
buf ( n417659 , n380401 );
nand ( n94865 , n417658 , n417659 );
buf ( n417661 , n94865 );
buf ( n417662 , n417661 );
nand ( n94868 , n94862 , n417662 );
buf ( n417664 , n94868 );
buf ( n417665 , n417664 );
xor ( n94871 , n417640 , n417665 );
buf ( n417667 , n58923 );
not ( n94873 , n417667 );
buf ( n417669 , n416367 );
not ( n94875 , n417669 );
or ( n94876 , n94873 , n94875 );
buf ( n417672 , n416613 );
buf ( n417673 , n414059 );
nand ( n94879 , n417672 , n417673 );
buf ( n417675 , n94879 );
buf ( n417676 , n417675 );
nand ( n94882 , n94876 , n417676 );
buf ( n417678 , n94882 );
buf ( n417679 , n417678 );
xor ( n94885 , n416785 , n416790 );
and ( n94886 , n94885 , n417129 );
and ( n94887 , n416785 , n416790 );
or ( n94888 , n94886 , n94887 );
buf ( n417684 , n94888 );
buf ( n417685 , n417684 );
xor ( n94891 , n417679 , n417685 );
xor ( n94892 , n93501 , n416061 );
xor ( n94893 , n94892 , n416078 );
buf ( n417689 , n94893 );
buf ( n417690 , n417689 );
xor ( n94896 , n94891 , n417690 );
buf ( n417692 , n94896 );
buf ( n417693 , n417692 );
xor ( n94899 , n94871 , n417693 );
buf ( n417695 , n94899 );
buf ( n417696 , n417695 );
and ( n94900 , n94844 , n417696 );
and ( n94901 , n417197 , n417635 );
or ( n94902 , n94900 , n94901 );
buf ( n417700 , n94902 );
not ( n94903 , n417700 );
xor ( n94904 , n417679 , n417685 );
and ( n94905 , n94904 , n417690 );
and ( n94906 , n417679 , n417685 );
or ( n94907 , n94905 , n94906 );
buf ( n417706 , n94907 );
buf ( n417707 , n380356 );
not ( n94910 , n417707 );
buf ( n417709 , n416741 );
not ( n94912 , n417709 );
or ( n94913 , n94910 , n94912 );
buf ( n417712 , n417654 );
buf ( n417713 , n380401 );
nand ( n94916 , n417712 , n417713 );
buf ( n417715 , n94916 );
buf ( n417716 , n417715 );
nand ( n94918 , n94913 , n417716 );
buf ( n417718 , n94918 );
buf ( n417719 , n417718 );
not ( n94921 , n417719 );
buf ( n417721 , n94921 );
and ( n94923 , n417706 , n417721 );
not ( n94924 , n417706 );
and ( n94925 , n94924 , n417718 );
or ( n94926 , n94923 , n94925 );
buf ( n417726 , n94926 );
xor ( n94928 , n416709 , n416712 );
xor ( n94929 , n94928 , n416717 );
buf ( n417729 , n94929 );
buf ( n417730 , n417729 );
not ( n94932 , n417730 );
buf ( n417732 , n94932 );
buf ( n417733 , n417732 );
and ( n94935 , n417726 , n417733 );
not ( n94936 , n417726 );
buf ( n417736 , n417729 );
and ( n94938 , n94936 , n417736 );
nor ( n94939 , n94935 , n94938 );
buf ( n417739 , n94939 );
buf ( n417740 , n417739 );
buf ( n417741 , n417664 );
buf ( n417742 , n417639 );
or ( n417743 , n417741 , n417742 );
buf ( n417744 , n417692 );
nand ( n417745 , n417743 , n417744 );
buf ( n417746 , n417745 );
buf ( n417747 , n417746 );
buf ( n417748 , n417664 );
buf ( n417749 , n417639 );
nand ( n94948 , n417748 , n417749 );
buf ( n94949 , n94948 );
buf ( n417752 , n94949 );
and ( n94951 , n417747 , n417752 );
buf ( n417754 , n94951 );
buf ( n417755 , n417754 );
nand ( n417756 , n417740 , n417755 );
buf ( n417757 , n417756 );
not ( n94956 , n417757 );
or ( n94957 , n94903 , n94956 );
buf ( n417760 , n417739 );
buf ( n417761 , n417754 );
or ( n417762 , n417760 , n417761 );
buf ( n417763 , n417762 );
nand ( n94962 , n94957 , n417763 );
buf ( n417765 , n94962 );
not ( n94964 , n417765 );
buf ( n417767 , n94964 );
buf ( n417768 , n417767 );
buf ( n417769 , n416754 );
not ( n94968 , n417769 );
buf ( n417771 , n416721 );
not ( n94970 , n417771 );
buf ( n417773 , n94192 );
not ( n94972 , n417773 );
and ( n94973 , n94970 , n94972 );
buf ( n417776 , n94192 );
buf ( n417777 , n416721 );
and ( n94976 , n417776 , n417777 );
nor ( n417779 , n94973 , n94976 );
buf ( n417780 , n417779 );
buf ( n417781 , n417780 );
not ( n94980 , n417781 );
or ( n417783 , n94968 , n94980 );
buf ( n417784 , n416754 );
buf ( n417785 , n417780 );
or ( n94984 , n417784 , n417785 );
nand ( n94985 , n417783 , n94984 );
buf ( n417788 , n94985 );
buf ( n417789 , n417788 );
buf ( n417790 , n417721 );
not ( n94989 , n417790 );
buf ( n417792 , n417732 );
not ( n417793 , n417792 );
or ( n94992 , n94989 , n417793 );
buf ( n417795 , n417706 );
nand ( n94994 , n94992 , n417795 );
buf ( n417797 , n94994 );
buf ( n417798 , n417797 );
buf ( n417799 , n417729 );
buf ( n417800 , n417718 );
nand ( n94999 , n417799 , n417800 );
buf ( n417802 , n94999 );
buf ( n417803 , n417802 );
nand ( n417804 , n417798 , n417803 );
buf ( n417805 , n417804 );
buf ( n417806 , n417805 );
nor ( n95005 , n417789 , n417806 );
buf ( n417808 , n95005 );
buf ( n417809 , n417808 );
or ( n95008 , n417768 , n417809 );
buf ( n417811 , n417788 );
buf ( n417812 , n417805 );
nand ( n95011 , n417811 , n417812 );
buf ( n417814 , n95011 );
buf ( n417815 , n417814 );
nand ( n95014 , n95008 , n417815 );
buf ( n417817 , n95014 );
not ( n95016 , n417817 );
or ( n95017 , n416770 , n95016 );
or ( n95018 , n416411 , n94210 );
nand ( n95019 , n95017 , n95018 );
not ( n417822 , n95019 );
xnor ( n417823 , n416277 , n416283 );
buf ( n417824 , n417823 );
buf ( n417825 , n416294 );
and ( n95023 , n417824 , n417825 );
not ( n95024 , n417824 );
buf ( n417828 , n416297 );
and ( n95026 , n95024 , n417828 );
nor ( n95027 , n95023 , n95026 );
buf ( n417831 , n95027 );
buf ( n417832 , n417831 );
buf ( n417833 , n416398 );
not ( n95031 , n417833 );
buf ( n417835 , n416318 );
not ( n95033 , n417835 );
or ( n95034 , n95031 , n95033 );
buf ( n417838 , n416392 );
nand ( n95036 , n95034 , n417838 );
buf ( n417840 , n95036 );
buf ( n417841 , n417840 );
buf ( n417842 , n416318 );
not ( n95038 , n417842 );
buf ( n417844 , n93839 );
nand ( n95040 , n95038 , n417844 );
buf ( n417846 , n95040 );
buf ( n417847 , n417846 );
and ( n95043 , n417841 , n417847 );
buf ( n417849 , n95043 );
buf ( n417850 , n417849 );
nand ( n95046 , n417832 , n417850 );
buf ( n417852 , n95046 );
not ( n95048 , n417852 );
or ( n95049 , n417822 , n95048 );
buf ( n417855 , n417831 );
buf ( n417856 , n417849 );
or ( n95051 , n417855 , n417856 );
buf ( n417858 , n95051 );
nand ( n95053 , n95049 , n417858 );
not ( n95054 , n95053 );
or ( n417861 , n416312 , n95054 );
buf ( n417862 , n416308 );
not ( n417863 , n417862 );
buf ( n417864 , n416303 );
nand ( n417865 , n417863 , n417864 );
buf ( n417866 , n417865 );
nand ( n417867 , n417861 , n417866 );
buf ( n417868 , n417867 );
nand ( n417869 , n416166 , n417868 );
buf ( n417870 , n417869 );
buf ( n417871 , n417870 );
buf ( n417872 , n416163 );
buf ( n417873 , n416158 );
or ( n417874 , n417872 , n417873 );
buf ( n417875 , n417874 );
buf ( n417876 , n417875 );
nand ( n417877 , n417871 , n417876 );
buf ( n417878 , n417877 );
not ( n417879 , n417878 );
or ( n417880 , n93390 , n417879 );
buf ( n417881 , n415823 );
buf ( n417882 , n415942 );
or ( n417883 , n417881 , n417882 );
buf ( n417884 , n417883 );
nand ( n417885 , n417880 , n417884 );
buf ( n417886 , n417885 );
nand ( n417887 , n93264 , n417886 );
buf ( n417888 , n417887 );
buf ( n417889 , n417888 );
buf ( n417890 , n415817 );
buf ( n417891 , n93182 );
or ( n417892 , n417890 , n417891 );
buf ( n417893 , n417892 );
buf ( n417894 , n417893 );
nand ( n417895 , n417889 , n417894 );
buf ( n417896 , n417895 );
buf ( n417897 , n417896 );
not ( n417898 , n417897 );
buf ( n417899 , n417898 );
buf ( n417900 , n417899 );
xor ( n417901 , n415787 , n415791 );
and ( n417902 , n417901 , n415805 );
and ( n417903 , n415787 , n415791 );
or ( n417904 , n417902 , n417903 );
buf ( n417905 , n417904 );
buf ( n417906 , n417905 );
buf ( n417907 , n414081 );
not ( n417908 , n417907 );
buf ( n417909 , n414110 );
not ( n417910 , n417909 );
or ( n417911 , n417908 , n417910 );
buf ( n417912 , n414078 );
buf ( n417913 , n414107 );
nand ( n417914 , n417912 , n417913 );
buf ( n417915 , n417914 );
buf ( n417916 , n417915 );
nand ( n417917 , n417911 , n417916 );
buf ( n417918 , n417917 );
buf ( n417919 , n417918 );
buf ( n417920 , n414070 );
buf ( n417921 , n417920 );
buf ( n417922 , n417921 );
buf ( n417923 , n417922 );
xor ( n417924 , n417919 , n417923 );
buf ( n417925 , n417924 );
buf ( n417926 , n417925 );
xor ( n417927 , n417906 , n417926 );
buf ( n417928 , n414196 );
buf ( n417929 , n414213 );
xor ( n417930 , n417928 , n417929 );
buf ( n417931 , n92503 );
xor ( n417932 , n417930 , n417931 );
buf ( n417933 , n417932 );
buf ( n417934 , n417933 );
xor ( n417935 , n417927 , n417934 );
buf ( n417936 , n417935 );
buf ( n417937 , n417936 );
buf ( n417938 , n93193 );
not ( n417939 , n417938 );
buf ( n417940 , n417939 );
buf ( n417941 , n417940 );
not ( n417942 , n417941 );
buf ( n417943 , n415810 );
not ( n417944 , n417943 );
or ( n417945 , n417942 , n417944 );
buf ( n417946 , n415771 );
not ( n417947 , n417946 );
buf ( n417948 , n417947 );
buf ( n417949 , n417948 );
nand ( n417950 , n417945 , n417949 );
buf ( n417951 , n417950 );
buf ( n417952 , n417951 );
buf ( n417953 , n415810 );
buf ( n417954 , n417940 );
or ( n417955 , n417953 , n417954 );
buf ( n417956 , n417955 );
buf ( n417957 , n417956 );
nand ( n417958 , n417952 , n417957 );
buf ( n417959 , n417958 );
buf ( n417960 , n417959 );
nor ( n417961 , n417937 , n417960 );
buf ( n417962 , n417961 );
buf ( n417963 , n417962 );
or ( n417964 , n417900 , n417963 );
buf ( n417965 , n417936 );
buf ( n417966 , n417959 );
nand ( n417967 , n417965 , n417966 );
buf ( n417968 , n417967 );
buf ( n417969 , n417968 );
nand ( n417970 , n417964 , n417969 );
buf ( n417971 , n417970 );
buf ( n417972 , n417971 );
xor ( n417973 , n417906 , n417926 );
and ( n417974 , n417973 , n417934 );
and ( n417975 , n417906 , n417926 );
or ( n417976 , n417974 , n417975 );
buf ( n417977 , n417976 );
not ( n417978 , n417977 );
xor ( n417979 , n91642 , n415067 );
and ( n417980 , n417979 , n414182 );
not ( n417981 , n417979 );
not ( n417982 , n414182 );
and ( n417983 , n417981 , n417982 );
nor ( n417984 , n417980 , n417983 );
nand ( n417985 , n417978 , n417984 );
buf ( n417986 , n417985 );
nand ( n417987 , n417972 , n417986 );
buf ( n417988 , n417987 );
buf ( n417989 , n417988 );
not ( n417990 , n417984 );
nand ( n417991 , n417990 , n417977 );
buf ( n417992 , n417991 );
nand ( n417993 , n417989 , n417992 );
buf ( n417994 , n417993 );
not ( n417995 , n417994 );
or ( n417996 , n415080 , n417995 );
buf ( n417997 , n92520 );
not ( n417998 , n417997 );
buf ( n417999 , n92515 );
nand ( n418000 , n417998 , n417999 );
buf ( n418001 , n418000 );
nand ( n418002 , n417996 , n418001 );
not ( n418003 , n418002 );
or ( n418004 , n414164 , n418003 );
not ( n418005 , n414162 );
nand ( n418006 , n418005 , n414149 );
nand ( n418007 , n418004 , n418006 );
buf ( n418008 , n418007 );
not ( n418009 , n418008 );
or ( n418010 , n413900 , n418009 );
buf ( n418011 , n413895 );
not ( n418012 , n418011 );
buf ( n418013 , n413883 );
nand ( n418014 , n418012 , n418013 );
buf ( n418015 , n418014 );
buf ( n418016 , n418015 );
nand ( n418017 , n418010 , n418016 );
buf ( n418018 , n418017 );
buf ( n418019 , n418018 );
and ( n418020 , n413612 , n418019 );
and ( n418021 , n413607 , n413611 );
or ( n418022 , n418020 , n418021 );
buf ( n418023 , n418022 );
buf ( n418024 , n418023 );
and ( n418025 , n90791 , n418024 );
and ( n418026 , n413327 , n413331 );
or ( n418027 , n418025 , n418026 );
buf ( n418028 , n418027 );
buf ( n418029 , n418028 );
and ( n418030 , n90539 , n418029 );
and ( n418031 , n413075 , n413079 );
or ( n418032 , n418030 , n418031 );
buf ( n418033 , n418032 );
buf ( n418034 , n418033 );
buf ( n418035 , n89919 );
buf ( n418036 , n411726 );
buf ( n418037 , n412428 );
or ( n418038 , n418036 , n418037 );
buf ( n418039 , n418038 );
buf ( n418040 , n418039 );
and ( n418041 , n418034 , n418035 , n418040 );
buf ( n418042 , n418041 );
buf ( n418043 , n418042 );
buf ( n418044 , n411278 );
nand ( n418045 , n418043 , n418044 );
buf ( n418046 , n418045 );
buf ( n418047 , n418046 );
nand ( n418048 , n412462 , n418047 );
buf ( n418049 , n418048 );
buf ( n418050 , n410790 );
buf ( n418051 , n410822 );
or ( n418052 , n418050 , n418051 );
buf ( n418053 , n418052 );
nand ( n418054 , n418049 , n418053 );
not ( n418055 , n418054 );
or ( n418056 , n88304 , n418055 );
xor ( n418057 , n407293 , n407318 );
and ( n418058 , n418057 , n407508 );
and ( n418059 , n407293 , n407318 );
or ( n418060 , n418058 , n418059 );
buf ( n418061 , n418060 );
buf ( n418062 , n418061 );
buf ( n418063 , n379890 );
not ( n418064 , n418063 );
buf ( n418065 , n83643 );
not ( n418066 , n418065 );
or ( n418067 , n418064 , n418066 );
buf ( n418068 , n83731 );
buf ( n418069 , n379916 );
nand ( n418070 , n418068 , n418069 );
buf ( n418071 , n418070 );
buf ( n418072 , n418071 );
nand ( n418073 , n418067 , n418072 );
buf ( n418074 , n418073 );
buf ( n418075 , n407457 );
not ( n418076 , n418075 );
buf ( n418077 , n407354 );
not ( n418078 , n418077 );
or ( n418079 , n418076 , n418078 );
buf ( n418080 , n407497 );
nand ( n418081 , n418079 , n418080 );
buf ( n418082 , n418081 );
buf ( n418083 , n407354 );
not ( n418084 , n418083 );
buf ( n418085 , n407454 );
nand ( n418086 , n418084 , n418085 );
buf ( n418087 , n418086 );
nand ( n418088 , n418082 , n418087 );
xor ( n418089 , n418074 , n418088 );
buf ( n418090 , n405008 );
buf ( n418091 , n405019 );
xor ( n418092 , n418090 , n418091 );
buf ( n418093 , n83237 );
xor ( n418094 , n418092 , n418093 );
buf ( n418095 , n418094 );
xnor ( n418096 , n418089 , n418095 );
buf ( n418097 , n418096 );
xor ( n418098 , n418062 , n418097 );
xor ( n418099 , n409159 , n409304 );
and ( n418100 , n418099 , n409376 );
and ( n418101 , n409159 , n409304 );
or ( n418102 , n418100 , n418101 );
buf ( n418103 , n418102 );
buf ( n418104 , n418103 );
xor ( n418105 , n418098 , n418104 );
buf ( n418106 , n418105 );
buf ( n418107 , n418106 );
xor ( n418108 , n409153 , n409379 );
and ( n418109 , n418108 , n409467 );
and ( n418110 , n409153 , n409379 );
or ( n418111 , n418109 , n418110 );
buf ( n418112 , n418111 );
buf ( n418113 , n418112 );
xor ( n418114 , n418107 , n418113 );
buf ( n418115 , n380356 );
not ( n418116 , n418115 );
buf ( n418117 , n380368 );
not ( n418118 , n418117 );
buf ( n418119 , n366077 );
not ( n418120 , n418119 );
or ( n418121 , n418118 , n418120 );
buf ( n418122 , n366078 );
buf ( n418123 , n384667 );
nand ( n418124 , n418122 , n418123 );
buf ( n418125 , n418124 );
buf ( n418126 , n418125 );
nand ( n418127 , n418121 , n418126 );
buf ( n418128 , n418127 );
buf ( n418129 , n418128 );
not ( n418130 , n418129 );
or ( n418131 , n418116 , n418130 );
buf ( n418132 , n407310 );
buf ( n418133 , n380404 );
nand ( n418134 , n418132 , n418133 );
buf ( n418135 , n418134 );
buf ( n418136 , n418135 );
nand ( n418137 , n418131 , n418136 );
buf ( n418138 , n418137 );
buf ( n418139 , n418138 );
buf ( n418140 , n405207 );
buf ( n418141 , n409320 );
or ( n418142 , n418140 , n418141 );
buf ( n418143 , n405217 );
buf ( n418144 , n398693 );
or ( n418145 , n418143 , n418144 );
nand ( n418146 , n418142 , n418145 );
buf ( n418147 , n418146 );
buf ( n418148 , n418147 );
xor ( n418149 , n409343 , n409356 );
and ( n418150 , n418149 , n409363 );
and ( n418151 , n409343 , n409356 );
or ( n418152 , n418150 , n418151 );
buf ( n418153 , n418152 );
buf ( n418154 , n418153 );
xor ( n418155 , n418148 , n418154 );
xor ( n418156 , n407469 , n407482 );
and ( n418157 , n418156 , n407495 );
and ( n418158 , n407469 , n407482 );
or ( n418159 , n418157 , n418158 );
buf ( n418160 , n418159 );
buf ( n418161 , n418160 );
xor ( n418162 , n418155 , n418161 );
buf ( n418163 , n418162 );
buf ( n418164 , n418163 );
xor ( n418165 , n418139 , n418164 );
xor ( n418166 , n86816 , n409366 );
and ( n418167 , n418166 , n409373 );
and ( n418168 , n86816 , n409366 );
or ( n418169 , n418167 , n418168 );
buf ( n418170 , n418169 );
buf ( n418171 , n418170 );
xor ( n418172 , n418165 , n418171 );
buf ( n418173 , n418172 );
buf ( n418174 , n418173 );
buf ( n418175 , n407510 );
buf ( n418176 , n407185 );
or ( n418177 , n418175 , n418176 );
buf ( n418178 , n407247 );
nand ( n418179 , n418177 , n418178 );
buf ( n418180 , n418179 );
buf ( n418181 , n418180 );
buf ( n418182 , n407510 );
buf ( n418183 , n407185 );
nand ( n418184 , n418182 , n418183 );
buf ( n418185 , n418184 );
buf ( n418186 , n418185 );
nand ( n418187 , n418181 , n418186 );
buf ( n418188 , n418187 );
buf ( n418189 , n418188 );
xor ( n418190 , n418174 , n418189 );
xnor ( n418191 , n405259 , n405273 );
xor ( n418192 , n405406 , n418191 );
buf ( n418193 , n418192 );
buf ( n418194 , n379263 );
not ( n418195 , n418194 );
buf ( n418196 , n404697 );
not ( n418197 , n418196 );
or ( n418198 , n418195 , n418197 );
buf ( n418199 , n407331 );
buf ( n418200 , n379299 );
nand ( n418201 , n418199 , n418200 );
buf ( n418202 , n418201 );
buf ( n418203 , n418202 );
nand ( n418204 , n418198 , n418203 );
buf ( n418205 , n418204 );
buf ( n418206 , n418205 );
xor ( n418207 , n418193 , n418206 );
xor ( n418208 , n407280 , n84953 );
and ( n418209 , n418208 , n407290 );
and ( n418210 , n407280 , n84953 );
or ( n418211 , n418209 , n418210 );
buf ( n418212 , n418211 );
buf ( n418213 , n418212 );
xor ( n418214 , n418207 , n418213 );
buf ( n418215 , n418214 );
buf ( n418216 , n418215 );
xor ( n418217 , n405719 , n407145 );
and ( n418218 , n418217 , n407183 );
and ( n418219 , n405719 , n407145 );
or ( n418220 , n418218 , n418219 );
buf ( n418221 , n418220 );
buf ( n418222 , n418221 );
xor ( n418223 , n418216 , n418222 );
xor ( n418224 , n404713 , n404750 );
xor ( n418225 , n418224 , n404768 );
buf ( n418226 , n418225 );
buf ( n418227 , n418226 );
buf ( n418228 , n58923 );
not ( n418229 , n418228 );
buf ( n418230 , n405610 );
not ( n418231 , n418230 );
or ( n418232 , n418229 , n418231 );
buf ( n418233 , n407175 );
buf ( n418234 , n58867 );
nand ( n418235 , n418233 , n418234 );
buf ( n418236 , n418235 );
buf ( n418237 , n418236 );
nand ( n418238 , n418232 , n418237 );
buf ( n418239 , n418238 );
buf ( n418240 , n418239 );
xor ( n418241 , n418227 , n418240 );
buf ( n418242 , n42266 );
buf ( n418243 , n379515 );
buf ( n418244 , n362426 );
and ( n418245 , n418243 , n418244 );
not ( n418246 , n418243 );
buf ( n418247 , n365773 );
and ( n418248 , n418246 , n418247 );
nor ( n418249 , n418245 , n418248 );
buf ( n418250 , n418249 );
buf ( n418251 , n418250 );
or ( n418252 , n418242 , n418251 );
buf ( n418253 , n405121 );
buf ( n418254 , n362388 );
or ( n418255 , n418253 , n418254 );
nand ( n418256 , n418252 , n418255 );
buf ( n418257 , n418256 );
buf ( n418258 , n418257 );
xor ( n418259 , n418241 , n418258 );
buf ( n418260 , n418259 );
buf ( n418261 , n418260 );
xor ( n418262 , n418223 , n418261 );
buf ( n418263 , n418262 );
buf ( n418264 , n418263 );
xor ( n418265 , n418190 , n418264 );
buf ( n418266 , n418265 );
buf ( n418267 , n418266 );
xor ( n418268 , n418114 , n418267 );
buf ( n418269 , n418268 );
buf ( n418270 , n418269 );
xor ( n418271 , n407512 , n409146 );
and ( n418272 , n418271 , n409470 );
and ( n418273 , n407512 , n409146 );
or ( n418274 , n418272 , n418273 );
buf ( n418275 , n418274 );
buf ( n418276 , n418275 );
nor ( n418277 , n418270 , n418276 );
buf ( n418278 , n418277 );
buf ( n418279 , n409472 );
buf ( n418280 , n410784 );
nor ( n418281 , n418279 , n418280 );
buf ( n418282 , n418281 );
nor ( n418283 , n418278 , n418282 );
nand ( n418284 , n418056 , n418283 );
buf ( n418285 , n418284 );
buf ( n418286 , n418269 );
buf ( n418287 , n418275 );
nand ( n418288 , n418286 , n418287 );
buf ( n418289 , n418288 );
buf ( n418290 , n418289 );
nand ( n418291 , n418285 , n418290 );
buf ( n418292 , n418291 );
buf ( n418293 , n418292 );
xor ( n418294 , n404672 , n404777 );
xnor ( n418295 , n418294 , n404675 );
xnor ( n418296 , n404816 , n404845 );
xnor ( n418297 , n418296 , n405130 );
xor ( n418298 , n418295 , n418297 );
buf ( n418299 , n418298 );
not ( n418300 , n418074 );
not ( n418301 , n418088 );
or ( n418302 , n418300 , n418301 );
buf ( n418303 , n418088 );
buf ( n418304 , n418074 );
nor ( n418305 , n418303 , n418304 );
buf ( n418306 , n418305 );
or ( n418307 , n418306 , n418095 );
nand ( n418308 , n418302 , n418307 );
buf ( n418309 , n418308 );
xor ( n418310 , n418227 , n418240 );
and ( n418311 , n418310 , n418258 );
and ( n418312 , n418227 , n418240 );
or ( n418313 , n418311 , n418312 );
buf ( n418314 , n418313 );
buf ( n418315 , n418314 );
xor ( n418316 , n418309 , n418315 );
xor ( n418317 , n405570 , n405595 );
xor ( n418318 , n418317 , n405621 );
buf ( n418319 , n418318 );
buf ( n418320 , n418319 );
and ( n418321 , n418316 , n418320 );
and ( n418322 , n418309 , n418315 );
or ( n418323 , n418321 , n418322 );
buf ( n418324 , n418323 );
buf ( n418325 , n418324 );
buf ( n418326 , n418325 );
buf ( n418327 , n418326 );
buf ( n418328 , n418327 );
xor ( n418329 , n418299 , n418328 );
buf ( n418330 , n418329 );
buf ( n418331 , n418330 );
xor ( n418332 , n418193 , n418206 );
and ( n418333 , n418332 , n418213 );
and ( n418334 , n418193 , n418206 );
or ( n418335 , n418333 , n418334 );
buf ( n418336 , n418335 );
buf ( n418337 , n418336 );
xor ( n418338 , n404683 , n404708 );
xor ( n418339 , n418338 , n404773 );
buf ( n418340 , n418339 );
buf ( n418341 , n418340 );
xor ( n418342 , n418337 , n418341 );
xor ( n418343 , n404851 , n405106 );
xor ( n418344 , n418343 , n405126 );
buf ( n418345 , n418344 );
buf ( n418346 , n418345 );
xor ( n418347 , n418342 , n418346 );
buf ( n418348 , n418347 );
buf ( n418349 , n418348 );
not ( n418350 , n418349 );
xor ( n418351 , n418309 , n418315 );
xor ( n418352 , n418351 , n418320 );
buf ( n418353 , n418352 );
buf ( n418354 , n418353 );
not ( n418355 , n418354 );
or ( n418356 , n418350 , n418355 );
xor ( n418357 , n418139 , n418164 );
and ( n418358 , n418357 , n418171 );
and ( n418359 , n418139 , n418164 );
or ( n418360 , n418358 , n418359 );
buf ( n418361 , n418360 );
buf ( n418362 , n418361 );
buf ( n418363 , n405228 );
not ( n418364 , n418363 );
xor ( n418365 , n405204 , n405417 );
buf ( n418366 , n418365 );
not ( n418367 , n418366 );
or ( n418368 , n418364 , n418367 );
buf ( n418369 , n418365 );
buf ( n418370 , n405228 );
or ( n418371 , n418369 , n418370 );
nand ( n418372 , n418368 , n418371 );
buf ( n418373 , n418372 );
buf ( n418374 , n418373 );
xor ( n418375 , n418148 , n418154 );
and ( n418376 , n418375 , n418161 );
and ( n418377 , n418148 , n418154 );
or ( n418378 , n418376 , n418377 );
buf ( n418379 , n418378 );
buf ( n418380 , n418379 );
xor ( n418381 , n418374 , n418380 );
buf ( n418382 , n418128 );
not ( n418383 , n418382 );
buf ( n418384 , n418383 );
buf ( n418385 , n418384 );
buf ( n418386 , n385064 );
or ( n418387 , n418385 , n418386 );
buf ( n418388 , n405556 );
buf ( n418389 , n384940 );
or ( n418390 , n418388 , n418389 );
nand ( n418391 , n418387 , n418390 );
buf ( n418392 , n418391 );
buf ( n418393 , n418392 );
xor ( n418394 , n418381 , n418393 );
buf ( n418395 , n418394 );
buf ( n418396 , n418395 );
xor ( n418397 , n418362 , n418396 );
xor ( n418398 , n418216 , n418222 );
and ( n418399 , n418398 , n418261 );
and ( n418400 , n418216 , n418222 );
or ( n418401 , n418399 , n418400 );
buf ( n418402 , n418401 );
buf ( n418403 , n418402 );
xor ( n418404 , n418397 , n418403 );
buf ( n418405 , n418404 );
buf ( n418406 , n418405 );
buf ( n418407 , n418353 );
not ( n418408 , n418407 );
not ( n418409 , n418348 );
buf ( n418410 , n418409 );
nand ( n418411 , n418408 , n418410 );
buf ( n418412 , n418411 );
buf ( n418413 , n418412 );
nand ( n418414 , n418406 , n418413 );
buf ( n418415 , n418414 );
buf ( n418416 , n418415 );
nand ( n418417 , n418356 , n418416 );
buf ( n418418 , n418417 );
buf ( n418419 , n418418 );
xor ( n418420 , n418331 , n418419 );
buf ( n418421 , n405632 );
buf ( n418422 , n405625 );
xor ( n418423 , n418421 , n418422 );
buf ( n418424 , n418423 );
buf ( n418425 , n418424 );
buf ( n418426 , n405636 );
and ( n418427 , n418425 , n418426 );
not ( n418428 , n418425 );
buf ( n418429 , n405546 );
and ( n418430 , n418428 , n418429 );
nor ( n418431 , n418427 , n418430 );
buf ( n418432 , n418431 );
buf ( n418433 , n418432 );
xor ( n418434 , n404534 , n82781 );
xor ( n418435 , n418434 , n404588 );
buf ( n418436 , n418435 );
buf ( n418437 , n418436 );
xor ( n418438 , n418374 , n418380 );
and ( n418439 , n418438 , n418393 );
and ( n418440 , n418374 , n418380 );
or ( n418441 , n418439 , n418440 );
buf ( n418442 , n418441 );
buf ( n418443 , n418442 );
xor ( n418444 , n418437 , n418443 );
xor ( n418445 , n418337 , n418341 );
and ( n418446 , n418445 , n418346 );
and ( n418447 , n418337 , n418341 );
or ( n418448 , n418446 , n418447 );
buf ( n418449 , n418448 );
buf ( n418450 , n418449 );
xor ( n418451 , n418444 , n418450 );
buf ( n418452 , n418451 );
buf ( n418453 , n418452 );
xor ( n418454 , n418433 , n418453 );
xor ( n418455 , n418362 , n418396 );
and ( n418456 , n418455 , n418403 );
and ( n418457 , n418362 , n418396 );
or ( n418458 , n418456 , n418457 );
buf ( n418459 , n418458 );
buf ( n418460 , n418459 );
xor ( n418461 , n418454 , n418460 );
buf ( n418462 , n418461 );
buf ( n418463 , n418462 );
xnor ( n418464 , n418420 , n418463 );
buf ( n418465 , n418464 );
buf ( n418466 , n418465 );
and ( n418467 , n418353 , n418348 );
not ( n418468 , n418353 );
and ( n418469 , n418468 , n418409 );
or ( n418470 , n418467 , n418469 );
xor ( n418471 , n418470 , n418405 );
xor ( n418472 , n418062 , n418097 );
and ( n418473 , n418472 , n418104 );
and ( n418474 , n418062 , n418097 );
or ( n418475 , n418473 , n418474 );
buf ( n418476 , n418475 );
not ( n418477 , n418476 );
nand ( n418478 , n418471 , n418477 );
buf ( n418479 , n418478 );
xor ( n418480 , n418174 , n418189 );
and ( n418481 , n418480 , n418264 );
and ( n418482 , n418174 , n418189 );
or ( n418483 , n418481 , n418482 );
buf ( n418484 , n418483 );
buf ( n418485 , n418484 );
buf ( n418486 , n418485 );
buf ( n418487 , n418486 );
buf ( n418488 , n418487 );
and ( n418489 , n418479 , n418488 );
nor ( n418490 , n418471 , n418477 );
buf ( n418491 , n418490 );
nor ( n418492 , n418489 , n418491 );
buf ( n418493 , n418492 );
buf ( n418494 , n418493 );
nand ( n418495 , n418466 , n418494 );
buf ( n418496 , n418495 );
buf ( n418497 , n418496 );
buf ( n418498 , n418484 );
buf ( n418499 , n418476 );
not ( n418500 , n418499 );
buf ( n418501 , n418500 );
buf ( n418502 , n418501 );
and ( n418503 , n418498 , n418502 );
not ( n418504 , n418498 );
buf ( n418505 , n418476 );
and ( n418506 , n418504 , n418505 );
nor ( n418507 , n418503 , n418506 );
buf ( n418508 , n418507 );
and ( n418509 , n418508 , n418471 );
not ( n418510 , n418508 );
not ( n418511 , n418471 );
and ( n418512 , n418510 , n418511 );
nor ( n418513 , n418509 , n418512 );
buf ( n418514 , n418513 );
not ( n418515 , n418514 );
buf ( n418516 , n418515 );
buf ( n418517 , n418516 );
xor ( n418518 , n418107 , n418113 );
and ( n418519 , n418518 , n418267 );
and ( n418520 , n418107 , n418113 );
or ( n418521 , n418519 , n418520 );
buf ( n418522 , n418521 );
buf ( n418523 , n418522 );
not ( n418524 , n418523 );
buf ( n418525 , n418524 );
buf ( n418526 , n418525 );
nand ( n418527 , n418517 , n418526 );
buf ( n418528 , n418527 );
buf ( n418529 , n418528 );
nand ( n418530 , n418293 , n418497 , n418529 );
buf ( n418531 , n418530 );
buf ( n418532 , n418531 );
buf ( n418533 , n418513 );
buf ( n418534 , n418522 );
nand ( n418535 , n418533 , n418534 );
buf ( n418536 , n418535 );
buf ( n418537 , n418536 );
not ( n418538 , n418537 );
buf ( n418539 , n418496 );
nand ( n418540 , n418538 , n418539 );
buf ( n418541 , n418540 );
buf ( n418542 , n418541 );
buf ( n418543 , n418465 );
not ( n418544 , n418543 );
buf ( n418545 , n418544 );
buf ( n418546 , n418545 );
buf ( n418547 , n418493 );
not ( n418548 , n418547 );
buf ( n418549 , n418548 );
buf ( n418550 , n418549 );
nand ( n418551 , n418546 , n418550 );
buf ( n418552 , n418551 );
buf ( n418553 , n418552 );
nand ( n418554 , n418532 , n418542 , n418553 );
buf ( n418555 , n418554 );
buf ( n418556 , n418555 );
xor ( n418557 , n405521 , n405649 );
xor ( n418558 , n418557 , n405654 );
buf ( n418559 , n418558 );
buf ( n418560 , n418559 );
not ( n418561 , n418560 );
not ( n418562 , n418295 );
not ( n418563 , n418297 );
and ( n418564 , n418562 , n418563 );
buf ( n418565 , n418295 );
buf ( n418566 , n418297 );
nand ( n418567 , n418565 , n418566 );
buf ( n418568 , n418567 );
and ( n418569 , n418324 , n418568 );
nor ( n418570 , n418564 , n418569 );
buf ( n418571 , n418570 );
not ( n418572 , n418571 );
buf ( n418573 , n418572 );
not ( n418574 , n418573 );
and ( n418575 , n83281 , n404786 );
not ( n418576 , n83281 );
and ( n418577 , n418576 , n404789 );
or ( n418578 , n418575 , n418577 );
buf ( n418579 , n418578 );
buf ( n418580 , n404658 );
and ( n418581 , n418579 , n418580 );
not ( n418582 , n418579 );
buf ( n418583 , n82880 );
and ( n418584 , n418582 , n418583 );
nor ( n418585 , n418581 , n418584 );
buf ( n418586 , n418585 );
buf ( n418587 , n418586 );
not ( n418588 , n418587 );
buf ( n418589 , n418588 );
not ( n418590 , n418589 );
or ( n418591 , n418574 , n418590 );
buf ( n418592 , n418570 );
not ( n418593 , n418592 );
buf ( n418594 , n418586 );
not ( n418595 , n418594 );
or ( n418596 , n418593 , n418595 );
xor ( n418597 , n418437 , n418443 );
and ( n418598 , n418597 , n418450 );
and ( n418599 , n418437 , n418443 );
or ( n418600 , n418598 , n418599 );
buf ( n418601 , n418600 );
buf ( n418602 , n418601 );
nand ( n418603 , n418596 , n418602 );
buf ( n418604 , n418603 );
nand ( n418605 , n418591 , n418604 );
not ( n418606 , n83285 );
or ( n418607 , n405448 , n405145 );
nand ( n418608 , n405145 , n405448 );
nand ( n418609 , n418607 , n418608 );
not ( n418610 , n418609 );
or ( n418611 , n418606 , n418610 );
or ( n418612 , n418609 , n83285 );
nand ( n418613 , n418611 , n418612 );
not ( n418614 , n418613 );
and ( n418615 , n418605 , n418614 );
not ( n418616 , n418605 );
and ( n418617 , n418616 , n418613 );
nor ( n418618 , n418615 , n418617 );
buf ( n418619 , n418618 );
not ( n418620 , n418619 );
buf ( n418621 , n418620 );
buf ( n418622 , n418621 );
not ( n418623 , n418622 );
or ( n418624 , n418561 , n418623 );
not ( n418625 , n418559 );
nand ( n418626 , n418625 , n418618 );
buf ( n418627 , n418626 );
nand ( n418628 , n418624 , n418627 );
buf ( n418629 , n418628 );
buf ( n418630 , n418629 );
not ( n418631 , n418630 );
buf ( n418632 , n418631 );
buf ( n418633 , n418632 );
buf ( n418634 , n405642 );
buf ( n418635 , n405532 );
xor ( n418636 , n418634 , n418635 );
buf ( n418637 , n405527 );
xor ( n418638 , n418636 , n418637 );
buf ( n418639 , n418638 );
buf ( n418640 , n418639 );
xor ( n418641 , n418433 , n418453 );
and ( n418642 , n418641 , n418460 );
and ( n418643 , n418433 , n418453 );
or ( n418644 , n418642 , n418643 );
buf ( n418645 , n418644 );
buf ( n418646 , n418645 );
xor ( n418647 , n418640 , n418646 );
buf ( n418648 , n418601 );
buf ( n418649 , n418573 );
xor ( n418650 , n418648 , n418649 );
buf ( n418651 , n418589 );
xor ( n418652 , n418650 , n418651 );
buf ( n418653 , n418652 );
buf ( n418654 , n418653 );
and ( n418655 , n418647 , n418654 );
and ( n418656 , n418640 , n418646 );
or ( n418657 , n418655 , n418656 );
buf ( n418658 , n418657 );
buf ( n418659 , n418658 );
not ( n418660 , n418659 );
buf ( n418661 , n418660 );
buf ( n418662 , n418661 );
nand ( n418663 , n418633 , n418662 );
buf ( n418664 , n418663 );
buf ( n418665 , n418664 );
xor ( n418666 , n418640 , n418646 );
xor ( n418667 , n418666 , n418654 );
buf ( n418668 , n418667 );
buf ( n418669 , n418668 );
not ( n418670 , n418669 );
buf ( n418671 , n418670 );
buf ( n418672 , n418671 );
buf ( n418673 , n418330 );
not ( n418674 , n418673 );
buf ( n418675 , n418418 );
not ( n418676 , n418675 );
or ( n418677 , n418674 , n418676 );
or ( n418678 , n418330 , n418418 );
nand ( n418679 , n418678 , n418462 );
buf ( n418680 , n418679 );
nand ( n418681 , n418677 , n418680 );
buf ( n418682 , n418681 );
buf ( n418683 , n418682 );
not ( n418684 , n418683 );
buf ( n418685 , n418684 );
buf ( n418686 , n418685 );
nand ( n418687 , n418672 , n418686 );
buf ( n418688 , n418687 );
buf ( n418689 , n418688 );
and ( n418690 , n418665 , n418689 );
buf ( n418691 , n418690 );
buf ( n418692 , n418691 );
buf ( n418693 , n405506 );
not ( n418694 , n418693 );
buf ( n418695 , n405658 );
not ( n418696 , n418695 );
buf ( n418697 , n418696 );
buf ( n418698 , n418697 );
not ( n418699 , n418698 );
or ( n418700 , n418694 , n418699 );
buf ( n418701 , n405511 );
buf ( n418702 , n405658 );
nand ( n418703 , n418701 , n418702 );
buf ( n418704 , n418703 );
buf ( n418705 , n418704 );
nand ( n418706 , n418700 , n418705 );
buf ( n418707 , n418706 );
buf ( n418708 , n418707 );
buf ( n418709 , n405499 );
and ( n418710 , n418708 , n418709 );
not ( n418711 , n418708 );
buf ( n418712 , n405502 );
and ( n418713 , n418711 , n418712 );
nor ( n418714 , n418710 , n418713 );
buf ( n418715 , n418714 );
buf ( n418716 , n418715 );
buf ( n418717 , n418559 );
not ( n418718 , n418717 );
buf ( n418719 , n418718 );
not ( n418720 , n418719 );
buf ( n418721 , n418613 );
buf ( n418722 , n418721 );
buf ( n418723 , n418722 );
not ( n418724 , n418723 );
and ( n418725 , n418720 , n418724 );
buf ( n418726 , n418719 );
buf ( n418727 , n418723 );
nand ( n418728 , n418726 , n418727 );
buf ( n418729 , n418728 );
and ( n418730 , n418729 , n418605 );
nor ( n418731 , n418725 , n418730 );
buf ( n418732 , n418731 );
nand ( n418733 , n418716 , n418732 );
buf ( n418734 , n418733 );
buf ( n418735 , n418734 );
nand ( n418736 , n418556 , n418692 , n418735 );
buf ( n418737 , n418736 );
buf ( n418738 , n418737 );
buf ( n418739 , n418629 );
buf ( n418740 , n418658 );
nand ( n418741 , n418739 , n418740 );
buf ( n418742 , n418741 );
buf ( n418743 , n418742 );
buf ( n418744 , n418668 );
buf ( n418745 , n418682 );
nand ( n418746 , n418744 , n418745 );
buf ( n418747 , n418746 );
buf ( n418748 , n418747 );
nand ( n418749 , n418743 , n418748 );
buf ( n418750 , n418749 );
buf ( n418751 , n418750 );
buf ( n418752 , n418664 );
and ( n418753 , n418751 , n418752 );
buf ( n418754 , n418753 );
buf ( n418755 , n418754 );
buf ( n418756 , n418734 );
nand ( n418757 , n418755 , n418756 );
buf ( n418758 , n418757 );
buf ( n418759 , n418758 );
or ( n418760 , n418715 , n418731 );
buf ( n418761 , n418760 );
nand ( n418762 , n418738 , n418759 , n418761 );
buf ( n418763 , n418762 );
buf ( n418764 , n418763 );
not ( n418765 , n418764 );
or ( n418766 , n405690 , n418765 );
buf ( n418767 , n405685 );
buf ( n418768 , n405493 );
buf ( n418769 , n405660 );
and ( n418770 , n418768 , n418769 );
buf ( n418771 , n418770 );
buf ( n418772 , n418771 );
nand ( n418773 , n418767 , n418772 );
buf ( n418774 , n418773 );
buf ( n418775 , n418774 );
or ( n418776 , n405668 , n405682 );
buf ( n418777 , n418776 );
and ( n418778 , n418775 , n418777 );
buf ( n418779 , n418778 );
buf ( n418780 , n418779 );
nand ( n418781 , n418766 , n418780 );
buf ( n418782 , n418781 );
not ( n418783 , n399723 );
not ( n418784 , n399731 );
or ( n418785 , n418783 , n418784 );
buf ( n418786 , n399696 );
buf ( n418787 , n399720 );
nand ( n418788 , n418786 , n418787 );
buf ( n418789 , n418788 );
nand ( n418790 , n418785 , n418789 );
xor ( n418791 , n418790 , n399682 );
not ( n418792 , n418791 );
xor ( n418793 , n398332 , n398598 );
xor ( n418794 , n418793 , n398776 );
buf ( n418795 , n418794 );
buf ( n418796 , n418795 );
not ( n418797 , n418796 );
buf ( n418798 , n418797 );
nand ( n418799 , n418792 , n418798 );
buf ( n418800 , n418799 );
buf ( n418801 , n404466 );
not ( n418802 , n418801 );
buf ( n418803 , n418802 );
buf ( n418804 , n418803 );
not ( n418805 , n418804 );
buf ( n418806 , n404479 );
not ( n418807 , n418806 );
or ( n418808 , n418805 , n418807 );
buf ( n418809 , n404466 );
not ( n418810 , n418809 );
buf ( n418811 , n404478 );
not ( n418812 , n418811 );
or ( n418813 , n418810 , n418812 );
buf ( n418814 , n404490 );
nand ( n418815 , n418813 , n418814 );
buf ( n418816 , n418815 );
buf ( n418817 , n418816 );
nand ( n418818 , n418808 , n418817 );
buf ( n418819 , n418818 );
buf ( n418820 , n418819 );
and ( n418821 , n418800 , n418820 );
not ( n418822 , n418791 );
nor ( n418823 , n418822 , n418798 );
buf ( n418824 , n418823 );
nor ( n418825 , n418821 , n418824 );
buf ( n418826 , n418825 );
and ( n418827 , n78431 , n77786 );
not ( n418828 , n78431 );
not ( n418829 , n77786 );
and ( n418830 , n418828 , n418829 );
nor ( n418831 , n418827 , n418830 );
not ( n418832 , n418831 );
or ( n418833 , n418832 , n399079 );
not ( n418834 , n399079 );
or ( n418835 , n418834 , n418831 );
nand ( n418836 , n418833 , n418835 );
nand ( n418837 , n418826 , n418836 );
not ( n418838 , n418837 );
buf ( n418839 , n418838 );
not ( n418840 , n418839 );
buf ( n418841 , n418840 );
buf ( n418842 , n404450 );
not ( n418843 , n418842 );
buf ( n418844 , n404506 );
not ( n418845 , n418844 );
or ( n418846 , n418843 , n418845 );
buf ( n418847 , n404456 );
not ( n418848 , n418847 );
buf ( n418849 , n404501 );
not ( n418850 , n418849 );
or ( n418851 , n418848 , n418850 );
buf ( n418852 , n404446 );
buf ( n418853 , n418852 );
nand ( n418854 , n418851 , n418853 );
buf ( n418855 , n418854 );
buf ( n418856 , n418855 );
nand ( n418857 , n418846 , n418856 );
buf ( n418858 , n418857 );
buf ( n418859 , n418858 );
not ( n418860 , n418819 );
xor ( n418861 , n418795 , n418860 );
xnor ( n418862 , n418861 , n418791 );
buf ( n418863 , n418862 );
nor ( n418864 , n418859 , n418863 );
buf ( n418865 , n418864 );
buf ( n418866 , n418865 );
not ( n418867 , n418866 );
buf ( n418868 , n418867 );
nand ( n418869 , n82759 , n418782 , n418841 , n418868 );
buf ( n418870 , n402508 );
buf ( n418871 , n403315 );
nand ( n418872 , n418870 , n418871 );
buf ( n418873 , n418872 );
buf ( n418874 , n418873 );
buf ( n418875 , n404436 );
not ( n418876 , n418875 );
buf ( n418877 , n418876 );
buf ( n418878 , n418877 );
buf ( n418879 , n404416 );
nand ( n418880 , n418878 , n418879 );
buf ( n418881 , n418880 );
buf ( n418882 , n418881 );
nand ( n418883 , n418874 , n418882 );
buf ( n418884 , n418883 );
buf ( n418885 , n418884 );
buf ( n418886 , n82756 );
buf ( n418887 , n403321 );
nand ( n418888 , n418885 , n418886 , n418887 );
buf ( n418889 , n418888 );
nor ( n418890 , n418836 , n418826 );
nor ( n418891 , n82749 , n82755 );
nor ( n418892 , n418890 , n418891 );
buf ( n418893 , n418862 );
buf ( n418894 , n418858 );
nand ( n418895 , n418893 , n418894 );
buf ( n418896 , n418895 );
nand ( n418897 , n418889 , n418892 , n418896 );
buf ( n418898 , n418890 );
not ( n418899 , n418898 );
buf ( n418900 , n418899 );
buf ( n418901 , n418900 );
buf ( n418902 , n418865 );
and ( n418903 , n418901 , n418902 );
buf ( n418904 , n418838 );
nor ( n418905 , n418903 , n418904 );
buf ( n418906 , n418905 );
nand ( n418907 , n418897 , n418906 );
nand ( n418908 , n418869 , n418907 );
not ( n418909 , n418908 );
or ( n418910 , n78652 , n418909 );
not ( n418911 , n399955 );
nand ( n418912 , n399073 , n399749 );
not ( n418913 , n418912 );
not ( n418914 , n418913 );
or ( n418915 , n418911 , n418914 );
or ( n418916 , n78649 , n399942 );
nand ( n418917 , n418915 , n418916 );
not ( n418918 , n418917 );
nand ( n418919 , n418910 , n418918 );
xor ( n418920 , n383405 , n383744 );
xor ( n418921 , n418920 , n383755 );
xor ( n418922 , n64698 , n385389 );
xor ( n418923 , n418922 , n385407 );
buf ( n418924 , n418923 );
nand ( n418925 , n418921 , n418924 );
buf ( n418926 , n418925 );
or ( n418927 , n418921 , n418924 );
xor ( n418928 , n399875 , n399879 );
and ( n418929 , n418928 , n399886 );
and ( n418930 , n399875 , n399879 );
or ( n418931 , n418929 , n418930 );
buf ( n418932 , n418931 );
nand ( n418933 , n418927 , n418932 );
buf ( n418934 , n418933 );
and ( n418935 , n418926 , n418934 );
buf ( n418936 , n418935 );
xor ( n418937 , n383396 , n383392 );
xnor ( n418938 , n418937 , n383758 );
and ( n418939 , n418936 , n418938 );
xor ( n418940 , n399753 , n399757 );
and ( n418941 , n418940 , n399771 );
and ( n418942 , n399753 , n399757 );
or ( n418943 , n418941 , n418942 );
buf ( n418944 , n418943 );
buf ( n418945 , n418944 );
buf ( n418946 , n399923 );
buf ( n418947 , n399917 );
or ( n418948 , n418946 , n418947 );
buf ( n418949 , n418948 );
buf ( n418950 , n418949 );
buf ( n418951 , n399930 );
and ( n418952 , n418950 , n418951 );
buf ( n418953 , n399923 );
buf ( n418954 , n399917 );
and ( n418955 , n418953 , n418954 );
buf ( n418956 , n418955 );
buf ( n418957 , n418956 );
nor ( n418958 , n418952 , n418957 );
buf ( n418959 , n418958 );
buf ( n418960 , n418959 );
xor ( n418961 , n418945 , n418960 );
buf ( n418962 , n385459 );
buf ( n418963 , n385542 );
xor ( n418964 , n418962 , n418963 );
buf ( n418965 , n385528 );
xnor ( n418966 , n418964 , n418965 );
buf ( n418967 , n418966 );
buf ( n418968 , n418967 );
and ( n418969 , n418961 , n418968 );
and ( n418970 , n418945 , n418960 );
or ( n418971 , n418969 , n418970 );
buf ( n418972 , n418971 );
or ( n418973 , n418939 , n418972 );
not ( n418974 , n418936 );
not ( n418975 , n418938 );
nand ( n418976 , n418974 , n418975 );
nand ( n418977 , n418973 , n418976 );
xor ( n418978 , n385412 , n385416 );
xor ( n418979 , n418978 , n385549 );
buf ( n418980 , n418979 );
buf ( n418981 , n418980 );
not ( n418982 , n418981 );
buf ( n418983 , n418982 );
buf ( n418984 , n418983 );
not ( n418985 , n418984 );
and ( n418986 , n385564 , n386170 );
not ( n418987 , n385564 );
not ( n418988 , n386170 );
and ( n418989 , n418987 , n418988 );
nor ( n418990 , n418986 , n418989 );
and ( n418991 , n418990 , n64918 );
not ( n418992 , n418990 );
and ( n418993 , n418992 , n385584 );
nor ( n418994 , n418991 , n418993 );
buf ( n418995 , n418994 );
not ( n418996 , n418995 );
or ( n418997 , n418985 , n418996 );
buf ( n418998 , n418932 );
buf ( n418999 , n418924 );
xor ( n419000 , n418998 , n418999 );
not ( n419001 , n418921 );
buf ( n419002 , n419001 );
xnor ( n419003 , n419000 , n419002 );
buf ( n419004 , n419003 );
not ( n419005 , n419004 );
xor ( n419006 , n385632 , n386164 );
buf ( n419007 , n385617 );
buf ( n419008 , n419007 );
buf ( n419009 , n419008 );
xor ( n419010 , n419006 , n419009 );
buf ( n419011 , n419010 );
not ( n419012 , n419011 );
not ( n419013 , n78533 );
not ( n419014 , n78536 );
and ( n419015 , n419013 , n419014 );
nand ( n419016 , n78533 , n78536 );
and ( n419017 , n399848 , n419016 );
nor ( n419018 , n419015 , n419017 );
buf ( n419019 , n419018 );
nand ( n419020 , n419012 , n419019 );
buf ( n419021 , n419020 );
not ( n419022 , n419021 );
or ( n419023 , n419005 , n419022 );
buf ( n419024 , n419018 );
not ( n419025 , n419024 );
buf ( n419026 , n419025 );
buf ( n419027 , n419026 );
buf ( n419028 , n419010 );
nand ( n419029 , n419027 , n419028 );
buf ( n419030 , n419029 );
nand ( n419031 , n419023 , n419030 );
buf ( n419032 , n419031 );
nand ( n419033 , n418997 , n419032 );
buf ( n419034 , n419033 );
buf ( n419035 , n419034 );
buf ( n419036 , n418994 );
not ( n419037 , n419036 );
buf ( n419038 , n418980 );
nand ( n419039 , n419037 , n419038 );
buf ( n419040 , n419039 );
buf ( n419041 , n419040 );
nand ( n419042 , n419035 , n419041 );
buf ( n419043 , n419042 );
buf ( n419044 , n419043 );
not ( n419045 , n419044 );
buf ( n419046 , n419045 );
and ( n419047 , n418977 , n419046 );
not ( n419048 , n418977 );
and ( n419049 , n419048 , n419043 );
nor ( n419050 , n419047 , n419049 );
xor ( n419051 , n386179 , n386180 );
buf ( n419052 , n419051 );
buf ( n419053 , n419052 );
buf ( n419054 , n386176 );
and ( n419055 , n419053 , n419054 );
not ( n419056 , n419053 );
buf ( n419057 , n386176 );
not ( n419058 , n419057 );
buf ( n419059 , n419058 );
buf ( n419060 , n419059 );
and ( n419061 , n419056 , n419060 );
nor ( n419062 , n419055 , n419061 );
buf ( n419063 , n419062 );
buf ( n419064 , n382391 );
buf ( n419065 , n61799 );
xor ( n419066 , n419064 , n419065 );
buf ( n419067 , n382385 );
xor ( n419068 , n419066 , n419067 );
buf ( n419069 , n419068 );
buf ( n419070 , n419069 );
xor ( n419071 , n382461 , n383385 );
xor ( n419072 , n419071 , n383761 );
buf ( n419073 , n419072 );
xor ( n419074 , n419070 , n419073 );
buf ( n419075 , n419074 );
xor ( n419076 , n419063 , n419075 );
xor ( n419077 , n419050 , n419076 );
and ( n419078 , n418936 , n418938 );
not ( n419079 , n418936 );
and ( n419080 , n419079 , n418975 );
nor ( n419081 , n419078 , n419080 );
xor ( n419082 , n419081 , n418972 );
buf ( n419083 , n419082 );
buf ( n419084 , n418983 );
not ( n419085 , n419084 );
buf ( n419086 , n418994 );
not ( n419087 , n419086 );
buf ( n419088 , n419087 );
buf ( n419089 , n419088 );
not ( n419090 , n419089 );
or ( n419091 , n419085 , n419090 );
buf ( n419092 , n418994 );
buf ( n419093 , n418980 );
nand ( n419094 , n419092 , n419093 );
buf ( n419095 , n419094 );
buf ( n419096 , n419095 );
nand ( n419097 , n419091 , n419096 );
buf ( n419098 , n419097 );
buf ( n419099 , n419098 );
buf ( n419100 , n419031 );
not ( n419101 , n419100 );
buf ( n419102 , n419101 );
buf ( n419103 , n419102 );
and ( n419104 , n419099 , n419103 );
not ( n419105 , n419099 );
buf ( n419106 , n419031 );
and ( n419107 , n419105 , n419106 );
nor ( n419108 , n419104 , n419107 );
buf ( n419109 , n419108 );
buf ( n419110 , n419109 );
xor ( n419111 , n419083 , n419110 );
buf ( n419112 , n399815 );
buf ( n419113 , n399794 );
not ( n419114 , n419113 );
buf ( n419115 , n419114 );
buf ( n419116 , n419115 );
buf ( n419117 , n399773 );
nand ( n419118 , n419116 , n419117 );
buf ( n419119 , n419118 );
buf ( n419120 , n419119 );
and ( n419121 , n419112 , n419120 );
buf ( n419122 , n399794 );
not ( n419123 , n419122 );
buf ( n419124 , n399773 );
nor ( n419125 , n419123 , n419124 );
buf ( n419126 , n419125 );
buf ( n419127 , n419126 );
nor ( n419128 , n419121 , n419127 );
buf ( n419129 , n419128 );
buf ( n419130 , n419129 );
xor ( n419131 , n399889 , n399913 );
and ( n419132 , n419131 , n399934 );
and ( n419133 , n399889 , n399913 );
or ( n419134 , n419132 , n419133 );
buf ( n419135 , n419134 );
buf ( n419136 , n419135 );
not ( n419137 , n419136 );
buf ( n419138 , n419137 );
buf ( n419139 , n419138 );
xor ( n419140 , n419130 , n419139 );
xor ( n419141 , n418945 , n418960 );
xor ( n419142 , n419141 , n418968 );
buf ( n419143 , n419142 );
buf ( n419144 , n419143 );
and ( n419145 , n419140 , n419144 );
and ( n419146 , n419130 , n419139 );
or ( n419147 , n419145 , n419146 );
buf ( n419148 , n419147 );
buf ( n419149 , n419148 );
and ( n419150 , n419111 , n419149 );
and ( n419151 , n419083 , n419110 );
or ( n419152 , n419150 , n419151 );
buf ( n419153 , n419152 );
nand ( n419154 , n419077 , n419153 );
xor ( n419155 , n419083 , n419110 );
xor ( n419156 , n419155 , n419149 );
buf ( n419157 , n419156 );
buf ( n419158 , n419010 );
buf ( n419159 , n419026 );
xor ( n419160 , n419158 , n419159 );
buf ( n419161 , n419004 );
xnor ( n419162 , n419160 , n419161 );
buf ( n419163 , n419162 );
xor ( n419164 , n399852 , n399864 );
and ( n419165 , n419164 , n399937 );
and ( n419166 , n399852 , n399864 );
or ( n419167 , n419165 , n419166 );
buf ( n419168 , n419167 );
buf ( n419169 , n419168 );
not ( n419170 , n419169 );
buf ( n419171 , n419170 );
xor ( n419172 , n419163 , n419171 );
xor ( n419173 , n419130 , n419139 );
xor ( n419174 , n419173 , n419144 );
buf ( n419175 , n419174 );
and ( n419176 , n419172 , n419175 );
and ( n419177 , n419163 , n419171 );
or ( n419178 , n419176 , n419177 );
nand ( n419179 , n419157 , n419178 );
not ( n419180 , n399939 );
buf ( n419181 , n78511 );
not ( n419182 , n419181 );
buf ( n419183 , n399822 );
not ( n419184 , n419183 );
buf ( n419185 , n419184 );
buf ( n419186 , n419185 );
nand ( n419187 , n419182 , n419186 );
buf ( n419188 , n419187 );
not ( n419189 , n419188 );
or ( n419190 , n419180 , n419189 );
buf ( n419191 , n419185 );
not ( n419192 , n419191 );
buf ( n419193 , n78511 );
nand ( n419194 , n419192 , n419193 );
buf ( n419195 , n419194 );
nand ( n419196 , n419190 , n419195 );
not ( n419197 , n419196 );
xor ( n419198 , n419163 , n419171 );
xor ( n419199 , n419198 , n419175 );
nand ( n419200 , n419197 , n419199 );
and ( n419201 , n419154 , n419179 , n419200 );
not ( n419202 , n419201 );
buf ( n419203 , n382409 );
not ( n419204 , n419203 );
buf ( n419205 , n382372 );
not ( n419206 , n419205 );
or ( n419207 , n419204 , n419206 );
buf ( n419208 , n382375 );
buf ( n419209 , n382406 );
nand ( n419210 , n419208 , n419209 );
buf ( n419211 , n419210 );
buf ( n419212 , n419211 );
nand ( n419213 , n419207 , n419212 );
buf ( n419214 , n419213 );
buf ( n419215 , n419214 );
buf ( n419216 , n383764 );
not ( n419217 , n419216 );
buf ( n419218 , n419217 );
buf ( n419219 , n419218 );
and ( n419220 , n419215 , n419219 );
not ( n419221 , n419215 );
buf ( n419222 , n383764 );
and ( n419223 , n419221 , n419222 );
nor ( n419224 , n419220 , n419223 );
buf ( n419225 , n419224 );
buf ( n419226 , n419225 );
xor ( n419227 , n385190 , n385197 );
xor ( n419228 , n419227 , n386186 );
buf ( n419229 , n419228 );
buf ( n419230 , n419229 );
xor ( n419231 , n419226 , n419230 );
buf ( n419232 , n419063 );
buf ( n419233 , n419072 );
buf ( n419234 , n419069 );
or ( n419235 , n419233 , n419234 );
buf ( n419236 , n419235 );
buf ( n419237 , n419236 );
and ( n419238 , n419232 , n419237 );
and ( n419239 , n419070 , n419073 );
buf ( n419240 , n419239 );
buf ( n419241 , n419240 );
nor ( n419242 , n419238 , n419241 );
buf ( n419243 , n419242 );
buf ( n419244 , n419243 );
and ( n419245 , n419231 , n419244 );
and ( n419246 , n419226 , n419230 );
or ( n419247 , n419245 , n419246 );
buf ( n419248 , n419247 );
not ( n419249 , n419248 );
not ( n419250 , n386190 );
not ( n419251 , n64538 );
and ( n419252 , n419250 , n419251 );
and ( n419253 , n386190 , n64538 );
nor ( n419254 , n419252 , n419253 );
not ( n419255 , n64531 );
and ( n419256 , n419254 , n419255 );
not ( n419257 , n419254 );
and ( n419258 , n419257 , n64531 );
nor ( n419259 , n419256 , n419258 );
not ( n419260 , n419259 );
or ( n419261 , n419249 , n419260 );
xor ( n419262 , n419226 , n419230 );
xor ( n419263 , n419262 , n419244 );
buf ( n419264 , n419263 );
not ( n419265 , n419076 );
not ( n419266 , n418977 );
nand ( n419267 , n419266 , n419046 );
not ( n419268 , n419267 );
or ( n419269 , n419265 , n419268 );
buf ( n419270 , n419046 );
not ( n419271 , n419270 );
buf ( n419272 , n418977 );
nand ( n419273 , n419271 , n419272 );
buf ( n419274 , n419273 );
nand ( n419275 , n419269 , n419274 );
not ( n419276 , n419275 );
nand ( n419277 , n419264 , n419276 );
nand ( n419278 , n419261 , n419277 );
nor ( n419279 , n419202 , n419278 );
and ( n419280 , n418919 , n419279 );
not ( n419281 , n419278 );
not ( n419282 , n419281 );
not ( n419283 , n419154 );
nor ( n419284 , n419197 , n419199 );
nand ( n419285 , n419284 , n419179 );
buf ( n419286 , n419285 );
buf ( n419287 , n419157 );
not ( n419288 , n419287 );
buf ( n419289 , n419288 );
not ( n419290 , n419178 );
nand ( n419291 , n419289 , n419290 );
buf ( n419292 , n419291 );
nand ( n419293 , n419286 , n419292 );
buf ( n419294 , n419293 );
not ( n419295 , n419294 );
or ( n419296 , n419283 , n419295 );
or ( n419297 , n419153 , n419077 );
nand ( n419298 , n419296 , n419297 );
not ( n419299 , n419298 );
or ( n419300 , n419282 , n419299 );
buf ( n419301 , n419264 );
not ( n419302 , n419301 );
buf ( n419303 , n419275 );
nand ( n419304 , n419302 , n419303 );
buf ( n419305 , n419304 );
nand ( n419306 , n419259 , n419248 );
buf ( n419307 , n419306 );
not ( n419308 , n419307 );
buf ( n419309 , n419308 );
nor ( n419310 , n419305 , n419309 );
buf ( n419311 , n419259 );
buf ( n419312 , n419248 );
or ( n419313 , n419311 , n419312 );
buf ( n419314 , n419313 );
not ( n419315 , n419314 );
nor ( n419316 , n419310 , n419315 );
nand ( n419317 , n419300 , n419316 );
nor ( n419318 , n419280 , n419317 );
buf ( n419319 , n374060 );
buf ( n419320 , n375849 );
nand ( n419321 , n419319 , n419320 );
buf ( n419322 , n419321 );
nor ( n419323 , n419318 , n419322 );
buf ( n419324 , n64524 );
not ( n419325 , n419324 );
buf ( n419326 , n386195 );
not ( n419327 , n419326 );
buf ( n419328 , n419327 );
buf ( n419329 , n419328 );
nand ( n419330 , n419325 , n419329 );
buf ( n419331 , n419330 );
nand ( n419332 , n419331 , n387093 );
not ( n419333 , n67818 );
not ( n419334 , n388709 );
or ( n419335 , n419333 , n419334 );
nand ( n419336 , n419335 , n67097 );
nor ( n419337 , n419332 , n419336 );
buf ( n419338 , n69484 );
buf ( n419339 , n72614 );
and ( n419340 , n419338 , n419339 );
buf ( n419341 , n419340 );
and ( n419342 , n393714 , n393636 );
and ( n419343 , n419337 , n419341 , n419342 );
nand ( n419344 , n393797 , n72761 );
nand ( n419345 , n72592 , n72600 );
nor ( n419346 , n419344 , n419345 );
buf ( n419347 , n71497 );
nand ( n419348 , n419343 , n419346 , n419347 );
not ( n419349 , n419348 );
and ( n419350 , n419323 , n419349 );
not ( n419351 , n375849 );
buf ( n419352 , n374052 );
not ( n419353 , n419352 );
buf ( n419354 , n373560 );
not ( n419355 , n419354 );
not ( n419356 , n373056 );
buf ( n419357 , n419356 );
not ( n419358 , n52818 );
buf ( n419359 , n419358 );
buf ( n419360 , n373080 );
not ( n419361 , n419360 );
buf ( n419362 , n419361 );
buf ( n419363 , n419362 );
nand ( n419364 , n419359 , n419363 );
buf ( n419365 , n419364 );
buf ( n419366 , n419365 );
or ( n419367 , n419357 , n419366 );
buf ( n419368 , n373053 );
not ( n419369 , n419368 );
buf ( n419370 , n373007 );
buf ( n419371 , n419370 );
buf ( n419372 , n419371 );
buf ( n419373 , n419372 );
nand ( n419374 , n419369 , n419373 );
buf ( n419375 , n419374 );
buf ( n419376 , n419375 );
nand ( n419377 , n419367 , n419376 );
buf ( n419378 , n419377 );
buf ( n419379 , n419378 );
not ( n419380 , n419379 );
or ( n419381 , n419355 , n419380 );
buf ( n419382 , n373537 );
buf ( n419383 , n373557 );
or ( n419384 , n419382 , n419383 );
buf ( n419385 , n419384 );
buf ( n419386 , n419385 );
nand ( n419387 , n419381 , n419386 );
buf ( n419388 , n419387 );
buf ( n419389 , n419388 );
not ( n419390 , n419389 );
or ( n419391 , n419353 , n419390 );
buf ( n419392 , n374046 );
buf ( n419393 , n53244 );
and ( n419394 , n419392 , n419393 );
buf ( n419395 , n419394 );
buf ( n419396 , n419395 );
not ( n419397 , n419396 );
buf ( n419398 , n419397 );
buf ( n419399 , n419398 );
not ( n419400 , n419399 );
buf ( n419401 , n374055 );
not ( n419402 , n419401 );
or ( n419403 , n419400 , n419402 );
buf ( n419404 , n371978 );
not ( n419405 , n419404 );
buf ( n419406 , n371997 );
nor ( n419407 , n419405 , n419406 );
buf ( n419408 , n419407 );
buf ( n419409 , n371330 );
buf ( n419410 , n371372 );
and ( n419411 , n419409 , n419410 );
buf ( n419412 , n419411 );
nor ( n419413 , n419408 , n419412 );
not ( n419414 , n419413 );
buf ( n419415 , n369164 );
buf ( n419416 , n370132 );
nand ( n419417 , n419415 , n419416 );
buf ( n419418 , n419417 );
not ( n419419 , n419418 );
nand ( n419420 , n372000 , n419419 );
not ( n419421 , n419420 );
or ( n419422 , n419414 , n419421 );
nor ( n419423 , n371974 , n371375 );
nand ( n419424 , n419422 , n419423 );
buf ( n419425 , n371973 );
buf ( n419426 , n371968 );
and ( n419427 , n419425 , n419426 );
buf ( n419428 , n419427 );
buf ( n419429 , n419428 );
buf ( n419430 , n419395 );
nor ( n419431 , n419429 , n419430 );
buf ( n419432 , n419431 );
nand ( n419433 , n419424 , n419432 );
buf ( n419434 , n419433 );
nand ( n419435 , n419403 , n419434 );
buf ( n419436 , n419435 );
buf ( n419437 , n419436 );
nand ( n419438 , n419391 , n419437 );
buf ( n419439 , n419438 );
not ( n419440 , n419439 );
or ( n419441 , n419351 , n419440 );
not ( n419442 , n375398 );
not ( n419443 , n55177 );
nor ( n419444 , n375520 , n375535 );
not ( n419445 , n419444 );
not ( n419446 , n375547 );
or ( n419447 , n419445 , n419446 );
buf ( n419448 , n375546 );
not ( n419449 , n419448 );
buf ( n419450 , n419449 );
buf ( n419451 , n419450 );
buf ( n419452 , n55212 );
not ( n419453 , n419452 );
buf ( n419454 , n419453 );
buf ( n419455 , n419454 );
nand ( n419456 , n419451 , n419455 );
buf ( n419457 , n419456 );
nand ( n419458 , n419447 , n419457 );
not ( n419459 , n419458 );
or ( n419460 , n419443 , n419459 );
buf ( n419461 , n55070 );
buf ( n419462 , n375501 );
nand ( n419463 , n419461 , n419462 );
buf ( n419464 , n419463 );
nand ( n419465 , n419460 , n419464 );
not ( n419466 , n419465 );
or ( n419467 , n419442 , n419466 );
or ( n419468 , n375274 , n55065 );
nand ( n419469 , n419467 , n419468 );
buf ( n419470 , n419469 );
buf ( n419471 , n375846 );
and ( n419472 , n419470 , n419471 );
buf ( n419473 , n375843 );
not ( n419474 , n419473 );
buf ( n419475 , n419474 );
buf ( n419476 , n419475 );
not ( n419477 , n419476 );
not ( n419478 , n375801 );
not ( n419479 , n55315 );
nand ( n419480 , n419479 , n55329 );
buf ( n419481 , n419480 );
not ( n419482 , n375816 );
buf ( n419483 , n419482 );
or ( n419484 , n419481 , n419483 );
buf ( n419485 , n375805 );
buf ( n419486 , n55483 );
or ( n419487 , n419485 , n419486 );
buf ( n419488 , n419487 );
buf ( n419489 , n419488 );
nand ( n419490 , n419484 , n419489 );
buf ( n419491 , n419490 );
not ( n419492 , n419491 );
or ( n419493 , n419478 , n419492 );
buf ( n419494 , n375754 );
buf ( n419495 , n375798 );
or ( n419496 , n419494 , n419495 );
buf ( n419497 , n419496 );
nand ( n419498 , n419493 , n419497 );
buf ( n419499 , n419498 );
not ( n419500 , n419499 );
or ( n419501 , n419477 , n419500 );
buf ( n419502 , n375836 );
buf ( n419503 , n375840 );
nand ( n419504 , n419502 , n419503 );
buf ( n419505 , n419504 );
buf ( n419506 , n419505 );
nand ( n419507 , n419501 , n419506 );
buf ( n419508 , n419507 );
buf ( n419509 , n419508 );
nor ( n419510 , n419472 , n419509 );
buf ( n419511 , n419510 );
nand ( n419512 , n419441 , n419511 );
nor ( n419513 , n419350 , n419512 );
nand ( n419514 , n72847 , n419513 );
buf ( n419515 , n419514 );
not ( n419516 , n419515 );
or ( n419517 , n364731 , n419516 );
not ( n419518 , n364147 );
buf ( n419519 , n363651 );
buf ( n419520 , n43127 );
nand ( n419521 , n419519 , n419520 );
buf ( n419522 , n419521 );
or ( n419523 , n419522 , n363914 );
nand ( n419524 , n363905 , n363911 );
nand ( n419525 , n419523 , n419524 );
not ( n419526 , n419525 );
or ( n419527 , n419518 , n419526 );
buf ( n419528 , n364140 );
not ( n419529 , n419528 );
buf ( n419530 , n364145 );
nand ( n419531 , n419529 , n419530 );
buf ( n419532 , n419531 );
nand ( n419533 , n419527 , n419532 );
and ( n419534 , n419533 , n364389 );
buf ( n419535 , n364154 );
buf ( n419536 , n364386 );
or ( n419537 , n419535 , n419536 );
buf ( n419538 , n419537 );
not ( n419539 , n419538 );
nor ( n419540 , n419534 , n419539 );
not ( n419541 , n44541 );
nor ( n419542 , n419541 , n364643 );
or ( n419543 , n364722 , n44560 );
nand ( n419544 , n419542 , n419543 );
or ( n419545 , n419540 , n419544 );
buf ( n419546 , n364539 );
not ( n419547 , n419546 );
buf ( n419548 , n419547 );
buf ( n419549 , n419548 );
buf ( n419550 , n44368 );
not ( n419551 , n419550 );
buf ( n419552 , n419551 );
buf ( n419553 , n419552 );
nand ( n419554 , n419549 , n419553 );
buf ( n419555 , n419554 );
buf ( n419556 , n364642 );
not ( n419557 , n419556 );
buf ( n419558 , n419557 );
or ( n419559 , n419555 , n419558 );
buf ( n419560 , n364634 );
buf ( n419561 , n44474 );
or ( n419562 , n419560 , n419561 );
buf ( n419563 , n419562 );
nand ( n419564 , n419559 , n419563 );
not ( n419565 , n419564 );
not ( n419566 , n44541 );
or ( n419567 , n419565 , n419566 );
buf ( n419568 , n44540 );
buf ( n419569 , n364649 );
or ( n419570 , n419568 , n419569 );
buf ( n419571 , n419570 );
nand ( n419572 , n419567 , n419571 );
and ( n419573 , n419572 , n419543 );
buf ( n419574 , n44560 );
buf ( n419575 , n364722 );
nand ( n419576 , n419574 , n419575 );
buf ( n419577 , n419576 );
not ( n419578 , n419577 );
nor ( n419579 , n419573 , n419578 );
nand ( n419580 , n419545 , n419579 );
buf ( n419581 , n419580 );
not ( n419582 , n419581 );
buf ( n419583 , n419582 );
nand ( n419584 , n419517 , n419583 );
buf ( n419585 , n419584 );
buf ( n419586 , n419585 );
not ( n419587 , n419586 );
or ( n419588 , n361494 , n419587 );
buf ( n419589 , n361486 );
not ( n419590 , n419589 );
buf ( n419591 , n361411 );
buf ( n419592 , n361378 );
nand ( n419593 , n419591 , n419592 );
buf ( n419594 , n419593 );
buf ( n419595 , n419594 );
buf ( n419596 , n41313 );
or ( n419597 , n419595 , n419596 );
buf ( n419598 , n41304 );
buf ( n419599 , n361449 );
nand ( n419600 , n419598 , n419599 );
buf ( n419601 , n419600 );
buf ( n419602 , n419601 );
nand ( n419603 , n419597 , n419602 );
buf ( n419604 , n419603 );
buf ( n419605 , n419604 );
not ( n419606 , n419605 );
or ( n419607 , n419590 , n419606 );
or ( n419608 , n361479 , n361483 );
buf ( n419609 , n419608 );
nand ( n419610 , n419607 , n419609 );
buf ( n419611 , n419610 );
buf ( n419612 , n419611 );
not ( n419613 , n419612 );
buf ( n419614 , n419613 );
buf ( n419615 , n419614 );
nand ( n419616 , n419588 , n419615 );
buf ( n419617 , n419616 );
buf ( n419618 , n419617 );
and ( n419619 , n419618 , n360796 );
not ( n419620 , n419618 );
and ( n419621 , n419620 , n360792 );
nor ( n419622 , n419619 , n419621 );
buf ( n419623 , n419622 );
buf ( n419624 , n364642 );
buf ( n419625 , n419563 );
nand ( n419626 , n419624 , n419625 );
buf ( n419627 , n419626 );
buf ( n419628 , n419627 );
buf ( n419629 , n419627 );
not ( n419630 , n419629 );
buf ( n419631 , n419630 );
buf ( n419632 , n419631 );
not ( n419633 , n364542 );
not ( n419634 , n364390 );
not ( n419635 , n419514 );
or ( n419636 , n419634 , n419635 );
buf ( n419637 , n419540 );
buf ( n419638 , n419637 );
nand ( n419639 , n419636 , n419638 );
not ( n419640 , n419639 );
or ( n419641 , n419633 , n419640 );
buf ( n419642 , n419555 );
buf ( n419643 , n419642 );
buf ( n419644 , n419643 );
nand ( n419645 , n419641 , n419644 );
buf ( n419646 , n419645 );
and ( n419647 , n419646 , n419632 );
not ( n419648 , n419646 );
and ( n419649 , n419648 , n419628 );
nor ( n419650 , n419647 , n419649 );
buf ( n419651 , n419650 );
buf ( n419652 , n419577 );
buf ( n419653 , n364726 );
nand ( n419654 , n419652 , n419653 );
buf ( n419655 , n419654 );
buf ( n419656 , n419655 );
buf ( n419657 , n419655 );
not ( n419658 , n419657 );
buf ( n419659 , n419658 );
buf ( n419660 , n419659 );
not ( n419661 , n419542 );
not ( n419662 , n419639 );
or ( n419663 , n419661 , n419662 );
buf ( n419664 , n419572 );
not ( n419665 , n419664 );
buf ( n419666 , n419665 );
nand ( n419667 , n419663 , n419666 );
buf ( n419668 , n419667 );
and ( n419669 , n419668 , n419660 );
not ( n419670 , n419668 );
and ( n419671 , n419670 , n419656 );
nor ( n419672 , n419669 , n419671 );
buf ( n419673 , n419672 );
buf ( n419674 , n361489 );
not ( n419675 , n419674 );
buf ( n419676 , n419608 );
nand ( n419677 , n419675 , n419676 );
buf ( n419678 , n419677 );
buf ( n419679 , n419678 );
buf ( n419680 , n419678 );
not ( n419681 , n419680 );
buf ( n419682 , n419681 );
buf ( n419683 , n419682 );
buf ( n419684 , n361458 );
not ( n419685 , n419684 );
buf ( n419686 , n419685 );
buf ( n419687 , n419686 );
not ( n419688 , n419687 );
buf ( n419689 , n419323 );
buf ( n419690 , n419689 );
buf ( n419691 , n419690 );
buf ( n419692 , n419349 );
nand ( n419693 , n419691 , n44564 , n419692 );
nand ( n419694 , n419512 , n44564 );
and ( n419695 , n419694 , n419582 );
not ( n419696 , n393853 );
not ( n419697 , n393773 );
or ( n419698 , n419696 , n419697 );
nor ( n419699 , n55520 , n364728 );
nand ( n419700 , n419698 , n419699 );
buf ( n419701 , n419700 );
nand ( n419702 , n419693 , n419695 , n419701 );
buf ( n419703 , n419702 );
not ( n419704 , n419703 );
or ( n419705 , n419688 , n419704 );
buf ( n419706 , n419604 );
not ( n419707 , n419706 );
buf ( n419708 , n419707 );
buf ( n419709 , n419708 );
nand ( n419710 , n419705 , n419709 );
buf ( n419711 , n419710 );
buf ( n419712 , n419711 );
and ( n419713 , n419712 , n419683 );
not ( n419714 , n419712 );
and ( n419715 , n419714 , n419679 );
nor ( n419716 , n419713 , n419715 );
buf ( n419717 , n419716 );
buf ( n419718 , n361414 );
buf ( n419719 , n419594 );
nand ( n419720 , n419718 , n419719 );
buf ( n419721 , n419720 );
buf ( n419722 , n419721 );
buf ( n419723 , n419721 );
not ( n419724 , n419723 );
buf ( n419725 , n419724 );
buf ( n419726 , n419725 );
buf ( n419727 , n419585 );
and ( n419728 , n419727 , n419726 );
not ( n419729 , n419727 );
and ( n419730 , n419729 , n419722 );
nor ( n419731 , n419728 , n419730 );
buf ( n419732 , n419731 );
buf ( n419733 , n419532 );
buf ( n419734 , n364147 );
nand ( n419735 , n419733 , n419734 );
buf ( n419736 , n419735 );
buf ( n419737 , n419736 );
buf ( n419738 , n419736 );
not ( n419739 , n419738 );
buf ( n419740 , n419739 );
buf ( n419741 , n419740 );
not ( n419742 , n363918 );
not ( n419743 , n419742 );
buf ( n419744 , n419514 );
not ( n419745 , n419744 );
or ( n419746 , n419743 , n419745 );
not ( n419747 , n419525 );
nand ( n419748 , n419746 , n419747 );
buf ( n419749 , n419748 );
and ( n419750 , n419749 , n419741 );
not ( n419751 , n419749 );
and ( n419752 , n419751 , n419737 );
nor ( n419753 , n419750 , n419752 );
buf ( n419754 , n419753 );
nand ( n419755 , n363917 , n419524 );
buf ( n419756 , n419755 );
buf ( n419757 , n419755 );
not ( n419758 , n419757 );
buf ( n419759 , n419758 );
buf ( n419760 , n419759 );
buf ( n419761 , n363654 );
not ( n419762 , n419761 );
buf ( n419763 , n419744 );
not ( n419764 , n419763 );
or ( n419765 , n419762 , n419764 );
buf ( n419766 , n419522 );
nand ( n419767 , n419765 , n419766 );
buf ( n419768 , n419767 );
buf ( n419769 , n419768 );
and ( n419770 , n419769 , n419760 );
not ( n419771 , n419769 );
and ( n419772 , n419771 , n419756 );
nor ( n419773 , n419770 , n419772 );
buf ( n419774 , n419773 );
buf ( n419775 , n393637 );
not ( n419776 , n419775 );
buf ( n419777 , n391981 );
buf ( n419778 , n419777 );
nand ( n419779 , n419776 , n419778 );
buf ( n419780 , n419779 );
buf ( n419781 , n419780 );
buf ( n419782 , n419780 );
not ( n419783 , n419782 );
buf ( n419784 , n419783 );
buf ( n419785 , n419784 );
buf ( n419786 , n419341 );
not ( n419787 , n419786 );
buf ( n419788 , n419787 );
buf ( n419789 , n419788 );
not ( n419790 , n419789 );
buf ( n419791 , n419790 );
buf ( n419792 , n419791 );
not ( n419793 , n419792 );
buf ( n419794 , n419337 );
not ( n419795 , n419794 );
buf ( n419796 , n419309 );
not ( n419797 , n419796 );
buf ( n419798 , n419797 );
not ( n419799 , n419798 );
buf ( n419800 , n419298 );
not ( n419801 , n419800 );
buf ( n419802 , n419801 );
not ( n419803 , n419802 );
buf ( n419804 , n419277 );
nand ( n419805 , n419803 , n419804 );
buf ( n419806 , n418908 );
buf ( n419807 , n419201 );
buf ( n419808 , n399956 );
nand ( n419809 , n419806 , n419804 , n419807 , n419808 );
nand ( n419810 , n419807 , n419804 , n418917 );
buf ( n419811 , n419305 );
nand ( n419812 , n419805 , n419809 , n419810 , n419811 );
not ( n419813 , n419812 );
or ( n419814 , n419799 , n419813 );
buf ( n419815 , n419314 );
buf ( n419816 , n419815 );
buf ( n419817 , n419816 );
nand ( n419818 , n419814 , n419817 );
not ( n419819 , n419818 );
or ( n419820 , n419795 , n419819 );
not ( n419821 , n386196 );
not ( n419822 , n419821 );
not ( n419823 , n67103 );
not ( n419824 , n419823 );
or ( n419825 , n419822 , n419824 );
buf ( n419826 , n387093 );
nand ( n419827 , n419825 , n419826 );
buf ( n419828 , n419827 );
buf ( n419829 , n67097 );
buf ( n419830 , n419829 );
not ( n419831 , n419830 );
buf ( n419832 , n419831 );
buf ( n419833 , n419832 );
or ( n419834 , n419828 , n419833 );
buf ( n419835 , n67080 );
or ( n419836 , n419835 , n67096 );
buf ( n419837 , n419836 );
nand ( n419838 , n419834 , n419837 );
buf ( n419839 , n419838 );
and ( n419840 , n419839 , n72622 );
not ( n419841 , n67814 );
nor ( n419842 , n419841 , n67818 );
buf ( n419843 , n419842 );
buf ( n419844 , n419843 );
buf ( n419845 , n419844 );
nor ( n419846 , n419840 , n419845 );
nand ( n419847 , n419820 , n419846 );
buf ( n419848 , n419847 );
not ( n419849 , n419848 );
or ( n419850 , n419793 , n419849 );
buf ( n419851 , n69486 );
buf ( n419852 , n419851 );
nand ( n419853 , n419850 , n419852 );
buf ( n419854 , n419853 );
buf ( n419855 , n419854 );
and ( n419856 , n419855 , n419785 );
not ( n419857 , n419855 );
and ( n419858 , n419857 , n419781 );
nor ( n419859 , n419856 , n419858 );
buf ( n419860 , n419859 );
buf ( n419861 , n393615 );
not ( n419862 , n419861 );
buf ( n419863 , n390428 );
buf ( n419864 , n419863 );
nand ( n419865 , n419862 , n419864 );
buf ( n419866 , n419865 );
buf ( n419867 , n419866 );
buf ( n419868 , n419866 );
not ( n419869 , n419868 );
buf ( n419870 , n419869 );
buf ( n419871 , n419870 );
buf ( n419872 , n393626 );
not ( n419873 , n419872 );
buf ( n419874 , n419847 );
not ( n419875 , n419874 );
or ( n419876 , n419873 , n419875 );
buf ( n419877 , n389596 );
buf ( n419878 , n419877 );
buf ( n419879 , n419878 );
buf ( n419880 , n419879 );
nand ( n419881 , n419876 , n419880 );
buf ( n419882 , n419881 );
buf ( n419883 , n419882 );
and ( n419884 , n419883 , n419871 );
not ( n419885 , n419883 );
and ( n419886 , n419885 , n419867 );
nor ( n419887 , n419884 , n419886 );
buf ( n419888 , n419887 );
buf ( n419889 , n419845 );
buf ( n419890 , n72622 );
not ( n419891 , n419890 );
buf ( n419892 , n419891 );
buf ( n419893 , n419892 );
or ( n419894 , n419889 , n419893 );
buf ( n419895 , n419894 );
buf ( n419896 , n419895 );
buf ( n419897 , n419895 );
not ( n419898 , n419897 );
buf ( n419899 , n419898 );
buf ( n419900 , n419899 );
buf ( n419901 , n419829 );
not ( n419902 , n419901 );
buf ( n419903 , n419332 );
not ( n419904 , n419903 );
buf ( n419905 , n419904 );
not ( n419906 , n419905 );
buf ( n419907 , n419812 );
buf ( n419908 , n419798 );
and ( n419909 , n419907 , n419908 );
buf ( n419910 , n419909 );
buf ( n419911 , n419910 );
not ( n419912 , n419911 );
or ( n419913 , n419906 , n419912 );
buf ( n419914 , n419827 );
not ( n419915 , n419914 );
buf ( n419916 , n419903 );
buf ( n419917 , n419817 );
nor ( n419918 , n419916 , n419917 );
buf ( n419919 , n419918 );
buf ( n419920 , n419919 );
nor ( n419921 , n419915 , n419920 );
buf ( n419922 , n419921 );
buf ( n419923 , n419922 );
nand ( n419924 , n419913 , n419923 );
buf ( n419925 , n419924 );
buf ( n419926 , n419925 );
not ( n419927 , n419926 );
or ( n419928 , n419902 , n419927 );
buf ( n419929 , n419836 );
nand ( n419930 , n419928 , n419929 );
buf ( n419931 , n419930 );
buf ( n419932 , n419931 );
and ( n419933 , n419932 , n419900 );
not ( n419934 , n419932 );
and ( n419935 , n419934 , n419896 );
nor ( n419936 , n419933 , n419935 );
buf ( n419937 , n419936 );
buf ( n419938 , n72816 );
buf ( n419939 , n419938 );
buf ( n419940 , n393599 );
nand ( n419941 , n419939 , n419940 );
buf ( n419942 , n419941 );
buf ( n419943 , n419941 );
not ( n419944 , n419943 );
buf ( n419945 , n419944 );
buf ( n419946 , n419945 );
not ( n419947 , n419344 );
not ( n419948 , n419947 );
not ( n419949 , n67823 );
not ( n419950 , n419949 );
buf ( n419951 , n69486 );
buf ( n419952 , n419777 );
nand ( n419953 , n419951 , n419952 );
buf ( n419954 , n419953 );
buf ( n419955 , n419954 );
not ( n419956 , n419955 );
buf ( n419957 , n419956 );
nand ( n419958 , n419950 , n419957 );
buf ( n419959 , n419788 );
buf ( n419960 , n419892 );
nor ( n419961 , n419959 , n419960 );
buf ( n419962 , n419961 );
not ( n419963 , n419962 );
nand ( n419964 , n419957 , n419963 );
buf ( n419965 , n419342 );
buf ( n419966 , n419965 );
buf ( n419967 , n419966 );
nand ( n419968 , n419958 , n419964 , n419967 );
buf ( n419969 , n419343 );
not ( n419970 , n419279 );
not ( n419971 , n399956 );
not ( n419972 , n418908 );
or ( n419973 , n419971 , n419972 );
nand ( n419974 , n419973 , n418918 );
not ( n419975 , n419974 );
or ( n419976 , n419970 , n419975 );
not ( n419977 , n419317 );
nand ( n419978 , n419976 , n419977 );
nand ( n419979 , n419969 , n419978 );
buf ( n419980 , n391967 );
nand ( n419981 , n70221 , n419980 );
not ( n419982 , n419981 );
not ( n419983 , n419982 );
nand ( n419984 , n419968 , n419979 , n419983 );
not ( n419985 , n419984 );
or ( n419986 , n419948 , n419985 );
not ( n419987 , n393839 );
nor ( n419988 , n72789 , n393792 );
nor ( n419989 , n419987 , n419988 );
nand ( n419990 , n419986 , n419989 );
buf ( n419991 , n419990 );
and ( n419992 , n419991 , n419946 );
not ( n419993 , n419991 );
and ( n419994 , n419993 , n419942 );
nor ( n419995 , n419992 , n419994 );
buf ( n419996 , n419995 );
xor ( n419997 , n360704 , n360758 );
and ( n419998 , n419997 , n360777 );
and ( n419999 , n360704 , n360758 );
or ( n420000 , n419998 , n419999 );
buf ( n420001 , n420000 );
buf ( n420002 , n40593 );
not ( n420003 , n420002 );
buf ( n420004 , n420003 );
buf ( n420005 , n362663 );
not ( n420006 , n420005 );
buf ( n420007 , n360168 );
not ( n420008 , n420007 );
buf ( n420009 , n420008 );
buf ( n420010 , n420009 );
not ( n420011 , n420010 );
or ( n420012 , n420006 , n420011 );
buf ( n420013 , n40603 );
nand ( n420014 , n420012 , n420013 );
buf ( n420015 , n420014 );
buf ( n420016 , n39891 );
not ( n420017 , n420016 );
buf ( n420018 , n359950 );
not ( n420019 , n420018 );
buf ( n420020 , n40092 );
not ( n420021 , n420020 );
or ( n420022 , n420019 , n420021 );
buf ( n420023 , n40093 );
buf ( n420024 , n359955 );
nand ( n420025 , n420023 , n420024 );
buf ( n420026 , n420025 );
buf ( n420027 , n420026 );
nand ( n420028 , n420022 , n420027 );
buf ( n420029 , n420028 );
buf ( n420030 , n420029 );
not ( n420031 , n420030 );
or ( n420032 , n420017 , n420031 );
buf ( n420033 , n360716 );
buf ( n420034 , n359919 );
nand ( n420035 , n420033 , n420034 );
buf ( n420036 , n420035 );
buf ( n420037 , n420036 );
nand ( n420038 , n420032 , n420037 );
buf ( n420039 , n420038 );
xor ( n420040 , n420015 , n420039 );
buf ( n420041 , n359815 );
not ( n420042 , n420041 );
buf ( n420043 , n360747 );
not ( n420044 , n420043 );
or ( n420045 , n420042 , n420044 );
buf ( n420046 , n359720 );
not ( n420047 , n420046 );
buf ( n420048 , n360138 );
not ( n420049 , n420048 );
or ( n420050 , n420047 , n420049 );
not ( n420051 , n360138 );
nand ( n420052 , n420051 , n359789 );
buf ( n420053 , n420052 );
nand ( n420054 , n420050 , n420053 );
buf ( n420055 , n420054 );
buf ( n420056 , n420055 );
buf ( n420057 , n39592 );
nand ( n420058 , n420056 , n420057 );
buf ( n420059 , n420058 );
buf ( n420060 , n420059 );
nand ( n420061 , n420045 , n420060 );
buf ( n420062 , n420061 );
xor ( n420063 , n420040 , n420062 );
xor ( n420064 , n420004 , n420063 );
xor ( n420065 , n360720 , n40611 );
and ( n420066 , n420065 , n360755 );
and ( n420067 , n360720 , n40611 );
or ( n420068 , n420066 , n420067 );
buf ( n420069 , n420068 );
xor ( n420070 , n420064 , n420069 );
nor ( n420071 , n420001 , n420070 );
not ( n420072 , n420071 );
buf ( n420073 , n420072 );
nand ( n420074 , n420001 , n420070 );
buf ( n420075 , n420074 );
nand ( n420076 , n420073 , n420075 );
buf ( n420077 , n420076 );
buf ( n420078 , n420077 );
buf ( n420079 , n420077 );
not ( n420080 , n420079 );
buf ( n420081 , n420080 );
buf ( n420082 , n420081 );
and ( n420083 , n361492 , n360788 );
buf ( n420084 , n420083 );
buf ( n420085 , n420084 );
not ( n420086 , n420085 );
buf ( n420087 , n419700 );
buf ( n420088 , n419694 );
buf ( n420089 , n419582 );
and ( n420090 , n420087 , n420088 , n420089 );
buf ( n420091 , n420090 );
buf ( n420092 , n420091 );
not ( n420093 , n420092 );
buf ( n420094 , n420093 );
buf ( n420095 , n420094 );
not ( n420096 , n420095 );
or ( n420097 , n420086 , n420096 );
nand ( n420098 , n44564 , n420084 );
not ( n420099 , n420098 );
and ( n420100 , n420099 , n419691 , n419692 );
buf ( n420101 , n360788 );
not ( n420102 , n420101 );
buf ( n420103 , n419611 );
not ( n420104 , n420103 );
or ( n420105 , n420102 , n420104 );
buf ( n420106 , n360782 );
nand ( n420107 , n420105 , n420106 );
buf ( n420108 , n420107 );
nor ( n420109 , n420100 , n420108 );
buf ( n420110 , n420109 );
nand ( n420111 , n420097 , n420110 );
buf ( n420112 , n420111 );
buf ( n420113 , n420112 );
and ( n420114 , n420113 , n420082 );
not ( n420115 , n420113 );
and ( n420116 , n420115 , n420078 );
nor ( n420117 , n420114 , n420116 );
buf ( n420118 , n420117 );
buf ( n420119 , n393791 );
not ( n420120 , n420119 );
buf ( n420121 , n393710 );
buf ( n420122 , n420121 );
nand ( n420123 , n420120 , n420122 );
buf ( n420124 , n420123 );
buf ( n420125 , n420124 );
buf ( n420126 , n420124 );
not ( n420127 , n420126 );
buf ( n420128 , n420127 );
buf ( n420129 , n420128 );
buf ( n420130 , n72772 );
not ( n420131 , n420130 );
not ( n420132 , n419969 );
not ( n420133 , n419978 );
or ( n420134 , n420132 , n420133 );
and ( n420135 , n419958 , n419964 , n419967 );
nor ( n420136 , n420135 , n419982 );
nand ( n420137 , n420134 , n420136 );
nand ( n420138 , n420137 , n72761 );
nand ( n420139 , n420131 , n420138 );
buf ( n420140 , n420139 );
and ( n420141 , n420140 , n420129 );
not ( n420142 , n420140 );
and ( n420143 , n420142 , n420125 );
nor ( n420144 , n420141 , n420143 );
buf ( n420145 , n420144 );
buf ( n420146 , n393839 );
buf ( n420147 , n72477 );
buf ( n420148 , n420147 );
nand ( n420149 , n420146 , n420148 );
buf ( n420150 , n420149 );
buf ( n420151 , n420150 );
buf ( n420152 , n420150 );
not ( n420153 , n420152 );
buf ( n420154 , n420153 );
buf ( n420155 , n420154 );
buf ( n420156 , n72761 );
buf ( n420157 , n420121 );
and ( n420158 , n420156 , n420157 );
buf ( n420159 , n420158 );
not ( n420160 , n420159 );
not ( n420161 , n420137 );
or ( n420162 , n420160 , n420161 );
buf ( n420163 , n420130 );
buf ( n420164 , n420121 );
and ( n420165 , n420163 , n420164 );
buf ( n420166 , n393791 );
nor ( n420167 , n420165 , n420166 );
buf ( n420168 , n420167 );
nand ( n420169 , n420162 , n420168 );
buf ( n420170 , n420169 );
and ( n420171 , n420170 , n420155 );
not ( n420172 , n420170 );
and ( n420173 , n420172 , n420151 );
nor ( n420174 , n420171 , n420173 );
buf ( n420175 , n420174 );
buf ( n420176 , n419408 );
not ( n420177 , n420176 );
buf ( n420178 , n420177 );
buf ( n420179 , n420178 );
buf ( n420180 , n372000 );
buf ( n420181 , n420180 );
nand ( n420182 , n420179 , n420181 );
buf ( n420183 , n420182 );
buf ( n420184 , n420183 );
buf ( n420185 , n420183 );
not ( n420186 , n420185 );
buf ( n420187 , n420186 );
buf ( n420188 , n420187 );
not ( n420189 , n49930 );
nand ( n420190 , n419349 , n419978 );
not ( n420191 , n393854 );
nand ( n420192 , n420190 , n420191 );
buf ( n420193 , n420192 );
not ( n420194 , n420193 );
or ( n420195 , n420189 , n420194 );
buf ( n420196 , n419418 );
nand ( n420197 , n420195 , n420196 );
buf ( n420198 , n420197 );
and ( n420199 , n420198 , n420188 );
not ( n420200 , n420198 );
and ( n420201 , n420200 , n420184 );
nor ( n420202 , n420199 , n420201 );
buf ( n420203 , n420202 );
not ( n420204 , n371974 );
buf ( n420205 , n419428 );
not ( n420206 , n420205 );
buf ( n420207 , n420206 );
nand ( n420208 , n420204 , n420207 );
buf ( n420209 , n420208 );
buf ( n420210 , n420208 );
not ( n420211 , n420210 );
buf ( n420212 , n420211 );
buf ( n420213 , n420212 );
and ( n420214 , n49930 , n371378 , n372000 );
buf ( n420215 , n420214 );
not ( n420216 , n420215 );
buf ( n420217 , n420193 );
not ( n420218 , n420217 );
or ( n420219 , n420216 , n420218 );
not ( n420220 , n372000 );
not ( n420221 , n419419 );
or ( n420222 , n420220 , n420221 );
nand ( n420223 , n420222 , n420178 );
buf ( n420224 , n420223 );
buf ( n420225 , n371378 );
buf ( n420226 , n420225 );
and ( n420227 , n420224 , n420226 );
buf ( n420228 , n371330 );
buf ( n420229 , n420228 );
buf ( n420230 , n371372 );
and ( n420231 , n420229 , n420230 );
buf ( n420232 , n420231 );
buf ( n420233 , n420232 );
nor ( n420234 , n420227 , n420233 );
buf ( n420235 , n420234 );
buf ( n420236 , n420235 );
nand ( n420237 , n420219 , n420236 );
buf ( n420238 , n420237 );
buf ( n420239 , n420238 );
and ( n420240 , n420239 , n420213 );
not ( n420241 , n420239 );
and ( n420242 , n420241 , n420209 );
nor ( n420243 , n420240 , n420242 );
buf ( n420244 , n420243 );
buf ( n420245 , n419154 );
buf ( n420246 , n419297 );
nand ( n420247 , n420245 , n420246 );
buf ( n420248 , n420247 );
buf ( n420249 , n420248 );
buf ( n420250 , n420248 );
not ( n420251 , n420250 );
buf ( n420252 , n420251 );
buf ( n420253 , n420252 );
buf ( n420254 , n419179 );
buf ( n420255 , n420254 );
not ( n420256 , n420255 );
not ( n420257 , n419200 );
buf ( n420258 , n399956 );
not ( n420259 , n420258 );
buf ( n420260 , n418908 );
buf ( n420261 , n420260 );
not ( n420262 , n420261 );
or ( n420263 , n420259 , n420262 );
buf ( n420264 , n418918 );
nand ( n420265 , n420263 , n420264 );
buf ( n420266 , n420265 );
not ( n420267 , n420266 );
or ( n420268 , n420257 , n420267 );
buf ( n420269 , n419284 );
buf ( n420270 , n420269 );
not ( n420271 , n420270 );
nand ( n420272 , n420268 , n420271 );
buf ( n420273 , n420272 );
not ( n420274 , n420273 );
or ( n420275 , n420256 , n420274 );
buf ( n420276 , n419291 );
nand ( n420277 , n420275 , n420276 );
buf ( n420278 , n420277 );
buf ( n420279 , n420278 );
and ( n420280 , n420279 , n420253 );
not ( n420281 , n420279 );
and ( n420282 , n420281 , n420249 );
nor ( n420283 , n420280 , n420282 );
buf ( n420284 , n420283 );
buf ( n420285 , n419823 );
buf ( n420286 , n419826 );
nand ( n420287 , n420285 , n420286 );
buf ( n420288 , n420287 );
buf ( n420289 , n420288 );
buf ( n420290 , n420288 );
not ( n420291 , n420290 );
buf ( n420292 , n420291 );
buf ( n420293 , n420292 );
buf ( n420294 , n419331 );
not ( n420295 , n420294 );
buf ( n420296 , n419978 );
not ( n420297 , n420296 );
or ( n420298 , n420295 , n420297 );
nand ( n420299 , n420298 , n419821 );
buf ( n420300 , n420299 );
and ( n420301 , n420300 , n420293 );
not ( n420302 , n420300 );
and ( n420303 , n420302 , n420289 );
nor ( n420304 , n420301 , n420303 );
buf ( n420305 , n420304 );
nand ( n420306 , n420294 , n419821 );
buf ( n420307 , n420306 );
buf ( n420308 , n420296 );
buf ( n420309 , n420306 );
buf ( n420310 , n420296 );
not ( n420311 , n420307 );
not ( n420312 , n420308 );
or ( n420313 , n420311 , n420312 );
or ( n420314 , n420309 , n420310 );
nand ( n420315 , n420313 , n420314 );
buf ( n420316 , n420315 );
buf ( n420317 , n419291 );
buf ( n420318 , n420254 );
nand ( n420319 , n420317 , n420318 );
buf ( n420320 , n420319 );
buf ( n420321 , n420320 );
buf ( n420322 , n420320 );
not ( n420323 , n420322 );
buf ( n420324 , n420323 );
buf ( n420325 , n420324 );
buf ( n420326 , n420272 );
and ( n420327 , n420326 , n420325 );
not ( n420328 , n420326 );
and ( n420329 , n420328 , n420321 );
nor ( n420330 , n420327 , n420329 );
buf ( n420331 , n420330 );
nand ( n420332 , n420271 , n419200 );
buf ( n420333 , n420332 );
buf ( n420334 , n420332 );
not ( n420335 , n420334 );
buf ( n420336 , n420335 );
buf ( n420337 , n420336 );
buf ( n420338 , n420266 );
and ( n420339 , n420338 , n420337 );
not ( n420340 , n420338 );
and ( n420341 , n420340 , n420333 );
nor ( n420342 , n420339 , n420341 );
buf ( n420343 , n420342 );
buf ( n420344 , n418916 );
buf ( n420345 , n399955 );
nand ( n420346 , n420344 , n420345 );
buf ( n420347 , n420346 );
buf ( n420348 , n420347 );
buf ( n420349 , n420347 );
not ( n420350 , n420349 );
buf ( n420351 , n420350 );
buf ( n420352 , n420351 );
not ( n420353 , n78445 );
not ( n420354 , n420260 );
or ( n420355 , n420353 , n420354 );
nand ( n420356 , n420355 , n418912 );
buf ( n420357 , n420356 );
and ( n420358 , n420357 , n420352 );
not ( n420359 , n420357 );
and ( n420360 , n420359 , n420348 );
nor ( n420361 , n420358 , n420360 );
buf ( n420362 , n420361 );
buf ( n420363 , n418900 );
buf ( n420364 , n418841 );
nand ( n420365 , n420363 , n420364 );
buf ( n420366 , n420365 );
buf ( n420367 , n420366 );
buf ( n420368 , n420366 );
not ( n420369 , n420368 );
buf ( n420370 , n420369 );
buf ( n420371 , n420370 );
buf ( n420372 , n418868 );
not ( n420373 , n420372 );
buf ( n420374 , n82759 );
not ( n420375 , n420374 );
buf ( n420376 , n418782 );
buf ( n420377 , n420376 );
buf ( n420378 , n420377 );
buf ( n420379 , n420378 );
not ( n420380 , n420379 );
or ( n420381 , n420375 , n420380 );
not ( n420382 , n418889 );
nor ( n420383 , n420382 , n418891 );
buf ( n420384 , n420383 );
nand ( n420385 , n420381 , n420384 );
buf ( n420386 , n420385 );
buf ( n420387 , n420386 );
not ( n420388 , n420387 );
or ( n420389 , n420373 , n420388 );
buf ( n420390 , n418896 );
nand ( n420391 , n420389 , n420390 );
buf ( n420392 , n420391 );
buf ( n420393 , n420392 );
and ( n420394 , n420393 , n420371 );
not ( n420395 , n420393 );
and ( n420396 , n420395 , n420367 );
nor ( n420397 , n420394 , n420396 );
buf ( n420398 , n420397 );
buf ( n420399 , n418896 );
buf ( n420400 , n418868 );
nand ( n420401 , n420399 , n420400 );
buf ( n420402 , n420401 );
buf ( n420403 , n420402 );
buf ( n420404 , n420402 );
not ( n420405 , n420404 );
buf ( n420406 , n420405 );
buf ( n420407 , n420406 );
buf ( n420408 , n420386 );
and ( n420409 , n420408 , n420407 );
not ( n420410 , n420408 );
and ( n420411 , n420410 , n420403 );
nor ( n420412 , n420409 , n420411 );
buf ( n420413 , n420412 );
not ( n420414 , n418891 );
nand ( n420415 , n420414 , n82756 );
buf ( n420416 , n420415 );
buf ( n420417 , n420415 );
not ( n420418 , n420417 );
buf ( n420419 , n420418 );
buf ( n420420 , n420419 );
buf ( n420421 , n404440 );
not ( n420422 , n420421 );
buf ( n420423 , n420378 );
not ( n420424 , n420423 );
or ( n420425 , n420422 , n420424 );
buf ( n420426 , n418884 );
buf ( n420427 , n403321 );
buf ( n420428 , n420427 );
nand ( n420429 , n420426 , n420428 );
buf ( n420430 , n420429 );
buf ( n420431 , n420430 );
nand ( n420432 , n420425 , n420431 );
buf ( n420433 , n420432 );
buf ( n420434 , n420433 );
and ( n420435 , n420434 , n420420 );
not ( n420436 , n420434 );
and ( n420437 , n420436 , n420416 );
nor ( n420438 , n420435 , n420437 );
buf ( n420439 , n420438 );
buf ( n420440 , n420427 );
buf ( n420441 , n418873 );
nand ( n420442 , n420440 , n420441 );
buf ( n420443 , n420442 );
buf ( n420444 , n420443 );
buf ( n420445 , n420443 );
not ( n420446 , n420445 );
buf ( n420447 , n420446 );
buf ( n420448 , n420447 );
buf ( n420449 , n82678 );
not ( n420450 , n420449 );
buf ( n420451 , n420378 );
not ( n420452 , n420451 );
or ( n420453 , n420450 , n420452 );
buf ( n420454 , n418881 );
buf ( n420455 , n420454 );
buf ( n420456 , n420455 );
buf ( n420457 , n420456 );
nand ( n420458 , n420453 , n420457 );
buf ( n420459 , n420458 );
buf ( n420460 , n420459 );
and ( n420461 , n420460 , n420448 );
not ( n420462 , n420460 );
and ( n420463 , n420462 , n420444 );
nor ( n420464 , n420461 , n420463 );
buf ( n420465 , n420464 );
buf ( n420466 , n420456 );
buf ( n420467 , n82678 );
nand ( n420468 , n420466 , n420467 );
buf ( n420469 , n420468 );
buf ( n420470 , n420469 );
buf ( n420471 , n420469 );
not ( n420472 , n420471 );
buf ( n420473 , n420472 );
buf ( n420474 , n420473 );
buf ( n420475 , n420378 );
and ( n420476 , n420475 , n420474 );
not ( n420477 , n420475 );
and ( n420478 , n420477 , n420470 );
nor ( n420479 , n420476 , n420478 );
buf ( n420480 , n420479 );
nand ( n420481 , n418776 , n405685 );
buf ( n420482 , n420481 );
buf ( n420483 , n420481 );
not ( n420484 , n420483 );
buf ( n420485 , n420484 );
buf ( n420486 , n420485 );
not ( n420487 , n405661 );
not ( n420488 , n418763 );
or ( n420489 , n420487 , n420488 );
not ( n420490 , n418771 );
nand ( n420491 , n420489 , n420490 );
buf ( n420492 , n420491 );
and ( n420493 , n420492 , n420486 );
not ( n420494 , n420492 );
and ( n420495 , n420494 , n420482 );
nor ( n420496 , n420493 , n420495 );
buf ( n420497 , n420496 );
buf ( n420498 , n418734 );
buf ( n420499 , n418760 );
nand ( n420500 , n420498 , n420499 );
buf ( n420501 , n420500 );
buf ( n420502 , n420501 );
buf ( n420503 , n420501 );
not ( n420504 , n420503 );
buf ( n420505 , n420504 );
buf ( n420506 , n420505 );
buf ( n420507 , n418691 );
not ( n420508 , n420507 );
buf ( n420509 , n418496 );
not ( n420510 , n420509 );
buf ( n420511 , n418528 );
not ( n420512 , n420511 );
buf ( n420513 , n418292 );
not ( n420514 , n420513 );
or ( n420515 , n420512 , n420514 );
buf ( n420516 , n418536 );
nand ( n420517 , n420515 , n420516 );
buf ( n420518 , n420517 );
buf ( n420519 , n420518 );
not ( n420520 , n420519 );
or ( n420521 , n420510 , n420520 );
buf ( n420522 , n418552 );
nand ( n420523 , n420521 , n420522 );
buf ( n420524 , n420523 );
buf ( n420525 , n420524 );
not ( n420526 , n420525 );
or ( n420527 , n420508 , n420526 );
buf ( n420528 , n418754 );
not ( n420529 , n420528 );
buf ( n420530 , n420529 );
buf ( n420531 , n420530 );
nand ( n420532 , n420527 , n420531 );
buf ( n420533 , n420532 );
buf ( n420534 , n420533 );
and ( n420535 , n420534 , n420506 );
not ( n420536 , n420534 );
and ( n420537 , n420536 , n420502 );
nor ( n420538 , n420535 , n420537 );
buf ( n420539 , n420538 );
buf ( n420540 , n418664 );
buf ( n420541 , n418742 );
nand ( n420542 , n420540 , n420541 );
buf ( n420543 , n420542 );
buf ( n420544 , n420543 );
buf ( n420545 , n420543 );
not ( n420546 , n420545 );
buf ( n420547 , n420546 );
buf ( n420548 , n420547 );
buf ( n420549 , n418688 );
not ( n420550 , n420549 );
buf ( n420551 , n420524 );
not ( n420552 , n420551 );
or ( n420553 , n420550 , n420552 );
buf ( n420554 , n418747 );
nand ( n420555 , n420553 , n420554 );
buf ( n420556 , n420555 );
buf ( n420557 , n420556 );
and ( n420558 , n420557 , n420548 );
not ( n420559 , n420557 );
and ( n420560 , n420559 , n420544 );
nor ( n420561 , n420558 , n420560 );
buf ( n420562 , n420561 );
buf ( n420563 , n418688 );
buf ( n420564 , n418747 );
nand ( n420565 , n420563 , n420564 );
buf ( n420566 , n420565 );
buf ( n420567 , n420566 );
buf ( n420568 , n420524 );
buf ( n420569 , n420566 );
buf ( n420570 , n420524 );
not ( n420571 , n420567 );
not ( n420572 , n420568 );
or ( n420573 , n420571 , n420572 );
or ( n420574 , n420569 , n420570 );
nand ( n420575 , n420573 , n420574 );
buf ( n420576 , n420575 );
buf ( n420577 , n89919 );
buf ( n420578 , n418039 );
not ( n420579 , n420578 );
buf ( n420580 , n418033 );
not ( n420581 , n420580 );
or ( n420582 , n420579 , n420581 );
buf ( n420583 , n412431 );
nand ( n420584 , n420582 , n420583 );
buf ( n420585 , n420584 );
buf ( n420586 , n420585 );
buf ( n420587 , n412456 );
buf ( n420588 , n420587 );
not ( n420589 , n420577 );
not ( n420590 , n420586 );
or ( n420591 , n420589 , n420590 );
nand ( n420592 , n420591 , n420588 );
buf ( n420593 , n420592 );
xor ( n420594 , n413075 , n413079 );
xor ( n420595 , n420594 , n418029 );
buf ( n420596 , n420595 );
xor ( n420597 , n413327 , n413331 );
xor ( n420598 , n420597 , n418024 );
buf ( n420599 , n420598 );
xor ( n420600 , n413607 , n413611 );
xor ( n420601 , n420600 , n418019 );
buf ( n420602 , n420601 );
buf ( n420603 , n418528 );
buf ( n420604 , n418536 );
nand ( n420605 , n420603 , n420604 );
buf ( n420606 , n420605 );
buf ( n420607 , n418015 );
buf ( n420608 , n413898 );
nand ( n420609 , n420607 , n420608 );
buf ( n420610 , n420609 );
buf ( n420611 , n420610 );
buf ( n420612 , n418007 );
buf ( n420613 , n420612 );
buf ( n420614 , n420613 );
buf ( n420615 , n420614 );
buf ( n420616 , n420614 );
buf ( n420617 , n420610 );
not ( n420618 , n420611 );
not ( n420619 , n420615 );
or ( n420620 , n420618 , n420619 );
or ( n420621 , n420616 , n420617 );
nand ( n420622 , n420620 , n420621 );
buf ( n420623 , n420622 );
not ( n420624 , n418282 );
buf ( n420625 , n420624 );
buf ( n420626 , n410787 );
nand ( n420627 , n420625 , n420626 );
buf ( n420628 , n420627 );
buf ( n420629 , n420628 );
not ( n420630 , n420629 );
buf ( n420631 , n420630 );
buf ( n420632 , n418053 );
buf ( n420633 , n410825 );
nand ( n420634 , n420632 , n420633 );
buf ( n420635 , n420634 );
buf ( n420636 , n411278 );
buf ( n420637 , n411284 );
nand ( n420638 , n420636 , n420637 );
buf ( n420639 , n420638 );
buf ( n420640 , n420587 );
buf ( n420641 , n89919 );
nand ( n420642 , n420640 , n420641 );
buf ( n420643 , n420642 );
buf ( n420644 , n412431 );
buf ( n420645 , n418039 );
nand ( n420646 , n420644 , n420645 );
buf ( n420647 , n420646 );
buf ( n420648 , n417896 );
buf ( n420649 , n417899 );
buf ( n420650 , n417962 );
not ( n420651 , n420650 );
buf ( n420652 , n417968 );
nand ( n420653 , n420651 , n420652 );
buf ( n420654 , n420653 );
buf ( n420655 , n420654 );
and ( n420656 , n420655 , n420649 );
not ( n420657 , n420655 );
and ( n420658 , n420657 , n420648 );
nor ( n420659 , n420656 , n420658 );
buf ( n420660 , n420659 );
buf ( n420661 , n419829 );
buf ( n420662 , n419836 );
nand ( n420663 , n420661 , n420662 );
buf ( n420664 , n420663 );
buf ( n420665 , n415079 );
buf ( n420666 , n418001 );
nand ( n420667 , n420665 , n420666 );
buf ( n420668 , n420667 );
buf ( n420669 , n393626 );
buf ( n420670 , n419879 );
nand ( n420671 , n420669 , n420670 );
buf ( n420672 , n420671 );
buf ( n420673 , n420672 );
not ( n420674 , n420673 );
buf ( n420675 , n420674 );
buf ( n420676 , n93182 );
buf ( n420677 , n415817 );
buf ( n420678 , n417893 );
not ( n420679 , n420676 );
not ( n420680 , n420677 );
or ( n420681 , n420679 , n420680 );
nand ( n420682 , n420681 , n420678 );
buf ( n420683 , n420682 );
buf ( n420684 , n417884 );
buf ( n420685 , n415945 );
nand ( n420686 , n420684 , n420685 );
buf ( n420687 , n420686 );
buf ( n420688 , n95053 );
buf ( n420689 , n417866 );
buf ( n420690 , n416311 );
nand ( n420691 , n420689 , n420690 );
buf ( n420692 , n420691 );
buf ( n420693 , n420692 );
buf ( n420694 , n420692 );
buf ( n420695 , n95053 );
not ( n420696 , n420688 );
not ( n420697 , n420693 );
or ( n420698 , n420696 , n420697 );
or ( n420699 , n420694 , n420695 );
nand ( n420700 , n420698 , n420699 );
buf ( n420701 , n420700 );
buf ( n420702 , n95019 );
buf ( n420703 , n417858 );
buf ( n420704 , n417852 );
nand ( n420705 , n420703 , n420704 );
buf ( n420706 , n420705 );
buf ( n420707 , n420706 );
buf ( n420708 , n420706 );
buf ( n420709 , n95019 );
not ( n420710 , n420702 );
not ( n420711 , n420707 );
or ( n420712 , n420710 , n420711 );
or ( n420713 , n420708 , n420709 );
nand ( n420714 , n420712 , n420713 );
buf ( n420715 , n420714 );
buf ( n420716 , n95018 );
buf ( n420717 , n416769 );
nand ( n420718 , n420716 , n420717 );
buf ( n420719 , n420718 );
buf ( n420720 , n420719 );
buf ( n420721 , n417817 );
buf ( n420722 , n417817 );
buf ( n420723 , n420719 );
not ( n420724 , n420720 );
not ( n420725 , n420721 );
or ( n420726 , n420724 , n420725 );
or ( n420727 , n420722 , n420723 );
nand ( n420728 , n420726 , n420727 );
buf ( n420729 , n420728 );
buf ( n420730 , n94962 );
buf ( n420731 , n417767 );
buf ( n420732 , n417808 );
not ( n420733 , n420732 );
buf ( n420734 , n417814 );
nand ( n420735 , n420733 , n420734 );
buf ( n420736 , n420735 );
buf ( n420737 , n420736 );
and ( n420738 , n420737 , n420731 );
not ( n420739 , n420737 );
and ( n420740 , n420739 , n420730 );
nor ( n420741 , n420738 , n420740 );
buf ( n420742 , n420741 );
not ( n420743 , n393774 );
buf ( n420744 , n72749 );
nand ( n420745 , n420743 , n420744 );
buf ( n420746 , n420745 );
not ( n420747 , n420746 );
buf ( n420748 , n420747 );
buf ( n420749 , n375549 );
buf ( n420750 , n420749 );
buf ( n420751 , n419439 );
buf ( n420752 , n420751 );
buf ( n420753 , n420752 );
buf ( n420754 , n420753 );
buf ( n420755 , n419469 );
not ( n420756 , n420755 );
buf ( n420757 , n420756 );
buf ( n420758 , n420757 );
not ( n420759 , n420750 );
not ( n420760 , n420754 );
or ( n420761 , n420759 , n420760 );
nand ( n420762 , n420761 , n420758 );
buf ( n420763 , n420762 );
buf ( n420764 , n72600 );
buf ( n420765 , n420764 );
buf ( n420766 , n72823 );
nand ( n420767 , n393803 , n393807 );
buf ( n420768 , n420767 );
not ( n420769 , n420765 );
not ( n420770 , n420766 );
or ( n420771 , n420769 , n420770 );
nand ( n420772 , n420771 , n420768 );
buf ( n420773 , n420772 );
buf ( n420774 , n417700 );
buf ( n420775 , n417757 );
buf ( n420776 , n417763 );
nand ( n420777 , n420775 , n420776 );
buf ( n420778 , n420777 );
buf ( n420779 , n420778 );
buf ( n420780 , n420778 );
buf ( n420781 , n417700 );
not ( n420782 , n420774 );
not ( n420783 , n420779 );
or ( n420784 , n420782 , n420783 );
or ( n420785 , n420780 , n420781 );
nand ( n420786 , n420784 , n420785 );
buf ( n420787 , n420786 );
buf ( n420788 , n393780 );
buf ( n420789 , n393768 );
buf ( n420790 , n420789 );
buf ( n420791 , n420790 );
nand ( n420792 , n420788 , n420791 );
buf ( n420793 , n420792 );
buf ( n420794 , n420793 );
not ( n420795 , n420794 );
buf ( n420796 , n420795 );
xor ( n420797 , n417197 , n417635 );
xor ( n420798 , n420797 , n417696 );
buf ( n420799 , n420798 );
nand ( n420800 , n393831 , n72808 );
buf ( n420801 , n420800 );
not ( n420802 , n420801 );
buf ( n420803 , n420802 );
buf ( n420804 , n419388 );
not ( n420805 , n420804 );
buf ( n420806 , n420805 );
buf ( n420807 , n420767 );
buf ( n420808 , n420764 );
nand ( n420809 , n420807 , n420808 );
buf ( n420810 , n420809 );
buf ( n420811 , n420810 );
not ( n420812 , n420811 );
buf ( n420813 , n420812 );
buf ( n420814 , n420223 );
not ( n420815 , n420814 );
buf ( n420816 , n420815 );
buf ( n420817 , n420196 );
buf ( n420818 , n49930 );
nand ( n420819 , n420817 , n420818 );
buf ( n420820 , n420819 );
buf ( n420821 , n417587 );
nand ( n420822 , n94817 , n94815 , n417625 );
nand ( n420823 , n94841 , n420822 );
buf ( n420824 , n420823 );
buf ( n420825 , n417587 );
buf ( n420826 , n420823 );
not ( n420827 , n420821 );
not ( n420828 , n420824 );
or ( n420829 , n420827 , n420828 );
or ( n420830 , n420825 , n420826 );
nand ( n420831 , n420829 , n420830 );
buf ( n420832 , n420831 );
not ( n420833 , n419356 );
buf ( n420834 , n420833 );
buf ( n420835 , n419375 );
nand ( n420836 , n420834 , n420835 );
buf ( n420837 , n420836 );
buf ( n420838 , n420837 );
not ( n420839 , n420838 );
buf ( n420840 , n420839 );
buf ( n420841 , n419398 );
buf ( n420842 , n374052 );
nand ( n420843 , n420841 , n420842 );
buf ( n420844 , n420843 );
buf ( n420845 , n420844 );
not ( n420846 , n420845 );
buf ( n420847 , n420846 );
buf ( n420848 , n373083 );
buf ( n420849 , n420848 );
buf ( n420850 , n420849 );
buf ( n420851 , n419365 );
buf ( n420852 , n420851 );
buf ( n420853 , n420852 );
buf ( n420854 , n419458 );
not ( n420855 , n420854 );
buf ( n420856 , n420855 );
xor ( n420857 , n417397 , n417573 );
xor ( n420858 , n420857 , n417578 );
buf ( n420859 , n420858 );
buf ( n420860 , n419464 );
buf ( n420861 , n55177 );
nand ( n420862 , n420860 , n420861 );
buf ( n420863 , n420862 );
buf ( n420864 , n420863 );
not ( n420865 , n420864 );
buf ( n420866 , n420865 );
buf ( n420867 , n375819 );
not ( n420868 , n420867 );
buf ( n420869 , n420868 );
buf ( n420870 , n419480 );
buf ( n420871 , n420870 );
buf ( n420872 , n55331 );
buf ( n420873 , n420872 );
nand ( n420874 , n420871 , n420873 );
buf ( n420875 , n420874 );
buf ( n420876 , n420875 );
not ( n420877 , n420876 );
buf ( n420878 , n420877 );
buf ( n420879 , n419497 );
buf ( n420880 , n375801 );
nand ( n420881 , n420879 , n420880 );
buf ( n420882 , n420881 );
buf ( n420883 , n419522 );
buf ( n420884 , n363654 );
nand ( n420885 , n420883 , n420884 );
buf ( n420886 , n420885 );
buf ( n420887 , n420108 );
buf ( n420888 , n359919 );
not ( n420889 , n420888 );
buf ( n420890 , n420029 );
not ( n420891 , n420890 );
or ( n420892 , n420889 , n420891 );
buf ( n420893 , n359950 );
not ( n420894 , n420893 );
buf ( n420895 , n359147 );
not ( n420896 , n420895 );
or ( n420897 , n420894 , n420896 );
buf ( n420898 , n360624 );
buf ( n420899 , n359955 );
nand ( n420900 , n420898 , n420899 );
buf ( n420901 , n420900 );
buf ( n420902 , n420901 );
nand ( n420903 , n420897 , n420902 );
buf ( n420904 , n420903 );
buf ( n420905 , n420904 );
buf ( n420906 , n39891 );
nand ( n420907 , n420905 , n420906 );
buf ( n420908 , n420907 );
buf ( n420909 , n420908 );
nand ( n420910 , n420892 , n420909 );
buf ( n420911 , n420910 );
not ( n420912 , n420911 );
buf ( n420913 , n39592 );
buf ( n420914 , n420913 );
not ( n420915 , n420914 );
buf ( n420916 , n359720 );
not ( n420917 , n420916 );
buf ( n420918 , n360116 );
buf ( n420919 , n420918 );
not ( n420920 , n420919 );
or ( n420921 , n420917 , n420920 );
buf ( n420922 , n360122 );
buf ( n420923 , n359789 );
nand ( n420924 , n420922 , n420923 );
buf ( n420925 , n420924 );
buf ( n420926 , n420925 );
nand ( n420927 , n420921 , n420926 );
buf ( n420928 , n420927 );
buf ( n420929 , n420928 );
not ( n420930 , n420929 );
or ( n420931 , n420915 , n420930 );
buf ( n420932 , n420055 );
buf ( n420933 , n359815 );
nand ( n420934 , n420932 , n420933 );
buf ( n420935 , n420934 );
buf ( n420936 , n420935 );
nand ( n420937 , n420931 , n420936 );
buf ( n420938 , n420937 );
buf ( n420939 , n420938 );
not ( n420940 , n420939 );
buf ( n420941 , n420940 );
not ( n420942 , n420941 );
or ( n420943 , n420912 , n420942 );
not ( n420944 , n420911 );
not ( n420945 , n420944 );
not ( n420946 , n420938 );
or ( n420947 , n420945 , n420946 );
not ( n420948 , n420015 );
not ( n420949 , n420039 );
or ( n420950 , n420948 , n420949 );
or ( n420951 , n420039 , n420015 );
nand ( n420952 , n420951 , n420062 );
nand ( n420953 , n420950 , n420952 );
nand ( n420954 , n420947 , n420953 );
nand ( n420955 , n420943 , n420954 );
not ( n420956 , n420955 );
buf ( n420957 , n359996 );
not ( n420958 , n420957 );
buf ( n420959 , n359919 );
not ( n420960 , n420959 );
buf ( n420961 , n420960 );
buf ( n420962 , n420961 );
not ( n420963 , n420962 );
or ( n420964 , n420958 , n420963 );
buf ( n420965 , n420904 );
nand ( n420966 , n420964 , n420965 );
buf ( n420967 , n420966 );
buf ( n420968 , n420967 );
buf ( n420969 , n420913 );
not ( n420970 , n420969 );
and ( n420971 , n40092 , n359720 );
not ( n420972 , n40092 );
and ( n420973 , n420972 , n359789 );
or ( n420974 , n420971 , n420973 );
buf ( n420975 , n420974 );
not ( n420976 , n420975 );
or ( n420977 , n420970 , n420976 );
buf ( n420978 , n420928 );
buf ( n420979 , n359815 );
nand ( n420980 , n420978 , n420979 );
buf ( n420981 , n420980 );
buf ( n420982 , n420981 );
nand ( n420983 , n420977 , n420982 );
buf ( n420984 , n420983 );
buf ( n420985 , n420984 );
xor ( n420986 , n420968 , n420985 );
buf ( n420987 , n420941 );
xor ( n420988 , n420986 , n420987 );
buf ( n420989 , n420988 );
nand ( n420990 , n420956 , n420989 );
buf ( n420991 , n420990 );
not ( n420992 , n420991 );
not ( n420993 , n420001 );
xor ( n420994 , n420953 , n420944 );
xnor ( n420995 , n420994 , n420941 );
not ( n420996 , n420004 );
not ( n420997 , n420069 );
or ( n420998 , n420996 , n420997 );
or ( n420999 , n420069 , n420004 );
nand ( n421000 , n420999 , n420063 );
nand ( n421001 , n420998 , n421000 );
nor ( n421002 , n420995 , n421001 );
not ( n421003 , n420070 );
or ( n421004 , n420993 , n421002 , n421003 );
nand ( n421005 , n421001 , n420995 );
nand ( n421006 , n421004 , n421005 );
buf ( n421007 , n421006 );
not ( n421008 , n421007 );
or ( n421009 , n420992 , n421008 );
not ( n421010 , n420989 );
nand ( n421011 , n421010 , n420955 );
buf ( n421012 , n421011 );
nand ( n421013 , n421009 , n421012 );
buf ( n421014 , n421013 );
buf ( n421015 , n421014 );
nor ( n421016 , n420887 , n421015 );
buf ( n421017 , n421016 );
buf ( n421018 , n94763 );
buf ( n421019 , n417563 );
not ( n421020 , n421019 );
buf ( n421021 , n417569 );
nand ( n421022 , n421020 , n421021 );
buf ( n421023 , n421022 );
buf ( n421024 , n421023 );
buf ( n421025 , n94763 );
buf ( n421026 , n421023 );
not ( n421027 , n421018 );
not ( n421028 , n421024 );
or ( n421029 , n421027 , n421028 );
or ( n421030 , n421025 , n421026 );
nand ( n421031 , n421029 , n421030 );
buf ( n421032 , n421031 );
buf ( n421033 , n420108 );
not ( n421034 , n421033 );
buf ( n421035 , n421034 );
buf ( n421036 , n419644 );
buf ( n421037 , n364542 );
nand ( n421038 , n421036 , n421037 );
buf ( n421039 , n421038 );
buf ( n421040 , n417428 );
buf ( n421041 , n417423 );
nand ( n421042 , n421040 , n421041 );
buf ( n421043 , n421042 );
buf ( n421044 , n421043 );
buf ( n421045 , n417538 );
buf ( n421046 , n417538 );
buf ( n421047 , n421043 );
not ( n421048 , n421044 );
not ( n421049 , n421045 );
or ( n421050 , n421048 , n421049 );
or ( n421051 , n421046 , n421047 );
nand ( n421052 , n421050 , n421051 );
buf ( n421053 , n421052 );
buf ( n421054 , n419601 );
buf ( n421055 , n361455 );
nand ( n421056 , n421054 , n421055 );
buf ( n421057 , n421056 );
xor ( n421058 , n417439 , n94740 );
xor ( n421059 , n421058 , n417534 );
buf ( n421060 , n421059 );
buf ( n421061 , n421014 );
not ( n421062 , n421061 );
buf ( n421063 , n421062 );
buf ( n421064 , n421002 );
buf ( n421065 , n421005 );
not ( n421066 , n421064 );
nand ( n421067 , n421066 , n421065 );
buf ( n421068 , n421067 );
xor ( n421069 , n417465 , n417504 );
xor ( n421070 , n421069 , n417516 );
buf ( n421071 , n421070 );
xor ( n421072 , n417467 , n417488 );
xor ( n421073 , n421072 , n417500 );
buf ( n421074 , n421073 );
buf ( n421075 , n420967 );
buf ( n421076 , n420938 );
buf ( n421077 , n420967 );
not ( n421078 , n421077 );
buf ( n421079 , n421078 );
buf ( n421080 , n421079 );
not ( n421081 , n421080 );
buf ( n421082 , n420941 );
not ( n421083 , n421082 );
or ( n421084 , n421081 , n421083 );
buf ( n421085 , n420984 );
nand ( n421086 , n421084 , n421085 );
buf ( n421087 , n421086 );
buf ( n421088 , n421087 );
not ( n421089 , n421075 );
not ( n421090 , n421076 );
or ( n421091 , n421089 , n421090 );
nand ( n421092 , n421091 , n421088 );
buf ( n421093 , n421092 );
buf ( n421094 , n420974 );
not ( n421095 , n421094 );
buf ( n421096 , n421095 );
buf ( n421097 , n421096 );
buf ( n421098 , n39707 );
or ( n421099 , n421097 , n421098 );
buf ( n421100 , n359147 );
buf ( n421101 , n359720 );
and ( n421102 , n421100 , n421101 );
not ( n421103 , n421100 );
buf ( n421104 , n359789 );
and ( n421105 , n421103 , n421104 );
nor ( n421106 , n421102 , n421105 );
buf ( n421107 , n421106 );
buf ( n421108 , n421107 );
buf ( n421109 , n361687 );
or ( n421110 , n421108 , n421109 );
nand ( n421111 , n421099 , n421110 );
buf ( n421112 , n421111 );
buf ( n421113 , n421112 );
not ( n421114 , n421113 );
buf ( n421115 , n421114 );
buf ( n421116 , n421115 );
buf ( n421117 , n39707 );
buf ( n421118 , n361687 );
and ( n421119 , n421117 , n421118 );
buf ( n421120 , n421107 );
nor ( n421121 , n421119 , n421120 );
buf ( n421122 , n421121 );
buf ( n421123 , n421122 );
nand ( n421124 , n421116 , n421123 );
buf ( n421125 , n421124 );
buf ( n421126 , n421125 );
buf ( n421127 , n421122 );
not ( n421128 , n421127 );
buf ( n421129 , n421112 );
nand ( n421130 , n421128 , n421129 );
buf ( n421131 , n421130 );
buf ( n421132 , n421131 );
nand ( n421133 , n421126 , n421132 );
buf ( n421134 , n421133 );
buf ( n421135 , n417235 );
buf ( n421136 , C0 );
buf ( n421137 , n421136 );
xor ( n421138 , n421135 , n421137 );
buf ( n421139 , n421138 );
buf ( n421140 , n420518 );
buf ( n421141 , n418552 );
buf ( n421142 , n418496 );
nand ( n421143 , n421141 , n421142 );
buf ( n421144 , n421143 );
buf ( n421145 , n421144 );
xnor ( n421146 , n421140 , n421145 );
buf ( n421147 , n421146 );
buf ( n421148 , n418292 );
buf ( n421149 , n420606 );
xnor ( n421150 , n421148 , n421149 );
buf ( n421151 , n421150 );
buf ( n421152 , n418049 );
buf ( n421153 , n420635 );
xnor ( n421154 , n421152 , n421153 );
buf ( n421155 , n421154 );
buf ( n421156 , n419968 );
buf ( n421157 , n419981 );
and ( n421158 , n421156 , n421157 );
buf ( n421159 , n421158 );
buf ( n421160 , n420593 );
buf ( n421161 , n420639 );
xnor ( n421162 , n421160 , n421161 );
buf ( n421163 , n421162 );
buf ( n421164 , n420585 );
buf ( n421165 , n420643 );
xnor ( n421166 , n421164 , n421165 );
buf ( n421167 , n421166 );
buf ( n421168 , n418033 );
buf ( n421169 , n420647 );
xnor ( n421170 , n421168 , n421169 );
buf ( n421171 , n421170 );
buf ( n421172 , n417994 );
buf ( n421173 , n420668 );
xnor ( n421174 , n421172 , n421173 );
buf ( n421175 , n421174 );
buf ( n421176 , n417971 );
nand ( n421177 , n417991 , n417985 );
buf ( n421178 , n421177 );
xnor ( n421179 , n421176 , n421178 );
buf ( n421180 , n421179 );
buf ( n421181 , n419925 );
buf ( n421182 , n420664 );
xnor ( n421183 , n421181 , n421182 );
buf ( n421184 , n421183 );
buf ( n421185 , n417885 );
buf ( n421186 , n420683 );
xnor ( n421187 , n421185 , n421186 );
buf ( n421188 , n421187 );
buf ( n421189 , n417878 );
buf ( n421190 , n420687 );
xnor ( n421191 , n421189 , n421190 );
buf ( n421192 , n421191 );
buf ( n421193 , n420193 );
buf ( n421194 , n420820 );
xnor ( n421195 , n421193 , n421194 );
buf ( n421196 , n421195 );
buf ( n421197 , n420232 );
buf ( n421198 , n420225 );
not ( n421199 , n421197 );
nand ( n421200 , n421199 , n421198 );
buf ( n421201 , n421200 );
xnor ( n421202 , n419744 , n420886 );
buf ( n421203 , n419444 );
buf ( n421204 , n421203 );
not ( n421205 , n421204 );
buf ( n421206 , n421205 );
buf ( n421207 , n419385 );
buf ( n421208 , n373560 );
nand ( n421209 , n421207 , n421208 );
buf ( n421210 , n421209 );
buf ( n421211 , n421206 );
buf ( n421212 , n375536 );
nand ( n421213 , n421211 , n421212 );
buf ( n421214 , n421213 );
buf ( n421215 , n373563 );
buf ( n421216 , n421215 );
not ( n421217 , n421216 );
buf ( n421218 , n421217 );
buf ( n421219 , n419491 );
buf ( n421220 , n372001 );
not ( n421221 , n420083 );
not ( n421222 , n419580 );
or ( n421223 , n421221 , n421222 );
nand ( n421224 , n421223 , n421035 );
not ( n421225 , n421224 );
not ( n421226 , n419482 );
and ( n421227 , n421226 , n420872 );
not ( n421228 , n420074 );
not ( n421229 , n420099 );
not ( n421230 , n419514 );
or ( n421231 , n421229 , n421230 );
nand ( n421232 , n421231 , n421225 );
nand ( n421233 , n421232 , n420072 );
not ( n421234 , n421233 );
or ( n421235 , n421228 , n421234 );
nand ( n421236 , n421235 , n421068 );
not ( n421237 , n420072 );
not ( n421238 , n421232 );
or ( n421239 , n421237 , n421238 );
not ( n421240 , n420074 );
nor ( n421241 , n421240 , n421068 );
nand ( n421242 , n421239 , n421241 );
nand ( n421243 , n421236 , n421242 );
buf ( n421244 , n419378 );
buf ( n421245 , n421244 );
or ( n421246 , n421245 , n421210 );
buf ( n421247 , n421220 );
not ( n421248 , n421247 );
buf ( n421249 , n420192 );
not ( n421250 , n421249 );
or ( n421251 , n421248 , n421250 );
buf ( n421252 , n419424 );
and ( n421253 , n421252 , n420207 );
buf ( n421254 , n421253 );
nand ( n421255 , n421251 , n421254 );
buf ( n421256 , n421255 );
or ( n421257 , n421246 , n421256 );
not ( n421258 , n421210 );
nand ( n421259 , n420833 , n420850 );
nor ( n421260 , n421258 , n421259 );
nand ( n421261 , n421260 , n421256 );
and ( n421262 , n421210 , n421245 );
not ( n421263 , n421259 );
nor ( n421264 , n421245 , n421210 , n421263 );
nor ( n421265 , n421262 , n421264 );
nand ( n421266 , n421257 , n421261 , n421265 );
not ( n421267 , n421201 );
nand ( n421268 , n420816 , n421267 );
or ( n421269 , n421268 , n420193 );
nand ( n421270 , n49930 , n420180 );
nor ( n421271 , n421267 , n421270 );
nand ( n421272 , n421271 , n420193 );
and ( n421273 , n420816 , n421267 , n421270 );
nor ( n421274 , n420816 , n421267 );
nor ( n421275 , n421273 , n421274 );
nand ( n421276 , n421269 , n421272 , n421275 );
not ( n421277 , n420990 );
nor ( n421278 , n421277 , n421002 , n420071 );
not ( n421279 , n421093 );
nand ( n421280 , n421279 , n421112 );
nand ( n421281 , n421278 , n421280 );
nor ( n421282 , n420098 , n421281 );
not ( n421283 , n421131 );
not ( n421284 , n421134 );
not ( n421285 , n420744 );
not ( n421286 , n419969 );
not ( n421287 , n419818 );
or ( n421288 , n421286 , n421287 );
nand ( n421289 , n421288 , n421159 );
not ( n421290 , n421289 );
or ( n421291 , n421285 , n421290 );
nand ( n421292 , n421291 , n420743 );
and ( n421293 , n421292 , n420796 );
not ( n421294 , n421292 );
and ( n421295 , n421294 , n420793 );
nor ( n421296 , n421293 , n421295 );
and ( n421297 , n420137 , n420748 );
not ( n421298 , n420137 );
and ( n421299 , n421298 , n420745 );
nor ( n421300 , n421297 , n421299 );
nand ( n421301 , n419818 , n419692 , n419699 );
not ( n421302 , n421301 );
not ( n421303 , n420091 );
or ( n421304 , n421302 , n421303 );
nand ( n421305 , n421304 , n361414 );
nand ( n421306 , n421093 , n421115 );
not ( n421307 , n421306 );
buf ( n421308 , n419498 );
nand ( n421309 , n419475 , n419505 );
nor ( n421310 , n421002 , n420071 );
not ( n421311 , n421310 );
not ( n421312 , n421232 );
or ( n421313 , n421311 , n421312 );
not ( n421314 , n421002 );
not ( n421315 , n420074 );
and ( n421316 , n421314 , n421315 );
not ( n421317 , n421005 );
nor ( n421318 , n421316 , n421317 );
nand ( n421319 , n421313 , n421318 );
nand ( n421320 , n420990 , n421011 );
not ( n421321 , n421320 );
and ( n421322 , n421319 , n421321 );
not ( n421323 , n421319 );
and ( n421324 , n421323 , n421320 );
nor ( n421325 , n421322 , n421324 );
and ( n421326 , n374060 , n420749 );
not ( n421327 , n419794 );
not ( n421328 , n419978 );
or ( n421329 , n421327 , n421328 );
nand ( n421330 , n421329 , n419846 );
nand ( n421331 , n419851 , n419777 );
or ( n421332 , n421330 , n421331 );
and ( n421333 , n419788 , n419851 , n419777 );
and ( n421334 , n419777 , n393637 );
nor ( n421335 , n421333 , n421334 );
nand ( n421336 , n421332 , n421335 );
nand ( n421337 , n419981 , n393714 );
and ( n421338 , n421336 , n421337 );
not ( n421339 , n421336 );
not ( n421340 , n421337 );
and ( n421341 , n421339 , n421340 );
nor ( n421342 , n421338 , n421341 );
and ( n421343 , n421280 , n421306 );
nand ( n421344 , n421017 , n421343 );
or ( n421345 , n421344 , n419702 );
not ( n421346 , n421278 );
nand ( n421347 , n421346 , n421063 );
not ( n421348 , n421347 );
not ( n421349 , n420084 );
nor ( n421350 , n421348 , n421349 , n421343 );
nand ( n421351 , n421350 , n419702 );
not ( n421352 , n421017 );
not ( n421353 , n421349 );
or ( n421354 , n421352 , n421353 );
nand ( n421355 , n421354 , n421347 );
and ( n421356 , n421355 , n421343 );
nor ( n421357 , n421348 , n421017 , n421343 );
nor ( n421358 , n421356 , n421357 );
nand ( n421359 , n421345 , n421351 , n421358 );
nand ( n421360 , n421226 , n419488 );
not ( n421361 , n421360 );
nand ( n421362 , n421361 , n420870 );
not ( n421363 , n420870 );
and ( n421364 , n421360 , n421363 );
nor ( n421365 , n421360 , n421363 , n420872 );
nor ( n421366 , n421364 , n421365 );
buf ( n421367 , n419346 );
not ( n421368 , n421367 );
not ( n421369 , n421289 );
or ( n421370 , n421368 , n421369 );
not ( n421371 , n419989 );
not ( n421372 , n419345 );
and ( n421373 , n421371 , n421372 );
nor ( n421374 , n421373 , n420773 );
nand ( n421375 , n421370 , n421374 );
nand ( n421376 , n419347 , n393814 );
not ( n421377 , n421376 );
and ( n421378 , n421375 , n421377 );
not ( n421379 , n421375 );
and ( n421380 , n421379 , n421376 );
nor ( n421381 , n421378 , n421380 );
and ( n421382 , n421330 , n420675 );
not ( n421383 , n421330 );
and ( n421384 , n421383 , n420672 );
nor ( n421385 , n421382 , n421384 );
not ( n421386 , n420763 );
not ( n421387 , n420190 );
not ( n421388 , n420191 );
or ( n421389 , n421387 , n421388 );
nand ( n421390 , n421389 , n421326 );
nand ( n421391 , n421386 , n421390 );
or ( n421392 , n421362 , n421391 );
and ( n421393 , n421360 , n420872 );
nand ( n421394 , n421393 , n421391 );
nand ( n421395 , n421392 , n421394 , n421366 );
and ( n421396 , n421391 , n420878 );
not ( n421397 , n421391 );
and ( n421398 , n421397 , n420875 );
nor ( n421399 , n421396 , n421398 );
and ( n421400 , n72808 , n419940 );
or ( n421401 , n421219 , n420882 );
or ( n421402 , n421401 , n421391 );
and ( n421403 , n421227 , n420882 );
nand ( n421404 , n421403 , n421391 );
not ( n421405 , n421227 );
not ( n421406 , n421401 );
and ( n421407 , n421405 , n421406 );
and ( n421408 , n420882 , n421219 );
nor ( n421409 , n421407 , n421408 );
nand ( n421410 , n421402 , n421404 , n421409 );
or ( n421411 , n421308 , n421309 );
not ( n421412 , n420749 );
buf ( n421413 , n374060 );
not ( n421414 , n421413 );
and ( n421415 , n393773 , n393853 );
nand ( n421416 , n421415 , n420190 );
not ( n421417 , n421416 );
or ( n421418 , n421414 , n421417 );
buf ( n421419 , n420753 );
not ( n421420 , n421419 );
buf ( n421421 , n421420 );
nand ( n421422 , n421418 , n421421 );
not ( n421423 , n421422 );
or ( n421424 , n421412 , n421423 );
nand ( n421425 , n421424 , n420757 );
or ( n421426 , n421411 , n421425 );
and ( n421427 , n420869 , n421309 );
nand ( n421428 , n421425 , n421427 );
and ( n421429 , n421309 , n421308 );
nor ( n421430 , n421308 , n421309 , n420869 );
nor ( n421431 , n421429 , n421430 );
nand ( n421432 , n421426 , n421428 , n421431 );
not ( n421433 , n419639 );
not ( n421434 , n421039 );
or ( n421435 , n421433 , n421434 );
or ( n421436 , n421039 , n419639 );
nand ( n421437 , n421435 , n421436 );
not ( n421438 , n421282 );
not ( n421439 , n419514 );
or ( n421440 , n421438 , n421439 );
nor ( n421441 , n421278 , n421307 );
nand ( n421442 , n421063 , n421441 );
nor ( n421443 , n421224 , n421307 );
nand ( n421444 , n421443 , n421063 );
or ( n421445 , n421307 , n421280 );
nand ( n421446 , n421442 , n421444 , n421445 );
nand ( n421447 , n421440 , n421446 );
or ( n421448 , n421447 , n421283 );
nand ( n421449 , n421448 , n421125 );
buf ( n421450 , n421449 );
and ( n421451 , n421447 , n421284 );
not ( n421452 , n421447 );
and ( n421453 , n421452 , n421134 );
nor ( n421454 , n421451 , n421453 );
not ( n421455 , n419594 );
not ( n421456 , n421305 );
or ( n421457 , n421455 , n421456 );
nand ( n421458 , n421457 , n421057 );
not ( n421459 , n419594 );
nor ( n421460 , n421459 , n421057 );
nand ( n421461 , n421460 , n421305 );
nand ( n421462 , n421458 , n421461 );
not ( n421463 , n420800 );
nand ( n421464 , n421463 , n419939 );
or ( n421465 , n421464 , n419990 );
not ( n421466 , n419940 );
nor ( n421467 , n421466 , n420803 );
nand ( n421468 , n421467 , n419990 );
not ( n421469 , n420803 );
not ( n421470 , n419939 );
and ( n421471 , n421469 , n421470 );
nor ( n421472 , n420800 , n419940 );
and ( n421473 , n421472 , n419939 );
nor ( n421474 , n421471 , n421473 );
nand ( n421475 , n421465 , n421468 , n421474 );
not ( n421476 , n420810 );
buf ( n421477 , n393835 );
nand ( n421478 , n421476 , n421477 );
or ( n421479 , n421478 , n419990 );
not ( n421480 , n421400 );
nor ( n421481 , n421480 , n420813 );
nand ( n421482 , n419990 , n421481 );
not ( n421483 , n420813 );
not ( n421484 , n421477 );
and ( n421485 , n421483 , n421484 );
not ( n421486 , n421477 );
nor ( n421487 , n420810 , n421400 , n421486 );
nor ( n421488 , n421485 , n421487 );
nand ( n421489 , n421479 , n421482 , n421488 );
not ( n421490 , n44479 );
not ( n421491 , n419639 );
or ( n421492 , n421490 , n421491 );
not ( n421493 , n419564 );
nand ( n421494 , n421492 , n421493 );
nand ( n421495 , n419571 , n44541 );
not ( n421496 , n421495 );
and ( n421497 , n421494 , n421496 );
not ( n421498 , n421494 );
and ( n421499 , n421498 , n421495 );
nor ( n421500 , n421497 , n421499 );
nor ( n421501 , n55218 , n375504 );
not ( n421502 , n421501 );
not ( n421503 , n421422 );
or ( n421504 , n421502 , n421503 );
not ( n421505 , n419465 );
nand ( n421506 , n421504 , n421505 );
nand ( n421507 , n419468 , n375398 );
not ( n421508 , n421507 );
and ( n421509 , n421506 , n421508 );
not ( n421510 , n421506 );
and ( n421511 , n421510 , n421507 );
nor ( n421512 , n421509 , n421511 );
not ( n421513 , n421214 );
not ( n421514 , n421413 );
not ( n421515 , n421416 );
or ( n421516 , n421514 , n421515 );
nand ( n421517 , n421516 , n421421 );
not ( n421518 , n375536 );
not ( n421519 , n421422 );
or ( n421520 , n421518 , n421519 );
nand ( n421521 , n421520 , n421206 );
nand ( n421522 , n375547 , n419457 );
not ( n421523 , n421522 );
and ( n421524 , n421521 , n421523 );
not ( n421525 , n421521 );
and ( n421526 , n421525 , n421522 );
nor ( n421527 , n421524 , n421526 );
nand ( n421528 , n420853 , n420850 );
not ( n421529 , n421528 );
and ( n421530 , n421256 , n421529 );
not ( n421531 , n421256 );
and ( n421532 , n421531 , n421528 );
nor ( n421533 , n421530 , n421532 );
not ( n421534 , n88302 );
nand ( n421535 , n421534 , n418054 );
nand ( n421536 , n78445 , n418912 );
not ( n421537 , n421536 );
not ( n421538 , n420260 );
or ( n421539 , n421537 , n421538 );
or ( n421540 , n421536 , n420260 );
nand ( n421541 , n421539 , n421540 );
xor ( n421542 , n352287 , n352288 );
xor ( n421543 , n421542 , n32526 );
buf ( n421544 , n421543 );
not ( n421545 , n32441 );
xor ( n421546 , n351031 , n351022 );
not ( n421547 , n421546 );
or ( n421548 , n421545 , n421547 );
or ( n421549 , n421546 , n32441 );
nand ( n421550 , n421548 , n421549 );
not ( n421551 , n416158 );
not ( n421552 , n416163 );
or ( n421553 , n421551 , n421552 );
nand ( n421554 , n421553 , n417875 );
not ( n421555 , n421554 );
not ( n421556 , n417867 );
or ( n421557 , n421555 , n421556 );
or ( n421558 , n417867 , n421554 );
nand ( n421559 , n421557 , n421558 );
not ( n421560 , n418002 );
nand ( n421561 , n418006 , n91612 );
not ( n421562 , n421561 );
or ( n421563 , n421560 , n421562 );
or ( n421564 , n418002 , n421561 );
nand ( n421565 , n421563 , n421564 );
nand ( n421566 , n421535 , n420624 );
not ( n421567 , n421566 );
not ( n421568 , n418289 );
nor ( n421569 , n421568 , n418278 );
not ( n421570 , n421569 );
or ( n421571 , n421567 , n421570 );
or ( n421572 , n421569 , n421566 );
nand ( n421573 , n421571 , n421572 );
xnor ( n421574 , n351116 , n351371 );
not ( n421575 , n421574 );
not ( n421576 , n32649 );
or ( n421577 , n421575 , n421576 );
or ( n421578 , n421574 , n32649 );
nand ( n421579 , n421577 , n421578 );
buf ( n421580 , n343235 );
buf ( n421581 , n343018 );
buf ( n421582 , n342430 );
xor ( n421583 , n421581 , n421582 );
buf ( n421584 , n421583 );
buf ( n421585 , n421584 );
xor ( n421586 , n421580 , n421585 );
buf ( n421587 , n421586 );
buf ( n421588 , n352831 );
buf ( n421589 , n352671 );
xor ( n421590 , n421588 , n421589 );
buf ( n421591 , n421590 );
buf ( n421592 , n343520 );
buf ( n421593 , n343354 );
xor ( n421594 , n421592 , n421593 );
buf ( n421595 , n421594 );
xor ( n421596 , n342940 , n343257 );
xor ( n421597 , n421596 , n343261 );
buf ( n421598 , n421597 );
xor ( n421599 , n342915 , n342916 );
xor ( n421600 , n421599 , n343266 );
buf ( n421601 , n421600 );
xor ( n421602 , n342887 , n343271 );
xor ( n421603 , n421602 , n343275 );
buf ( n421604 , n421603 );
xor ( n421605 , n342860 , n342885 );
xor ( n421606 , n421605 , n343280 );
buf ( n421607 , n421606 );
xor ( n421608 , n417386 , n94698 );
xor ( n421609 , n421608 , n417583 );
buf ( n421610 , n421609 );
xor ( n421611 , n343093 , n343094 );
buf ( n421612 , n421611 );
xor ( n421613 , n343090 , n343091 );
xor ( n421614 , n421613 , n343097 );
buf ( n421615 , n421614 );
xnor ( n421616 , n351130 , n351354 );
not ( n421617 , n420844 );
nand ( n421618 , n421617 , n420806 );
or ( n421619 , n421256 , n421618 );
not ( n421620 , n421218 );
nor ( n421621 , n421620 , n420847 );
nand ( n421622 , n421256 , n421621 );
not ( n421623 , n420847 );
not ( n421624 , n420806 );
and ( n421625 , n421623 , n421624 );
nor ( n421626 , n421618 , n421218 );
nor ( n421627 , n421625 , n421626 );
nand ( n421628 , n421619 , n421622 , n421627 );
not ( n421629 , n55218 );
not ( n421630 , n43984 );
not ( n421631 , n419744 );
or ( n421632 , n421630 , n421631 );
not ( n421633 , n419533 );
nand ( n421634 , n421632 , n421633 );
nand ( n421635 , n419538 , n364389 );
not ( n421636 , n421635 );
and ( n421637 , n421634 , n421636 );
not ( n421638 , n421634 );
and ( n421639 , n421638 , n421635 );
nor ( n421640 , n421637 , n421639 );
nand ( n421641 , n419808 , n419806 , n419807 );
nand ( n421642 , n419807 , n418917 );
xor ( n421643 , n343086 , n343107 );
xor ( n421644 , n421643 , n343109 );
buf ( n421645 , n421644 );
buf ( n421646 , n421422 );
and ( n421647 , n421646 , n421513 );
not ( n421648 , n421646 );
and ( n421649 , n421648 , n421214 );
nor ( n421650 , n421647 , n421649 );
not ( n421651 , n421517 );
not ( n421652 , n420856 );
nor ( n421653 , n420863 , n421652 );
nand ( n421654 , n421651 , n421653 );
not ( n421655 , n421629 );
nor ( n421656 , n421655 , n420866 );
nand ( n421657 , n421517 , n421656 );
not ( n421658 , n420866 );
not ( n421659 , n420856 );
and ( n421660 , n421658 , n421659 );
nor ( n421661 , n420863 , n421652 , n421629 );
nor ( n421662 , n421660 , n421661 );
nand ( n421663 , n421654 , n421657 , n421662 );
not ( n421664 , n420837 );
nand ( n421665 , n421664 , n420853 );
or ( n421666 , n421256 , n421665 );
not ( n421667 , n420850 );
nor ( n421668 , n421667 , n420840 );
nand ( n421669 , n421256 , n421668 );
not ( n421670 , n420840 );
not ( n421671 , n420853 );
and ( n421672 , n421670 , n421671 );
not ( n421673 , n420853 );
nor ( n421674 , n420837 , n421673 , n420850 );
nor ( n421675 , n421672 , n421674 );
nand ( n421676 , n421666 , n421669 , n421675 );
buf ( n421677 , n420628 );
buf ( n421678 , n420631 );
buf ( n421679 , n410825 );
buf ( n421680 , n418054 );
nand ( n421681 , n421679 , n421680 );
buf ( n421682 , n421681 );
buf ( n421683 , n421682 );
and ( n421684 , n421683 , n421678 );
not ( n421685 , n421683 );
and ( n421686 , n421685 , n421677 );
nor ( n421687 , n421684 , n421686 );
buf ( n421688 , n421687 );
buf ( n421689 , n419817 );
buf ( n421690 , n419798 );
nand ( n421691 , n421689 , n421690 );
buf ( n421692 , n421691 );
buf ( n421693 , n421692 );
buf ( n421694 , n421692 );
not ( n421695 , n421694 );
buf ( n421696 , n421695 );
buf ( n421697 , n421696 );
buf ( n421698 , n419812 );
and ( n421699 , n421698 , n421697 );
not ( n421700 , n421698 );
and ( n421701 , n421700 , n421693 );
nor ( n421702 , n421699 , n421701 );
buf ( n421703 , n421702 );
nand ( n421704 , n419811 , n419804 );
not ( n421705 , n421704 );
not ( n421706 , n419803 );
nand ( n421707 , n421706 , n421641 , n421642 );
not ( n421708 , n421707 );
or ( n421709 , n421705 , n421708 );
or ( n421710 , n421704 , n421707 );
nand ( n421711 , n421709 , n421710 );
nand ( n421712 , n420490 , n405661 );
not ( n421713 , n421712 );
buf ( n421714 , n418763 );
not ( n421715 , n421714 );
or ( n421716 , n421713 , n421715 );
or ( n421717 , n421712 , n421714 );
nand ( n421718 , n421716 , n421717 );
xnor ( n421719 , n421616 , n32530 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
