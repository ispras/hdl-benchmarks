`define DC_CST_INIT 0 
`define DC_CST_LOOKUP 1 
`define DC_CST_FILL 2 
`define DC_CST_WPFILL 3 
`define DC_CST_WPWB 4 
`define DC_CST_WPDATA 5 
`define DC_CST_RPFILL 6 
`define DC_CST_RPWB 7 
`define DC_CST_RPDATA 8 
`define DC_CST_UCPROBE 9 
`define DC_CST_UCWAIT 10 
`define DC_CST_WAIT 11 
`define DC_CST_RPALGN 12 
`define DC_CST_RPDVAL 13 
`define DC_CST_QUIET 14 
`define DC_CST_MISS 15 
`define DC_CST_GNTRAM 16 
`define DC_CST_LAST 16 
`define DC_CST_CLEAR_VECT 17'd0 
`define DC_CST_RESET_VECT 17'd1 

`define DC_IST_RESET 0 
`define DC_IST_WRITE 1 
`define DC_IST_WAIT 2 
`define DC_IST_IDLE 3 
`define DC_IST_LAST 3 
`define DC_IST_CLEAR_VECT 4'd0 
`define DC_IST_RESET_VECT 4'd1 

`define IC_CST_INIT 0 
`define IC_CST_LOOKUP 1 
`define IC_CST_WB 2 
`define IC_CST_FILL 3 
`define IC_CST_UCWAIT 4 
`define IC_CST_GNTRAM 5 
`define IC_CST_LAST 5 
`define IC_CST_RESET_VECT 6'd1 

`define IC_IST_RESET 0 
`define IC_IST_WRITE 1 
`define IC_IST_WAIT 2 
`define IC_IST_IDLE 3 
`define IC_IST_LAST 3 
`define IC_IST_RESET_VECT 4'd1 
