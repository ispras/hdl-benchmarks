module mul_11_21_11(a, b, c);
  input [10:0] a;
  input [20:0] b;
  output [10:0] c;
  assign c = a * b;
endmodule
